
module first_nns_comb_W7_N256 ( q, DB, min_val_out );
  input [6:0] q;
  input [1791:0] DB;
  output [6:0] min_val_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121;

  XOR U1793 ( .A(DB[1791]), .B(n1), .Z(min_val_out[6]) );
  AND U1794 ( .A(n2), .B(n3), .Z(n1) );
  XOR U1795 ( .A(n4), .B(n5), .Z(n3) );
  XOR U1796 ( .A(DB[1791]), .B(DB[1784]), .Z(n5) );
  AND U1797 ( .A(n6), .B(n7), .Z(n4) );
  XOR U1798 ( .A(n8), .B(n9), .Z(n7) );
  XOR U1799 ( .A(DB[1784]), .B(DB[1777]), .Z(n9) );
  AND U1800 ( .A(n10), .B(n11), .Z(n8) );
  XOR U1801 ( .A(n12), .B(n13), .Z(n11) );
  XOR U1802 ( .A(DB[1777]), .B(DB[1770]), .Z(n13) );
  AND U1803 ( .A(n14), .B(n15), .Z(n12) );
  XOR U1804 ( .A(n16), .B(n17), .Z(n15) );
  XOR U1805 ( .A(DB[1770]), .B(DB[1763]), .Z(n17) );
  AND U1806 ( .A(n18), .B(n19), .Z(n16) );
  XOR U1807 ( .A(n20), .B(n21), .Z(n19) );
  XOR U1808 ( .A(DB[1763]), .B(DB[1756]), .Z(n21) );
  AND U1809 ( .A(n22), .B(n23), .Z(n20) );
  XOR U1810 ( .A(n24), .B(n25), .Z(n23) );
  XOR U1811 ( .A(DB[1756]), .B(DB[1749]), .Z(n25) );
  AND U1812 ( .A(n26), .B(n27), .Z(n24) );
  XOR U1813 ( .A(n28), .B(n29), .Z(n27) );
  XOR U1814 ( .A(DB[1749]), .B(DB[1742]), .Z(n29) );
  AND U1815 ( .A(n30), .B(n31), .Z(n28) );
  XOR U1816 ( .A(n32), .B(n33), .Z(n31) );
  XOR U1817 ( .A(DB[1742]), .B(DB[1735]), .Z(n33) );
  AND U1818 ( .A(n34), .B(n35), .Z(n32) );
  XOR U1819 ( .A(n36), .B(n37), .Z(n35) );
  XOR U1820 ( .A(DB[1735]), .B(DB[1728]), .Z(n37) );
  AND U1821 ( .A(n38), .B(n39), .Z(n36) );
  XOR U1822 ( .A(n40), .B(n41), .Z(n39) );
  XOR U1823 ( .A(DB[1728]), .B(DB[1721]), .Z(n41) );
  AND U1824 ( .A(n42), .B(n43), .Z(n40) );
  XOR U1825 ( .A(n44), .B(n45), .Z(n43) );
  XOR U1826 ( .A(DB[1721]), .B(DB[1714]), .Z(n45) );
  AND U1827 ( .A(n46), .B(n47), .Z(n44) );
  XOR U1828 ( .A(n48), .B(n49), .Z(n47) );
  XOR U1829 ( .A(DB[1714]), .B(DB[1707]), .Z(n49) );
  AND U1830 ( .A(n50), .B(n51), .Z(n48) );
  XOR U1831 ( .A(n52), .B(n53), .Z(n51) );
  XOR U1832 ( .A(DB[1707]), .B(DB[1700]), .Z(n53) );
  AND U1833 ( .A(n54), .B(n55), .Z(n52) );
  XOR U1834 ( .A(n56), .B(n57), .Z(n55) );
  XOR U1835 ( .A(DB[1700]), .B(DB[1693]), .Z(n57) );
  AND U1836 ( .A(n58), .B(n59), .Z(n56) );
  XOR U1837 ( .A(n60), .B(n61), .Z(n59) );
  XOR U1838 ( .A(DB[1693]), .B(DB[1686]), .Z(n61) );
  AND U1839 ( .A(n62), .B(n63), .Z(n60) );
  XOR U1840 ( .A(n64), .B(n65), .Z(n63) );
  XOR U1841 ( .A(DB[1686]), .B(DB[1679]), .Z(n65) );
  AND U1842 ( .A(n66), .B(n67), .Z(n64) );
  XOR U1843 ( .A(n68), .B(n69), .Z(n67) );
  XOR U1844 ( .A(DB[1679]), .B(DB[1672]), .Z(n69) );
  AND U1845 ( .A(n70), .B(n71), .Z(n68) );
  XOR U1846 ( .A(n72), .B(n73), .Z(n71) );
  XOR U1847 ( .A(DB[1672]), .B(DB[1665]), .Z(n73) );
  AND U1848 ( .A(n74), .B(n75), .Z(n72) );
  XOR U1849 ( .A(n76), .B(n77), .Z(n75) );
  XOR U1850 ( .A(DB[1665]), .B(DB[1658]), .Z(n77) );
  AND U1851 ( .A(n78), .B(n79), .Z(n76) );
  XOR U1852 ( .A(n80), .B(n81), .Z(n79) );
  XOR U1853 ( .A(DB[1658]), .B(DB[1651]), .Z(n81) );
  AND U1854 ( .A(n82), .B(n83), .Z(n80) );
  XOR U1855 ( .A(n84), .B(n85), .Z(n83) );
  XOR U1856 ( .A(DB[1651]), .B(DB[1644]), .Z(n85) );
  AND U1857 ( .A(n86), .B(n87), .Z(n84) );
  XOR U1858 ( .A(n88), .B(n89), .Z(n87) );
  XOR U1859 ( .A(DB[1644]), .B(DB[1637]), .Z(n89) );
  AND U1860 ( .A(n90), .B(n91), .Z(n88) );
  XOR U1861 ( .A(n92), .B(n93), .Z(n91) );
  XOR U1862 ( .A(DB[1637]), .B(DB[1630]), .Z(n93) );
  AND U1863 ( .A(n94), .B(n95), .Z(n92) );
  XOR U1864 ( .A(n96), .B(n97), .Z(n95) );
  XOR U1865 ( .A(DB[1630]), .B(DB[1623]), .Z(n97) );
  AND U1866 ( .A(n98), .B(n99), .Z(n96) );
  XOR U1867 ( .A(n100), .B(n101), .Z(n99) );
  XOR U1868 ( .A(DB[1623]), .B(DB[1616]), .Z(n101) );
  AND U1869 ( .A(n102), .B(n103), .Z(n100) );
  XOR U1870 ( .A(n104), .B(n105), .Z(n103) );
  XOR U1871 ( .A(DB[1616]), .B(DB[1609]), .Z(n105) );
  AND U1872 ( .A(n106), .B(n107), .Z(n104) );
  XOR U1873 ( .A(n108), .B(n109), .Z(n107) );
  XOR U1874 ( .A(DB[1609]), .B(DB[1602]), .Z(n109) );
  AND U1875 ( .A(n110), .B(n111), .Z(n108) );
  XOR U1876 ( .A(n112), .B(n113), .Z(n111) );
  XOR U1877 ( .A(DB[1602]), .B(DB[1595]), .Z(n113) );
  AND U1878 ( .A(n114), .B(n115), .Z(n112) );
  XOR U1879 ( .A(n116), .B(n117), .Z(n115) );
  XOR U1880 ( .A(DB[1595]), .B(DB[1588]), .Z(n117) );
  AND U1881 ( .A(n118), .B(n119), .Z(n116) );
  XOR U1882 ( .A(n120), .B(n121), .Z(n119) );
  XOR U1883 ( .A(DB[1588]), .B(DB[1581]), .Z(n121) );
  AND U1884 ( .A(n122), .B(n123), .Z(n120) );
  XOR U1885 ( .A(n124), .B(n125), .Z(n123) );
  XOR U1886 ( .A(DB[1581]), .B(DB[1574]), .Z(n125) );
  AND U1887 ( .A(n126), .B(n127), .Z(n124) );
  XOR U1888 ( .A(n128), .B(n129), .Z(n127) );
  XOR U1889 ( .A(DB[1574]), .B(DB[1567]), .Z(n129) );
  AND U1890 ( .A(n130), .B(n131), .Z(n128) );
  XOR U1891 ( .A(n132), .B(n133), .Z(n131) );
  XOR U1892 ( .A(DB[1567]), .B(DB[1560]), .Z(n133) );
  AND U1893 ( .A(n134), .B(n135), .Z(n132) );
  XOR U1894 ( .A(n136), .B(n137), .Z(n135) );
  XOR U1895 ( .A(DB[1560]), .B(DB[1553]), .Z(n137) );
  AND U1896 ( .A(n138), .B(n139), .Z(n136) );
  XOR U1897 ( .A(n140), .B(n141), .Z(n139) );
  XOR U1898 ( .A(DB[1553]), .B(DB[1546]), .Z(n141) );
  AND U1899 ( .A(n142), .B(n143), .Z(n140) );
  XOR U1900 ( .A(n144), .B(n145), .Z(n143) );
  XOR U1901 ( .A(DB[1546]), .B(DB[1539]), .Z(n145) );
  AND U1902 ( .A(n146), .B(n147), .Z(n144) );
  XOR U1903 ( .A(n148), .B(n149), .Z(n147) );
  XOR U1904 ( .A(DB[1539]), .B(DB[1532]), .Z(n149) );
  AND U1905 ( .A(n150), .B(n151), .Z(n148) );
  XOR U1906 ( .A(n152), .B(n153), .Z(n151) );
  XOR U1907 ( .A(DB[1532]), .B(DB[1525]), .Z(n153) );
  AND U1908 ( .A(n154), .B(n155), .Z(n152) );
  XOR U1909 ( .A(n156), .B(n157), .Z(n155) );
  XOR U1910 ( .A(DB[1525]), .B(DB[1518]), .Z(n157) );
  AND U1911 ( .A(n158), .B(n159), .Z(n156) );
  XOR U1912 ( .A(n160), .B(n161), .Z(n159) );
  XOR U1913 ( .A(DB[1518]), .B(DB[1511]), .Z(n161) );
  AND U1914 ( .A(n162), .B(n163), .Z(n160) );
  XOR U1915 ( .A(n164), .B(n165), .Z(n163) );
  XOR U1916 ( .A(DB[1511]), .B(DB[1504]), .Z(n165) );
  AND U1917 ( .A(n166), .B(n167), .Z(n164) );
  XOR U1918 ( .A(n168), .B(n169), .Z(n167) );
  XOR U1919 ( .A(DB[1504]), .B(DB[1497]), .Z(n169) );
  AND U1920 ( .A(n170), .B(n171), .Z(n168) );
  XOR U1921 ( .A(n172), .B(n173), .Z(n171) );
  XOR U1922 ( .A(DB[1497]), .B(DB[1490]), .Z(n173) );
  AND U1923 ( .A(n174), .B(n175), .Z(n172) );
  XOR U1924 ( .A(n176), .B(n177), .Z(n175) );
  XOR U1925 ( .A(DB[1490]), .B(DB[1483]), .Z(n177) );
  AND U1926 ( .A(n178), .B(n179), .Z(n176) );
  XOR U1927 ( .A(n180), .B(n181), .Z(n179) );
  XOR U1928 ( .A(DB[1483]), .B(DB[1476]), .Z(n181) );
  AND U1929 ( .A(n182), .B(n183), .Z(n180) );
  XOR U1930 ( .A(n184), .B(n185), .Z(n183) );
  XOR U1931 ( .A(DB[1476]), .B(DB[1469]), .Z(n185) );
  AND U1932 ( .A(n186), .B(n187), .Z(n184) );
  XOR U1933 ( .A(n188), .B(n189), .Z(n187) );
  XOR U1934 ( .A(DB[1469]), .B(DB[1462]), .Z(n189) );
  AND U1935 ( .A(n190), .B(n191), .Z(n188) );
  XOR U1936 ( .A(n192), .B(n193), .Z(n191) );
  XOR U1937 ( .A(DB[1462]), .B(DB[1455]), .Z(n193) );
  AND U1938 ( .A(n194), .B(n195), .Z(n192) );
  XOR U1939 ( .A(n196), .B(n197), .Z(n195) );
  XOR U1940 ( .A(DB[1455]), .B(DB[1448]), .Z(n197) );
  AND U1941 ( .A(n198), .B(n199), .Z(n196) );
  XOR U1942 ( .A(n200), .B(n201), .Z(n199) );
  XOR U1943 ( .A(DB[1448]), .B(DB[1441]), .Z(n201) );
  AND U1944 ( .A(n202), .B(n203), .Z(n200) );
  XOR U1945 ( .A(n204), .B(n205), .Z(n203) );
  XOR U1946 ( .A(DB[1441]), .B(DB[1434]), .Z(n205) );
  AND U1947 ( .A(n206), .B(n207), .Z(n204) );
  XOR U1948 ( .A(n208), .B(n209), .Z(n207) );
  XOR U1949 ( .A(DB[1434]), .B(DB[1427]), .Z(n209) );
  AND U1950 ( .A(n210), .B(n211), .Z(n208) );
  XOR U1951 ( .A(n212), .B(n213), .Z(n211) );
  XOR U1952 ( .A(DB[1427]), .B(DB[1420]), .Z(n213) );
  AND U1953 ( .A(n214), .B(n215), .Z(n212) );
  XOR U1954 ( .A(n216), .B(n217), .Z(n215) );
  XOR U1955 ( .A(DB[1420]), .B(DB[1413]), .Z(n217) );
  AND U1956 ( .A(n218), .B(n219), .Z(n216) );
  XOR U1957 ( .A(n220), .B(n221), .Z(n219) );
  XOR U1958 ( .A(DB[1413]), .B(DB[1406]), .Z(n221) );
  AND U1959 ( .A(n222), .B(n223), .Z(n220) );
  XOR U1960 ( .A(n224), .B(n225), .Z(n223) );
  XOR U1961 ( .A(DB[1406]), .B(DB[1399]), .Z(n225) );
  AND U1962 ( .A(n226), .B(n227), .Z(n224) );
  XOR U1963 ( .A(n228), .B(n229), .Z(n227) );
  XOR U1964 ( .A(DB[1399]), .B(DB[1392]), .Z(n229) );
  AND U1965 ( .A(n230), .B(n231), .Z(n228) );
  XOR U1966 ( .A(n232), .B(n233), .Z(n231) );
  XOR U1967 ( .A(DB[1392]), .B(DB[1385]), .Z(n233) );
  AND U1968 ( .A(n234), .B(n235), .Z(n232) );
  XOR U1969 ( .A(n236), .B(n237), .Z(n235) );
  XOR U1970 ( .A(DB[1385]), .B(DB[1378]), .Z(n237) );
  AND U1971 ( .A(n238), .B(n239), .Z(n236) );
  XOR U1972 ( .A(n240), .B(n241), .Z(n239) );
  XOR U1973 ( .A(DB[1378]), .B(DB[1371]), .Z(n241) );
  AND U1974 ( .A(n242), .B(n243), .Z(n240) );
  XOR U1975 ( .A(n244), .B(n245), .Z(n243) );
  XOR U1976 ( .A(DB[1371]), .B(DB[1364]), .Z(n245) );
  AND U1977 ( .A(n246), .B(n247), .Z(n244) );
  XOR U1978 ( .A(n248), .B(n249), .Z(n247) );
  XOR U1979 ( .A(DB[1364]), .B(DB[1357]), .Z(n249) );
  AND U1980 ( .A(n250), .B(n251), .Z(n248) );
  XOR U1981 ( .A(n252), .B(n253), .Z(n251) );
  XOR U1982 ( .A(DB[1357]), .B(DB[1350]), .Z(n253) );
  AND U1983 ( .A(n254), .B(n255), .Z(n252) );
  XOR U1984 ( .A(n256), .B(n257), .Z(n255) );
  XOR U1985 ( .A(DB[1350]), .B(DB[1343]), .Z(n257) );
  AND U1986 ( .A(n258), .B(n259), .Z(n256) );
  XOR U1987 ( .A(n260), .B(n261), .Z(n259) );
  XOR U1988 ( .A(DB[1343]), .B(DB[1336]), .Z(n261) );
  AND U1989 ( .A(n262), .B(n263), .Z(n260) );
  XOR U1990 ( .A(n264), .B(n265), .Z(n263) );
  XOR U1991 ( .A(DB[1336]), .B(DB[1329]), .Z(n265) );
  AND U1992 ( .A(n266), .B(n267), .Z(n264) );
  XOR U1993 ( .A(n268), .B(n269), .Z(n267) );
  XOR U1994 ( .A(DB[1329]), .B(DB[1322]), .Z(n269) );
  AND U1995 ( .A(n270), .B(n271), .Z(n268) );
  XOR U1996 ( .A(n272), .B(n273), .Z(n271) );
  XOR U1997 ( .A(DB[1322]), .B(DB[1315]), .Z(n273) );
  AND U1998 ( .A(n274), .B(n275), .Z(n272) );
  XOR U1999 ( .A(n276), .B(n277), .Z(n275) );
  XOR U2000 ( .A(DB[1315]), .B(DB[1308]), .Z(n277) );
  AND U2001 ( .A(n278), .B(n279), .Z(n276) );
  XOR U2002 ( .A(n280), .B(n281), .Z(n279) );
  XOR U2003 ( .A(DB[1308]), .B(DB[1301]), .Z(n281) );
  AND U2004 ( .A(n282), .B(n283), .Z(n280) );
  XOR U2005 ( .A(n284), .B(n285), .Z(n283) );
  XOR U2006 ( .A(DB[1301]), .B(DB[1294]), .Z(n285) );
  AND U2007 ( .A(n286), .B(n287), .Z(n284) );
  XOR U2008 ( .A(n288), .B(n289), .Z(n287) );
  XOR U2009 ( .A(DB[1294]), .B(DB[1287]), .Z(n289) );
  AND U2010 ( .A(n290), .B(n291), .Z(n288) );
  XOR U2011 ( .A(n292), .B(n293), .Z(n291) );
  XOR U2012 ( .A(DB[1287]), .B(DB[1280]), .Z(n293) );
  AND U2013 ( .A(n294), .B(n295), .Z(n292) );
  XOR U2014 ( .A(n296), .B(n297), .Z(n295) );
  XOR U2015 ( .A(DB[1280]), .B(DB[1273]), .Z(n297) );
  AND U2016 ( .A(n298), .B(n299), .Z(n296) );
  XOR U2017 ( .A(n300), .B(n301), .Z(n299) );
  XOR U2018 ( .A(DB[1273]), .B(DB[1266]), .Z(n301) );
  AND U2019 ( .A(n302), .B(n303), .Z(n300) );
  XOR U2020 ( .A(n304), .B(n305), .Z(n303) );
  XOR U2021 ( .A(DB[1266]), .B(DB[1259]), .Z(n305) );
  AND U2022 ( .A(n306), .B(n307), .Z(n304) );
  XOR U2023 ( .A(n308), .B(n309), .Z(n307) );
  XOR U2024 ( .A(DB[1259]), .B(DB[1252]), .Z(n309) );
  AND U2025 ( .A(n310), .B(n311), .Z(n308) );
  XOR U2026 ( .A(n312), .B(n313), .Z(n311) );
  XOR U2027 ( .A(DB[1252]), .B(DB[1245]), .Z(n313) );
  AND U2028 ( .A(n314), .B(n315), .Z(n312) );
  XOR U2029 ( .A(n316), .B(n317), .Z(n315) );
  XOR U2030 ( .A(DB[1245]), .B(DB[1238]), .Z(n317) );
  AND U2031 ( .A(n318), .B(n319), .Z(n316) );
  XOR U2032 ( .A(n320), .B(n321), .Z(n319) );
  XOR U2033 ( .A(DB[1238]), .B(DB[1231]), .Z(n321) );
  AND U2034 ( .A(n322), .B(n323), .Z(n320) );
  XOR U2035 ( .A(n324), .B(n325), .Z(n323) );
  XOR U2036 ( .A(DB[1231]), .B(DB[1224]), .Z(n325) );
  AND U2037 ( .A(n326), .B(n327), .Z(n324) );
  XOR U2038 ( .A(n328), .B(n329), .Z(n327) );
  XOR U2039 ( .A(DB[1224]), .B(DB[1217]), .Z(n329) );
  AND U2040 ( .A(n330), .B(n331), .Z(n328) );
  XOR U2041 ( .A(n332), .B(n333), .Z(n331) );
  XOR U2042 ( .A(DB[1217]), .B(DB[1210]), .Z(n333) );
  AND U2043 ( .A(n334), .B(n335), .Z(n332) );
  XOR U2044 ( .A(n336), .B(n337), .Z(n335) );
  XOR U2045 ( .A(DB[1210]), .B(DB[1203]), .Z(n337) );
  AND U2046 ( .A(n338), .B(n339), .Z(n336) );
  XOR U2047 ( .A(n340), .B(n341), .Z(n339) );
  XOR U2048 ( .A(DB[1203]), .B(DB[1196]), .Z(n341) );
  AND U2049 ( .A(n342), .B(n343), .Z(n340) );
  XOR U2050 ( .A(n344), .B(n345), .Z(n343) );
  XOR U2051 ( .A(DB[1196]), .B(DB[1189]), .Z(n345) );
  AND U2052 ( .A(n346), .B(n347), .Z(n344) );
  XOR U2053 ( .A(n348), .B(n349), .Z(n347) );
  XOR U2054 ( .A(DB[1189]), .B(DB[1182]), .Z(n349) );
  AND U2055 ( .A(n350), .B(n351), .Z(n348) );
  XOR U2056 ( .A(n352), .B(n353), .Z(n351) );
  XOR U2057 ( .A(DB[1182]), .B(DB[1175]), .Z(n353) );
  AND U2058 ( .A(n354), .B(n355), .Z(n352) );
  XOR U2059 ( .A(n356), .B(n357), .Z(n355) );
  XOR U2060 ( .A(DB[1175]), .B(DB[1168]), .Z(n357) );
  AND U2061 ( .A(n358), .B(n359), .Z(n356) );
  XOR U2062 ( .A(n360), .B(n361), .Z(n359) );
  XOR U2063 ( .A(DB[1168]), .B(DB[1161]), .Z(n361) );
  AND U2064 ( .A(n362), .B(n363), .Z(n360) );
  XOR U2065 ( .A(n364), .B(n365), .Z(n363) );
  XOR U2066 ( .A(DB[1161]), .B(DB[1154]), .Z(n365) );
  AND U2067 ( .A(n366), .B(n367), .Z(n364) );
  XOR U2068 ( .A(n368), .B(n369), .Z(n367) );
  XOR U2069 ( .A(DB[1154]), .B(DB[1147]), .Z(n369) );
  AND U2070 ( .A(n370), .B(n371), .Z(n368) );
  XOR U2071 ( .A(n372), .B(n373), .Z(n371) );
  XOR U2072 ( .A(DB[1147]), .B(DB[1140]), .Z(n373) );
  AND U2073 ( .A(n374), .B(n375), .Z(n372) );
  XOR U2074 ( .A(n376), .B(n377), .Z(n375) );
  XOR U2075 ( .A(DB[1140]), .B(DB[1133]), .Z(n377) );
  AND U2076 ( .A(n378), .B(n379), .Z(n376) );
  XOR U2077 ( .A(n380), .B(n381), .Z(n379) );
  XOR U2078 ( .A(DB[1133]), .B(DB[1126]), .Z(n381) );
  AND U2079 ( .A(n382), .B(n383), .Z(n380) );
  XOR U2080 ( .A(n384), .B(n385), .Z(n383) );
  XOR U2081 ( .A(DB[1126]), .B(DB[1119]), .Z(n385) );
  AND U2082 ( .A(n386), .B(n387), .Z(n384) );
  XOR U2083 ( .A(n388), .B(n389), .Z(n387) );
  XOR U2084 ( .A(DB[1119]), .B(DB[1112]), .Z(n389) );
  AND U2085 ( .A(n390), .B(n391), .Z(n388) );
  XOR U2086 ( .A(n392), .B(n393), .Z(n391) );
  XOR U2087 ( .A(DB[1112]), .B(DB[1105]), .Z(n393) );
  AND U2088 ( .A(n394), .B(n395), .Z(n392) );
  XOR U2089 ( .A(n396), .B(n397), .Z(n395) );
  XOR U2090 ( .A(DB[1105]), .B(DB[1098]), .Z(n397) );
  AND U2091 ( .A(n398), .B(n399), .Z(n396) );
  XOR U2092 ( .A(n400), .B(n401), .Z(n399) );
  XOR U2093 ( .A(DB[1098]), .B(DB[1091]), .Z(n401) );
  AND U2094 ( .A(n402), .B(n403), .Z(n400) );
  XOR U2095 ( .A(n404), .B(n405), .Z(n403) );
  XOR U2096 ( .A(DB[1091]), .B(DB[1084]), .Z(n405) );
  AND U2097 ( .A(n406), .B(n407), .Z(n404) );
  XOR U2098 ( .A(n408), .B(n409), .Z(n407) );
  XOR U2099 ( .A(DB[1084]), .B(DB[1077]), .Z(n409) );
  AND U2100 ( .A(n410), .B(n411), .Z(n408) );
  XOR U2101 ( .A(n412), .B(n413), .Z(n411) );
  XOR U2102 ( .A(DB[1077]), .B(DB[1070]), .Z(n413) );
  AND U2103 ( .A(n414), .B(n415), .Z(n412) );
  XOR U2104 ( .A(n416), .B(n417), .Z(n415) );
  XOR U2105 ( .A(DB[1070]), .B(DB[1063]), .Z(n417) );
  AND U2106 ( .A(n418), .B(n419), .Z(n416) );
  XOR U2107 ( .A(n420), .B(n421), .Z(n419) );
  XOR U2108 ( .A(DB[1063]), .B(DB[1056]), .Z(n421) );
  AND U2109 ( .A(n422), .B(n423), .Z(n420) );
  XOR U2110 ( .A(n424), .B(n425), .Z(n423) );
  XOR U2111 ( .A(DB[1056]), .B(DB[1049]), .Z(n425) );
  AND U2112 ( .A(n426), .B(n427), .Z(n424) );
  XOR U2113 ( .A(n428), .B(n429), .Z(n427) );
  XOR U2114 ( .A(DB[1049]), .B(DB[1042]), .Z(n429) );
  AND U2115 ( .A(n430), .B(n431), .Z(n428) );
  XOR U2116 ( .A(n432), .B(n433), .Z(n431) );
  XOR U2117 ( .A(DB[1042]), .B(DB[1035]), .Z(n433) );
  AND U2118 ( .A(n434), .B(n435), .Z(n432) );
  XOR U2119 ( .A(n436), .B(n437), .Z(n435) );
  XOR U2120 ( .A(DB[1035]), .B(DB[1028]), .Z(n437) );
  AND U2121 ( .A(n438), .B(n439), .Z(n436) );
  XOR U2122 ( .A(n440), .B(n441), .Z(n439) );
  XOR U2123 ( .A(DB[1028]), .B(DB[1021]), .Z(n441) );
  AND U2124 ( .A(n442), .B(n443), .Z(n440) );
  XOR U2125 ( .A(n444), .B(n445), .Z(n443) );
  XOR U2126 ( .A(DB[1021]), .B(DB[1014]), .Z(n445) );
  AND U2127 ( .A(n446), .B(n447), .Z(n444) );
  XOR U2128 ( .A(n448), .B(n449), .Z(n447) );
  XOR U2129 ( .A(DB[1014]), .B(DB[1007]), .Z(n449) );
  AND U2130 ( .A(n450), .B(n451), .Z(n448) );
  XOR U2131 ( .A(n452), .B(n453), .Z(n451) );
  XOR U2132 ( .A(DB[1007]), .B(DB[1000]), .Z(n453) );
  AND U2133 ( .A(n454), .B(n455), .Z(n452) );
  XOR U2134 ( .A(n456), .B(n457), .Z(n455) );
  XOR U2135 ( .A(DB[993]), .B(DB[1000]), .Z(n457) );
  AND U2136 ( .A(n458), .B(n459), .Z(n456) );
  XOR U2137 ( .A(n460), .B(n461), .Z(n459) );
  XOR U2138 ( .A(DB[993]), .B(DB[986]), .Z(n461) );
  AND U2139 ( .A(n462), .B(n463), .Z(n460) );
  XOR U2140 ( .A(n464), .B(n465), .Z(n463) );
  XOR U2141 ( .A(DB[986]), .B(DB[979]), .Z(n465) );
  AND U2142 ( .A(n466), .B(n467), .Z(n464) );
  XOR U2143 ( .A(n468), .B(n469), .Z(n467) );
  XOR U2144 ( .A(DB[979]), .B(DB[972]), .Z(n469) );
  AND U2145 ( .A(n470), .B(n471), .Z(n468) );
  XOR U2146 ( .A(n472), .B(n473), .Z(n471) );
  XOR U2147 ( .A(DB[972]), .B(DB[965]), .Z(n473) );
  AND U2148 ( .A(n474), .B(n475), .Z(n472) );
  XOR U2149 ( .A(n476), .B(n477), .Z(n475) );
  XOR U2150 ( .A(DB[965]), .B(DB[958]), .Z(n477) );
  AND U2151 ( .A(n478), .B(n479), .Z(n476) );
  XOR U2152 ( .A(n480), .B(n481), .Z(n479) );
  XOR U2153 ( .A(DB[958]), .B(DB[951]), .Z(n481) );
  AND U2154 ( .A(n482), .B(n483), .Z(n480) );
  XOR U2155 ( .A(n484), .B(n485), .Z(n483) );
  XOR U2156 ( .A(DB[951]), .B(DB[944]), .Z(n485) );
  AND U2157 ( .A(n486), .B(n487), .Z(n484) );
  XOR U2158 ( .A(n488), .B(n489), .Z(n487) );
  XOR U2159 ( .A(DB[944]), .B(DB[937]), .Z(n489) );
  AND U2160 ( .A(n490), .B(n491), .Z(n488) );
  XOR U2161 ( .A(n492), .B(n493), .Z(n491) );
  XOR U2162 ( .A(DB[937]), .B(DB[930]), .Z(n493) );
  AND U2163 ( .A(n494), .B(n495), .Z(n492) );
  XOR U2164 ( .A(n496), .B(n497), .Z(n495) );
  XOR U2165 ( .A(DB[930]), .B(DB[923]), .Z(n497) );
  AND U2166 ( .A(n498), .B(n499), .Z(n496) );
  XOR U2167 ( .A(n500), .B(n501), .Z(n499) );
  XOR U2168 ( .A(DB[923]), .B(DB[916]), .Z(n501) );
  AND U2169 ( .A(n502), .B(n503), .Z(n500) );
  XOR U2170 ( .A(n504), .B(n505), .Z(n503) );
  XOR U2171 ( .A(DB[916]), .B(DB[909]), .Z(n505) );
  AND U2172 ( .A(n506), .B(n507), .Z(n504) );
  XOR U2173 ( .A(n508), .B(n509), .Z(n507) );
  XOR U2174 ( .A(DB[909]), .B(DB[902]), .Z(n509) );
  AND U2175 ( .A(n510), .B(n511), .Z(n508) );
  XOR U2176 ( .A(n512), .B(n513), .Z(n511) );
  XOR U2177 ( .A(DB[902]), .B(DB[895]), .Z(n513) );
  AND U2178 ( .A(n514), .B(n515), .Z(n512) );
  XOR U2179 ( .A(n516), .B(n517), .Z(n515) );
  XOR U2180 ( .A(DB[895]), .B(DB[888]), .Z(n517) );
  AND U2181 ( .A(n518), .B(n519), .Z(n516) );
  XOR U2182 ( .A(n520), .B(n521), .Z(n519) );
  XOR U2183 ( .A(DB[888]), .B(DB[881]), .Z(n521) );
  AND U2184 ( .A(n522), .B(n523), .Z(n520) );
  XOR U2185 ( .A(n524), .B(n525), .Z(n523) );
  XOR U2186 ( .A(DB[881]), .B(DB[874]), .Z(n525) );
  AND U2187 ( .A(n526), .B(n527), .Z(n524) );
  XOR U2188 ( .A(n528), .B(n529), .Z(n527) );
  XOR U2189 ( .A(DB[874]), .B(DB[867]), .Z(n529) );
  AND U2190 ( .A(n530), .B(n531), .Z(n528) );
  XOR U2191 ( .A(n532), .B(n533), .Z(n531) );
  XOR U2192 ( .A(DB[867]), .B(DB[860]), .Z(n533) );
  AND U2193 ( .A(n534), .B(n535), .Z(n532) );
  XOR U2194 ( .A(n536), .B(n537), .Z(n535) );
  XOR U2195 ( .A(DB[860]), .B(DB[853]), .Z(n537) );
  AND U2196 ( .A(n538), .B(n539), .Z(n536) );
  XOR U2197 ( .A(n540), .B(n541), .Z(n539) );
  XOR U2198 ( .A(DB[853]), .B(DB[846]), .Z(n541) );
  AND U2199 ( .A(n542), .B(n543), .Z(n540) );
  XOR U2200 ( .A(n544), .B(n545), .Z(n543) );
  XOR U2201 ( .A(DB[846]), .B(DB[839]), .Z(n545) );
  AND U2202 ( .A(n546), .B(n547), .Z(n544) );
  XOR U2203 ( .A(n548), .B(n549), .Z(n547) );
  XOR U2204 ( .A(DB[839]), .B(DB[832]), .Z(n549) );
  AND U2205 ( .A(n550), .B(n551), .Z(n548) );
  XOR U2206 ( .A(n552), .B(n553), .Z(n551) );
  XOR U2207 ( .A(DB[832]), .B(DB[825]), .Z(n553) );
  AND U2208 ( .A(n554), .B(n555), .Z(n552) );
  XOR U2209 ( .A(n556), .B(n557), .Z(n555) );
  XOR U2210 ( .A(DB[825]), .B(DB[818]), .Z(n557) );
  AND U2211 ( .A(n558), .B(n559), .Z(n556) );
  XOR U2212 ( .A(n560), .B(n561), .Z(n559) );
  XOR U2213 ( .A(DB[818]), .B(DB[811]), .Z(n561) );
  AND U2214 ( .A(n562), .B(n563), .Z(n560) );
  XOR U2215 ( .A(n564), .B(n565), .Z(n563) );
  XOR U2216 ( .A(DB[811]), .B(DB[804]), .Z(n565) );
  AND U2217 ( .A(n566), .B(n567), .Z(n564) );
  XOR U2218 ( .A(n568), .B(n569), .Z(n567) );
  XOR U2219 ( .A(DB[804]), .B(DB[797]), .Z(n569) );
  AND U2220 ( .A(n570), .B(n571), .Z(n568) );
  XOR U2221 ( .A(n572), .B(n573), .Z(n571) );
  XOR U2222 ( .A(DB[797]), .B(DB[790]), .Z(n573) );
  AND U2223 ( .A(n574), .B(n575), .Z(n572) );
  XOR U2224 ( .A(n576), .B(n577), .Z(n575) );
  XOR U2225 ( .A(DB[790]), .B(DB[783]), .Z(n577) );
  AND U2226 ( .A(n578), .B(n579), .Z(n576) );
  XOR U2227 ( .A(n580), .B(n581), .Z(n579) );
  XOR U2228 ( .A(DB[783]), .B(DB[776]), .Z(n581) );
  AND U2229 ( .A(n582), .B(n583), .Z(n580) );
  XOR U2230 ( .A(n584), .B(n585), .Z(n583) );
  XOR U2231 ( .A(DB[776]), .B(DB[769]), .Z(n585) );
  AND U2232 ( .A(n586), .B(n587), .Z(n584) );
  XOR U2233 ( .A(n588), .B(n589), .Z(n587) );
  XOR U2234 ( .A(DB[769]), .B(DB[762]), .Z(n589) );
  AND U2235 ( .A(n590), .B(n591), .Z(n588) );
  XOR U2236 ( .A(n592), .B(n593), .Z(n591) );
  XOR U2237 ( .A(DB[762]), .B(DB[755]), .Z(n593) );
  AND U2238 ( .A(n594), .B(n595), .Z(n592) );
  XOR U2239 ( .A(n596), .B(n597), .Z(n595) );
  XOR U2240 ( .A(DB[755]), .B(DB[748]), .Z(n597) );
  AND U2241 ( .A(n598), .B(n599), .Z(n596) );
  XOR U2242 ( .A(n600), .B(n601), .Z(n599) );
  XOR U2243 ( .A(DB[748]), .B(DB[741]), .Z(n601) );
  AND U2244 ( .A(n602), .B(n603), .Z(n600) );
  XOR U2245 ( .A(n604), .B(n605), .Z(n603) );
  XOR U2246 ( .A(DB[741]), .B(DB[734]), .Z(n605) );
  AND U2247 ( .A(n606), .B(n607), .Z(n604) );
  XOR U2248 ( .A(n608), .B(n609), .Z(n607) );
  XOR U2249 ( .A(DB[734]), .B(DB[727]), .Z(n609) );
  AND U2250 ( .A(n610), .B(n611), .Z(n608) );
  XOR U2251 ( .A(n612), .B(n613), .Z(n611) );
  XOR U2252 ( .A(DB[727]), .B(DB[720]), .Z(n613) );
  AND U2253 ( .A(n614), .B(n615), .Z(n612) );
  XOR U2254 ( .A(n616), .B(n617), .Z(n615) );
  XOR U2255 ( .A(DB[720]), .B(DB[713]), .Z(n617) );
  AND U2256 ( .A(n618), .B(n619), .Z(n616) );
  XOR U2257 ( .A(n620), .B(n621), .Z(n619) );
  XOR U2258 ( .A(DB[713]), .B(DB[706]), .Z(n621) );
  AND U2259 ( .A(n622), .B(n623), .Z(n620) );
  XOR U2260 ( .A(n624), .B(n625), .Z(n623) );
  XOR U2261 ( .A(DB[706]), .B(DB[699]), .Z(n625) );
  AND U2262 ( .A(n626), .B(n627), .Z(n624) );
  XOR U2263 ( .A(n628), .B(n629), .Z(n627) );
  XOR U2264 ( .A(DB[699]), .B(DB[692]), .Z(n629) );
  AND U2265 ( .A(n630), .B(n631), .Z(n628) );
  XOR U2266 ( .A(n632), .B(n633), .Z(n631) );
  XOR U2267 ( .A(DB[692]), .B(DB[685]), .Z(n633) );
  AND U2268 ( .A(n634), .B(n635), .Z(n632) );
  XOR U2269 ( .A(n636), .B(n637), .Z(n635) );
  XOR U2270 ( .A(DB[685]), .B(DB[678]), .Z(n637) );
  AND U2271 ( .A(n638), .B(n639), .Z(n636) );
  XOR U2272 ( .A(n640), .B(n641), .Z(n639) );
  XOR U2273 ( .A(DB[678]), .B(DB[671]), .Z(n641) );
  AND U2274 ( .A(n642), .B(n643), .Z(n640) );
  XOR U2275 ( .A(n644), .B(n645), .Z(n643) );
  XOR U2276 ( .A(DB[671]), .B(DB[664]), .Z(n645) );
  AND U2277 ( .A(n646), .B(n647), .Z(n644) );
  XOR U2278 ( .A(n648), .B(n649), .Z(n647) );
  XOR U2279 ( .A(DB[664]), .B(DB[657]), .Z(n649) );
  AND U2280 ( .A(n650), .B(n651), .Z(n648) );
  XOR U2281 ( .A(n652), .B(n653), .Z(n651) );
  XOR U2282 ( .A(DB[657]), .B(DB[650]), .Z(n653) );
  AND U2283 ( .A(n654), .B(n655), .Z(n652) );
  XOR U2284 ( .A(n656), .B(n657), .Z(n655) );
  XOR U2285 ( .A(DB[650]), .B(DB[643]), .Z(n657) );
  AND U2286 ( .A(n658), .B(n659), .Z(n656) );
  XOR U2287 ( .A(n660), .B(n661), .Z(n659) );
  XOR U2288 ( .A(DB[643]), .B(DB[636]), .Z(n661) );
  AND U2289 ( .A(n662), .B(n663), .Z(n660) );
  XOR U2290 ( .A(n664), .B(n665), .Z(n663) );
  XOR U2291 ( .A(DB[636]), .B(DB[629]), .Z(n665) );
  AND U2292 ( .A(n666), .B(n667), .Z(n664) );
  XOR U2293 ( .A(n668), .B(n669), .Z(n667) );
  XOR U2294 ( .A(DB[629]), .B(DB[622]), .Z(n669) );
  AND U2295 ( .A(n670), .B(n671), .Z(n668) );
  XOR U2296 ( .A(n672), .B(n673), .Z(n671) );
  XOR U2297 ( .A(DB[622]), .B(DB[615]), .Z(n673) );
  AND U2298 ( .A(n674), .B(n675), .Z(n672) );
  XOR U2299 ( .A(n676), .B(n677), .Z(n675) );
  XOR U2300 ( .A(DB[615]), .B(DB[608]), .Z(n677) );
  AND U2301 ( .A(n678), .B(n679), .Z(n676) );
  XOR U2302 ( .A(n680), .B(n681), .Z(n679) );
  XOR U2303 ( .A(DB[608]), .B(DB[601]), .Z(n681) );
  AND U2304 ( .A(n682), .B(n683), .Z(n680) );
  XOR U2305 ( .A(n684), .B(n685), .Z(n683) );
  XOR U2306 ( .A(DB[601]), .B(DB[594]), .Z(n685) );
  AND U2307 ( .A(n686), .B(n687), .Z(n684) );
  XOR U2308 ( .A(n688), .B(n689), .Z(n687) );
  XOR U2309 ( .A(DB[594]), .B(DB[587]), .Z(n689) );
  AND U2310 ( .A(n690), .B(n691), .Z(n688) );
  XOR U2311 ( .A(n692), .B(n693), .Z(n691) );
  XOR U2312 ( .A(DB[587]), .B(DB[580]), .Z(n693) );
  AND U2313 ( .A(n694), .B(n695), .Z(n692) );
  XOR U2314 ( .A(n696), .B(n697), .Z(n695) );
  XOR U2315 ( .A(DB[580]), .B(DB[573]), .Z(n697) );
  AND U2316 ( .A(n698), .B(n699), .Z(n696) );
  XOR U2317 ( .A(n700), .B(n701), .Z(n699) );
  XOR U2318 ( .A(DB[573]), .B(DB[566]), .Z(n701) );
  AND U2319 ( .A(n702), .B(n703), .Z(n700) );
  XOR U2320 ( .A(n704), .B(n705), .Z(n703) );
  XOR U2321 ( .A(DB[566]), .B(DB[559]), .Z(n705) );
  AND U2322 ( .A(n706), .B(n707), .Z(n704) );
  XOR U2323 ( .A(n708), .B(n709), .Z(n707) );
  XOR U2324 ( .A(DB[559]), .B(DB[552]), .Z(n709) );
  AND U2325 ( .A(n710), .B(n711), .Z(n708) );
  XOR U2326 ( .A(n712), .B(n713), .Z(n711) );
  XOR U2327 ( .A(DB[552]), .B(DB[545]), .Z(n713) );
  AND U2328 ( .A(n714), .B(n715), .Z(n712) );
  XOR U2329 ( .A(n716), .B(n717), .Z(n715) );
  XOR U2330 ( .A(DB[545]), .B(DB[538]), .Z(n717) );
  AND U2331 ( .A(n718), .B(n719), .Z(n716) );
  XOR U2332 ( .A(n720), .B(n721), .Z(n719) );
  XOR U2333 ( .A(DB[538]), .B(DB[531]), .Z(n721) );
  AND U2334 ( .A(n722), .B(n723), .Z(n720) );
  XOR U2335 ( .A(n724), .B(n725), .Z(n723) );
  XOR U2336 ( .A(DB[531]), .B(DB[524]), .Z(n725) );
  AND U2337 ( .A(n726), .B(n727), .Z(n724) );
  XOR U2338 ( .A(n728), .B(n729), .Z(n727) );
  XOR U2339 ( .A(DB[524]), .B(DB[517]), .Z(n729) );
  AND U2340 ( .A(n730), .B(n731), .Z(n728) );
  XOR U2341 ( .A(n732), .B(n733), .Z(n731) );
  XOR U2342 ( .A(DB[517]), .B(DB[510]), .Z(n733) );
  AND U2343 ( .A(n734), .B(n735), .Z(n732) );
  XOR U2344 ( .A(n736), .B(n737), .Z(n735) );
  XOR U2345 ( .A(DB[510]), .B(DB[503]), .Z(n737) );
  AND U2346 ( .A(n738), .B(n739), .Z(n736) );
  XOR U2347 ( .A(n740), .B(n741), .Z(n739) );
  XOR U2348 ( .A(DB[503]), .B(DB[496]), .Z(n741) );
  AND U2349 ( .A(n742), .B(n743), .Z(n740) );
  XOR U2350 ( .A(n744), .B(n745), .Z(n743) );
  XOR U2351 ( .A(DB[496]), .B(DB[489]), .Z(n745) );
  AND U2352 ( .A(n746), .B(n747), .Z(n744) );
  XOR U2353 ( .A(n748), .B(n749), .Z(n747) );
  XOR U2354 ( .A(DB[489]), .B(DB[482]), .Z(n749) );
  AND U2355 ( .A(n750), .B(n751), .Z(n748) );
  XOR U2356 ( .A(n752), .B(n753), .Z(n751) );
  XOR U2357 ( .A(DB[482]), .B(DB[475]), .Z(n753) );
  AND U2358 ( .A(n754), .B(n755), .Z(n752) );
  XOR U2359 ( .A(n756), .B(n757), .Z(n755) );
  XOR U2360 ( .A(DB[475]), .B(DB[468]), .Z(n757) );
  AND U2361 ( .A(n758), .B(n759), .Z(n756) );
  XOR U2362 ( .A(n760), .B(n761), .Z(n759) );
  XOR U2363 ( .A(DB[468]), .B(DB[461]), .Z(n761) );
  AND U2364 ( .A(n762), .B(n763), .Z(n760) );
  XOR U2365 ( .A(n764), .B(n765), .Z(n763) );
  XOR U2366 ( .A(DB[461]), .B(DB[454]), .Z(n765) );
  AND U2367 ( .A(n766), .B(n767), .Z(n764) );
  XOR U2368 ( .A(n768), .B(n769), .Z(n767) );
  XOR U2369 ( .A(DB[454]), .B(DB[447]), .Z(n769) );
  AND U2370 ( .A(n770), .B(n771), .Z(n768) );
  XOR U2371 ( .A(n772), .B(n773), .Z(n771) );
  XOR U2372 ( .A(DB[447]), .B(DB[440]), .Z(n773) );
  AND U2373 ( .A(n774), .B(n775), .Z(n772) );
  XOR U2374 ( .A(n776), .B(n777), .Z(n775) );
  XOR U2375 ( .A(DB[440]), .B(DB[433]), .Z(n777) );
  AND U2376 ( .A(n778), .B(n779), .Z(n776) );
  XOR U2377 ( .A(n780), .B(n781), .Z(n779) );
  XOR U2378 ( .A(DB[433]), .B(DB[426]), .Z(n781) );
  AND U2379 ( .A(n782), .B(n783), .Z(n780) );
  XOR U2380 ( .A(n784), .B(n785), .Z(n783) );
  XOR U2381 ( .A(DB[426]), .B(DB[419]), .Z(n785) );
  AND U2382 ( .A(n786), .B(n787), .Z(n784) );
  XOR U2383 ( .A(n788), .B(n789), .Z(n787) );
  XOR U2384 ( .A(DB[419]), .B(DB[412]), .Z(n789) );
  AND U2385 ( .A(n790), .B(n791), .Z(n788) );
  XOR U2386 ( .A(n792), .B(n793), .Z(n791) );
  XOR U2387 ( .A(DB[412]), .B(DB[405]), .Z(n793) );
  AND U2388 ( .A(n794), .B(n795), .Z(n792) );
  XOR U2389 ( .A(n796), .B(n797), .Z(n795) );
  XOR U2390 ( .A(DB[405]), .B(DB[398]), .Z(n797) );
  AND U2391 ( .A(n798), .B(n799), .Z(n796) );
  XOR U2392 ( .A(n800), .B(n801), .Z(n799) );
  XOR U2393 ( .A(DB[398]), .B(DB[391]), .Z(n801) );
  AND U2394 ( .A(n802), .B(n803), .Z(n800) );
  XOR U2395 ( .A(n804), .B(n805), .Z(n803) );
  XOR U2396 ( .A(DB[391]), .B(DB[384]), .Z(n805) );
  AND U2397 ( .A(n806), .B(n807), .Z(n804) );
  XOR U2398 ( .A(n808), .B(n809), .Z(n807) );
  XOR U2399 ( .A(DB[384]), .B(DB[377]), .Z(n809) );
  AND U2400 ( .A(n810), .B(n811), .Z(n808) );
  XOR U2401 ( .A(n812), .B(n813), .Z(n811) );
  XOR U2402 ( .A(DB[377]), .B(DB[370]), .Z(n813) );
  AND U2403 ( .A(n814), .B(n815), .Z(n812) );
  XOR U2404 ( .A(n816), .B(n817), .Z(n815) );
  XOR U2405 ( .A(DB[370]), .B(DB[363]), .Z(n817) );
  AND U2406 ( .A(n818), .B(n819), .Z(n816) );
  XOR U2407 ( .A(n820), .B(n821), .Z(n819) );
  XOR U2408 ( .A(DB[363]), .B(DB[356]), .Z(n821) );
  AND U2409 ( .A(n822), .B(n823), .Z(n820) );
  XOR U2410 ( .A(n824), .B(n825), .Z(n823) );
  XOR U2411 ( .A(DB[356]), .B(DB[349]), .Z(n825) );
  AND U2412 ( .A(n826), .B(n827), .Z(n824) );
  XOR U2413 ( .A(n828), .B(n829), .Z(n827) );
  XOR U2414 ( .A(DB[349]), .B(DB[342]), .Z(n829) );
  AND U2415 ( .A(n830), .B(n831), .Z(n828) );
  XOR U2416 ( .A(n832), .B(n833), .Z(n831) );
  XOR U2417 ( .A(DB[342]), .B(DB[335]), .Z(n833) );
  AND U2418 ( .A(n834), .B(n835), .Z(n832) );
  XOR U2419 ( .A(n836), .B(n837), .Z(n835) );
  XOR U2420 ( .A(DB[335]), .B(DB[328]), .Z(n837) );
  AND U2421 ( .A(n838), .B(n839), .Z(n836) );
  XOR U2422 ( .A(n840), .B(n841), .Z(n839) );
  XOR U2423 ( .A(DB[328]), .B(DB[321]), .Z(n841) );
  AND U2424 ( .A(n842), .B(n843), .Z(n840) );
  XOR U2425 ( .A(n844), .B(n845), .Z(n843) );
  XOR U2426 ( .A(DB[321]), .B(DB[314]), .Z(n845) );
  AND U2427 ( .A(n846), .B(n847), .Z(n844) );
  XOR U2428 ( .A(n848), .B(n849), .Z(n847) );
  XOR U2429 ( .A(DB[314]), .B(DB[307]), .Z(n849) );
  AND U2430 ( .A(n850), .B(n851), .Z(n848) );
  XOR U2431 ( .A(n852), .B(n853), .Z(n851) );
  XOR U2432 ( .A(DB[307]), .B(DB[300]), .Z(n853) );
  AND U2433 ( .A(n854), .B(n855), .Z(n852) );
  XOR U2434 ( .A(n856), .B(n857), .Z(n855) );
  XOR U2435 ( .A(DB[300]), .B(DB[293]), .Z(n857) );
  AND U2436 ( .A(n858), .B(n859), .Z(n856) );
  XOR U2437 ( .A(n860), .B(n861), .Z(n859) );
  XOR U2438 ( .A(DB[293]), .B(DB[286]), .Z(n861) );
  AND U2439 ( .A(n862), .B(n863), .Z(n860) );
  XOR U2440 ( .A(n864), .B(n865), .Z(n863) );
  XOR U2441 ( .A(DB[286]), .B(DB[279]), .Z(n865) );
  AND U2442 ( .A(n866), .B(n867), .Z(n864) );
  XOR U2443 ( .A(n868), .B(n869), .Z(n867) );
  XOR U2444 ( .A(DB[279]), .B(DB[272]), .Z(n869) );
  AND U2445 ( .A(n870), .B(n871), .Z(n868) );
  XOR U2446 ( .A(n872), .B(n873), .Z(n871) );
  XOR U2447 ( .A(DB[272]), .B(DB[265]), .Z(n873) );
  AND U2448 ( .A(n874), .B(n875), .Z(n872) );
  XOR U2449 ( .A(n876), .B(n877), .Z(n875) );
  XOR U2450 ( .A(DB[265]), .B(DB[258]), .Z(n877) );
  AND U2451 ( .A(n878), .B(n879), .Z(n876) );
  XOR U2452 ( .A(n880), .B(n881), .Z(n879) );
  XOR U2453 ( .A(DB[258]), .B(DB[251]), .Z(n881) );
  AND U2454 ( .A(n882), .B(n883), .Z(n880) );
  XOR U2455 ( .A(n884), .B(n885), .Z(n883) );
  XOR U2456 ( .A(DB[251]), .B(DB[244]), .Z(n885) );
  AND U2457 ( .A(n886), .B(n887), .Z(n884) );
  XOR U2458 ( .A(n888), .B(n889), .Z(n887) );
  XOR U2459 ( .A(DB[244]), .B(DB[237]), .Z(n889) );
  AND U2460 ( .A(n890), .B(n891), .Z(n888) );
  XOR U2461 ( .A(n892), .B(n893), .Z(n891) );
  XOR U2462 ( .A(DB[237]), .B(DB[230]), .Z(n893) );
  AND U2463 ( .A(n894), .B(n895), .Z(n892) );
  XOR U2464 ( .A(n896), .B(n897), .Z(n895) );
  XOR U2465 ( .A(DB[230]), .B(DB[223]), .Z(n897) );
  AND U2466 ( .A(n898), .B(n899), .Z(n896) );
  XOR U2467 ( .A(n900), .B(n901), .Z(n899) );
  XOR U2468 ( .A(DB[223]), .B(DB[216]), .Z(n901) );
  AND U2469 ( .A(n902), .B(n903), .Z(n900) );
  XOR U2470 ( .A(n904), .B(n905), .Z(n903) );
  XOR U2471 ( .A(DB[216]), .B(DB[209]), .Z(n905) );
  AND U2472 ( .A(n906), .B(n907), .Z(n904) );
  XOR U2473 ( .A(n908), .B(n909), .Z(n907) );
  XOR U2474 ( .A(DB[209]), .B(DB[202]), .Z(n909) );
  AND U2475 ( .A(n910), .B(n911), .Z(n908) );
  XOR U2476 ( .A(n912), .B(n913), .Z(n911) );
  XOR U2477 ( .A(DB[202]), .B(DB[195]), .Z(n913) );
  AND U2478 ( .A(n914), .B(n915), .Z(n912) );
  XOR U2479 ( .A(n916), .B(n917), .Z(n915) );
  XOR U2480 ( .A(DB[195]), .B(DB[188]), .Z(n917) );
  AND U2481 ( .A(n918), .B(n919), .Z(n916) );
  XOR U2482 ( .A(n920), .B(n921), .Z(n919) );
  XOR U2483 ( .A(DB[188]), .B(DB[181]), .Z(n921) );
  AND U2484 ( .A(n922), .B(n923), .Z(n920) );
  XOR U2485 ( .A(n924), .B(n925), .Z(n923) );
  XOR U2486 ( .A(DB[181]), .B(DB[174]), .Z(n925) );
  AND U2487 ( .A(n926), .B(n927), .Z(n924) );
  XOR U2488 ( .A(n928), .B(n929), .Z(n927) );
  XOR U2489 ( .A(DB[174]), .B(DB[167]), .Z(n929) );
  AND U2490 ( .A(n930), .B(n931), .Z(n928) );
  XOR U2491 ( .A(n932), .B(n933), .Z(n931) );
  XOR U2492 ( .A(DB[167]), .B(DB[160]), .Z(n933) );
  AND U2493 ( .A(n934), .B(n935), .Z(n932) );
  XOR U2494 ( .A(n936), .B(n937), .Z(n935) );
  XOR U2495 ( .A(DB[160]), .B(DB[153]), .Z(n937) );
  AND U2496 ( .A(n938), .B(n939), .Z(n936) );
  XOR U2497 ( .A(n940), .B(n941), .Z(n939) );
  XOR U2498 ( .A(DB[153]), .B(DB[146]), .Z(n941) );
  AND U2499 ( .A(n942), .B(n943), .Z(n940) );
  XOR U2500 ( .A(n944), .B(n945), .Z(n943) );
  XOR U2501 ( .A(DB[146]), .B(DB[139]), .Z(n945) );
  AND U2502 ( .A(n946), .B(n947), .Z(n944) );
  XOR U2503 ( .A(n948), .B(n949), .Z(n947) );
  XOR U2504 ( .A(DB[139]), .B(DB[132]), .Z(n949) );
  AND U2505 ( .A(n950), .B(n951), .Z(n948) );
  XOR U2506 ( .A(n952), .B(n953), .Z(n951) );
  XOR U2507 ( .A(DB[132]), .B(DB[125]), .Z(n953) );
  AND U2508 ( .A(n954), .B(n955), .Z(n952) );
  XOR U2509 ( .A(n956), .B(n957), .Z(n955) );
  XOR U2510 ( .A(DB[125]), .B(DB[118]), .Z(n957) );
  AND U2511 ( .A(n958), .B(n959), .Z(n956) );
  XOR U2512 ( .A(n960), .B(n961), .Z(n959) );
  XOR U2513 ( .A(DB[118]), .B(DB[111]), .Z(n961) );
  AND U2514 ( .A(n962), .B(n963), .Z(n960) );
  XOR U2515 ( .A(n964), .B(n965), .Z(n963) );
  XOR U2516 ( .A(DB[111]), .B(DB[104]), .Z(n965) );
  AND U2517 ( .A(n966), .B(n967), .Z(n964) );
  XOR U2518 ( .A(n968), .B(n969), .Z(n967) );
  XOR U2519 ( .A(DB[97]), .B(DB[104]), .Z(n969) );
  AND U2520 ( .A(n970), .B(n971), .Z(n968) );
  XOR U2521 ( .A(n972), .B(n973), .Z(n971) );
  XOR U2522 ( .A(DB[97]), .B(DB[90]), .Z(n973) );
  AND U2523 ( .A(n974), .B(n975), .Z(n972) );
  XOR U2524 ( .A(n976), .B(n977), .Z(n975) );
  XOR U2525 ( .A(DB[90]), .B(DB[83]), .Z(n977) );
  AND U2526 ( .A(n978), .B(n979), .Z(n976) );
  XOR U2527 ( .A(n980), .B(n981), .Z(n979) );
  XOR U2528 ( .A(DB[83]), .B(DB[76]), .Z(n981) );
  AND U2529 ( .A(n982), .B(n983), .Z(n980) );
  XOR U2530 ( .A(n984), .B(n985), .Z(n983) );
  XOR U2531 ( .A(DB[76]), .B(DB[69]), .Z(n985) );
  AND U2532 ( .A(n986), .B(n987), .Z(n984) );
  XOR U2533 ( .A(n988), .B(n989), .Z(n987) );
  XOR U2534 ( .A(DB[69]), .B(DB[62]), .Z(n989) );
  AND U2535 ( .A(n990), .B(n991), .Z(n988) );
  XOR U2536 ( .A(n992), .B(n993), .Z(n991) );
  XOR U2537 ( .A(DB[62]), .B(DB[55]), .Z(n993) );
  AND U2538 ( .A(n994), .B(n995), .Z(n992) );
  XOR U2539 ( .A(n996), .B(n997), .Z(n995) );
  XOR U2540 ( .A(DB[55]), .B(DB[48]), .Z(n997) );
  AND U2541 ( .A(n998), .B(n999), .Z(n996) );
  XOR U2542 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U2543 ( .A(DB[48]), .B(DB[41]), .Z(n1001) );
  AND U2544 ( .A(n1002), .B(n1003), .Z(n1000) );
  XOR U2545 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U2546 ( .A(DB[41]), .B(DB[34]), .Z(n1005) );
  AND U2547 ( .A(n1006), .B(n1007), .Z(n1004) );
  XOR U2548 ( .A(n1008), .B(n1009), .Z(n1007) );
  XOR U2549 ( .A(DB[34]), .B(DB[27]), .Z(n1009) );
  AND U2550 ( .A(n1010), .B(n1011), .Z(n1008) );
  XOR U2551 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR U2552 ( .A(DB[27]), .B(DB[20]), .Z(n1013) );
  AND U2553 ( .A(n1014), .B(n1015), .Z(n1012) );
  XOR U2554 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U2555 ( .A(DB[20]), .B(DB[13]), .Z(n1017) );
  AND U2556 ( .A(n1018), .B(n1019), .Z(n1016) );
  XOR U2557 ( .A(DB[6]), .B(DB[13]), .Z(n1019) );
  XOR U2558 ( .A(DB[1790]), .B(n1020), .Z(min_val_out[5]) );
  AND U2559 ( .A(n2), .B(n1021), .Z(n1020) );
  XOR U2560 ( .A(n1022), .B(n1023), .Z(n1021) );
  XOR U2561 ( .A(DB[1790]), .B(DB[1783]), .Z(n1023) );
  AND U2562 ( .A(n6), .B(n1024), .Z(n1022) );
  XOR U2563 ( .A(n1025), .B(n1026), .Z(n1024) );
  XOR U2564 ( .A(DB[1783]), .B(DB[1776]), .Z(n1026) );
  AND U2565 ( .A(n10), .B(n1027), .Z(n1025) );
  XOR U2566 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U2567 ( .A(DB[1776]), .B(DB[1769]), .Z(n1029) );
  AND U2568 ( .A(n14), .B(n1030), .Z(n1028) );
  XOR U2569 ( .A(n1031), .B(n1032), .Z(n1030) );
  XOR U2570 ( .A(DB[1769]), .B(DB[1762]), .Z(n1032) );
  AND U2571 ( .A(n18), .B(n1033), .Z(n1031) );
  XOR U2572 ( .A(n1034), .B(n1035), .Z(n1033) );
  XOR U2573 ( .A(DB[1762]), .B(DB[1755]), .Z(n1035) );
  AND U2574 ( .A(n22), .B(n1036), .Z(n1034) );
  XOR U2575 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U2576 ( .A(DB[1755]), .B(DB[1748]), .Z(n1038) );
  AND U2577 ( .A(n26), .B(n1039), .Z(n1037) );
  XOR U2578 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U2579 ( .A(DB[1748]), .B(DB[1741]), .Z(n1041) );
  AND U2580 ( .A(n30), .B(n1042), .Z(n1040) );
  XOR U2581 ( .A(n1043), .B(n1044), .Z(n1042) );
  XOR U2582 ( .A(DB[1741]), .B(DB[1734]), .Z(n1044) );
  AND U2583 ( .A(n34), .B(n1045), .Z(n1043) );
  XOR U2584 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U2585 ( .A(DB[1734]), .B(DB[1727]), .Z(n1047) );
  AND U2586 ( .A(n38), .B(n1048), .Z(n1046) );
  XOR U2587 ( .A(n1049), .B(n1050), .Z(n1048) );
  XOR U2588 ( .A(DB[1727]), .B(DB[1720]), .Z(n1050) );
  AND U2589 ( .A(n42), .B(n1051), .Z(n1049) );
  XOR U2590 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR U2591 ( .A(DB[1720]), .B(DB[1713]), .Z(n1053) );
  AND U2592 ( .A(n46), .B(n1054), .Z(n1052) );
  XOR U2593 ( .A(n1055), .B(n1056), .Z(n1054) );
  XOR U2594 ( .A(DB[1713]), .B(DB[1706]), .Z(n1056) );
  AND U2595 ( .A(n50), .B(n1057), .Z(n1055) );
  XOR U2596 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U2597 ( .A(DB[1706]), .B(DB[1699]), .Z(n1059) );
  AND U2598 ( .A(n54), .B(n1060), .Z(n1058) );
  XOR U2599 ( .A(n1061), .B(n1062), .Z(n1060) );
  XOR U2600 ( .A(DB[1699]), .B(DB[1692]), .Z(n1062) );
  AND U2601 ( .A(n58), .B(n1063), .Z(n1061) );
  XOR U2602 ( .A(n1064), .B(n1065), .Z(n1063) );
  XOR U2603 ( .A(DB[1692]), .B(DB[1685]), .Z(n1065) );
  AND U2604 ( .A(n62), .B(n1066), .Z(n1064) );
  XOR U2605 ( .A(n1067), .B(n1068), .Z(n1066) );
  XOR U2606 ( .A(DB[1685]), .B(DB[1678]), .Z(n1068) );
  AND U2607 ( .A(n66), .B(n1069), .Z(n1067) );
  XOR U2608 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U2609 ( .A(DB[1678]), .B(DB[1671]), .Z(n1071) );
  AND U2610 ( .A(n70), .B(n1072), .Z(n1070) );
  XOR U2611 ( .A(n1073), .B(n1074), .Z(n1072) );
  XOR U2612 ( .A(DB[1671]), .B(DB[1664]), .Z(n1074) );
  AND U2613 ( .A(n74), .B(n1075), .Z(n1073) );
  XOR U2614 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U2615 ( .A(DB[1664]), .B(DB[1657]), .Z(n1077) );
  AND U2616 ( .A(n78), .B(n1078), .Z(n1076) );
  XOR U2617 ( .A(n1079), .B(n1080), .Z(n1078) );
  XOR U2618 ( .A(DB[1657]), .B(DB[1650]), .Z(n1080) );
  AND U2619 ( .A(n82), .B(n1081), .Z(n1079) );
  XOR U2620 ( .A(n1082), .B(n1083), .Z(n1081) );
  XOR U2621 ( .A(DB[1650]), .B(DB[1643]), .Z(n1083) );
  AND U2622 ( .A(n86), .B(n1084), .Z(n1082) );
  XOR U2623 ( .A(n1085), .B(n1086), .Z(n1084) );
  XOR U2624 ( .A(DB[1643]), .B(DB[1636]), .Z(n1086) );
  AND U2625 ( .A(n90), .B(n1087), .Z(n1085) );
  XOR U2626 ( .A(n1088), .B(n1089), .Z(n1087) );
  XOR U2627 ( .A(DB[1636]), .B(DB[1629]), .Z(n1089) );
  AND U2628 ( .A(n94), .B(n1090), .Z(n1088) );
  XOR U2629 ( .A(n1091), .B(n1092), .Z(n1090) );
  XOR U2630 ( .A(DB[1629]), .B(DB[1622]), .Z(n1092) );
  AND U2631 ( .A(n98), .B(n1093), .Z(n1091) );
  XOR U2632 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U2633 ( .A(DB[1622]), .B(DB[1615]), .Z(n1095) );
  AND U2634 ( .A(n102), .B(n1096), .Z(n1094) );
  XOR U2635 ( .A(n1097), .B(n1098), .Z(n1096) );
  XOR U2636 ( .A(DB[1615]), .B(DB[1608]), .Z(n1098) );
  AND U2637 ( .A(n106), .B(n1099), .Z(n1097) );
  XOR U2638 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U2639 ( .A(DB[1608]), .B(DB[1601]), .Z(n1101) );
  AND U2640 ( .A(n110), .B(n1102), .Z(n1100) );
  XOR U2641 ( .A(n1103), .B(n1104), .Z(n1102) );
  XOR U2642 ( .A(DB[1601]), .B(DB[1594]), .Z(n1104) );
  AND U2643 ( .A(n114), .B(n1105), .Z(n1103) );
  XOR U2644 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U2645 ( .A(DB[1594]), .B(DB[1587]), .Z(n1107) );
  AND U2646 ( .A(n118), .B(n1108), .Z(n1106) );
  XOR U2647 ( .A(n1109), .B(n1110), .Z(n1108) );
  XOR U2648 ( .A(DB[1587]), .B(DB[1580]), .Z(n1110) );
  AND U2649 ( .A(n122), .B(n1111), .Z(n1109) );
  XOR U2650 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR U2651 ( .A(DB[1580]), .B(DB[1573]), .Z(n1113) );
  AND U2652 ( .A(n126), .B(n1114), .Z(n1112) );
  XOR U2653 ( .A(n1115), .B(n1116), .Z(n1114) );
  XOR U2654 ( .A(DB[1573]), .B(DB[1566]), .Z(n1116) );
  AND U2655 ( .A(n130), .B(n1117), .Z(n1115) );
  XOR U2656 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U2657 ( .A(DB[1566]), .B(DB[1559]), .Z(n1119) );
  AND U2658 ( .A(n134), .B(n1120), .Z(n1118) );
  XOR U2659 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U2660 ( .A(DB[1559]), .B(DB[1552]), .Z(n1122) );
  AND U2661 ( .A(n138), .B(n1123), .Z(n1121) );
  XOR U2662 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U2663 ( .A(DB[1552]), .B(DB[1545]), .Z(n1125) );
  AND U2664 ( .A(n142), .B(n1126), .Z(n1124) );
  XOR U2665 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U2666 ( .A(DB[1545]), .B(DB[1538]), .Z(n1128) );
  AND U2667 ( .A(n146), .B(n1129), .Z(n1127) );
  XOR U2668 ( .A(n1130), .B(n1131), .Z(n1129) );
  XOR U2669 ( .A(DB[1538]), .B(DB[1531]), .Z(n1131) );
  AND U2670 ( .A(n150), .B(n1132), .Z(n1130) );
  XOR U2671 ( .A(n1133), .B(n1134), .Z(n1132) );
  XOR U2672 ( .A(DB[1531]), .B(DB[1524]), .Z(n1134) );
  AND U2673 ( .A(n154), .B(n1135), .Z(n1133) );
  XOR U2674 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U2675 ( .A(DB[1524]), .B(DB[1517]), .Z(n1137) );
  AND U2676 ( .A(n158), .B(n1138), .Z(n1136) );
  XOR U2677 ( .A(n1139), .B(n1140), .Z(n1138) );
  XOR U2678 ( .A(DB[1517]), .B(DB[1510]), .Z(n1140) );
  AND U2679 ( .A(n162), .B(n1141), .Z(n1139) );
  XOR U2680 ( .A(n1142), .B(n1143), .Z(n1141) );
  XOR U2681 ( .A(DB[1510]), .B(DB[1503]), .Z(n1143) );
  AND U2682 ( .A(n166), .B(n1144), .Z(n1142) );
  XOR U2683 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U2684 ( .A(DB[1503]), .B(DB[1496]), .Z(n1146) );
  AND U2685 ( .A(n170), .B(n1147), .Z(n1145) );
  XOR U2686 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U2687 ( .A(DB[1496]), .B(DB[1489]), .Z(n1149) );
  AND U2688 ( .A(n174), .B(n1150), .Z(n1148) );
  XOR U2689 ( .A(n1151), .B(n1152), .Z(n1150) );
  XOR U2690 ( .A(DB[1489]), .B(DB[1482]), .Z(n1152) );
  AND U2691 ( .A(n178), .B(n1153), .Z(n1151) );
  XOR U2692 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U2693 ( .A(DB[1482]), .B(DB[1475]), .Z(n1155) );
  AND U2694 ( .A(n182), .B(n1156), .Z(n1154) );
  XOR U2695 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U2696 ( .A(DB[1475]), .B(DB[1468]), .Z(n1158) );
  AND U2697 ( .A(n186), .B(n1159), .Z(n1157) );
  XOR U2698 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U2699 ( .A(DB[1468]), .B(DB[1461]), .Z(n1161) );
  AND U2700 ( .A(n190), .B(n1162), .Z(n1160) );
  XOR U2701 ( .A(n1163), .B(n1164), .Z(n1162) );
  XOR U2702 ( .A(DB[1461]), .B(DB[1454]), .Z(n1164) );
  AND U2703 ( .A(n194), .B(n1165), .Z(n1163) );
  XOR U2704 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U2705 ( .A(DB[1454]), .B(DB[1447]), .Z(n1167) );
  AND U2706 ( .A(n198), .B(n1168), .Z(n1166) );
  XOR U2707 ( .A(n1169), .B(n1170), .Z(n1168) );
  XOR U2708 ( .A(DB[1447]), .B(DB[1440]), .Z(n1170) );
  AND U2709 ( .A(n202), .B(n1171), .Z(n1169) );
  XOR U2710 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U2711 ( .A(DB[1440]), .B(DB[1433]), .Z(n1173) );
  AND U2712 ( .A(n206), .B(n1174), .Z(n1172) );
  XOR U2713 ( .A(n1175), .B(n1176), .Z(n1174) );
  XOR U2714 ( .A(DB[1433]), .B(DB[1426]), .Z(n1176) );
  AND U2715 ( .A(n210), .B(n1177), .Z(n1175) );
  XOR U2716 ( .A(n1178), .B(n1179), .Z(n1177) );
  XOR U2717 ( .A(DB[1426]), .B(DB[1419]), .Z(n1179) );
  AND U2718 ( .A(n214), .B(n1180), .Z(n1178) );
  XOR U2719 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U2720 ( .A(DB[1419]), .B(DB[1412]), .Z(n1182) );
  AND U2721 ( .A(n218), .B(n1183), .Z(n1181) );
  XOR U2722 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U2723 ( .A(DB[1412]), .B(DB[1405]), .Z(n1185) );
  AND U2724 ( .A(n222), .B(n1186), .Z(n1184) );
  XOR U2725 ( .A(n1187), .B(n1188), .Z(n1186) );
  XOR U2726 ( .A(DB[1405]), .B(DB[1398]), .Z(n1188) );
  AND U2727 ( .A(n226), .B(n1189), .Z(n1187) );
  XOR U2728 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U2729 ( .A(DB[1398]), .B(DB[1391]), .Z(n1191) );
  AND U2730 ( .A(n230), .B(n1192), .Z(n1190) );
  XOR U2731 ( .A(n1193), .B(n1194), .Z(n1192) );
  XOR U2732 ( .A(DB[1391]), .B(DB[1384]), .Z(n1194) );
  AND U2733 ( .A(n234), .B(n1195), .Z(n1193) );
  XOR U2734 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR U2735 ( .A(DB[1384]), .B(DB[1377]), .Z(n1197) );
  AND U2736 ( .A(n238), .B(n1198), .Z(n1196) );
  XOR U2737 ( .A(n1199), .B(n1200), .Z(n1198) );
  XOR U2738 ( .A(DB[1377]), .B(DB[1370]), .Z(n1200) );
  AND U2739 ( .A(n242), .B(n1201), .Z(n1199) );
  XOR U2740 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U2741 ( .A(DB[1370]), .B(DB[1363]), .Z(n1203) );
  AND U2742 ( .A(n246), .B(n1204), .Z(n1202) );
  XOR U2743 ( .A(n1205), .B(n1206), .Z(n1204) );
  XOR U2744 ( .A(DB[1363]), .B(DB[1356]), .Z(n1206) );
  AND U2745 ( .A(n250), .B(n1207), .Z(n1205) );
  XOR U2746 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U2747 ( .A(DB[1356]), .B(DB[1349]), .Z(n1209) );
  AND U2748 ( .A(n254), .B(n1210), .Z(n1208) );
  XOR U2749 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U2750 ( .A(DB[1349]), .B(DB[1342]), .Z(n1212) );
  AND U2751 ( .A(n258), .B(n1213), .Z(n1211) );
  XOR U2752 ( .A(n1214), .B(n1215), .Z(n1213) );
  XOR U2753 ( .A(DB[1342]), .B(DB[1335]), .Z(n1215) );
  AND U2754 ( .A(n262), .B(n1216), .Z(n1214) );
  XOR U2755 ( .A(n1217), .B(n1218), .Z(n1216) );
  XOR U2756 ( .A(DB[1335]), .B(DB[1328]), .Z(n1218) );
  AND U2757 ( .A(n266), .B(n1219), .Z(n1217) );
  XOR U2758 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U2759 ( .A(DB[1328]), .B(DB[1321]), .Z(n1221) );
  AND U2760 ( .A(n270), .B(n1222), .Z(n1220) );
  XOR U2761 ( .A(n1223), .B(n1224), .Z(n1222) );
  XOR U2762 ( .A(DB[1321]), .B(DB[1314]), .Z(n1224) );
  AND U2763 ( .A(n274), .B(n1225), .Z(n1223) );
  XOR U2764 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U2765 ( .A(DB[1314]), .B(DB[1307]), .Z(n1227) );
  AND U2766 ( .A(n278), .B(n1228), .Z(n1226) );
  XOR U2767 ( .A(n1229), .B(n1230), .Z(n1228) );
  XOR U2768 ( .A(DB[1307]), .B(DB[1300]), .Z(n1230) );
  AND U2769 ( .A(n282), .B(n1231), .Z(n1229) );
  XOR U2770 ( .A(n1232), .B(n1233), .Z(n1231) );
  XOR U2771 ( .A(DB[1300]), .B(DB[1293]), .Z(n1233) );
  AND U2772 ( .A(n286), .B(n1234), .Z(n1232) );
  XOR U2773 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U2774 ( .A(DB[1293]), .B(DB[1286]), .Z(n1236) );
  AND U2775 ( .A(n290), .B(n1237), .Z(n1235) );
  XOR U2776 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U2777 ( .A(DB[1286]), .B(DB[1279]), .Z(n1239) );
  AND U2778 ( .A(n294), .B(n1240), .Z(n1238) );
  XOR U2779 ( .A(n1241), .B(n1242), .Z(n1240) );
  XOR U2780 ( .A(DB[1279]), .B(DB[1272]), .Z(n1242) );
  AND U2781 ( .A(n298), .B(n1243), .Z(n1241) );
  XOR U2782 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U2783 ( .A(DB[1272]), .B(DB[1265]), .Z(n1245) );
  AND U2784 ( .A(n302), .B(n1246), .Z(n1244) );
  XOR U2785 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U2786 ( .A(DB[1265]), .B(DB[1258]), .Z(n1248) );
  AND U2787 ( .A(n306), .B(n1249), .Z(n1247) );
  XOR U2788 ( .A(n1250), .B(n1251), .Z(n1249) );
  XOR U2789 ( .A(DB[1258]), .B(DB[1251]), .Z(n1251) );
  AND U2790 ( .A(n310), .B(n1252), .Z(n1250) );
  XOR U2791 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U2792 ( .A(DB[1251]), .B(DB[1244]), .Z(n1254) );
  AND U2793 ( .A(n314), .B(n1255), .Z(n1253) );
  XOR U2794 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U2795 ( .A(DB[1244]), .B(DB[1237]), .Z(n1257) );
  AND U2796 ( .A(n318), .B(n1258), .Z(n1256) );
  XOR U2797 ( .A(n1259), .B(n1260), .Z(n1258) );
  XOR U2798 ( .A(DB[1237]), .B(DB[1230]), .Z(n1260) );
  AND U2799 ( .A(n322), .B(n1261), .Z(n1259) );
  XOR U2800 ( .A(n1262), .B(n1263), .Z(n1261) );
  XOR U2801 ( .A(DB[1230]), .B(DB[1223]), .Z(n1263) );
  AND U2802 ( .A(n326), .B(n1264), .Z(n1262) );
  XOR U2803 ( .A(n1265), .B(n1266), .Z(n1264) );
  XOR U2804 ( .A(DB[1223]), .B(DB[1216]), .Z(n1266) );
  AND U2805 ( .A(n330), .B(n1267), .Z(n1265) );
  XOR U2806 ( .A(n1268), .B(n1269), .Z(n1267) );
  XOR U2807 ( .A(DB[1216]), .B(DB[1209]), .Z(n1269) );
  AND U2808 ( .A(n334), .B(n1270), .Z(n1268) );
  XOR U2809 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U2810 ( .A(DB[1209]), .B(DB[1202]), .Z(n1272) );
  AND U2811 ( .A(n338), .B(n1273), .Z(n1271) );
  XOR U2812 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U2813 ( .A(DB[1202]), .B(DB[1195]), .Z(n1275) );
  AND U2814 ( .A(n342), .B(n1276), .Z(n1274) );
  XOR U2815 ( .A(n1277), .B(n1278), .Z(n1276) );
  XOR U2816 ( .A(DB[1195]), .B(DB[1188]), .Z(n1278) );
  AND U2817 ( .A(n346), .B(n1279), .Z(n1277) );
  XOR U2818 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U2819 ( .A(DB[1188]), .B(DB[1181]), .Z(n1281) );
  AND U2820 ( .A(n350), .B(n1282), .Z(n1280) );
  XOR U2821 ( .A(n1283), .B(n1284), .Z(n1282) );
  XOR U2822 ( .A(DB[1181]), .B(DB[1174]), .Z(n1284) );
  AND U2823 ( .A(n354), .B(n1285), .Z(n1283) );
  XOR U2824 ( .A(n1286), .B(n1287), .Z(n1285) );
  XOR U2825 ( .A(DB[1174]), .B(DB[1167]), .Z(n1287) );
  AND U2826 ( .A(n358), .B(n1288), .Z(n1286) );
  XOR U2827 ( .A(n1289), .B(n1290), .Z(n1288) );
  XOR U2828 ( .A(DB[1167]), .B(DB[1160]), .Z(n1290) );
  AND U2829 ( .A(n362), .B(n1291), .Z(n1289) );
  XOR U2830 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U2831 ( .A(DB[1160]), .B(DB[1153]), .Z(n1293) );
  AND U2832 ( .A(n366), .B(n1294), .Z(n1292) );
  XOR U2833 ( .A(n1295), .B(n1296), .Z(n1294) );
  XOR U2834 ( .A(DB[1153]), .B(DB[1146]), .Z(n1296) );
  AND U2835 ( .A(n370), .B(n1297), .Z(n1295) );
  XOR U2836 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U2837 ( .A(DB[1146]), .B(DB[1139]), .Z(n1299) );
  AND U2838 ( .A(n374), .B(n1300), .Z(n1298) );
  XOR U2839 ( .A(n1301), .B(n1302), .Z(n1300) );
  XOR U2840 ( .A(DB[1139]), .B(DB[1132]), .Z(n1302) );
  AND U2841 ( .A(n378), .B(n1303), .Z(n1301) );
  XOR U2842 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U2843 ( .A(DB[1132]), .B(DB[1125]), .Z(n1305) );
  AND U2844 ( .A(n382), .B(n1306), .Z(n1304) );
  XOR U2845 ( .A(n1307), .B(n1308), .Z(n1306) );
  XOR U2846 ( .A(DB[1125]), .B(DB[1118]), .Z(n1308) );
  AND U2847 ( .A(n386), .B(n1309), .Z(n1307) );
  XOR U2848 ( .A(n1310), .B(n1311), .Z(n1309) );
  XOR U2849 ( .A(DB[1118]), .B(DB[1111]), .Z(n1311) );
  AND U2850 ( .A(n390), .B(n1312), .Z(n1310) );
  XOR U2851 ( .A(n1313), .B(n1314), .Z(n1312) );
  XOR U2852 ( .A(DB[1111]), .B(DB[1104]), .Z(n1314) );
  AND U2853 ( .A(n394), .B(n1315), .Z(n1313) );
  XOR U2854 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U2855 ( .A(DB[1104]), .B(DB[1097]), .Z(n1317) );
  AND U2856 ( .A(n398), .B(n1318), .Z(n1316) );
  XOR U2857 ( .A(n1319), .B(n1320), .Z(n1318) );
  XOR U2858 ( .A(DB[1097]), .B(DB[1090]), .Z(n1320) );
  AND U2859 ( .A(n402), .B(n1321), .Z(n1319) );
  XOR U2860 ( .A(n1322), .B(n1323), .Z(n1321) );
  XOR U2861 ( .A(DB[1090]), .B(DB[1083]), .Z(n1323) );
  AND U2862 ( .A(n406), .B(n1324), .Z(n1322) );
  XOR U2863 ( .A(n1325), .B(n1326), .Z(n1324) );
  XOR U2864 ( .A(DB[1083]), .B(DB[1076]), .Z(n1326) );
  AND U2865 ( .A(n410), .B(n1327), .Z(n1325) );
  XOR U2866 ( .A(n1328), .B(n1329), .Z(n1327) );
  XOR U2867 ( .A(DB[1076]), .B(DB[1069]), .Z(n1329) );
  AND U2868 ( .A(n414), .B(n1330), .Z(n1328) );
  XOR U2869 ( .A(n1331), .B(n1332), .Z(n1330) );
  XOR U2870 ( .A(DB[1069]), .B(DB[1062]), .Z(n1332) );
  AND U2871 ( .A(n418), .B(n1333), .Z(n1331) );
  XOR U2872 ( .A(n1334), .B(n1335), .Z(n1333) );
  XOR U2873 ( .A(DB[1062]), .B(DB[1055]), .Z(n1335) );
  AND U2874 ( .A(n422), .B(n1336), .Z(n1334) );
  XOR U2875 ( .A(n1337), .B(n1338), .Z(n1336) );
  XOR U2876 ( .A(DB[1055]), .B(DB[1048]), .Z(n1338) );
  AND U2877 ( .A(n426), .B(n1339), .Z(n1337) );
  XOR U2878 ( .A(n1340), .B(n1341), .Z(n1339) );
  XOR U2879 ( .A(DB[1048]), .B(DB[1041]), .Z(n1341) );
  AND U2880 ( .A(n430), .B(n1342), .Z(n1340) );
  XOR U2881 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U2882 ( .A(DB[1041]), .B(DB[1034]), .Z(n1344) );
  AND U2883 ( .A(n434), .B(n1345), .Z(n1343) );
  XOR U2884 ( .A(n1346), .B(n1347), .Z(n1345) );
  XOR U2885 ( .A(DB[1034]), .B(DB[1027]), .Z(n1347) );
  AND U2886 ( .A(n438), .B(n1348), .Z(n1346) );
  XOR U2887 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U2888 ( .A(DB[1027]), .B(DB[1020]), .Z(n1350) );
  AND U2889 ( .A(n442), .B(n1351), .Z(n1349) );
  XOR U2890 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR U2891 ( .A(DB[1020]), .B(DB[1013]), .Z(n1353) );
  AND U2892 ( .A(n446), .B(n1354), .Z(n1352) );
  XOR U2893 ( .A(n1355), .B(n1356), .Z(n1354) );
  XOR U2894 ( .A(DB[1013]), .B(DB[1006]), .Z(n1356) );
  AND U2895 ( .A(n450), .B(n1357), .Z(n1355) );
  XOR U2896 ( .A(n1358), .B(n1359), .Z(n1357) );
  XOR U2897 ( .A(DB[999]), .B(DB[1006]), .Z(n1359) );
  AND U2898 ( .A(n454), .B(n1360), .Z(n1358) );
  XOR U2899 ( .A(n1361), .B(n1362), .Z(n1360) );
  XOR U2900 ( .A(DB[999]), .B(DB[992]), .Z(n1362) );
  AND U2901 ( .A(n458), .B(n1363), .Z(n1361) );
  XOR U2902 ( .A(n1364), .B(n1365), .Z(n1363) );
  XOR U2903 ( .A(DB[992]), .B(DB[985]), .Z(n1365) );
  AND U2904 ( .A(n462), .B(n1366), .Z(n1364) );
  XOR U2905 ( .A(n1367), .B(n1368), .Z(n1366) );
  XOR U2906 ( .A(DB[985]), .B(DB[978]), .Z(n1368) );
  AND U2907 ( .A(n466), .B(n1369), .Z(n1367) );
  XOR U2908 ( .A(n1370), .B(n1371), .Z(n1369) );
  XOR U2909 ( .A(DB[978]), .B(DB[971]), .Z(n1371) );
  AND U2910 ( .A(n470), .B(n1372), .Z(n1370) );
  XOR U2911 ( .A(n1373), .B(n1374), .Z(n1372) );
  XOR U2912 ( .A(DB[971]), .B(DB[964]), .Z(n1374) );
  AND U2913 ( .A(n474), .B(n1375), .Z(n1373) );
  XOR U2914 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U2915 ( .A(DB[964]), .B(DB[957]), .Z(n1377) );
  AND U2916 ( .A(n478), .B(n1378), .Z(n1376) );
  XOR U2917 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U2918 ( .A(DB[957]), .B(DB[950]), .Z(n1380) );
  AND U2919 ( .A(n482), .B(n1381), .Z(n1379) );
  XOR U2920 ( .A(n1382), .B(n1383), .Z(n1381) );
  XOR U2921 ( .A(DB[950]), .B(DB[943]), .Z(n1383) );
  AND U2922 ( .A(n486), .B(n1384), .Z(n1382) );
  XOR U2923 ( .A(n1385), .B(n1386), .Z(n1384) );
  XOR U2924 ( .A(DB[943]), .B(DB[936]), .Z(n1386) );
  AND U2925 ( .A(n490), .B(n1387), .Z(n1385) );
  XOR U2926 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U2927 ( .A(DB[936]), .B(DB[929]), .Z(n1389) );
  AND U2928 ( .A(n494), .B(n1390), .Z(n1388) );
  XOR U2929 ( .A(n1391), .B(n1392), .Z(n1390) );
  XOR U2930 ( .A(DB[929]), .B(DB[922]), .Z(n1392) );
  AND U2931 ( .A(n498), .B(n1393), .Z(n1391) );
  XOR U2932 ( .A(n1394), .B(n1395), .Z(n1393) );
  XOR U2933 ( .A(DB[922]), .B(DB[915]), .Z(n1395) );
  AND U2934 ( .A(n502), .B(n1396), .Z(n1394) );
  XOR U2935 ( .A(n1397), .B(n1398), .Z(n1396) );
  XOR U2936 ( .A(DB[915]), .B(DB[908]), .Z(n1398) );
  AND U2937 ( .A(n506), .B(n1399), .Z(n1397) );
  XOR U2938 ( .A(n1400), .B(n1401), .Z(n1399) );
  XOR U2939 ( .A(DB[908]), .B(DB[901]), .Z(n1401) );
  AND U2940 ( .A(n510), .B(n1402), .Z(n1400) );
  XOR U2941 ( .A(n1403), .B(n1404), .Z(n1402) );
  XOR U2942 ( .A(DB[901]), .B(DB[894]), .Z(n1404) );
  AND U2943 ( .A(n514), .B(n1405), .Z(n1403) );
  XOR U2944 ( .A(n1406), .B(n1407), .Z(n1405) );
  XOR U2945 ( .A(DB[894]), .B(DB[887]), .Z(n1407) );
  AND U2946 ( .A(n518), .B(n1408), .Z(n1406) );
  XOR U2947 ( .A(n1409), .B(n1410), .Z(n1408) );
  XOR U2948 ( .A(DB[887]), .B(DB[880]), .Z(n1410) );
  AND U2949 ( .A(n522), .B(n1411), .Z(n1409) );
  XOR U2950 ( .A(n1412), .B(n1413), .Z(n1411) );
  XOR U2951 ( .A(DB[880]), .B(DB[873]), .Z(n1413) );
  AND U2952 ( .A(n526), .B(n1414), .Z(n1412) );
  XOR U2953 ( .A(n1415), .B(n1416), .Z(n1414) );
  XOR U2954 ( .A(DB[873]), .B(DB[866]), .Z(n1416) );
  AND U2955 ( .A(n530), .B(n1417), .Z(n1415) );
  XOR U2956 ( .A(n1418), .B(n1419), .Z(n1417) );
  XOR U2957 ( .A(DB[866]), .B(DB[859]), .Z(n1419) );
  AND U2958 ( .A(n534), .B(n1420), .Z(n1418) );
  XOR U2959 ( .A(n1421), .B(n1422), .Z(n1420) );
  XOR U2960 ( .A(DB[859]), .B(DB[852]), .Z(n1422) );
  AND U2961 ( .A(n538), .B(n1423), .Z(n1421) );
  XOR U2962 ( .A(n1424), .B(n1425), .Z(n1423) );
  XOR U2963 ( .A(DB[852]), .B(DB[845]), .Z(n1425) );
  AND U2964 ( .A(n542), .B(n1426), .Z(n1424) );
  XOR U2965 ( .A(n1427), .B(n1428), .Z(n1426) );
  XOR U2966 ( .A(DB[845]), .B(DB[838]), .Z(n1428) );
  AND U2967 ( .A(n546), .B(n1429), .Z(n1427) );
  XOR U2968 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U2969 ( .A(DB[838]), .B(DB[831]), .Z(n1431) );
  AND U2970 ( .A(n550), .B(n1432), .Z(n1430) );
  XOR U2971 ( .A(n1433), .B(n1434), .Z(n1432) );
  XOR U2972 ( .A(DB[831]), .B(DB[824]), .Z(n1434) );
  AND U2973 ( .A(n554), .B(n1435), .Z(n1433) );
  XOR U2974 ( .A(n1436), .B(n1437), .Z(n1435) );
  XOR U2975 ( .A(DB[824]), .B(DB[817]), .Z(n1437) );
  AND U2976 ( .A(n558), .B(n1438), .Z(n1436) );
  XOR U2977 ( .A(n1439), .B(n1440), .Z(n1438) );
  XOR U2978 ( .A(DB[817]), .B(DB[810]), .Z(n1440) );
  AND U2979 ( .A(n562), .B(n1441), .Z(n1439) );
  XOR U2980 ( .A(n1442), .B(n1443), .Z(n1441) );
  XOR U2981 ( .A(DB[810]), .B(DB[803]), .Z(n1443) );
  AND U2982 ( .A(n566), .B(n1444), .Z(n1442) );
  XOR U2983 ( .A(n1445), .B(n1446), .Z(n1444) );
  XOR U2984 ( .A(DB[803]), .B(DB[796]), .Z(n1446) );
  AND U2985 ( .A(n570), .B(n1447), .Z(n1445) );
  XOR U2986 ( .A(n1448), .B(n1449), .Z(n1447) );
  XOR U2987 ( .A(DB[796]), .B(DB[789]), .Z(n1449) );
  AND U2988 ( .A(n574), .B(n1450), .Z(n1448) );
  XOR U2989 ( .A(n1451), .B(n1452), .Z(n1450) );
  XOR U2990 ( .A(DB[789]), .B(DB[782]), .Z(n1452) );
  AND U2991 ( .A(n578), .B(n1453), .Z(n1451) );
  XOR U2992 ( .A(n1454), .B(n1455), .Z(n1453) );
  XOR U2993 ( .A(DB[782]), .B(DB[775]), .Z(n1455) );
  AND U2994 ( .A(n582), .B(n1456), .Z(n1454) );
  XOR U2995 ( .A(n1457), .B(n1458), .Z(n1456) );
  XOR U2996 ( .A(DB[775]), .B(DB[768]), .Z(n1458) );
  AND U2997 ( .A(n586), .B(n1459), .Z(n1457) );
  XOR U2998 ( .A(n1460), .B(n1461), .Z(n1459) );
  XOR U2999 ( .A(DB[768]), .B(DB[761]), .Z(n1461) );
  AND U3000 ( .A(n590), .B(n1462), .Z(n1460) );
  XOR U3001 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U3002 ( .A(DB[761]), .B(DB[754]), .Z(n1464) );
  AND U3003 ( .A(n594), .B(n1465), .Z(n1463) );
  XOR U3004 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U3005 ( .A(DB[754]), .B(DB[747]), .Z(n1467) );
  AND U3006 ( .A(n598), .B(n1468), .Z(n1466) );
  XOR U3007 ( .A(n1469), .B(n1470), .Z(n1468) );
  XOR U3008 ( .A(DB[747]), .B(DB[740]), .Z(n1470) );
  AND U3009 ( .A(n602), .B(n1471), .Z(n1469) );
  XOR U3010 ( .A(n1472), .B(n1473), .Z(n1471) );
  XOR U3011 ( .A(DB[740]), .B(DB[733]), .Z(n1473) );
  AND U3012 ( .A(n606), .B(n1474), .Z(n1472) );
  XOR U3013 ( .A(n1475), .B(n1476), .Z(n1474) );
  XOR U3014 ( .A(DB[733]), .B(DB[726]), .Z(n1476) );
  AND U3015 ( .A(n610), .B(n1477), .Z(n1475) );
  XOR U3016 ( .A(n1478), .B(n1479), .Z(n1477) );
  XOR U3017 ( .A(DB[726]), .B(DB[719]), .Z(n1479) );
  AND U3018 ( .A(n614), .B(n1480), .Z(n1478) );
  XOR U3019 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U3020 ( .A(DB[719]), .B(DB[712]), .Z(n1482) );
  AND U3021 ( .A(n618), .B(n1483), .Z(n1481) );
  XOR U3022 ( .A(n1484), .B(n1485), .Z(n1483) );
  XOR U3023 ( .A(DB[712]), .B(DB[705]), .Z(n1485) );
  AND U3024 ( .A(n622), .B(n1486), .Z(n1484) );
  XOR U3025 ( .A(n1487), .B(n1488), .Z(n1486) );
  XOR U3026 ( .A(DB[705]), .B(DB[698]), .Z(n1488) );
  AND U3027 ( .A(n626), .B(n1489), .Z(n1487) );
  XOR U3028 ( .A(n1490), .B(n1491), .Z(n1489) );
  XOR U3029 ( .A(DB[698]), .B(DB[691]), .Z(n1491) );
  AND U3030 ( .A(n630), .B(n1492), .Z(n1490) );
  XOR U3031 ( .A(n1493), .B(n1494), .Z(n1492) );
  XOR U3032 ( .A(DB[691]), .B(DB[684]), .Z(n1494) );
  AND U3033 ( .A(n634), .B(n1495), .Z(n1493) );
  XOR U3034 ( .A(n1496), .B(n1497), .Z(n1495) );
  XOR U3035 ( .A(DB[684]), .B(DB[677]), .Z(n1497) );
  AND U3036 ( .A(n638), .B(n1498), .Z(n1496) );
  XOR U3037 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U3038 ( .A(DB[677]), .B(DB[670]), .Z(n1500) );
  AND U3039 ( .A(n642), .B(n1501), .Z(n1499) );
  XOR U3040 ( .A(n1502), .B(n1503), .Z(n1501) );
  XOR U3041 ( .A(DB[670]), .B(DB[663]), .Z(n1503) );
  AND U3042 ( .A(n646), .B(n1504), .Z(n1502) );
  XOR U3043 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U3044 ( .A(DB[663]), .B(DB[656]), .Z(n1506) );
  AND U3045 ( .A(n650), .B(n1507), .Z(n1505) );
  XOR U3046 ( .A(n1508), .B(n1509), .Z(n1507) );
  XOR U3047 ( .A(DB[656]), .B(DB[649]), .Z(n1509) );
  AND U3048 ( .A(n654), .B(n1510), .Z(n1508) );
  XOR U3049 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U3050 ( .A(DB[649]), .B(DB[642]), .Z(n1512) );
  AND U3051 ( .A(n658), .B(n1513), .Z(n1511) );
  XOR U3052 ( .A(n1514), .B(n1515), .Z(n1513) );
  XOR U3053 ( .A(DB[642]), .B(DB[635]), .Z(n1515) );
  AND U3054 ( .A(n662), .B(n1516), .Z(n1514) );
  XOR U3055 ( .A(n1517), .B(n1518), .Z(n1516) );
  XOR U3056 ( .A(DB[635]), .B(DB[628]), .Z(n1518) );
  AND U3057 ( .A(n666), .B(n1519), .Z(n1517) );
  XOR U3058 ( .A(n1520), .B(n1521), .Z(n1519) );
  XOR U3059 ( .A(DB[628]), .B(DB[621]), .Z(n1521) );
  AND U3060 ( .A(n670), .B(n1522), .Z(n1520) );
  XOR U3061 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U3062 ( .A(DB[621]), .B(DB[614]), .Z(n1524) );
  AND U3063 ( .A(n674), .B(n1525), .Z(n1523) );
  XOR U3064 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U3065 ( .A(DB[614]), .B(DB[607]), .Z(n1527) );
  AND U3066 ( .A(n678), .B(n1528), .Z(n1526) );
  XOR U3067 ( .A(n1529), .B(n1530), .Z(n1528) );
  XOR U3068 ( .A(DB[607]), .B(DB[600]), .Z(n1530) );
  AND U3069 ( .A(n682), .B(n1531), .Z(n1529) );
  XOR U3070 ( .A(n1532), .B(n1533), .Z(n1531) );
  XOR U3071 ( .A(DB[600]), .B(DB[593]), .Z(n1533) );
  AND U3072 ( .A(n686), .B(n1534), .Z(n1532) );
  XOR U3073 ( .A(n1535), .B(n1536), .Z(n1534) );
  XOR U3074 ( .A(DB[593]), .B(DB[586]), .Z(n1536) );
  AND U3075 ( .A(n690), .B(n1537), .Z(n1535) );
  XOR U3076 ( .A(n1538), .B(n1539), .Z(n1537) );
  XOR U3077 ( .A(DB[586]), .B(DB[579]), .Z(n1539) );
  AND U3078 ( .A(n694), .B(n1540), .Z(n1538) );
  XOR U3079 ( .A(n1541), .B(n1542), .Z(n1540) );
  XOR U3080 ( .A(DB[579]), .B(DB[572]), .Z(n1542) );
  AND U3081 ( .A(n698), .B(n1543), .Z(n1541) );
  XOR U3082 ( .A(n1544), .B(n1545), .Z(n1543) );
  XOR U3083 ( .A(DB[572]), .B(DB[565]), .Z(n1545) );
  AND U3084 ( .A(n702), .B(n1546), .Z(n1544) );
  XOR U3085 ( .A(n1547), .B(n1548), .Z(n1546) );
  XOR U3086 ( .A(DB[565]), .B(DB[558]), .Z(n1548) );
  AND U3087 ( .A(n706), .B(n1549), .Z(n1547) );
  XOR U3088 ( .A(n1550), .B(n1551), .Z(n1549) );
  XOR U3089 ( .A(DB[558]), .B(DB[551]), .Z(n1551) );
  AND U3090 ( .A(n710), .B(n1552), .Z(n1550) );
  XOR U3091 ( .A(n1553), .B(n1554), .Z(n1552) );
  XOR U3092 ( .A(DB[551]), .B(DB[544]), .Z(n1554) );
  AND U3093 ( .A(n714), .B(n1555), .Z(n1553) );
  XOR U3094 ( .A(n1556), .B(n1557), .Z(n1555) );
  XOR U3095 ( .A(DB[544]), .B(DB[537]), .Z(n1557) );
  AND U3096 ( .A(n718), .B(n1558), .Z(n1556) );
  XOR U3097 ( .A(n1559), .B(n1560), .Z(n1558) );
  XOR U3098 ( .A(DB[537]), .B(DB[530]), .Z(n1560) );
  AND U3099 ( .A(n722), .B(n1561), .Z(n1559) );
  XOR U3100 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U3101 ( .A(DB[530]), .B(DB[523]), .Z(n1563) );
  AND U3102 ( .A(n726), .B(n1564), .Z(n1562) );
  XOR U3103 ( .A(n1565), .B(n1566), .Z(n1564) );
  XOR U3104 ( .A(DB[523]), .B(DB[516]), .Z(n1566) );
  AND U3105 ( .A(n730), .B(n1567), .Z(n1565) );
  XOR U3106 ( .A(n1568), .B(n1569), .Z(n1567) );
  XOR U3107 ( .A(DB[516]), .B(DB[509]), .Z(n1569) );
  AND U3108 ( .A(n734), .B(n1570), .Z(n1568) );
  XOR U3109 ( .A(n1571), .B(n1572), .Z(n1570) );
  XOR U3110 ( .A(DB[509]), .B(DB[502]), .Z(n1572) );
  AND U3111 ( .A(n738), .B(n1573), .Z(n1571) );
  XOR U3112 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U3113 ( .A(DB[502]), .B(DB[495]), .Z(n1575) );
  AND U3114 ( .A(n742), .B(n1576), .Z(n1574) );
  XOR U3115 ( .A(n1577), .B(n1578), .Z(n1576) );
  XOR U3116 ( .A(DB[495]), .B(DB[488]), .Z(n1578) );
  AND U3117 ( .A(n746), .B(n1579), .Z(n1577) );
  XOR U3118 ( .A(n1580), .B(n1581), .Z(n1579) );
  XOR U3119 ( .A(DB[488]), .B(DB[481]), .Z(n1581) );
  AND U3120 ( .A(n750), .B(n1582), .Z(n1580) );
  XOR U3121 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U3122 ( .A(DB[481]), .B(DB[474]), .Z(n1584) );
  AND U3123 ( .A(n754), .B(n1585), .Z(n1583) );
  XOR U3124 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U3125 ( .A(DB[474]), .B(DB[467]), .Z(n1587) );
  AND U3126 ( .A(n758), .B(n1588), .Z(n1586) );
  XOR U3127 ( .A(n1589), .B(n1590), .Z(n1588) );
  XOR U3128 ( .A(DB[467]), .B(DB[460]), .Z(n1590) );
  AND U3129 ( .A(n762), .B(n1591), .Z(n1589) );
  XOR U3130 ( .A(n1592), .B(n1593), .Z(n1591) );
  XOR U3131 ( .A(DB[460]), .B(DB[453]), .Z(n1593) );
  AND U3132 ( .A(n766), .B(n1594), .Z(n1592) );
  XOR U3133 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U3134 ( .A(DB[453]), .B(DB[446]), .Z(n1596) );
  AND U3135 ( .A(n770), .B(n1597), .Z(n1595) );
  XOR U3136 ( .A(n1598), .B(n1599), .Z(n1597) );
  XOR U3137 ( .A(DB[446]), .B(DB[439]), .Z(n1599) );
  AND U3138 ( .A(n774), .B(n1600), .Z(n1598) );
  XOR U3139 ( .A(n1601), .B(n1602), .Z(n1600) );
  XOR U3140 ( .A(DB[439]), .B(DB[432]), .Z(n1602) );
  AND U3141 ( .A(n778), .B(n1603), .Z(n1601) );
  XOR U3142 ( .A(n1604), .B(n1605), .Z(n1603) );
  XOR U3143 ( .A(DB[432]), .B(DB[425]), .Z(n1605) );
  AND U3144 ( .A(n782), .B(n1606), .Z(n1604) );
  XOR U3145 ( .A(n1607), .B(n1608), .Z(n1606) );
  XOR U3146 ( .A(DB[425]), .B(DB[418]), .Z(n1608) );
  AND U3147 ( .A(n786), .B(n1609), .Z(n1607) );
  XOR U3148 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U3149 ( .A(DB[418]), .B(DB[411]), .Z(n1611) );
  AND U3150 ( .A(n790), .B(n1612), .Z(n1610) );
  XOR U3151 ( .A(n1613), .B(n1614), .Z(n1612) );
  XOR U3152 ( .A(DB[411]), .B(DB[404]), .Z(n1614) );
  AND U3153 ( .A(n794), .B(n1615), .Z(n1613) );
  XOR U3154 ( .A(n1616), .B(n1617), .Z(n1615) );
  XOR U3155 ( .A(DB[404]), .B(DB[397]), .Z(n1617) );
  AND U3156 ( .A(n798), .B(n1618), .Z(n1616) );
  XOR U3157 ( .A(n1619), .B(n1620), .Z(n1618) );
  XOR U3158 ( .A(DB[397]), .B(DB[390]), .Z(n1620) );
  AND U3159 ( .A(n802), .B(n1621), .Z(n1619) );
  XOR U3160 ( .A(n1622), .B(n1623), .Z(n1621) );
  XOR U3161 ( .A(DB[390]), .B(DB[383]), .Z(n1623) );
  AND U3162 ( .A(n806), .B(n1624), .Z(n1622) );
  XOR U3163 ( .A(n1625), .B(n1626), .Z(n1624) );
  XOR U3164 ( .A(DB[383]), .B(DB[376]), .Z(n1626) );
  AND U3165 ( .A(n810), .B(n1627), .Z(n1625) );
  XOR U3166 ( .A(n1628), .B(n1629), .Z(n1627) );
  XOR U3167 ( .A(DB[376]), .B(DB[369]), .Z(n1629) );
  AND U3168 ( .A(n814), .B(n1630), .Z(n1628) );
  XOR U3169 ( .A(n1631), .B(n1632), .Z(n1630) );
  XOR U3170 ( .A(DB[369]), .B(DB[362]), .Z(n1632) );
  AND U3171 ( .A(n818), .B(n1633), .Z(n1631) );
  XOR U3172 ( .A(n1634), .B(n1635), .Z(n1633) );
  XOR U3173 ( .A(DB[362]), .B(DB[355]), .Z(n1635) );
  AND U3174 ( .A(n822), .B(n1636), .Z(n1634) );
  XOR U3175 ( .A(n1637), .B(n1638), .Z(n1636) );
  XOR U3176 ( .A(DB[355]), .B(DB[348]), .Z(n1638) );
  AND U3177 ( .A(n826), .B(n1639), .Z(n1637) );
  XOR U3178 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U3179 ( .A(DB[348]), .B(DB[341]), .Z(n1641) );
  AND U3180 ( .A(n830), .B(n1642), .Z(n1640) );
  XOR U3181 ( .A(n1643), .B(n1644), .Z(n1642) );
  XOR U3182 ( .A(DB[341]), .B(DB[334]), .Z(n1644) );
  AND U3183 ( .A(n834), .B(n1645), .Z(n1643) );
  XOR U3184 ( .A(n1646), .B(n1647), .Z(n1645) );
  XOR U3185 ( .A(DB[334]), .B(DB[327]), .Z(n1647) );
  AND U3186 ( .A(n838), .B(n1648), .Z(n1646) );
  XOR U3187 ( .A(n1649), .B(n1650), .Z(n1648) );
  XOR U3188 ( .A(DB[327]), .B(DB[320]), .Z(n1650) );
  AND U3189 ( .A(n842), .B(n1651), .Z(n1649) );
  XOR U3190 ( .A(n1652), .B(n1653), .Z(n1651) );
  XOR U3191 ( .A(DB[320]), .B(DB[313]), .Z(n1653) );
  AND U3192 ( .A(n846), .B(n1654), .Z(n1652) );
  XOR U3193 ( .A(n1655), .B(n1656), .Z(n1654) );
  XOR U3194 ( .A(DB[313]), .B(DB[306]), .Z(n1656) );
  AND U3195 ( .A(n850), .B(n1657), .Z(n1655) );
  XOR U3196 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U3197 ( .A(DB[306]), .B(DB[299]), .Z(n1659) );
  AND U3198 ( .A(n854), .B(n1660), .Z(n1658) );
  XOR U3199 ( .A(n1661), .B(n1662), .Z(n1660) );
  XOR U3200 ( .A(DB[299]), .B(DB[292]), .Z(n1662) );
  AND U3201 ( .A(n858), .B(n1663), .Z(n1661) );
  XOR U3202 ( .A(n1664), .B(n1665), .Z(n1663) );
  XOR U3203 ( .A(DB[292]), .B(DB[285]), .Z(n1665) );
  AND U3204 ( .A(n862), .B(n1666), .Z(n1664) );
  XOR U3205 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U3206 ( .A(DB[285]), .B(DB[278]), .Z(n1668) );
  AND U3207 ( .A(n866), .B(n1669), .Z(n1667) );
  XOR U3208 ( .A(n1670), .B(n1671), .Z(n1669) );
  XOR U3209 ( .A(DB[278]), .B(DB[271]), .Z(n1671) );
  AND U3210 ( .A(n870), .B(n1672), .Z(n1670) );
  XOR U3211 ( .A(n1673), .B(n1674), .Z(n1672) );
  XOR U3212 ( .A(DB[271]), .B(DB[264]), .Z(n1674) );
  AND U3213 ( .A(n874), .B(n1675), .Z(n1673) );
  XOR U3214 ( .A(n1676), .B(n1677), .Z(n1675) );
  XOR U3215 ( .A(DB[264]), .B(DB[257]), .Z(n1677) );
  AND U3216 ( .A(n878), .B(n1678), .Z(n1676) );
  XOR U3217 ( .A(n1679), .B(n1680), .Z(n1678) );
  XOR U3218 ( .A(DB[257]), .B(DB[250]), .Z(n1680) );
  AND U3219 ( .A(n882), .B(n1681), .Z(n1679) );
  XOR U3220 ( .A(n1682), .B(n1683), .Z(n1681) );
  XOR U3221 ( .A(DB[250]), .B(DB[243]), .Z(n1683) );
  AND U3222 ( .A(n886), .B(n1684), .Z(n1682) );
  XOR U3223 ( .A(n1685), .B(n1686), .Z(n1684) );
  XOR U3224 ( .A(DB[243]), .B(DB[236]), .Z(n1686) );
  AND U3225 ( .A(n890), .B(n1687), .Z(n1685) );
  XOR U3226 ( .A(n1688), .B(n1689), .Z(n1687) );
  XOR U3227 ( .A(DB[236]), .B(DB[229]), .Z(n1689) );
  AND U3228 ( .A(n894), .B(n1690), .Z(n1688) );
  XOR U3229 ( .A(n1691), .B(n1692), .Z(n1690) );
  XOR U3230 ( .A(DB[229]), .B(DB[222]), .Z(n1692) );
  AND U3231 ( .A(n898), .B(n1693), .Z(n1691) );
  XOR U3232 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U3233 ( .A(DB[222]), .B(DB[215]), .Z(n1695) );
  AND U3234 ( .A(n902), .B(n1696), .Z(n1694) );
  XOR U3235 ( .A(n1697), .B(n1698), .Z(n1696) );
  XOR U3236 ( .A(DB[215]), .B(DB[208]), .Z(n1698) );
  AND U3237 ( .A(n906), .B(n1699), .Z(n1697) );
  XOR U3238 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U3239 ( .A(DB[208]), .B(DB[201]), .Z(n1701) );
  AND U3240 ( .A(n910), .B(n1702), .Z(n1700) );
  XOR U3241 ( .A(n1703), .B(n1704), .Z(n1702) );
  XOR U3242 ( .A(DB[201]), .B(DB[194]), .Z(n1704) );
  AND U3243 ( .A(n914), .B(n1705), .Z(n1703) );
  XOR U3244 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U3245 ( .A(DB[194]), .B(DB[187]), .Z(n1707) );
  AND U3246 ( .A(n918), .B(n1708), .Z(n1706) );
  XOR U3247 ( .A(n1709), .B(n1710), .Z(n1708) );
  XOR U3248 ( .A(DB[187]), .B(DB[180]), .Z(n1710) );
  AND U3249 ( .A(n922), .B(n1711), .Z(n1709) );
  XOR U3250 ( .A(n1712), .B(n1713), .Z(n1711) );
  XOR U3251 ( .A(DB[180]), .B(DB[173]), .Z(n1713) );
  AND U3252 ( .A(n926), .B(n1714), .Z(n1712) );
  XOR U3253 ( .A(n1715), .B(n1716), .Z(n1714) );
  XOR U3254 ( .A(DB[173]), .B(DB[166]), .Z(n1716) );
  AND U3255 ( .A(n930), .B(n1717), .Z(n1715) );
  XOR U3256 ( .A(n1718), .B(n1719), .Z(n1717) );
  XOR U3257 ( .A(DB[166]), .B(DB[159]), .Z(n1719) );
  AND U3258 ( .A(n934), .B(n1720), .Z(n1718) );
  XOR U3259 ( .A(n1721), .B(n1722), .Z(n1720) );
  XOR U3260 ( .A(DB[159]), .B(DB[152]), .Z(n1722) );
  AND U3261 ( .A(n938), .B(n1723), .Z(n1721) );
  XOR U3262 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U3263 ( .A(DB[152]), .B(DB[145]), .Z(n1725) );
  AND U3264 ( .A(n942), .B(n1726), .Z(n1724) );
  XOR U3265 ( .A(n1727), .B(n1728), .Z(n1726) );
  XOR U3266 ( .A(DB[145]), .B(DB[138]), .Z(n1728) );
  AND U3267 ( .A(n946), .B(n1729), .Z(n1727) );
  XOR U3268 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U3269 ( .A(DB[138]), .B(DB[131]), .Z(n1731) );
  AND U3270 ( .A(n950), .B(n1732), .Z(n1730) );
  XOR U3271 ( .A(n1733), .B(n1734), .Z(n1732) );
  XOR U3272 ( .A(DB[131]), .B(DB[124]), .Z(n1734) );
  AND U3273 ( .A(n954), .B(n1735), .Z(n1733) );
  XOR U3274 ( .A(n1736), .B(n1737), .Z(n1735) );
  XOR U3275 ( .A(DB[124]), .B(DB[117]), .Z(n1737) );
  AND U3276 ( .A(n958), .B(n1738), .Z(n1736) );
  XOR U3277 ( .A(n1739), .B(n1740), .Z(n1738) );
  XOR U3278 ( .A(DB[117]), .B(DB[110]), .Z(n1740) );
  AND U3279 ( .A(n962), .B(n1741), .Z(n1739) );
  XOR U3280 ( .A(n1742), .B(n1743), .Z(n1741) );
  XOR U3281 ( .A(DB[110]), .B(DB[103]), .Z(n1743) );
  AND U3282 ( .A(n966), .B(n1744), .Z(n1742) );
  XOR U3283 ( .A(n1745), .B(n1746), .Z(n1744) );
  XOR U3284 ( .A(DB[96]), .B(DB[103]), .Z(n1746) );
  AND U3285 ( .A(n970), .B(n1747), .Z(n1745) );
  XOR U3286 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U3287 ( .A(DB[96]), .B(DB[89]), .Z(n1749) );
  AND U3288 ( .A(n974), .B(n1750), .Z(n1748) );
  XOR U3289 ( .A(n1751), .B(n1752), .Z(n1750) );
  XOR U3290 ( .A(DB[89]), .B(DB[82]), .Z(n1752) );
  AND U3291 ( .A(n978), .B(n1753), .Z(n1751) );
  XOR U3292 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U3293 ( .A(DB[82]), .B(DB[75]), .Z(n1755) );
  AND U3294 ( .A(n982), .B(n1756), .Z(n1754) );
  XOR U3295 ( .A(n1757), .B(n1758), .Z(n1756) );
  XOR U3296 ( .A(DB[75]), .B(DB[68]), .Z(n1758) );
  AND U3297 ( .A(n986), .B(n1759), .Z(n1757) );
  XOR U3298 ( .A(n1760), .B(n1761), .Z(n1759) );
  XOR U3299 ( .A(DB[68]), .B(DB[61]), .Z(n1761) );
  AND U3300 ( .A(n990), .B(n1762), .Z(n1760) );
  XOR U3301 ( .A(n1763), .B(n1764), .Z(n1762) );
  XOR U3302 ( .A(DB[61]), .B(DB[54]), .Z(n1764) );
  AND U3303 ( .A(n994), .B(n1765), .Z(n1763) );
  XOR U3304 ( .A(n1766), .B(n1767), .Z(n1765) );
  XOR U3305 ( .A(DB[54]), .B(DB[47]), .Z(n1767) );
  AND U3306 ( .A(n998), .B(n1768), .Z(n1766) );
  XOR U3307 ( .A(n1769), .B(n1770), .Z(n1768) );
  XOR U3308 ( .A(DB[47]), .B(DB[40]), .Z(n1770) );
  AND U3309 ( .A(n1002), .B(n1771), .Z(n1769) );
  XOR U3310 ( .A(n1772), .B(n1773), .Z(n1771) );
  XOR U3311 ( .A(DB[40]), .B(DB[33]), .Z(n1773) );
  AND U3312 ( .A(n1006), .B(n1774), .Z(n1772) );
  XOR U3313 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U3314 ( .A(DB[33]), .B(DB[26]), .Z(n1776) );
  AND U3315 ( .A(n1010), .B(n1777), .Z(n1775) );
  XOR U3316 ( .A(n1778), .B(n1779), .Z(n1777) );
  XOR U3317 ( .A(DB[26]), .B(DB[19]), .Z(n1779) );
  AND U3318 ( .A(n1014), .B(n1780), .Z(n1778) );
  XOR U3319 ( .A(n1781), .B(n1782), .Z(n1780) );
  XOR U3320 ( .A(DB[19]), .B(DB[12]), .Z(n1782) );
  AND U3321 ( .A(n1018), .B(n1783), .Z(n1781) );
  XOR U3322 ( .A(DB[5]), .B(DB[12]), .Z(n1783) );
  XOR U3323 ( .A(DB[1789]), .B(n1784), .Z(min_val_out[4]) );
  AND U3324 ( .A(n2), .B(n1785), .Z(n1784) );
  XOR U3325 ( .A(n1786), .B(n1787), .Z(n1785) );
  XOR U3326 ( .A(DB[1789]), .B(DB[1782]), .Z(n1787) );
  AND U3327 ( .A(n6), .B(n1788), .Z(n1786) );
  XOR U3328 ( .A(n1789), .B(n1790), .Z(n1788) );
  XOR U3329 ( .A(DB[1782]), .B(DB[1775]), .Z(n1790) );
  AND U3330 ( .A(n10), .B(n1791), .Z(n1789) );
  XOR U3331 ( .A(n1792), .B(n1793), .Z(n1791) );
  XOR U3332 ( .A(DB[1775]), .B(DB[1768]), .Z(n1793) );
  AND U3333 ( .A(n14), .B(n1794), .Z(n1792) );
  XOR U3334 ( .A(n1795), .B(n1796), .Z(n1794) );
  XOR U3335 ( .A(DB[1768]), .B(DB[1761]), .Z(n1796) );
  AND U3336 ( .A(n18), .B(n1797), .Z(n1795) );
  XOR U3337 ( .A(n1798), .B(n1799), .Z(n1797) );
  XOR U3338 ( .A(DB[1761]), .B(DB[1754]), .Z(n1799) );
  AND U3339 ( .A(n22), .B(n1800), .Z(n1798) );
  XOR U3340 ( .A(n1801), .B(n1802), .Z(n1800) );
  XOR U3341 ( .A(DB[1754]), .B(DB[1747]), .Z(n1802) );
  AND U3342 ( .A(n26), .B(n1803), .Z(n1801) );
  XOR U3343 ( .A(n1804), .B(n1805), .Z(n1803) );
  XOR U3344 ( .A(DB[1747]), .B(DB[1740]), .Z(n1805) );
  AND U3345 ( .A(n30), .B(n1806), .Z(n1804) );
  XOR U3346 ( .A(n1807), .B(n1808), .Z(n1806) );
  XOR U3347 ( .A(DB[1740]), .B(DB[1733]), .Z(n1808) );
  AND U3348 ( .A(n34), .B(n1809), .Z(n1807) );
  XOR U3349 ( .A(n1810), .B(n1811), .Z(n1809) );
  XOR U3350 ( .A(DB[1733]), .B(DB[1726]), .Z(n1811) );
  AND U3351 ( .A(n38), .B(n1812), .Z(n1810) );
  XOR U3352 ( .A(n1813), .B(n1814), .Z(n1812) );
  XOR U3353 ( .A(DB[1726]), .B(DB[1719]), .Z(n1814) );
  AND U3354 ( .A(n42), .B(n1815), .Z(n1813) );
  XOR U3355 ( .A(n1816), .B(n1817), .Z(n1815) );
  XOR U3356 ( .A(DB[1719]), .B(DB[1712]), .Z(n1817) );
  AND U3357 ( .A(n46), .B(n1818), .Z(n1816) );
  XOR U3358 ( .A(n1819), .B(n1820), .Z(n1818) );
  XOR U3359 ( .A(DB[1712]), .B(DB[1705]), .Z(n1820) );
  AND U3360 ( .A(n50), .B(n1821), .Z(n1819) );
  XOR U3361 ( .A(n1822), .B(n1823), .Z(n1821) );
  XOR U3362 ( .A(DB[1705]), .B(DB[1698]), .Z(n1823) );
  AND U3363 ( .A(n54), .B(n1824), .Z(n1822) );
  XOR U3364 ( .A(n1825), .B(n1826), .Z(n1824) );
  XOR U3365 ( .A(DB[1698]), .B(DB[1691]), .Z(n1826) );
  AND U3366 ( .A(n58), .B(n1827), .Z(n1825) );
  XOR U3367 ( .A(n1828), .B(n1829), .Z(n1827) );
  XOR U3368 ( .A(DB[1691]), .B(DB[1684]), .Z(n1829) );
  AND U3369 ( .A(n62), .B(n1830), .Z(n1828) );
  XOR U3370 ( .A(n1831), .B(n1832), .Z(n1830) );
  XOR U3371 ( .A(DB[1684]), .B(DB[1677]), .Z(n1832) );
  AND U3372 ( .A(n66), .B(n1833), .Z(n1831) );
  XOR U3373 ( .A(n1834), .B(n1835), .Z(n1833) );
  XOR U3374 ( .A(DB[1677]), .B(DB[1670]), .Z(n1835) );
  AND U3375 ( .A(n70), .B(n1836), .Z(n1834) );
  XOR U3376 ( .A(n1837), .B(n1838), .Z(n1836) );
  XOR U3377 ( .A(DB[1670]), .B(DB[1663]), .Z(n1838) );
  AND U3378 ( .A(n74), .B(n1839), .Z(n1837) );
  XOR U3379 ( .A(n1840), .B(n1841), .Z(n1839) );
  XOR U3380 ( .A(DB[1663]), .B(DB[1656]), .Z(n1841) );
  AND U3381 ( .A(n78), .B(n1842), .Z(n1840) );
  XOR U3382 ( .A(n1843), .B(n1844), .Z(n1842) );
  XOR U3383 ( .A(DB[1656]), .B(DB[1649]), .Z(n1844) );
  AND U3384 ( .A(n82), .B(n1845), .Z(n1843) );
  XOR U3385 ( .A(n1846), .B(n1847), .Z(n1845) );
  XOR U3386 ( .A(DB[1649]), .B(DB[1642]), .Z(n1847) );
  AND U3387 ( .A(n86), .B(n1848), .Z(n1846) );
  XOR U3388 ( .A(n1849), .B(n1850), .Z(n1848) );
  XOR U3389 ( .A(DB[1642]), .B(DB[1635]), .Z(n1850) );
  AND U3390 ( .A(n90), .B(n1851), .Z(n1849) );
  XOR U3391 ( .A(n1852), .B(n1853), .Z(n1851) );
  XOR U3392 ( .A(DB[1635]), .B(DB[1628]), .Z(n1853) );
  AND U3393 ( .A(n94), .B(n1854), .Z(n1852) );
  XOR U3394 ( .A(n1855), .B(n1856), .Z(n1854) );
  XOR U3395 ( .A(DB[1628]), .B(DB[1621]), .Z(n1856) );
  AND U3396 ( .A(n98), .B(n1857), .Z(n1855) );
  XOR U3397 ( .A(n1858), .B(n1859), .Z(n1857) );
  XOR U3398 ( .A(DB[1621]), .B(DB[1614]), .Z(n1859) );
  AND U3399 ( .A(n102), .B(n1860), .Z(n1858) );
  XOR U3400 ( .A(n1861), .B(n1862), .Z(n1860) );
  XOR U3401 ( .A(DB[1614]), .B(DB[1607]), .Z(n1862) );
  AND U3402 ( .A(n106), .B(n1863), .Z(n1861) );
  XOR U3403 ( .A(n1864), .B(n1865), .Z(n1863) );
  XOR U3404 ( .A(DB[1607]), .B(DB[1600]), .Z(n1865) );
  AND U3405 ( .A(n110), .B(n1866), .Z(n1864) );
  XOR U3406 ( .A(n1867), .B(n1868), .Z(n1866) );
  XOR U3407 ( .A(DB[1600]), .B(DB[1593]), .Z(n1868) );
  AND U3408 ( .A(n114), .B(n1869), .Z(n1867) );
  XOR U3409 ( .A(n1870), .B(n1871), .Z(n1869) );
  XOR U3410 ( .A(DB[1593]), .B(DB[1586]), .Z(n1871) );
  AND U3411 ( .A(n118), .B(n1872), .Z(n1870) );
  XOR U3412 ( .A(n1873), .B(n1874), .Z(n1872) );
  XOR U3413 ( .A(DB[1586]), .B(DB[1579]), .Z(n1874) );
  AND U3414 ( .A(n122), .B(n1875), .Z(n1873) );
  XOR U3415 ( .A(n1876), .B(n1877), .Z(n1875) );
  XOR U3416 ( .A(DB[1579]), .B(DB[1572]), .Z(n1877) );
  AND U3417 ( .A(n126), .B(n1878), .Z(n1876) );
  XOR U3418 ( .A(n1879), .B(n1880), .Z(n1878) );
  XOR U3419 ( .A(DB[1572]), .B(DB[1565]), .Z(n1880) );
  AND U3420 ( .A(n130), .B(n1881), .Z(n1879) );
  XOR U3421 ( .A(n1882), .B(n1883), .Z(n1881) );
  XOR U3422 ( .A(DB[1565]), .B(DB[1558]), .Z(n1883) );
  AND U3423 ( .A(n134), .B(n1884), .Z(n1882) );
  XOR U3424 ( .A(n1885), .B(n1886), .Z(n1884) );
  XOR U3425 ( .A(DB[1558]), .B(DB[1551]), .Z(n1886) );
  AND U3426 ( .A(n138), .B(n1887), .Z(n1885) );
  XOR U3427 ( .A(n1888), .B(n1889), .Z(n1887) );
  XOR U3428 ( .A(DB[1551]), .B(DB[1544]), .Z(n1889) );
  AND U3429 ( .A(n142), .B(n1890), .Z(n1888) );
  XOR U3430 ( .A(n1891), .B(n1892), .Z(n1890) );
  XOR U3431 ( .A(DB[1544]), .B(DB[1537]), .Z(n1892) );
  AND U3432 ( .A(n146), .B(n1893), .Z(n1891) );
  XOR U3433 ( .A(n1894), .B(n1895), .Z(n1893) );
  XOR U3434 ( .A(DB[1537]), .B(DB[1530]), .Z(n1895) );
  AND U3435 ( .A(n150), .B(n1896), .Z(n1894) );
  XOR U3436 ( .A(n1897), .B(n1898), .Z(n1896) );
  XOR U3437 ( .A(DB[1530]), .B(DB[1523]), .Z(n1898) );
  AND U3438 ( .A(n154), .B(n1899), .Z(n1897) );
  XOR U3439 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U3440 ( .A(DB[1523]), .B(DB[1516]), .Z(n1901) );
  AND U3441 ( .A(n158), .B(n1902), .Z(n1900) );
  XOR U3442 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U3443 ( .A(DB[1516]), .B(DB[1509]), .Z(n1904) );
  AND U3444 ( .A(n162), .B(n1905), .Z(n1903) );
  XOR U3445 ( .A(n1906), .B(n1907), .Z(n1905) );
  XOR U3446 ( .A(DB[1509]), .B(DB[1502]), .Z(n1907) );
  AND U3447 ( .A(n166), .B(n1908), .Z(n1906) );
  XOR U3448 ( .A(n1909), .B(n1910), .Z(n1908) );
  XOR U3449 ( .A(DB[1502]), .B(DB[1495]), .Z(n1910) );
  AND U3450 ( .A(n170), .B(n1911), .Z(n1909) );
  XOR U3451 ( .A(n1912), .B(n1913), .Z(n1911) );
  XOR U3452 ( .A(DB[1495]), .B(DB[1488]), .Z(n1913) );
  AND U3453 ( .A(n174), .B(n1914), .Z(n1912) );
  XOR U3454 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR U3455 ( .A(DB[1488]), .B(DB[1481]), .Z(n1916) );
  AND U3456 ( .A(n178), .B(n1917), .Z(n1915) );
  XOR U3457 ( .A(n1918), .B(n1919), .Z(n1917) );
  XOR U3458 ( .A(DB[1481]), .B(DB[1474]), .Z(n1919) );
  AND U3459 ( .A(n182), .B(n1920), .Z(n1918) );
  XOR U3460 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U3461 ( .A(DB[1474]), .B(DB[1467]), .Z(n1922) );
  AND U3462 ( .A(n186), .B(n1923), .Z(n1921) );
  XOR U3463 ( .A(n1924), .B(n1925), .Z(n1923) );
  XOR U3464 ( .A(DB[1467]), .B(DB[1460]), .Z(n1925) );
  AND U3465 ( .A(n190), .B(n1926), .Z(n1924) );
  XOR U3466 ( .A(n1927), .B(n1928), .Z(n1926) );
  XOR U3467 ( .A(DB[1460]), .B(DB[1453]), .Z(n1928) );
  AND U3468 ( .A(n194), .B(n1929), .Z(n1927) );
  XOR U3469 ( .A(n1930), .B(n1931), .Z(n1929) );
  XOR U3470 ( .A(DB[1453]), .B(DB[1446]), .Z(n1931) );
  AND U3471 ( .A(n198), .B(n1932), .Z(n1930) );
  XOR U3472 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U3473 ( .A(DB[1446]), .B(DB[1439]), .Z(n1934) );
  AND U3474 ( .A(n202), .B(n1935), .Z(n1933) );
  XOR U3475 ( .A(n1936), .B(n1937), .Z(n1935) );
  XOR U3476 ( .A(DB[1439]), .B(DB[1432]), .Z(n1937) );
  AND U3477 ( .A(n206), .B(n1938), .Z(n1936) );
  XOR U3478 ( .A(n1939), .B(n1940), .Z(n1938) );
  XOR U3479 ( .A(DB[1432]), .B(DB[1425]), .Z(n1940) );
  AND U3480 ( .A(n210), .B(n1941), .Z(n1939) );
  XOR U3481 ( .A(n1942), .B(n1943), .Z(n1941) );
  XOR U3482 ( .A(DB[1425]), .B(DB[1418]), .Z(n1943) );
  AND U3483 ( .A(n214), .B(n1944), .Z(n1942) );
  XOR U3484 ( .A(n1945), .B(n1946), .Z(n1944) );
  XOR U3485 ( .A(DB[1418]), .B(DB[1411]), .Z(n1946) );
  AND U3486 ( .A(n218), .B(n1947), .Z(n1945) );
  XOR U3487 ( .A(n1948), .B(n1949), .Z(n1947) );
  XOR U3488 ( .A(DB[1411]), .B(DB[1404]), .Z(n1949) );
  AND U3489 ( .A(n222), .B(n1950), .Z(n1948) );
  XOR U3490 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U3491 ( .A(DB[1404]), .B(DB[1397]), .Z(n1952) );
  AND U3492 ( .A(n226), .B(n1953), .Z(n1951) );
  XOR U3493 ( .A(n1954), .B(n1955), .Z(n1953) );
  XOR U3494 ( .A(DB[1397]), .B(DB[1390]), .Z(n1955) );
  AND U3495 ( .A(n230), .B(n1956), .Z(n1954) );
  XOR U3496 ( .A(n1957), .B(n1958), .Z(n1956) );
  XOR U3497 ( .A(DB[1390]), .B(DB[1383]), .Z(n1958) );
  AND U3498 ( .A(n234), .B(n1959), .Z(n1957) );
  XOR U3499 ( .A(n1960), .B(n1961), .Z(n1959) );
  XOR U3500 ( .A(DB[1383]), .B(DB[1376]), .Z(n1961) );
  AND U3501 ( .A(n238), .B(n1962), .Z(n1960) );
  XOR U3502 ( .A(n1963), .B(n1964), .Z(n1962) );
  XOR U3503 ( .A(DB[1376]), .B(DB[1369]), .Z(n1964) );
  AND U3504 ( .A(n242), .B(n1965), .Z(n1963) );
  XOR U3505 ( .A(n1966), .B(n1967), .Z(n1965) );
  XOR U3506 ( .A(DB[1369]), .B(DB[1362]), .Z(n1967) );
  AND U3507 ( .A(n246), .B(n1968), .Z(n1966) );
  XOR U3508 ( .A(n1969), .B(n1970), .Z(n1968) );
  XOR U3509 ( .A(DB[1362]), .B(DB[1355]), .Z(n1970) );
  AND U3510 ( .A(n250), .B(n1971), .Z(n1969) );
  XOR U3511 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR U3512 ( .A(DB[1355]), .B(DB[1348]), .Z(n1973) );
  AND U3513 ( .A(n254), .B(n1974), .Z(n1972) );
  XOR U3514 ( .A(n1975), .B(n1976), .Z(n1974) );
  XOR U3515 ( .A(DB[1348]), .B(DB[1341]), .Z(n1976) );
  AND U3516 ( .A(n258), .B(n1977), .Z(n1975) );
  XOR U3517 ( .A(n1978), .B(n1979), .Z(n1977) );
  XOR U3518 ( .A(DB[1341]), .B(DB[1334]), .Z(n1979) );
  AND U3519 ( .A(n262), .B(n1980), .Z(n1978) );
  XOR U3520 ( .A(n1981), .B(n1982), .Z(n1980) );
  XOR U3521 ( .A(DB[1334]), .B(DB[1327]), .Z(n1982) );
  AND U3522 ( .A(n266), .B(n1983), .Z(n1981) );
  XOR U3523 ( .A(n1984), .B(n1985), .Z(n1983) );
  XOR U3524 ( .A(DB[1327]), .B(DB[1320]), .Z(n1985) );
  AND U3525 ( .A(n270), .B(n1986), .Z(n1984) );
  XOR U3526 ( .A(n1987), .B(n1988), .Z(n1986) );
  XOR U3527 ( .A(DB[1320]), .B(DB[1313]), .Z(n1988) );
  AND U3528 ( .A(n274), .B(n1989), .Z(n1987) );
  XOR U3529 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U3530 ( .A(DB[1313]), .B(DB[1306]), .Z(n1991) );
  AND U3531 ( .A(n278), .B(n1992), .Z(n1990) );
  XOR U3532 ( .A(n1993), .B(n1994), .Z(n1992) );
  XOR U3533 ( .A(DB[1306]), .B(DB[1299]), .Z(n1994) );
  AND U3534 ( .A(n282), .B(n1995), .Z(n1993) );
  XOR U3535 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U3536 ( .A(DB[1299]), .B(DB[1292]), .Z(n1997) );
  AND U3537 ( .A(n286), .B(n1998), .Z(n1996) );
  XOR U3538 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR U3539 ( .A(DB[1292]), .B(DB[1285]), .Z(n2000) );
  AND U3540 ( .A(n290), .B(n2001), .Z(n1999) );
  XOR U3541 ( .A(n2002), .B(n2003), .Z(n2001) );
  XOR U3542 ( .A(DB[1285]), .B(DB[1278]), .Z(n2003) );
  AND U3543 ( .A(n294), .B(n2004), .Z(n2002) );
  XOR U3544 ( .A(n2005), .B(n2006), .Z(n2004) );
  XOR U3545 ( .A(DB[1278]), .B(DB[1271]), .Z(n2006) );
  AND U3546 ( .A(n298), .B(n2007), .Z(n2005) );
  XOR U3547 ( .A(n2008), .B(n2009), .Z(n2007) );
  XOR U3548 ( .A(DB[1271]), .B(DB[1264]), .Z(n2009) );
  AND U3549 ( .A(n302), .B(n2010), .Z(n2008) );
  XOR U3550 ( .A(n2011), .B(n2012), .Z(n2010) );
  XOR U3551 ( .A(DB[1264]), .B(DB[1257]), .Z(n2012) );
  AND U3552 ( .A(n306), .B(n2013), .Z(n2011) );
  XOR U3553 ( .A(n2014), .B(n2015), .Z(n2013) );
  XOR U3554 ( .A(DB[1257]), .B(DB[1250]), .Z(n2015) );
  AND U3555 ( .A(n310), .B(n2016), .Z(n2014) );
  XOR U3556 ( .A(n2017), .B(n2018), .Z(n2016) );
  XOR U3557 ( .A(DB[1250]), .B(DB[1243]), .Z(n2018) );
  AND U3558 ( .A(n314), .B(n2019), .Z(n2017) );
  XOR U3559 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U3560 ( .A(DB[1243]), .B(DB[1236]), .Z(n2021) );
  AND U3561 ( .A(n318), .B(n2022), .Z(n2020) );
  XOR U3562 ( .A(n2023), .B(n2024), .Z(n2022) );
  XOR U3563 ( .A(DB[1236]), .B(DB[1229]), .Z(n2024) );
  AND U3564 ( .A(n322), .B(n2025), .Z(n2023) );
  XOR U3565 ( .A(n2026), .B(n2027), .Z(n2025) );
  XOR U3566 ( .A(DB[1229]), .B(DB[1222]), .Z(n2027) );
  AND U3567 ( .A(n326), .B(n2028), .Z(n2026) );
  XOR U3568 ( .A(n2029), .B(n2030), .Z(n2028) );
  XOR U3569 ( .A(DB[1222]), .B(DB[1215]), .Z(n2030) );
  AND U3570 ( .A(n330), .B(n2031), .Z(n2029) );
  XOR U3571 ( .A(n2032), .B(n2033), .Z(n2031) );
  XOR U3572 ( .A(DB[1215]), .B(DB[1208]), .Z(n2033) );
  AND U3573 ( .A(n334), .B(n2034), .Z(n2032) );
  XOR U3574 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U3575 ( .A(DB[1208]), .B(DB[1201]), .Z(n2036) );
  AND U3576 ( .A(n338), .B(n2037), .Z(n2035) );
  XOR U3577 ( .A(n2038), .B(n2039), .Z(n2037) );
  XOR U3578 ( .A(DB[1201]), .B(DB[1194]), .Z(n2039) );
  AND U3579 ( .A(n342), .B(n2040), .Z(n2038) );
  XOR U3580 ( .A(n2041), .B(n2042), .Z(n2040) );
  XOR U3581 ( .A(DB[1194]), .B(DB[1187]), .Z(n2042) );
  AND U3582 ( .A(n346), .B(n2043), .Z(n2041) );
  XOR U3583 ( .A(n2044), .B(n2045), .Z(n2043) );
  XOR U3584 ( .A(DB[1187]), .B(DB[1180]), .Z(n2045) );
  AND U3585 ( .A(n350), .B(n2046), .Z(n2044) );
  XOR U3586 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U3587 ( .A(DB[1180]), .B(DB[1173]), .Z(n2048) );
  AND U3588 ( .A(n354), .B(n2049), .Z(n2047) );
  XOR U3589 ( .A(n2050), .B(n2051), .Z(n2049) );
  XOR U3590 ( .A(DB[1173]), .B(DB[1166]), .Z(n2051) );
  AND U3591 ( .A(n358), .B(n2052), .Z(n2050) );
  XOR U3592 ( .A(n2053), .B(n2054), .Z(n2052) );
  XOR U3593 ( .A(DB[1166]), .B(DB[1159]), .Z(n2054) );
  AND U3594 ( .A(n362), .B(n2055), .Z(n2053) );
  XOR U3595 ( .A(n2056), .B(n2057), .Z(n2055) );
  XOR U3596 ( .A(DB[1159]), .B(DB[1152]), .Z(n2057) );
  AND U3597 ( .A(n366), .B(n2058), .Z(n2056) );
  XOR U3598 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U3599 ( .A(DB[1152]), .B(DB[1145]), .Z(n2060) );
  AND U3600 ( .A(n370), .B(n2061), .Z(n2059) );
  XOR U3601 ( .A(n2062), .B(n2063), .Z(n2061) );
  XOR U3602 ( .A(DB[1145]), .B(DB[1138]), .Z(n2063) );
  AND U3603 ( .A(n374), .B(n2064), .Z(n2062) );
  XOR U3604 ( .A(n2065), .B(n2066), .Z(n2064) );
  XOR U3605 ( .A(DB[1138]), .B(DB[1131]), .Z(n2066) );
  AND U3606 ( .A(n378), .B(n2067), .Z(n2065) );
  XOR U3607 ( .A(n2068), .B(n2069), .Z(n2067) );
  XOR U3608 ( .A(DB[1131]), .B(DB[1124]), .Z(n2069) );
  AND U3609 ( .A(n382), .B(n2070), .Z(n2068) );
  XOR U3610 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U3611 ( .A(DB[1124]), .B(DB[1117]), .Z(n2072) );
  AND U3612 ( .A(n386), .B(n2073), .Z(n2071) );
  XOR U3613 ( .A(n2074), .B(n2075), .Z(n2073) );
  XOR U3614 ( .A(DB[1117]), .B(DB[1110]), .Z(n2075) );
  AND U3615 ( .A(n390), .B(n2076), .Z(n2074) );
  XOR U3616 ( .A(n2077), .B(n2078), .Z(n2076) );
  XOR U3617 ( .A(DB[1110]), .B(DB[1103]), .Z(n2078) );
  AND U3618 ( .A(n394), .B(n2079), .Z(n2077) );
  XOR U3619 ( .A(n2080), .B(n2081), .Z(n2079) );
  XOR U3620 ( .A(DB[1103]), .B(DB[1096]), .Z(n2081) );
  AND U3621 ( .A(n398), .B(n2082), .Z(n2080) );
  XOR U3622 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U3623 ( .A(DB[1096]), .B(DB[1089]), .Z(n2084) );
  AND U3624 ( .A(n402), .B(n2085), .Z(n2083) );
  XOR U3625 ( .A(n2086), .B(n2087), .Z(n2085) );
  XOR U3626 ( .A(DB[1089]), .B(DB[1082]), .Z(n2087) );
  AND U3627 ( .A(n406), .B(n2088), .Z(n2086) );
  XOR U3628 ( .A(n2089), .B(n2090), .Z(n2088) );
  XOR U3629 ( .A(DB[1082]), .B(DB[1075]), .Z(n2090) );
  AND U3630 ( .A(n410), .B(n2091), .Z(n2089) );
  XOR U3631 ( .A(n2092), .B(n2093), .Z(n2091) );
  XOR U3632 ( .A(DB[1075]), .B(DB[1068]), .Z(n2093) );
  AND U3633 ( .A(n414), .B(n2094), .Z(n2092) );
  XOR U3634 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U3635 ( .A(DB[1068]), .B(DB[1061]), .Z(n2096) );
  AND U3636 ( .A(n418), .B(n2097), .Z(n2095) );
  XOR U3637 ( .A(n2098), .B(n2099), .Z(n2097) );
  XOR U3638 ( .A(DB[1061]), .B(DB[1054]), .Z(n2099) );
  AND U3639 ( .A(n422), .B(n2100), .Z(n2098) );
  XOR U3640 ( .A(n2101), .B(n2102), .Z(n2100) );
  XOR U3641 ( .A(DB[1054]), .B(DB[1047]), .Z(n2102) );
  AND U3642 ( .A(n426), .B(n2103), .Z(n2101) );
  XOR U3643 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR U3644 ( .A(DB[1047]), .B(DB[1040]), .Z(n2105) );
  AND U3645 ( .A(n430), .B(n2106), .Z(n2104) );
  XOR U3646 ( .A(n2107), .B(n2108), .Z(n2106) );
  XOR U3647 ( .A(DB[1040]), .B(DB[1033]), .Z(n2108) );
  AND U3648 ( .A(n434), .B(n2109), .Z(n2107) );
  XOR U3649 ( .A(n2110), .B(n2111), .Z(n2109) );
  XOR U3650 ( .A(DB[1033]), .B(DB[1026]), .Z(n2111) );
  AND U3651 ( .A(n438), .B(n2112), .Z(n2110) );
  XOR U3652 ( .A(n2113), .B(n2114), .Z(n2112) );
  XOR U3653 ( .A(DB[1026]), .B(DB[1019]), .Z(n2114) );
  AND U3654 ( .A(n442), .B(n2115), .Z(n2113) );
  XOR U3655 ( .A(n2116), .B(n2117), .Z(n2115) );
  XOR U3656 ( .A(DB[1019]), .B(DB[1012]), .Z(n2117) );
  AND U3657 ( .A(n446), .B(n2118), .Z(n2116) );
  XOR U3658 ( .A(n2119), .B(n2120), .Z(n2118) );
  XOR U3659 ( .A(DB[1012]), .B(DB[1005]), .Z(n2120) );
  AND U3660 ( .A(n450), .B(n2121), .Z(n2119) );
  XOR U3661 ( .A(n2122), .B(n2123), .Z(n2121) );
  XOR U3662 ( .A(DB[998]), .B(DB[1005]), .Z(n2123) );
  AND U3663 ( .A(n454), .B(n2124), .Z(n2122) );
  XOR U3664 ( .A(n2125), .B(n2126), .Z(n2124) );
  XOR U3665 ( .A(DB[998]), .B(DB[991]), .Z(n2126) );
  AND U3666 ( .A(n458), .B(n2127), .Z(n2125) );
  XOR U3667 ( .A(n2128), .B(n2129), .Z(n2127) );
  XOR U3668 ( .A(DB[991]), .B(DB[984]), .Z(n2129) );
  AND U3669 ( .A(n462), .B(n2130), .Z(n2128) );
  XOR U3670 ( .A(n2131), .B(n2132), .Z(n2130) );
  XOR U3671 ( .A(DB[984]), .B(DB[977]), .Z(n2132) );
  AND U3672 ( .A(n466), .B(n2133), .Z(n2131) );
  XOR U3673 ( .A(n2134), .B(n2135), .Z(n2133) );
  XOR U3674 ( .A(DB[977]), .B(DB[970]), .Z(n2135) );
  AND U3675 ( .A(n470), .B(n2136), .Z(n2134) );
  XOR U3676 ( .A(n2137), .B(n2138), .Z(n2136) );
  XOR U3677 ( .A(DB[970]), .B(DB[963]), .Z(n2138) );
  AND U3678 ( .A(n474), .B(n2139), .Z(n2137) );
  XOR U3679 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U3680 ( .A(DB[963]), .B(DB[956]), .Z(n2141) );
  AND U3681 ( .A(n478), .B(n2142), .Z(n2140) );
  XOR U3682 ( .A(n2143), .B(n2144), .Z(n2142) );
  XOR U3683 ( .A(DB[956]), .B(DB[949]), .Z(n2144) );
  AND U3684 ( .A(n482), .B(n2145), .Z(n2143) );
  XOR U3685 ( .A(n2146), .B(n2147), .Z(n2145) );
  XOR U3686 ( .A(DB[949]), .B(DB[942]), .Z(n2147) );
  AND U3687 ( .A(n486), .B(n2148), .Z(n2146) );
  XOR U3688 ( .A(n2149), .B(n2150), .Z(n2148) );
  XOR U3689 ( .A(DB[942]), .B(DB[935]), .Z(n2150) );
  AND U3690 ( .A(n490), .B(n2151), .Z(n2149) );
  XOR U3691 ( .A(n2152), .B(n2153), .Z(n2151) );
  XOR U3692 ( .A(DB[935]), .B(DB[928]), .Z(n2153) );
  AND U3693 ( .A(n494), .B(n2154), .Z(n2152) );
  XOR U3694 ( .A(n2155), .B(n2156), .Z(n2154) );
  XOR U3695 ( .A(DB[928]), .B(DB[921]), .Z(n2156) );
  AND U3696 ( .A(n498), .B(n2157), .Z(n2155) );
  XOR U3697 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U3698 ( .A(DB[921]), .B(DB[914]), .Z(n2159) );
  AND U3699 ( .A(n502), .B(n2160), .Z(n2158) );
  XOR U3700 ( .A(n2161), .B(n2162), .Z(n2160) );
  XOR U3701 ( .A(DB[914]), .B(DB[907]), .Z(n2162) );
  AND U3702 ( .A(n506), .B(n2163), .Z(n2161) );
  XOR U3703 ( .A(n2164), .B(n2165), .Z(n2163) );
  XOR U3704 ( .A(DB[907]), .B(DB[900]), .Z(n2165) );
  AND U3705 ( .A(n510), .B(n2166), .Z(n2164) );
  XOR U3706 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U3707 ( .A(DB[900]), .B(DB[893]), .Z(n2168) );
  AND U3708 ( .A(n514), .B(n2169), .Z(n2167) );
  XOR U3709 ( .A(n2170), .B(n2171), .Z(n2169) );
  XOR U3710 ( .A(DB[893]), .B(DB[886]), .Z(n2171) );
  AND U3711 ( .A(n518), .B(n2172), .Z(n2170) );
  XOR U3712 ( .A(n2173), .B(n2174), .Z(n2172) );
  XOR U3713 ( .A(DB[886]), .B(DB[879]), .Z(n2174) );
  AND U3714 ( .A(n522), .B(n2175), .Z(n2173) );
  XOR U3715 ( .A(n2176), .B(n2177), .Z(n2175) );
  XOR U3716 ( .A(DB[879]), .B(DB[872]), .Z(n2177) );
  AND U3717 ( .A(n526), .B(n2178), .Z(n2176) );
  XOR U3718 ( .A(n2179), .B(n2180), .Z(n2178) );
  XOR U3719 ( .A(DB[872]), .B(DB[865]), .Z(n2180) );
  AND U3720 ( .A(n530), .B(n2181), .Z(n2179) );
  XOR U3721 ( .A(n2182), .B(n2183), .Z(n2181) );
  XOR U3722 ( .A(DB[865]), .B(DB[858]), .Z(n2183) );
  AND U3723 ( .A(n534), .B(n2184), .Z(n2182) );
  XOR U3724 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U3725 ( .A(DB[858]), .B(DB[851]), .Z(n2186) );
  AND U3726 ( .A(n538), .B(n2187), .Z(n2185) );
  XOR U3727 ( .A(n2188), .B(n2189), .Z(n2187) );
  XOR U3728 ( .A(DB[851]), .B(DB[844]), .Z(n2189) );
  AND U3729 ( .A(n542), .B(n2190), .Z(n2188) );
  XOR U3730 ( .A(n2191), .B(n2192), .Z(n2190) );
  XOR U3731 ( .A(DB[844]), .B(DB[837]), .Z(n2192) );
  AND U3732 ( .A(n546), .B(n2193), .Z(n2191) );
  XOR U3733 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U3734 ( .A(DB[837]), .B(DB[830]), .Z(n2195) );
  AND U3735 ( .A(n550), .B(n2196), .Z(n2194) );
  XOR U3736 ( .A(n2197), .B(n2198), .Z(n2196) );
  XOR U3737 ( .A(DB[830]), .B(DB[823]), .Z(n2198) );
  AND U3738 ( .A(n554), .B(n2199), .Z(n2197) );
  XOR U3739 ( .A(n2200), .B(n2201), .Z(n2199) );
  XOR U3740 ( .A(DB[823]), .B(DB[816]), .Z(n2201) );
  AND U3741 ( .A(n558), .B(n2202), .Z(n2200) );
  XOR U3742 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR U3743 ( .A(DB[816]), .B(DB[809]), .Z(n2204) );
  AND U3744 ( .A(n562), .B(n2205), .Z(n2203) );
  XOR U3745 ( .A(n2206), .B(n2207), .Z(n2205) );
  XOR U3746 ( .A(DB[809]), .B(DB[802]), .Z(n2207) );
  AND U3747 ( .A(n566), .B(n2208), .Z(n2206) );
  XOR U3748 ( .A(n2209), .B(n2210), .Z(n2208) );
  XOR U3749 ( .A(DB[802]), .B(DB[795]), .Z(n2210) );
  AND U3750 ( .A(n570), .B(n2211), .Z(n2209) );
  XOR U3751 ( .A(n2212), .B(n2213), .Z(n2211) );
  XOR U3752 ( .A(DB[795]), .B(DB[788]), .Z(n2213) );
  AND U3753 ( .A(n574), .B(n2214), .Z(n2212) );
  XOR U3754 ( .A(n2215), .B(n2216), .Z(n2214) );
  XOR U3755 ( .A(DB[788]), .B(DB[781]), .Z(n2216) );
  AND U3756 ( .A(n578), .B(n2217), .Z(n2215) );
  XOR U3757 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U3758 ( .A(DB[781]), .B(DB[774]), .Z(n2219) );
  AND U3759 ( .A(n582), .B(n2220), .Z(n2218) );
  XOR U3760 ( .A(n2221), .B(n2222), .Z(n2220) );
  XOR U3761 ( .A(DB[774]), .B(DB[767]), .Z(n2222) );
  AND U3762 ( .A(n586), .B(n2223), .Z(n2221) );
  XOR U3763 ( .A(n2224), .B(n2225), .Z(n2223) );
  XOR U3764 ( .A(DB[767]), .B(DB[760]), .Z(n2225) );
  AND U3765 ( .A(n590), .B(n2226), .Z(n2224) );
  XOR U3766 ( .A(n2227), .B(n2228), .Z(n2226) );
  XOR U3767 ( .A(DB[760]), .B(DB[753]), .Z(n2228) );
  AND U3768 ( .A(n594), .B(n2229), .Z(n2227) );
  XOR U3769 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U3770 ( .A(DB[753]), .B(DB[746]), .Z(n2231) );
  AND U3771 ( .A(n598), .B(n2232), .Z(n2230) );
  XOR U3772 ( .A(n2233), .B(n2234), .Z(n2232) );
  XOR U3773 ( .A(DB[746]), .B(DB[739]), .Z(n2234) );
  AND U3774 ( .A(n602), .B(n2235), .Z(n2233) );
  XOR U3775 ( .A(n2236), .B(n2237), .Z(n2235) );
  XOR U3776 ( .A(DB[739]), .B(DB[732]), .Z(n2237) );
  AND U3777 ( .A(n606), .B(n2238), .Z(n2236) );
  XOR U3778 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U3779 ( .A(DB[732]), .B(DB[725]), .Z(n2240) );
  AND U3780 ( .A(n610), .B(n2241), .Z(n2239) );
  XOR U3781 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U3782 ( .A(DB[725]), .B(DB[718]), .Z(n2243) );
  AND U3783 ( .A(n614), .B(n2244), .Z(n2242) );
  XOR U3784 ( .A(n2245), .B(n2246), .Z(n2244) );
  XOR U3785 ( .A(DB[718]), .B(DB[711]), .Z(n2246) );
  AND U3786 ( .A(n618), .B(n2247), .Z(n2245) );
  XOR U3787 ( .A(n2248), .B(n2249), .Z(n2247) );
  XOR U3788 ( .A(DB[711]), .B(DB[704]), .Z(n2249) );
  AND U3789 ( .A(n622), .B(n2250), .Z(n2248) );
  XOR U3790 ( .A(n2251), .B(n2252), .Z(n2250) );
  XOR U3791 ( .A(DB[704]), .B(DB[697]), .Z(n2252) );
  AND U3792 ( .A(n626), .B(n2253), .Z(n2251) );
  XOR U3793 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR U3794 ( .A(DB[697]), .B(DB[690]), .Z(n2255) );
  AND U3795 ( .A(n630), .B(n2256), .Z(n2254) );
  XOR U3796 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U3797 ( .A(DB[690]), .B(DB[683]), .Z(n2258) );
  AND U3798 ( .A(n634), .B(n2259), .Z(n2257) );
  XOR U3799 ( .A(n2260), .B(n2261), .Z(n2259) );
  XOR U3800 ( .A(DB[683]), .B(DB[676]), .Z(n2261) );
  AND U3801 ( .A(n638), .B(n2262), .Z(n2260) );
  XOR U3802 ( .A(n2263), .B(n2264), .Z(n2262) );
  XOR U3803 ( .A(DB[676]), .B(DB[669]), .Z(n2264) );
  AND U3804 ( .A(n642), .B(n2265), .Z(n2263) );
  XOR U3805 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U3806 ( .A(DB[669]), .B(DB[662]), .Z(n2267) );
  AND U3807 ( .A(n646), .B(n2268), .Z(n2266) );
  XOR U3808 ( .A(n2269), .B(n2270), .Z(n2268) );
  XOR U3809 ( .A(DB[662]), .B(DB[655]), .Z(n2270) );
  AND U3810 ( .A(n650), .B(n2271), .Z(n2269) );
  XOR U3811 ( .A(n2272), .B(n2273), .Z(n2271) );
  XOR U3812 ( .A(DB[655]), .B(DB[648]), .Z(n2273) );
  AND U3813 ( .A(n654), .B(n2274), .Z(n2272) );
  XOR U3814 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U3815 ( .A(DB[648]), .B(DB[641]), .Z(n2276) );
  AND U3816 ( .A(n658), .B(n2277), .Z(n2275) );
  XOR U3817 ( .A(n2278), .B(n2279), .Z(n2277) );
  XOR U3818 ( .A(DB[641]), .B(DB[634]), .Z(n2279) );
  AND U3819 ( .A(n662), .B(n2280), .Z(n2278) );
  XOR U3820 ( .A(n2281), .B(n2282), .Z(n2280) );
  XOR U3821 ( .A(DB[634]), .B(DB[627]), .Z(n2282) );
  AND U3822 ( .A(n666), .B(n2283), .Z(n2281) );
  XOR U3823 ( .A(n2284), .B(n2285), .Z(n2283) );
  XOR U3824 ( .A(DB[627]), .B(DB[620]), .Z(n2285) );
  AND U3825 ( .A(n670), .B(n2286), .Z(n2284) );
  XOR U3826 ( .A(n2287), .B(n2288), .Z(n2286) );
  XOR U3827 ( .A(DB[620]), .B(DB[613]), .Z(n2288) );
  AND U3828 ( .A(n674), .B(n2289), .Z(n2287) );
  XOR U3829 ( .A(n2290), .B(n2291), .Z(n2289) );
  XOR U3830 ( .A(DB[613]), .B(DB[606]), .Z(n2291) );
  AND U3831 ( .A(n678), .B(n2292), .Z(n2290) );
  XOR U3832 ( .A(n2293), .B(n2294), .Z(n2292) );
  XOR U3833 ( .A(DB[606]), .B(DB[599]), .Z(n2294) );
  AND U3834 ( .A(n682), .B(n2295), .Z(n2293) );
  XOR U3835 ( .A(n2296), .B(n2297), .Z(n2295) );
  XOR U3836 ( .A(DB[599]), .B(DB[592]), .Z(n2297) );
  AND U3837 ( .A(n686), .B(n2298), .Z(n2296) );
  XOR U3838 ( .A(n2299), .B(n2300), .Z(n2298) );
  XOR U3839 ( .A(DB[592]), .B(DB[585]), .Z(n2300) );
  AND U3840 ( .A(n690), .B(n2301), .Z(n2299) );
  XOR U3841 ( .A(n2302), .B(n2303), .Z(n2301) );
  XOR U3842 ( .A(DB[585]), .B(DB[578]), .Z(n2303) );
  AND U3843 ( .A(n694), .B(n2304), .Z(n2302) );
  XOR U3844 ( .A(n2305), .B(n2306), .Z(n2304) );
  XOR U3845 ( .A(DB[578]), .B(DB[571]), .Z(n2306) );
  AND U3846 ( .A(n698), .B(n2307), .Z(n2305) );
  XOR U3847 ( .A(n2308), .B(n2309), .Z(n2307) );
  XOR U3848 ( .A(DB[571]), .B(DB[564]), .Z(n2309) );
  AND U3849 ( .A(n702), .B(n2310), .Z(n2308) );
  XOR U3850 ( .A(n2311), .B(n2312), .Z(n2310) );
  XOR U3851 ( .A(DB[564]), .B(DB[557]), .Z(n2312) );
  AND U3852 ( .A(n706), .B(n2313), .Z(n2311) );
  XOR U3853 ( .A(n2314), .B(n2315), .Z(n2313) );
  XOR U3854 ( .A(DB[557]), .B(DB[550]), .Z(n2315) );
  AND U3855 ( .A(n710), .B(n2316), .Z(n2314) );
  XOR U3856 ( .A(n2317), .B(n2318), .Z(n2316) );
  XOR U3857 ( .A(DB[550]), .B(DB[543]), .Z(n2318) );
  AND U3858 ( .A(n714), .B(n2319), .Z(n2317) );
  XOR U3859 ( .A(n2320), .B(n2321), .Z(n2319) );
  XOR U3860 ( .A(DB[543]), .B(DB[536]), .Z(n2321) );
  AND U3861 ( .A(n718), .B(n2322), .Z(n2320) );
  XOR U3862 ( .A(n2323), .B(n2324), .Z(n2322) );
  XOR U3863 ( .A(DB[536]), .B(DB[529]), .Z(n2324) );
  AND U3864 ( .A(n722), .B(n2325), .Z(n2323) );
  XOR U3865 ( .A(n2326), .B(n2327), .Z(n2325) );
  XOR U3866 ( .A(DB[529]), .B(DB[522]), .Z(n2327) );
  AND U3867 ( .A(n726), .B(n2328), .Z(n2326) );
  XOR U3868 ( .A(n2329), .B(n2330), .Z(n2328) );
  XOR U3869 ( .A(DB[522]), .B(DB[515]), .Z(n2330) );
  AND U3870 ( .A(n730), .B(n2331), .Z(n2329) );
  XOR U3871 ( .A(n2332), .B(n2333), .Z(n2331) );
  XOR U3872 ( .A(DB[515]), .B(DB[508]), .Z(n2333) );
  AND U3873 ( .A(n734), .B(n2334), .Z(n2332) );
  XOR U3874 ( .A(n2335), .B(n2336), .Z(n2334) );
  XOR U3875 ( .A(DB[508]), .B(DB[501]), .Z(n2336) );
  AND U3876 ( .A(n738), .B(n2337), .Z(n2335) );
  XOR U3877 ( .A(n2338), .B(n2339), .Z(n2337) );
  XOR U3878 ( .A(DB[501]), .B(DB[494]), .Z(n2339) );
  AND U3879 ( .A(n742), .B(n2340), .Z(n2338) );
  XOR U3880 ( .A(n2341), .B(n2342), .Z(n2340) );
  XOR U3881 ( .A(DB[494]), .B(DB[487]), .Z(n2342) );
  AND U3882 ( .A(n746), .B(n2343), .Z(n2341) );
  XOR U3883 ( .A(n2344), .B(n2345), .Z(n2343) );
  XOR U3884 ( .A(DB[487]), .B(DB[480]), .Z(n2345) );
  AND U3885 ( .A(n750), .B(n2346), .Z(n2344) );
  XOR U3886 ( .A(n2347), .B(n2348), .Z(n2346) );
  XOR U3887 ( .A(DB[480]), .B(DB[473]), .Z(n2348) );
  AND U3888 ( .A(n754), .B(n2349), .Z(n2347) );
  XOR U3889 ( .A(n2350), .B(n2351), .Z(n2349) );
  XOR U3890 ( .A(DB[473]), .B(DB[466]), .Z(n2351) );
  AND U3891 ( .A(n758), .B(n2352), .Z(n2350) );
  XOR U3892 ( .A(n2353), .B(n2354), .Z(n2352) );
  XOR U3893 ( .A(DB[466]), .B(DB[459]), .Z(n2354) );
  AND U3894 ( .A(n762), .B(n2355), .Z(n2353) );
  XOR U3895 ( .A(n2356), .B(n2357), .Z(n2355) );
  XOR U3896 ( .A(DB[459]), .B(DB[452]), .Z(n2357) );
  AND U3897 ( .A(n766), .B(n2358), .Z(n2356) );
  XOR U3898 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U3899 ( .A(DB[452]), .B(DB[445]), .Z(n2360) );
  AND U3900 ( .A(n770), .B(n2361), .Z(n2359) );
  XOR U3901 ( .A(n2362), .B(n2363), .Z(n2361) );
  XOR U3902 ( .A(DB[445]), .B(DB[438]), .Z(n2363) );
  AND U3903 ( .A(n774), .B(n2364), .Z(n2362) );
  XOR U3904 ( .A(n2365), .B(n2366), .Z(n2364) );
  XOR U3905 ( .A(DB[438]), .B(DB[431]), .Z(n2366) );
  AND U3906 ( .A(n778), .B(n2367), .Z(n2365) );
  XOR U3907 ( .A(n2368), .B(n2369), .Z(n2367) );
  XOR U3908 ( .A(DB[431]), .B(DB[424]), .Z(n2369) );
  AND U3909 ( .A(n782), .B(n2370), .Z(n2368) );
  XOR U3910 ( .A(n2371), .B(n2372), .Z(n2370) );
  XOR U3911 ( .A(DB[424]), .B(DB[417]), .Z(n2372) );
  AND U3912 ( .A(n786), .B(n2373), .Z(n2371) );
  XOR U3913 ( .A(n2374), .B(n2375), .Z(n2373) );
  XOR U3914 ( .A(DB[417]), .B(DB[410]), .Z(n2375) );
  AND U3915 ( .A(n790), .B(n2376), .Z(n2374) );
  XOR U3916 ( .A(n2377), .B(n2378), .Z(n2376) );
  XOR U3917 ( .A(DB[410]), .B(DB[403]), .Z(n2378) );
  AND U3918 ( .A(n794), .B(n2379), .Z(n2377) );
  XOR U3919 ( .A(n2380), .B(n2381), .Z(n2379) );
  XOR U3920 ( .A(DB[403]), .B(DB[396]), .Z(n2381) );
  AND U3921 ( .A(n798), .B(n2382), .Z(n2380) );
  XOR U3922 ( .A(n2383), .B(n2384), .Z(n2382) );
  XOR U3923 ( .A(DB[396]), .B(DB[389]), .Z(n2384) );
  AND U3924 ( .A(n802), .B(n2385), .Z(n2383) );
  XOR U3925 ( .A(n2386), .B(n2387), .Z(n2385) );
  XOR U3926 ( .A(DB[389]), .B(DB[382]), .Z(n2387) );
  AND U3927 ( .A(n806), .B(n2388), .Z(n2386) );
  XOR U3928 ( .A(n2389), .B(n2390), .Z(n2388) );
  XOR U3929 ( .A(DB[382]), .B(DB[375]), .Z(n2390) );
  AND U3930 ( .A(n810), .B(n2391), .Z(n2389) );
  XOR U3931 ( .A(n2392), .B(n2393), .Z(n2391) );
  XOR U3932 ( .A(DB[375]), .B(DB[368]), .Z(n2393) );
  AND U3933 ( .A(n814), .B(n2394), .Z(n2392) );
  XOR U3934 ( .A(n2395), .B(n2396), .Z(n2394) );
  XOR U3935 ( .A(DB[368]), .B(DB[361]), .Z(n2396) );
  AND U3936 ( .A(n818), .B(n2397), .Z(n2395) );
  XOR U3937 ( .A(n2398), .B(n2399), .Z(n2397) );
  XOR U3938 ( .A(DB[361]), .B(DB[354]), .Z(n2399) );
  AND U3939 ( .A(n822), .B(n2400), .Z(n2398) );
  XOR U3940 ( .A(n2401), .B(n2402), .Z(n2400) );
  XOR U3941 ( .A(DB[354]), .B(DB[347]), .Z(n2402) );
  AND U3942 ( .A(n826), .B(n2403), .Z(n2401) );
  XOR U3943 ( .A(n2404), .B(n2405), .Z(n2403) );
  XOR U3944 ( .A(DB[347]), .B(DB[340]), .Z(n2405) );
  AND U3945 ( .A(n830), .B(n2406), .Z(n2404) );
  XOR U3946 ( .A(n2407), .B(n2408), .Z(n2406) );
  XOR U3947 ( .A(DB[340]), .B(DB[333]), .Z(n2408) );
  AND U3948 ( .A(n834), .B(n2409), .Z(n2407) );
  XOR U3949 ( .A(n2410), .B(n2411), .Z(n2409) );
  XOR U3950 ( .A(DB[333]), .B(DB[326]), .Z(n2411) );
  AND U3951 ( .A(n838), .B(n2412), .Z(n2410) );
  XOR U3952 ( .A(n2413), .B(n2414), .Z(n2412) );
  XOR U3953 ( .A(DB[326]), .B(DB[319]), .Z(n2414) );
  AND U3954 ( .A(n842), .B(n2415), .Z(n2413) );
  XOR U3955 ( .A(n2416), .B(n2417), .Z(n2415) );
  XOR U3956 ( .A(DB[319]), .B(DB[312]), .Z(n2417) );
  AND U3957 ( .A(n846), .B(n2418), .Z(n2416) );
  XOR U3958 ( .A(n2419), .B(n2420), .Z(n2418) );
  XOR U3959 ( .A(DB[312]), .B(DB[305]), .Z(n2420) );
  AND U3960 ( .A(n850), .B(n2421), .Z(n2419) );
  XOR U3961 ( .A(n2422), .B(n2423), .Z(n2421) );
  XOR U3962 ( .A(DB[305]), .B(DB[298]), .Z(n2423) );
  AND U3963 ( .A(n854), .B(n2424), .Z(n2422) );
  XOR U3964 ( .A(n2425), .B(n2426), .Z(n2424) );
  XOR U3965 ( .A(DB[298]), .B(DB[291]), .Z(n2426) );
  AND U3966 ( .A(n858), .B(n2427), .Z(n2425) );
  XOR U3967 ( .A(n2428), .B(n2429), .Z(n2427) );
  XOR U3968 ( .A(DB[291]), .B(DB[284]), .Z(n2429) );
  AND U3969 ( .A(n862), .B(n2430), .Z(n2428) );
  XOR U3970 ( .A(n2431), .B(n2432), .Z(n2430) );
  XOR U3971 ( .A(DB[284]), .B(DB[277]), .Z(n2432) );
  AND U3972 ( .A(n866), .B(n2433), .Z(n2431) );
  XOR U3973 ( .A(n2434), .B(n2435), .Z(n2433) );
  XOR U3974 ( .A(DB[277]), .B(DB[270]), .Z(n2435) );
  AND U3975 ( .A(n870), .B(n2436), .Z(n2434) );
  XOR U3976 ( .A(n2437), .B(n2438), .Z(n2436) );
  XOR U3977 ( .A(DB[270]), .B(DB[263]), .Z(n2438) );
  AND U3978 ( .A(n874), .B(n2439), .Z(n2437) );
  XOR U3979 ( .A(n2440), .B(n2441), .Z(n2439) );
  XOR U3980 ( .A(DB[263]), .B(DB[256]), .Z(n2441) );
  AND U3981 ( .A(n878), .B(n2442), .Z(n2440) );
  XOR U3982 ( .A(n2443), .B(n2444), .Z(n2442) );
  XOR U3983 ( .A(DB[256]), .B(DB[249]), .Z(n2444) );
  AND U3984 ( .A(n882), .B(n2445), .Z(n2443) );
  XOR U3985 ( .A(n2446), .B(n2447), .Z(n2445) );
  XOR U3986 ( .A(DB[249]), .B(DB[242]), .Z(n2447) );
  AND U3987 ( .A(n886), .B(n2448), .Z(n2446) );
  XOR U3988 ( .A(n2449), .B(n2450), .Z(n2448) );
  XOR U3989 ( .A(DB[242]), .B(DB[235]), .Z(n2450) );
  AND U3990 ( .A(n890), .B(n2451), .Z(n2449) );
  XOR U3991 ( .A(n2452), .B(n2453), .Z(n2451) );
  XOR U3992 ( .A(DB[235]), .B(DB[228]), .Z(n2453) );
  AND U3993 ( .A(n894), .B(n2454), .Z(n2452) );
  XOR U3994 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U3995 ( .A(DB[228]), .B(DB[221]), .Z(n2456) );
  AND U3996 ( .A(n898), .B(n2457), .Z(n2455) );
  XOR U3997 ( .A(n2458), .B(n2459), .Z(n2457) );
  XOR U3998 ( .A(DB[221]), .B(DB[214]), .Z(n2459) );
  AND U3999 ( .A(n902), .B(n2460), .Z(n2458) );
  XOR U4000 ( .A(n2461), .B(n2462), .Z(n2460) );
  XOR U4001 ( .A(DB[214]), .B(DB[207]), .Z(n2462) );
  AND U4002 ( .A(n906), .B(n2463), .Z(n2461) );
  XOR U4003 ( .A(n2464), .B(n2465), .Z(n2463) );
  XOR U4004 ( .A(DB[207]), .B(DB[200]), .Z(n2465) );
  AND U4005 ( .A(n910), .B(n2466), .Z(n2464) );
  XOR U4006 ( .A(n2467), .B(n2468), .Z(n2466) );
  XOR U4007 ( .A(DB[200]), .B(DB[193]), .Z(n2468) );
  AND U4008 ( .A(n914), .B(n2469), .Z(n2467) );
  XOR U4009 ( .A(n2470), .B(n2471), .Z(n2469) );
  XOR U4010 ( .A(DB[193]), .B(DB[186]), .Z(n2471) );
  AND U4011 ( .A(n918), .B(n2472), .Z(n2470) );
  XOR U4012 ( .A(n2473), .B(n2474), .Z(n2472) );
  XOR U4013 ( .A(DB[186]), .B(DB[179]), .Z(n2474) );
  AND U4014 ( .A(n922), .B(n2475), .Z(n2473) );
  XOR U4015 ( .A(n2476), .B(n2477), .Z(n2475) );
  XOR U4016 ( .A(DB[179]), .B(DB[172]), .Z(n2477) );
  AND U4017 ( .A(n926), .B(n2478), .Z(n2476) );
  XOR U4018 ( .A(n2479), .B(n2480), .Z(n2478) );
  XOR U4019 ( .A(DB[172]), .B(DB[165]), .Z(n2480) );
  AND U4020 ( .A(n930), .B(n2481), .Z(n2479) );
  XOR U4021 ( .A(n2482), .B(n2483), .Z(n2481) );
  XOR U4022 ( .A(DB[165]), .B(DB[158]), .Z(n2483) );
  AND U4023 ( .A(n934), .B(n2484), .Z(n2482) );
  XOR U4024 ( .A(n2485), .B(n2486), .Z(n2484) );
  XOR U4025 ( .A(DB[158]), .B(DB[151]), .Z(n2486) );
  AND U4026 ( .A(n938), .B(n2487), .Z(n2485) );
  XOR U4027 ( .A(n2488), .B(n2489), .Z(n2487) );
  XOR U4028 ( .A(DB[151]), .B(DB[144]), .Z(n2489) );
  AND U4029 ( .A(n942), .B(n2490), .Z(n2488) );
  XOR U4030 ( .A(n2491), .B(n2492), .Z(n2490) );
  XOR U4031 ( .A(DB[144]), .B(DB[137]), .Z(n2492) );
  AND U4032 ( .A(n946), .B(n2493), .Z(n2491) );
  XOR U4033 ( .A(n2494), .B(n2495), .Z(n2493) );
  XOR U4034 ( .A(DB[137]), .B(DB[130]), .Z(n2495) );
  AND U4035 ( .A(n950), .B(n2496), .Z(n2494) );
  XOR U4036 ( .A(n2497), .B(n2498), .Z(n2496) );
  XOR U4037 ( .A(DB[130]), .B(DB[123]), .Z(n2498) );
  AND U4038 ( .A(n954), .B(n2499), .Z(n2497) );
  XOR U4039 ( .A(n2500), .B(n2501), .Z(n2499) );
  XOR U4040 ( .A(DB[123]), .B(DB[116]), .Z(n2501) );
  AND U4041 ( .A(n958), .B(n2502), .Z(n2500) );
  XOR U4042 ( .A(n2503), .B(n2504), .Z(n2502) );
  XOR U4043 ( .A(DB[116]), .B(DB[109]), .Z(n2504) );
  AND U4044 ( .A(n962), .B(n2505), .Z(n2503) );
  XOR U4045 ( .A(n2506), .B(n2507), .Z(n2505) );
  XOR U4046 ( .A(DB[109]), .B(DB[102]), .Z(n2507) );
  AND U4047 ( .A(n966), .B(n2508), .Z(n2506) );
  XOR U4048 ( .A(n2509), .B(n2510), .Z(n2508) );
  XOR U4049 ( .A(DB[95]), .B(DB[102]), .Z(n2510) );
  AND U4050 ( .A(n970), .B(n2511), .Z(n2509) );
  XOR U4051 ( .A(n2512), .B(n2513), .Z(n2511) );
  XOR U4052 ( .A(DB[95]), .B(DB[88]), .Z(n2513) );
  AND U4053 ( .A(n974), .B(n2514), .Z(n2512) );
  XOR U4054 ( .A(n2515), .B(n2516), .Z(n2514) );
  XOR U4055 ( .A(DB[88]), .B(DB[81]), .Z(n2516) );
  AND U4056 ( .A(n978), .B(n2517), .Z(n2515) );
  XOR U4057 ( .A(n2518), .B(n2519), .Z(n2517) );
  XOR U4058 ( .A(DB[81]), .B(DB[74]), .Z(n2519) );
  AND U4059 ( .A(n982), .B(n2520), .Z(n2518) );
  XOR U4060 ( .A(n2521), .B(n2522), .Z(n2520) );
  XOR U4061 ( .A(DB[74]), .B(DB[67]), .Z(n2522) );
  AND U4062 ( .A(n986), .B(n2523), .Z(n2521) );
  XOR U4063 ( .A(n2524), .B(n2525), .Z(n2523) );
  XOR U4064 ( .A(DB[67]), .B(DB[60]), .Z(n2525) );
  AND U4065 ( .A(n990), .B(n2526), .Z(n2524) );
  XOR U4066 ( .A(n2527), .B(n2528), .Z(n2526) );
  XOR U4067 ( .A(DB[60]), .B(DB[53]), .Z(n2528) );
  AND U4068 ( .A(n994), .B(n2529), .Z(n2527) );
  XOR U4069 ( .A(n2530), .B(n2531), .Z(n2529) );
  XOR U4070 ( .A(DB[53]), .B(DB[46]), .Z(n2531) );
  AND U4071 ( .A(n998), .B(n2532), .Z(n2530) );
  XOR U4072 ( .A(n2533), .B(n2534), .Z(n2532) );
  XOR U4073 ( .A(DB[46]), .B(DB[39]), .Z(n2534) );
  AND U4074 ( .A(n1002), .B(n2535), .Z(n2533) );
  XOR U4075 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR U4076 ( .A(DB[39]), .B(DB[32]), .Z(n2537) );
  AND U4077 ( .A(n1006), .B(n2538), .Z(n2536) );
  XOR U4078 ( .A(n2539), .B(n2540), .Z(n2538) );
  XOR U4079 ( .A(DB[32]), .B(DB[25]), .Z(n2540) );
  AND U4080 ( .A(n1010), .B(n2541), .Z(n2539) );
  XOR U4081 ( .A(n2542), .B(n2543), .Z(n2541) );
  XOR U4082 ( .A(DB[25]), .B(DB[18]), .Z(n2543) );
  AND U4083 ( .A(n1014), .B(n2544), .Z(n2542) );
  XOR U4084 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U4085 ( .A(DB[18]), .B(DB[11]), .Z(n2546) );
  AND U4086 ( .A(n1018), .B(n2547), .Z(n2545) );
  XOR U4087 ( .A(DB[4]), .B(DB[11]), .Z(n2547) );
  XOR U4088 ( .A(DB[1788]), .B(n2548), .Z(min_val_out[3]) );
  AND U4089 ( .A(n2), .B(n2549), .Z(n2548) );
  XOR U4090 ( .A(n2550), .B(n2551), .Z(n2549) );
  XOR U4091 ( .A(DB[1788]), .B(DB[1781]), .Z(n2551) );
  AND U4092 ( .A(n6), .B(n2552), .Z(n2550) );
  XOR U4093 ( .A(n2553), .B(n2554), .Z(n2552) );
  XOR U4094 ( .A(DB[1781]), .B(DB[1774]), .Z(n2554) );
  AND U4095 ( .A(n10), .B(n2555), .Z(n2553) );
  XOR U4096 ( .A(n2556), .B(n2557), .Z(n2555) );
  XOR U4097 ( .A(DB[1774]), .B(DB[1767]), .Z(n2557) );
  AND U4098 ( .A(n14), .B(n2558), .Z(n2556) );
  XOR U4099 ( .A(n2559), .B(n2560), .Z(n2558) );
  XOR U4100 ( .A(DB[1767]), .B(DB[1760]), .Z(n2560) );
  AND U4101 ( .A(n18), .B(n2561), .Z(n2559) );
  XOR U4102 ( .A(n2562), .B(n2563), .Z(n2561) );
  XOR U4103 ( .A(DB[1760]), .B(DB[1753]), .Z(n2563) );
  AND U4104 ( .A(n22), .B(n2564), .Z(n2562) );
  XOR U4105 ( .A(n2565), .B(n2566), .Z(n2564) );
  XOR U4106 ( .A(DB[1753]), .B(DB[1746]), .Z(n2566) );
  AND U4107 ( .A(n26), .B(n2567), .Z(n2565) );
  XOR U4108 ( .A(n2568), .B(n2569), .Z(n2567) );
  XOR U4109 ( .A(DB[1746]), .B(DB[1739]), .Z(n2569) );
  AND U4110 ( .A(n30), .B(n2570), .Z(n2568) );
  XOR U4111 ( .A(n2571), .B(n2572), .Z(n2570) );
  XOR U4112 ( .A(DB[1739]), .B(DB[1732]), .Z(n2572) );
  AND U4113 ( .A(n34), .B(n2573), .Z(n2571) );
  XOR U4114 ( .A(n2574), .B(n2575), .Z(n2573) );
  XOR U4115 ( .A(DB[1732]), .B(DB[1725]), .Z(n2575) );
  AND U4116 ( .A(n38), .B(n2576), .Z(n2574) );
  XOR U4117 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR U4118 ( .A(DB[1725]), .B(DB[1718]), .Z(n2578) );
  AND U4119 ( .A(n42), .B(n2579), .Z(n2577) );
  XOR U4120 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U4121 ( .A(DB[1718]), .B(DB[1711]), .Z(n2581) );
  AND U4122 ( .A(n46), .B(n2582), .Z(n2580) );
  XOR U4123 ( .A(n2583), .B(n2584), .Z(n2582) );
  XOR U4124 ( .A(DB[1711]), .B(DB[1704]), .Z(n2584) );
  AND U4125 ( .A(n50), .B(n2585), .Z(n2583) );
  XOR U4126 ( .A(n2586), .B(n2587), .Z(n2585) );
  XOR U4127 ( .A(DB[1704]), .B(DB[1697]), .Z(n2587) );
  AND U4128 ( .A(n54), .B(n2588), .Z(n2586) );
  XOR U4129 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR U4130 ( .A(DB[1697]), .B(DB[1690]), .Z(n2590) );
  AND U4131 ( .A(n58), .B(n2591), .Z(n2589) );
  XOR U4132 ( .A(n2592), .B(n2593), .Z(n2591) );
  XOR U4133 ( .A(DB[1690]), .B(DB[1683]), .Z(n2593) );
  AND U4134 ( .A(n62), .B(n2594), .Z(n2592) );
  XOR U4135 ( .A(n2595), .B(n2596), .Z(n2594) );
  XOR U4136 ( .A(DB[1683]), .B(DB[1676]), .Z(n2596) );
  AND U4137 ( .A(n66), .B(n2597), .Z(n2595) );
  XOR U4138 ( .A(n2598), .B(n2599), .Z(n2597) );
  XOR U4139 ( .A(DB[1676]), .B(DB[1669]), .Z(n2599) );
  AND U4140 ( .A(n70), .B(n2600), .Z(n2598) );
  XOR U4141 ( .A(n2601), .B(n2602), .Z(n2600) );
  XOR U4142 ( .A(DB[1669]), .B(DB[1662]), .Z(n2602) );
  AND U4143 ( .A(n74), .B(n2603), .Z(n2601) );
  XOR U4144 ( .A(n2604), .B(n2605), .Z(n2603) );
  XOR U4145 ( .A(DB[1662]), .B(DB[1655]), .Z(n2605) );
  AND U4146 ( .A(n78), .B(n2606), .Z(n2604) );
  XOR U4147 ( .A(n2607), .B(n2608), .Z(n2606) );
  XOR U4148 ( .A(DB[1655]), .B(DB[1648]), .Z(n2608) );
  AND U4149 ( .A(n82), .B(n2609), .Z(n2607) );
  XOR U4150 ( .A(n2610), .B(n2611), .Z(n2609) );
  XOR U4151 ( .A(DB[1648]), .B(DB[1641]), .Z(n2611) );
  AND U4152 ( .A(n86), .B(n2612), .Z(n2610) );
  XOR U4153 ( .A(n2613), .B(n2614), .Z(n2612) );
  XOR U4154 ( .A(DB[1641]), .B(DB[1634]), .Z(n2614) );
  AND U4155 ( .A(n90), .B(n2615), .Z(n2613) );
  XOR U4156 ( .A(n2616), .B(n2617), .Z(n2615) );
  XOR U4157 ( .A(DB[1634]), .B(DB[1627]), .Z(n2617) );
  AND U4158 ( .A(n94), .B(n2618), .Z(n2616) );
  XOR U4159 ( .A(n2619), .B(n2620), .Z(n2618) );
  XOR U4160 ( .A(DB[1627]), .B(DB[1620]), .Z(n2620) );
  AND U4161 ( .A(n98), .B(n2621), .Z(n2619) );
  XOR U4162 ( .A(n2622), .B(n2623), .Z(n2621) );
  XOR U4163 ( .A(DB[1620]), .B(DB[1613]), .Z(n2623) );
  AND U4164 ( .A(n102), .B(n2624), .Z(n2622) );
  XOR U4165 ( .A(n2625), .B(n2626), .Z(n2624) );
  XOR U4166 ( .A(DB[1613]), .B(DB[1606]), .Z(n2626) );
  AND U4167 ( .A(n106), .B(n2627), .Z(n2625) );
  XOR U4168 ( .A(n2628), .B(n2629), .Z(n2627) );
  XOR U4169 ( .A(DB[1606]), .B(DB[1599]), .Z(n2629) );
  AND U4170 ( .A(n110), .B(n2630), .Z(n2628) );
  XOR U4171 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U4172 ( .A(DB[1599]), .B(DB[1592]), .Z(n2632) );
  AND U4173 ( .A(n114), .B(n2633), .Z(n2631) );
  XOR U4174 ( .A(n2634), .B(n2635), .Z(n2633) );
  XOR U4175 ( .A(DB[1592]), .B(DB[1585]), .Z(n2635) );
  AND U4176 ( .A(n118), .B(n2636), .Z(n2634) );
  XOR U4177 ( .A(n2637), .B(n2638), .Z(n2636) );
  XOR U4178 ( .A(DB[1585]), .B(DB[1578]), .Z(n2638) );
  AND U4179 ( .A(n122), .B(n2639), .Z(n2637) );
  XOR U4180 ( .A(n2640), .B(n2641), .Z(n2639) );
  XOR U4181 ( .A(DB[1578]), .B(DB[1571]), .Z(n2641) );
  AND U4182 ( .A(n126), .B(n2642), .Z(n2640) );
  XOR U4183 ( .A(n2643), .B(n2644), .Z(n2642) );
  XOR U4184 ( .A(DB[1571]), .B(DB[1564]), .Z(n2644) );
  AND U4185 ( .A(n130), .B(n2645), .Z(n2643) );
  XOR U4186 ( .A(n2646), .B(n2647), .Z(n2645) );
  XOR U4187 ( .A(DB[1564]), .B(DB[1557]), .Z(n2647) );
  AND U4188 ( .A(n134), .B(n2648), .Z(n2646) );
  XOR U4189 ( .A(n2649), .B(n2650), .Z(n2648) );
  XOR U4190 ( .A(DB[1557]), .B(DB[1550]), .Z(n2650) );
  AND U4191 ( .A(n138), .B(n2651), .Z(n2649) );
  XOR U4192 ( .A(n2652), .B(n2653), .Z(n2651) );
  XOR U4193 ( .A(DB[1550]), .B(DB[1543]), .Z(n2653) );
  AND U4194 ( .A(n142), .B(n2654), .Z(n2652) );
  XOR U4195 ( .A(n2655), .B(n2656), .Z(n2654) );
  XOR U4196 ( .A(DB[1543]), .B(DB[1536]), .Z(n2656) );
  AND U4197 ( .A(n146), .B(n2657), .Z(n2655) );
  XOR U4198 ( .A(n2658), .B(n2659), .Z(n2657) );
  XOR U4199 ( .A(DB[1536]), .B(DB[1529]), .Z(n2659) );
  AND U4200 ( .A(n150), .B(n2660), .Z(n2658) );
  XOR U4201 ( .A(n2661), .B(n2662), .Z(n2660) );
  XOR U4202 ( .A(DB[1529]), .B(DB[1522]), .Z(n2662) );
  AND U4203 ( .A(n154), .B(n2663), .Z(n2661) );
  XOR U4204 ( .A(n2664), .B(n2665), .Z(n2663) );
  XOR U4205 ( .A(DB[1522]), .B(DB[1515]), .Z(n2665) );
  AND U4206 ( .A(n158), .B(n2666), .Z(n2664) );
  XOR U4207 ( .A(n2667), .B(n2668), .Z(n2666) );
  XOR U4208 ( .A(DB[1515]), .B(DB[1508]), .Z(n2668) );
  AND U4209 ( .A(n162), .B(n2669), .Z(n2667) );
  XOR U4210 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR U4211 ( .A(DB[1508]), .B(DB[1501]), .Z(n2671) );
  AND U4212 ( .A(n166), .B(n2672), .Z(n2670) );
  XOR U4213 ( .A(n2673), .B(n2674), .Z(n2672) );
  XOR U4214 ( .A(DB[1501]), .B(DB[1494]), .Z(n2674) );
  AND U4215 ( .A(n170), .B(n2675), .Z(n2673) );
  XOR U4216 ( .A(n2676), .B(n2677), .Z(n2675) );
  XOR U4217 ( .A(DB[1494]), .B(DB[1487]), .Z(n2677) );
  AND U4218 ( .A(n174), .B(n2678), .Z(n2676) );
  XOR U4219 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR U4220 ( .A(DB[1487]), .B(DB[1480]), .Z(n2680) );
  AND U4221 ( .A(n178), .B(n2681), .Z(n2679) );
  XOR U4222 ( .A(n2682), .B(n2683), .Z(n2681) );
  XOR U4223 ( .A(DB[1480]), .B(DB[1473]), .Z(n2683) );
  AND U4224 ( .A(n182), .B(n2684), .Z(n2682) );
  XOR U4225 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR U4226 ( .A(DB[1473]), .B(DB[1466]), .Z(n2686) );
  AND U4227 ( .A(n186), .B(n2687), .Z(n2685) );
  XOR U4228 ( .A(n2688), .B(n2689), .Z(n2687) );
  XOR U4229 ( .A(DB[1466]), .B(DB[1459]), .Z(n2689) );
  AND U4230 ( .A(n190), .B(n2690), .Z(n2688) );
  XOR U4231 ( .A(n2691), .B(n2692), .Z(n2690) );
  XOR U4232 ( .A(DB[1459]), .B(DB[1452]), .Z(n2692) );
  AND U4233 ( .A(n194), .B(n2693), .Z(n2691) );
  XOR U4234 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR U4235 ( .A(DB[1452]), .B(DB[1445]), .Z(n2695) );
  AND U4236 ( .A(n198), .B(n2696), .Z(n2694) );
  XOR U4237 ( .A(n2697), .B(n2698), .Z(n2696) );
  XOR U4238 ( .A(DB[1445]), .B(DB[1438]), .Z(n2698) );
  AND U4239 ( .A(n202), .B(n2699), .Z(n2697) );
  XOR U4240 ( .A(n2700), .B(n2701), .Z(n2699) );
  XOR U4241 ( .A(DB[1438]), .B(DB[1431]), .Z(n2701) );
  AND U4242 ( .A(n206), .B(n2702), .Z(n2700) );
  XOR U4243 ( .A(n2703), .B(n2704), .Z(n2702) );
  XOR U4244 ( .A(DB[1431]), .B(DB[1424]), .Z(n2704) );
  AND U4245 ( .A(n210), .B(n2705), .Z(n2703) );
  XOR U4246 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U4247 ( .A(DB[1424]), .B(DB[1417]), .Z(n2707) );
  AND U4248 ( .A(n214), .B(n2708), .Z(n2706) );
  XOR U4249 ( .A(n2709), .B(n2710), .Z(n2708) );
  XOR U4250 ( .A(DB[1417]), .B(DB[1410]), .Z(n2710) );
  AND U4251 ( .A(n218), .B(n2711), .Z(n2709) );
  XOR U4252 ( .A(n2712), .B(n2713), .Z(n2711) );
  XOR U4253 ( .A(DB[1410]), .B(DB[1403]), .Z(n2713) );
  AND U4254 ( .A(n222), .B(n2714), .Z(n2712) );
  XOR U4255 ( .A(n2715), .B(n2716), .Z(n2714) );
  XOR U4256 ( .A(DB[1403]), .B(DB[1396]), .Z(n2716) );
  AND U4257 ( .A(n226), .B(n2717), .Z(n2715) );
  XOR U4258 ( .A(n2718), .B(n2719), .Z(n2717) );
  XOR U4259 ( .A(DB[1396]), .B(DB[1389]), .Z(n2719) );
  AND U4260 ( .A(n230), .B(n2720), .Z(n2718) );
  XOR U4261 ( .A(n2721), .B(n2722), .Z(n2720) );
  XOR U4262 ( .A(DB[1389]), .B(DB[1382]), .Z(n2722) );
  AND U4263 ( .A(n234), .B(n2723), .Z(n2721) );
  XOR U4264 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR U4265 ( .A(DB[1382]), .B(DB[1375]), .Z(n2725) );
  AND U4266 ( .A(n238), .B(n2726), .Z(n2724) );
  XOR U4267 ( .A(n2727), .B(n2728), .Z(n2726) );
  XOR U4268 ( .A(DB[1375]), .B(DB[1368]), .Z(n2728) );
  AND U4269 ( .A(n242), .B(n2729), .Z(n2727) );
  XOR U4270 ( .A(n2730), .B(n2731), .Z(n2729) );
  XOR U4271 ( .A(DB[1368]), .B(DB[1361]), .Z(n2731) );
  AND U4272 ( .A(n246), .B(n2732), .Z(n2730) );
  XOR U4273 ( .A(n2733), .B(n2734), .Z(n2732) );
  XOR U4274 ( .A(DB[1361]), .B(DB[1354]), .Z(n2734) );
  AND U4275 ( .A(n250), .B(n2735), .Z(n2733) );
  XOR U4276 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR U4277 ( .A(DB[1354]), .B(DB[1347]), .Z(n2737) );
  AND U4278 ( .A(n254), .B(n2738), .Z(n2736) );
  XOR U4279 ( .A(n2739), .B(n2740), .Z(n2738) );
  XOR U4280 ( .A(DB[1347]), .B(DB[1340]), .Z(n2740) );
  AND U4281 ( .A(n258), .B(n2741), .Z(n2739) );
  XOR U4282 ( .A(n2742), .B(n2743), .Z(n2741) );
  XOR U4283 ( .A(DB[1340]), .B(DB[1333]), .Z(n2743) );
  AND U4284 ( .A(n262), .B(n2744), .Z(n2742) );
  XOR U4285 ( .A(n2745), .B(n2746), .Z(n2744) );
  XOR U4286 ( .A(DB[1333]), .B(DB[1326]), .Z(n2746) );
  AND U4287 ( .A(n266), .B(n2747), .Z(n2745) );
  XOR U4288 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR U4289 ( .A(DB[1326]), .B(DB[1319]), .Z(n2749) );
  AND U4290 ( .A(n270), .B(n2750), .Z(n2748) );
  XOR U4291 ( .A(n2751), .B(n2752), .Z(n2750) );
  XOR U4292 ( .A(DB[1319]), .B(DB[1312]), .Z(n2752) );
  AND U4293 ( .A(n274), .B(n2753), .Z(n2751) );
  XOR U4294 ( .A(n2754), .B(n2755), .Z(n2753) );
  XOR U4295 ( .A(DB[1312]), .B(DB[1305]), .Z(n2755) );
  AND U4296 ( .A(n278), .B(n2756), .Z(n2754) );
  XOR U4297 ( .A(n2757), .B(n2758), .Z(n2756) );
  XOR U4298 ( .A(DB[1305]), .B(DB[1298]), .Z(n2758) );
  AND U4299 ( .A(n282), .B(n2759), .Z(n2757) );
  XOR U4300 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U4301 ( .A(DB[1298]), .B(DB[1291]), .Z(n2761) );
  AND U4302 ( .A(n286), .B(n2762), .Z(n2760) );
  XOR U4303 ( .A(n2763), .B(n2764), .Z(n2762) );
  XOR U4304 ( .A(DB[1291]), .B(DB[1284]), .Z(n2764) );
  AND U4305 ( .A(n290), .B(n2765), .Z(n2763) );
  XOR U4306 ( .A(n2766), .B(n2767), .Z(n2765) );
  XOR U4307 ( .A(DB[1284]), .B(DB[1277]), .Z(n2767) );
  AND U4308 ( .A(n294), .B(n2768), .Z(n2766) );
  XOR U4309 ( .A(n2769), .B(n2770), .Z(n2768) );
  XOR U4310 ( .A(DB[1277]), .B(DB[1270]), .Z(n2770) );
  AND U4311 ( .A(n298), .B(n2771), .Z(n2769) );
  XOR U4312 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U4313 ( .A(DB[1270]), .B(DB[1263]), .Z(n2773) );
  AND U4314 ( .A(n302), .B(n2774), .Z(n2772) );
  XOR U4315 ( .A(n2775), .B(n2776), .Z(n2774) );
  XOR U4316 ( .A(DB[1263]), .B(DB[1256]), .Z(n2776) );
  AND U4317 ( .A(n306), .B(n2777), .Z(n2775) );
  XOR U4318 ( .A(n2778), .B(n2779), .Z(n2777) );
  XOR U4319 ( .A(DB[1256]), .B(DB[1249]), .Z(n2779) );
  AND U4320 ( .A(n310), .B(n2780), .Z(n2778) );
  XOR U4321 ( .A(n2781), .B(n2782), .Z(n2780) );
  XOR U4322 ( .A(DB[1249]), .B(DB[1242]), .Z(n2782) );
  AND U4323 ( .A(n314), .B(n2783), .Z(n2781) );
  XOR U4324 ( .A(n2784), .B(n2785), .Z(n2783) );
  XOR U4325 ( .A(DB[1242]), .B(DB[1235]), .Z(n2785) );
  AND U4326 ( .A(n318), .B(n2786), .Z(n2784) );
  XOR U4327 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U4328 ( .A(DB[1235]), .B(DB[1228]), .Z(n2788) );
  AND U4329 ( .A(n322), .B(n2789), .Z(n2787) );
  XOR U4330 ( .A(n2790), .B(n2791), .Z(n2789) );
  XOR U4331 ( .A(DB[1228]), .B(DB[1221]), .Z(n2791) );
  AND U4332 ( .A(n326), .B(n2792), .Z(n2790) );
  XOR U4333 ( .A(n2793), .B(n2794), .Z(n2792) );
  XOR U4334 ( .A(DB[1221]), .B(DB[1214]), .Z(n2794) );
  AND U4335 ( .A(n330), .B(n2795), .Z(n2793) );
  XOR U4336 ( .A(n2796), .B(n2797), .Z(n2795) );
  XOR U4337 ( .A(DB[1214]), .B(DB[1207]), .Z(n2797) );
  AND U4338 ( .A(n334), .B(n2798), .Z(n2796) );
  XOR U4339 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR U4340 ( .A(DB[1207]), .B(DB[1200]), .Z(n2800) );
  AND U4341 ( .A(n338), .B(n2801), .Z(n2799) );
  XOR U4342 ( .A(n2802), .B(n2803), .Z(n2801) );
  XOR U4343 ( .A(DB[1200]), .B(DB[1193]), .Z(n2803) );
  AND U4344 ( .A(n342), .B(n2804), .Z(n2802) );
  XOR U4345 ( .A(n2805), .B(n2806), .Z(n2804) );
  XOR U4346 ( .A(DB[1193]), .B(DB[1186]), .Z(n2806) );
  AND U4347 ( .A(n346), .B(n2807), .Z(n2805) );
  XOR U4348 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U4349 ( .A(DB[1186]), .B(DB[1179]), .Z(n2809) );
  AND U4350 ( .A(n350), .B(n2810), .Z(n2808) );
  XOR U4351 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR U4352 ( .A(DB[1179]), .B(DB[1172]), .Z(n2812) );
  AND U4353 ( .A(n354), .B(n2813), .Z(n2811) );
  XOR U4354 ( .A(n2814), .B(n2815), .Z(n2813) );
  XOR U4355 ( .A(DB[1172]), .B(DB[1165]), .Z(n2815) );
  AND U4356 ( .A(n358), .B(n2816), .Z(n2814) );
  XOR U4357 ( .A(n2817), .B(n2818), .Z(n2816) );
  XOR U4358 ( .A(DB[1165]), .B(DB[1158]), .Z(n2818) );
  AND U4359 ( .A(n362), .B(n2819), .Z(n2817) );
  XOR U4360 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U4361 ( .A(DB[1158]), .B(DB[1151]), .Z(n2821) );
  AND U4362 ( .A(n366), .B(n2822), .Z(n2820) );
  XOR U4363 ( .A(n2823), .B(n2824), .Z(n2822) );
  XOR U4364 ( .A(DB[1151]), .B(DB[1144]), .Z(n2824) );
  AND U4365 ( .A(n370), .B(n2825), .Z(n2823) );
  XOR U4366 ( .A(n2826), .B(n2827), .Z(n2825) );
  XOR U4367 ( .A(DB[1144]), .B(DB[1137]), .Z(n2827) );
  AND U4368 ( .A(n374), .B(n2828), .Z(n2826) );
  XOR U4369 ( .A(n2829), .B(n2830), .Z(n2828) );
  XOR U4370 ( .A(DB[1137]), .B(DB[1130]), .Z(n2830) );
  AND U4371 ( .A(n378), .B(n2831), .Z(n2829) );
  XOR U4372 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U4373 ( .A(DB[1130]), .B(DB[1123]), .Z(n2833) );
  AND U4374 ( .A(n382), .B(n2834), .Z(n2832) );
  XOR U4375 ( .A(n2835), .B(n2836), .Z(n2834) );
  XOR U4376 ( .A(DB[1123]), .B(DB[1116]), .Z(n2836) );
  AND U4377 ( .A(n386), .B(n2837), .Z(n2835) );
  XOR U4378 ( .A(n2838), .B(n2839), .Z(n2837) );
  XOR U4379 ( .A(DB[1116]), .B(DB[1109]), .Z(n2839) );
  AND U4380 ( .A(n390), .B(n2840), .Z(n2838) );
  XOR U4381 ( .A(n2841), .B(n2842), .Z(n2840) );
  XOR U4382 ( .A(DB[1109]), .B(DB[1102]), .Z(n2842) );
  AND U4383 ( .A(n394), .B(n2843), .Z(n2841) );
  XOR U4384 ( .A(n2844), .B(n2845), .Z(n2843) );
  XOR U4385 ( .A(DB[1102]), .B(DB[1095]), .Z(n2845) );
  AND U4386 ( .A(n398), .B(n2846), .Z(n2844) );
  XOR U4387 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U4388 ( .A(DB[1095]), .B(DB[1088]), .Z(n2848) );
  AND U4389 ( .A(n402), .B(n2849), .Z(n2847) );
  XOR U4390 ( .A(n2850), .B(n2851), .Z(n2849) );
  XOR U4391 ( .A(DB[1088]), .B(DB[1081]), .Z(n2851) );
  AND U4392 ( .A(n406), .B(n2852), .Z(n2850) );
  XOR U4393 ( .A(n2853), .B(n2854), .Z(n2852) );
  XOR U4394 ( .A(DB[1081]), .B(DB[1074]), .Z(n2854) );
  AND U4395 ( .A(n410), .B(n2855), .Z(n2853) );
  XOR U4396 ( .A(n2856), .B(n2857), .Z(n2855) );
  XOR U4397 ( .A(DB[1074]), .B(DB[1067]), .Z(n2857) );
  AND U4398 ( .A(n414), .B(n2858), .Z(n2856) );
  XOR U4399 ( .A(n2859), .B(n2860), .Z(n2858) );
  XOR U4400 ( .A(DB[1067]), .B(DB[1060]), .Z(n2860) );
  AND U4401 ( .A(n418), .B(n2861), .Z(n2859) );
  XOR U4402 ( .A(n2862), .B(n2863), .Z(n2861) );
  XOR U4403 ( .A(DB[1060]), .B(DB[1053]), .Z(n2863) );
  AND U4404 ( .A(n422), .B(n2864), .Z(n2862) );
  XOR U4405 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR U4406 ( .A(DB[1053]), .B(DB[1046]), .Z(n2866) );
  AND U4407 ( .A(n426), .B(n2867), .Z(n2865) );
  XOR U4408 ( .A(n2868), .B(n2869), .Z(n2867) );
  XOR U4409 ( .A(DB[1046]), .B(DB[1039]), .Z(n2869) );
  AND U4410 ( .A(n430), .B(n2870), .Z(n2868) );
  XOR U4411 ( .A(n2871), .B(n2872), .Z(n2870) );
  XOR U4412 ( .A(DB[1039]), .B(DB[1032]), .Z(n2872) );
  AND U4413 ( .A(n434), .B(n2873), .Z(n2871) );
  XOR U4414 ( .A(n2874), .B(n2875), .Z(n2873) );
  XOR U4415 ( .A(DB[1032]), .B(DB[1025]), .Z(n2875) );
  AND U4416 ( .A(n438), .B(n2876), .Z(n2874) );
  XOR U4417 ( .A(n2877), .B(n2878), .Z(n2876) );
  XOR U4418 ( .A(DB[1025]), .B(DB[1018]), .Z(n2878) );
  AND U4419 ( .A(n442), .B(n2879), .Z(n2877) );
  XOR U4420 ( .A(n2880), .B(n2881), .Z(n2879) );
  XOR U4421 ( .A(DB[1018]), .B(DB[1011]), .Z(n2881) );
  AND U4422 ( .A(n446), .B(n2882), .Z(n2880) );
  XOR U4423 ( .A(n2883), .B(n2884), .Z(n2882) );
  XOR U4424 ( .A(DB[1011]), .B(DB[1004]), .Z(n2884) );
  AND U4425 ( .A(n450), .B(n2885), .Z(n2883) );
  XOR U4426 ( .A(n2886), .B(n2887), .Z(n2885) );
  XOR U4427 ( .A(DB[997]), .B(DB[1004]), .Z(n2887) );
  AND U4428 ( .A(n454), .B(n2888), .Z(n2886) );
  XOR U4429 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR U4430 ( .A(DB[997]), .B(DB[990]), .Z(n2890) );
  AND U4431 ( .A(n458), .B(n2891), .Z(n2889) );
  XOR U4432 ( .A(n2892), .B(n2893), .Z(n2891) );
  XOR U4433 ( .A(DB[990]), .B(DB[983]), .Z(n2893) );
  AND U4434 ( .A(n462), .B(n2894), .Z(n2892) );
  XOR U4435 ( .A(n2895), .B(n2896), .Z(n2894) );
  XOR U4436 ( .A(DB[983]), .B(DB[976]), .Z(n2896) );
  AND U4437 ( .A(n466), .B(n2897), .Z(n2895) );
  XOR U4438 ( .A(n2898), .B(n2899), .Z(n2897) );
  XOR U4439 ( .A(DB[976]), .B(DB[969]), .Z(n2899) );
  AND U4440 ( .A(n470), .B(n2900), .Z(n2898) );
  XOR U4441 ( .A(n2901), .B(n2902), .Z(n2900) );
  XOR U4442 ( .A(DB[969]), .B(DB[962]), .Z(n2902) );
  AND U4443 ( .A(n474), .B(n2903), .Z(n2901) );
  XOR U4444 ( .A(n2904), .B(n2905), .Z(n2903) );
  XOR U4445 ( .A(DB[962]), .B(DB[955]), .Z(n2905) );
  AND U4446 ( .A(n478), .B(n2906), .Z(n2904) );
  XOR U4447 ( .A(n2907), .B(n2908), .Z(n2906) );
  XOR U4448 ( .A(DB[955]), .B(DB[948]), .Z(n2908) );
  AND U4449 ( .A(n482), .B(n2909), .Z(n2907) );
  XOR U4450 ( .A(n2910), .B(n2911), .Z(n2909) );
  XOR U4451 ( .A(DB[948]), .B(DB[941]), .Z(n2911) );
  AND U4452 ( .A(n486), .B(n2912), .Z(n2910) );
  XOR U4453 ( .A(n2913), .B(n2914), .Z(n2912) );
  XOR U4454 ( .A(DB[941]), .B(DB[934]), .Z(n2914) );
  AND U4455 ( .A(n490), .B(n2915), .Z(n2913) );
  XOR U4456 ( .A(n2916), .B(n2917), .Z(n2915) );
  XOR U4457 ( .A(DB[934]), .B(DB[927]), .Z(n2917) );
  AND U4458 ( .A(n494), .B(n2918), .Z(n2916) );
  XOR U4459 ( .A(n2919), .B(n2920), .Z(n2918) );
  XOR U4460 ( .A(DB[927]), .B(DB[920]), .Z(n2920) );
  AND U4461 ( .A(n498), .B(n2921), .Z(n2919) );
  XOR U4462 ( .A(n2922), .B(n2923), .Z(n2921) );
  XOR U4463 ( .A(DB[920]), .B(DB[913]), .Z(n2923) );
  AND U4464 ( .A(n502), .B(n2924), .Z(n2922) );
  XOR U4465 ( .A(n2925), .B(n2926), .Z(n2924) );
  XOR U4466 ( .A(DB[913]), .B(DB[906]), .Z(n2926) );
  AND U4467 ( .A(n506), .B(n2927), .Z(n2925) );
  XOR U4468 ( .A(n2928), .B(n2929), .Z(n2927) );
  XOR U4469 ( .A(DB[906]), .B(DB[899]), .Z(n2929) );
  AND U4470 ( .A(n510), .B(n2930), .Z(n2928) );
  XOR U4471 ( .A(n2931), .B(n2932), .Z(n2930) );
  XOR U4472 ( .A(DB[899]), .B(DB[892]), .Z(n2932) );
  AND U4473 ( .A(n514), .B(n2933), .Z(n2931) );
  XOR U4474 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR U4475 ( .A(DB[892]), .B(DB[885]), .Z(n2935) );
  AND U4476 ( .A(n518), .B(n2936), .Z(n2934) );
  XOR U4477 ( .A(n2937), .B(n2938), .Z(n2936) );
  XOR U4478 ( .A(DB[885]), .B(DB[878]), .Z(n2938) );
  AND U4479 ( .A(n522), .B(n2939), .Z(n2937) );
  XOR U4480 ( .A(n2940), .B(n2941), .Z(n2939) );
  XOR U4481 ( .A(DB[878]), .B(DB[871]), .Z(n2941) );
  AND U4482 ( .A(n526), .B(n2942), .Z(n2940) );
  XOR U4483 ( .A(n2943), .B(n2944), .Z(n2942) );
  XOR U4484 ( .A(DB[871]), .B(DB[864]), .Z(n2944) );
  AND U4485 ( .A(n530), .B(n2945), .Z(n2943) );
  XOR U4486 ( .A(n2946), .B(n2947), .Z(n2945) );
  XOR U4487 ( .A(DB[864]), .B(DB[857]), .Z(n2947) );
  AND U4488 ( .A(n534), .B(n2948), .Z(n2946) );
  XOR U4489 ( .A(n2949), .B(n2950), .Z(n2948) );
  XOR U4490 ( .A(DB[857]), .B(DB[850]), .Z(n2950) );
  AND U4491 ( .A(n538), .B(n2951), .Z(n2949) );
  XOR U4492 ( .A(n2952), .B(n2953), .Z(n2951) );
  XOR U4493 ( .A(DB[850]), .B(DB[843]), .Z(n2953) );
  AND U4494 ( .A(n542), .B(n2954), .Z(n2952) );
  XOR U4495 ( .A(n2955), .B(n2956), .Z(n2954) );
  XOR U4496 ( .A(DB[843]), .B(DB[836]), .Z(n2956) );
  AND U4497 ( .A(n546), .B(n2957), .Z(n2955) );
  XOR U4498 ( .A(n2958), .B(n2959), .Z(n2957) );
  XOR U4499 ( .A(DB[836]), .B(DB[829]), .Z(n2959) );
  AND U4500 ( .A(n550), .B(n2960), .Z(n2958) );
  XOR U4501 ( .A(n2961), .B(n2962), .Z(n2960) );
  XOR U4502 ( .A(DB[829]), .B(DB[822]), .Z(n2962) );
  AND U4503 ( .A(n554), .B(n2963), .Z(n2961) );
  XOR U4504 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR U4505 ( .A(DB[822]), .B(DB[815]), .Z(n2965) );
  AND U4506 ( .A(n558), .B(n2966), .Z(n2964) );
  XOR U4507 ( .A(n2967), .B(n2968), .Z(n2966) );
  XOR U4508 ( .A(DB[815]), .B(DB[808]), .Z(n2968) );
  AND U4509 ( .A(n562), .B(n2969), .Z(n2967) );
  XOR U4510 ( .A(n2970), .B(n2971), .Z(n2969) );
  XOR U4511 ( .A(DB[808]), .B(DB[801]), .Z(n2971) );
  AND U4512 ( .A(n566), .B(n2972), .Z(n2970) );
  XOR U4513 ( .A(n2973), .B(n2974), .Z(n2972) );
  XOR U4514 ( .A(DB[801]), .B(DB[794]), .Z(n2974) );
  AND U4515 ( .A(n570), .B(n2975), .Z(n2973) );
  XOR U4516 ( .A(n2976), .B(n2977), .Z(n2975) );
  XOR U4517 ( .A(DB[794]), .B(DB[787]), .Z(n2977) );
  AND U4518 ( .A(n574), .B(n2978), .Z(n2976) );
  XOR U4519 ( .A(n2979), .B(n2980), .Z(n2978) );
  XOR U4520 ( .A(DB[787]), .B(DB[780]), .Z(n2980) );
  AND U4521 ( .A(n578), .B(n2981), .Z(n2979) );
  XOR U4522 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR U4523 ( .A(DB[780]), .B(DB[773]), .Z(n2983) );
  AND U4524 ( .A(n582), .B(n2984), .Z(n2982) );
  XOR U4525 ( .A(n2985), .B(n2986), .Z(n2984) );
  XOR U4526 ( .A(DB[773]), .B(DB[766]), .Z(n2986) );
  AND U4527 ( .A(n586), .B(n2987), .Z(n2985) );
  XOR U4528 ( .A(n2988), .B(n2989), .Z(n2987) );
  XOR U4529 ( .A(DB[766]), .B(DB[759]), .Z(n2989) );
  AND U4530 ( .A(n590), .B(n2990), .Z(n2988) );
  XOR U4531 ( .A(n2991), .B(n2992), .Z(n2990) );
  XOR U4532 ( .A(DB[759]), .B(DB[752]), .Z(n2992) );
  AND U4533 ( .A(n594), .B(n2993), .Z(n2991) );
  XOR U4534 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U4535 ( .A(DB[752]), .B(DB[745]), .Z(n2995) );
  AND U4536 ( .A(n598), .B(n2996), .Z(n2994) );
  XOR U4537 ( .A(n2997), .B(n2998), .Z(n2996) );
  XOR U4538 ( .A(DB[745]), .B(DB[738]), .Z(n2998) );
  AND U4539 ( .A(n602), .B(n2999), .Z(n2997) );
  XOR U4540 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U4541 ( .A(DB[738]), .B(DB[731]), .Z(n3001) );
  AND U4542 ( .A(n606), .B(n3002), .Z(n3000) );
  XOR U4543 ( .A(n3003), .B(n3004), .Z(n3002) );
  XOR U4544 ( .A(DB[731]), .B(DB[724]), .Z(n3004) );
  AND U4545 ( .A(n610), .B(n3005), .Z(n3003) );
  XOR U4546 ( .A(n3006), .B(n3007), .Z(n3005) );
  XOR U4547 ( .A(DB[724]), .B(DB[717]), .Z(n3007) );
  AND U4548 ( .A(n614), .B(n3008), .Z(n3006) );
  XOR U4549 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR U4550 ( .A(DB[717]), .B(DB[710]), .Z(n3010) );
  AND U4551 ( .A(n618), .B(n3011), .Z(n3009) );
  XOR U4552 ( .A(n3012), .B(n3013), .Z(n3011) );
  XOR U4553 ( .A(DB[710]), .B(DB[703]), .Z(n3013) );
  AND U4554 ( .A(n622), .B(n3014), .Z(n3012) );
  XOR U4555 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U4556 ( .A(DB[703]), .B(DB[696]), .Z(n3016) );
  AND U4557 ( .A(n626), .B(n3017), .Z(n3015) );
  XOR U4558 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U4559 ( .A(DB[696]), .B(DB[689]), .Z(n3019) );
  AND U4560 ( .A(n630), .B(n3020), .Z(n3018) );
  XOR U4561 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR U4562 ( .A(DB[689]), .B(DB[682]), .Z(n3022) );
  AND U4563 ( .A(n634), .B(n3023), .Z(n3021) );
  XOR U4564 ( .A(n3024), .B(n3025), .Z(n3023) );
  XOR U4565 ( .A(DB[682]), .B(DB[675]), .Z(n3025) );
  AND U4566 ( .A(n638), .B(n3026), .Z(n3024) );
  XOR U4567 ( .A(n3027), .B(n3028), .Z(n3026) );
  XOR U4568 ( .A(DB[675]), .B(DB[668]), .Z(n3028) );
  AND U4569 ( .A(n642), .B(n3029), .Z(n3027) );
  XOR U4570 ( .A(n3030), .B(n3031), .Z(n3029) );
  XOR U4571 ( .A(DB[668]), .B(DB[661]), .Z(n3031) );
  AND U4572 ( .A(n646), .B(n3032), .Z(n3030) );
  XOR U4573 ( .A(n3033), .B(n3034), .Z(n3032) );
  XOR U4574 ( .A(DB[661]), .B(DB[654]), .Z(n3034) );
  AND U4575 ( .A(n650), .B(n3035), .Z(n3033) );
  XOR U4576 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U4577 ( .A(DB[654]), .B(DB[647]), .Z(n3037) );
  AND U4578 ( .A(n654), .B(n3038), .Z(n3036) );
  XOR U4579 ( .A(n3039), .B(n3040), .Z(n3038) );
  XOR U4580 ( .A(DB[647]), .B(DB[640]), .Z(n3040) );
  AND U4581 ( .A(n658), .B(n3041), .Z(n3039) );
  XOR U4582 ( .A(n3042), .B(n3043), .Z(n3041) );
  XOR U4583 ( .A(DB[640]), .B(DB[633]), .Z(n3043) );
  AND U4584 ( .A(n662), .B(n3044), .Z(n3042) );
  XOR U4585 ( .A(n3045), .B(n3046), .Z(n3044) );
  XOR U4586 ( .A(DB[633]), .B(DB[626]), .Z(n3046) );
  AND U4587 ( .A(n666), .B(n3047), .Z(n3045) );
  XOR U4588 ( .A(n3048), .B(n3049), .Z(n3047) );
  XOR U4589 ( .A(DB[626]), .B(DB[619]), .Z(n3049) );
  AND U4590 ( .A(n670), .B(n3050), .Z(n3048) );
  XOR U4591 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U4592 ( .A(DB[619]), .B(DB[612]), .Z(n3052) );
  AND U4593 ( .A(n674), .B(n3053), .Z(n3051) );
  XOR U4594 ( .A(n3054), .B(n3055), .Z(n3053) );
  XOR U4595 ( .A(DB[612]), .B(DB[605]), .Z(n3055) );
  AND U4596 ( .A(n678), .B(n3056), .Z(n3054) );
  XOR U4597 ( .A(n3057), .B(n3058), .Z(n3056) );
  XOR U4598 ( .A(DB[605]), .B(DB[598]), .Z(n3058) );
  AND U4599 ( .A(n682), .B(n3059), .Z(n3057) );
  XOR U4600 ( .A(n3060), .B(n3061), .Z(n3059) );
  XOR U4601 ( .A(DB[598]), .B(DB[591]), .Z(n3061) );
  AND U4602 ( .A(n686), .B(n3062), .Z(n3060) );
  XOR U4603 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR U4604 ( .A(DB[591]), .B(DB[584]), .Z(n3064) );
  AND U4605 ( .A(n690), .B(n3065), .Z(n3063) );
  XOR U4606 ( .A(n3066), .B(n3067), .Z(n3065) );
  XOR U4607 ( .A(DB[584]), .B(DB[577]), .Z(n3067) );
  AND U4608 ( .A(n694), .B(n3068), .Z(n3066) );
  XOR U4609 ( .A(n3069), .B(n3070), .Z(n3068) );
  XOR U4610 ( .A(DB[577]), .B(DB[570]), .Z(n3070) );
  AND U4611 ( .A(n698), .B(n3071), .Z(n3069) );
  XOR U4612 ( .A(n3072), .B(n3073), .Z(n3071) );
  XOR U4613 ( .A(DB[570]), .B(DB[563]), .Z(n3073) );
  AND U4614 ( .A(n702), .B(n3074), .Z(n3072) );
  XOR U4615 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR U4616 ( .A(DB[563]), .B(DB[556]), .Z(n3076) );
  AND U4617 ( .A(n706), .B(n3077), .Z(n3075) );
  XOR U4618 ( .A(n3078), .B(n3079), .Z(n3077) );
  XOR U4619 ( .A(DB[556]), .B(DB[549]), .Z(n3079) );
  AND U4620 ( .A(n710), .B(n3080), .Z(n3078) );
  XOR U4621 ( .A(n3081), .B(n3082), .Z(n3080) );
  XOR U4622 ( .A(DB[549]), .B(DB[542]), .Z(n3082) );
  AND U4623 ( .A(n714), .B(n3083), .Z(n3081) );
  XOR U4624 ( .A(n3084), .B(n3085), .Z(n3083) );
  XOR U4625 ( .A(DB[542]), .B(DB[535]), .Z(n3085) );
  AND U4626 ( .A(n718), .B(n3086), .Z(n3084) );
  XOR U4627 ( .A(n3087), .B(n3088), .Z(n3086) );
  XOR U4628 ( .A(DB[535]), .B(DB[528]), .Z(n3088) );
  AND U4629 ( .A(n722), .B(n3089), .Z(n3087) );
  XOR U4630 ( .A(n3090), .B(n3091), .Z(n3089) );
  XOR U4631 ( .A(DB[528]), .B(DB[521]), .Z(n3091) );
  AND U4632 ( .A(n726), .B(n3092), .Z(n3090) );
  XOR U4633 ( .A(n3093), .B(n3094), .Z(n3092) );
  XOR U4634 ( .A(DB[521]), .B(DB[514]), .Z(n3094) );
  AND U4635 ( .A(n730), .B(n3095), .Z(n3093) );
  XOR U4636 ( .A(n3096), .B(n3097), .Z(n3095) );
  XOR U4637 ( .A(DB[514]), .B(DB[507]), .Z(n3097) );
  AND U4638 ( .A(n734), .B(n3098), .Z(n3096) );
  XOR U4639 ( .A(n3099), .B(n3100), .Z(n3098) );
  XOR U4640 ( .A(DB[507]), .B(DB[500]), .Z(n3100) );
  AND U4641 ( .A(n738), .B(n3101), .Z(n3099) );
  XOR U4642 ( .A(n3102), .B(n3103), .Z(n3101) );
  XOR U4643 ( .A(DB[500]), .B(DB[493]), .Z(n3103) );
  AND U4644 ( .A(n742), .B(n3104), .Z(n3102) );
  XOR U4645 ( .A(n3105), .B(n3106), .Z(n3104) );
  XOR U4646 ( .A(DB[493]), .B(DB[486]), .Z(n3106) );
  AND U4647 ( .A(n746), .B(n3107), .Z(n3105) );
  XOR U4648 ( .A(n3108), .B(n3109), .Z(n3107) );
  XOR U4649 ( .A(DB[486]), .B(DB[479]), .Z(n3109) );
  AND U4650 ( .A(n750), .B(n3110), .Z(n3108) );
  XOR U4651 ( .A(n3111), .B(n3112), .Z(n3110) );
  XOR U4652 ( .A(DB[479]), .B(DB[472]), .Z(n3112) );
  AND U4653 ( .A(n754), .B(n3113), .Z(n3111) );
  XOR U4654 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR U4655 ( .A(DB[472]), .B(DB[465]), .Z(n3115) );
  AND U4656 ( .A(n758), .B(n3116), .Z(n3114) );
  XOR U4657 ( .A(n3117), .B(n3118), .Z(n3116) );
  XOR U4658 ( .A(DB[465]), .B(DB[458]), .Z(n3118) );
  AND U4659 ( .A(n762), .B(n3119), .Z(n3117) );
  XOR U4660 ( .A(n3120), .B(n3121), .Z(n3119) );
  XOR U4661 ( .A(DB[458]), .B(DB[451]), .Z(n3121) );
  AND U4662 ( .A(n766), .B(n3122), .Z(n3120) );
  XOR U4663 ( .A(n3123), .B(n3124), .Z(n3122) );
  XOR U4664 ( .A(DB[451]), .B(DB[444]), .Z(n3124) );
  AND U4665 ( .A(n770), .B(n3125), .Z(n3123) );
  XOR U4666 ( .A(n3126), .B(n3127), .Z(n3125) );
  XOR U4667 ( .A(DB[444]), .B(DB[437]), .Z(n3127) );
  AND U4668 ( .A(n774), .B(n3128), .Z(n3126) );
  XOR U4669 ( .A(n3129), .B(n3130), .Z(n3128) );
  XOR U4670 ( .A(DB[437]), .B(DB[430]), .Z(n3130) );
  AND U4671 ( .A(n778), .B(n3131), .Z(n3129) );
  XOR U4672 ( .A(n3132), .B(n3133), .Z(n3131) );
  XOR U4673 ( .A(DB[430]), .B(DB[423]), .Z(n3133) );
  AND U4674 ( .A(n782), .B(n3134), .Z(n3132) );
  XOR U4675 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U4676 ( .A(DB[423]), .B(DB[416]), .Z(n3136) );
  AND U4677 ( .A(n786), .B(n3137), .Z(n3135) );
  XOR U4678 ( .A(n3138), .B(n3139), .Z(n3137) );
  XOR U4679 ( .A(DB[416]), .B(DB[409]), .Z(n3139) );
  AND U4680 ( .A(n790), .B(n3140), .Z(n3138) );
  XOR U4681 ( .A(n3141), .B(n3142), .Z(n3140) );
  XOR U4682 ( .A(DB[409]), .B(DB[402]), .Z(n3142) );
  AND U4683 ( .A(n794), .B(n3143), .Z(n3141) );
  XOR U4684 ( .A(n3144), .B(n3145), .Z(n3143) );
  XOR U4685 ( .A(DB[402]), .B(DB[395]), .Z(n3145) );
  AND U4686 ( .A(n798), .B(n3146), .Z(n3144) );
  XOR U4687 ( .A(n3147), .B(n3148), .Z(n3146) );
  XOR U4688 ( .A(DB[395]), .B(DB[388]), .Z(n3148) );
  AND U4689 ( .A(n802), .B(n3149), .Z(n3147) );
  XOR U4690 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U4691 ( .A(DB[388]), .B(DB[381]), .Z(n3151) );
  AND U4692 ( .A(n806), .B(n3152), .Z(n3150) );
  XOR U4693 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U4694 ( .A(DB[381]), .B(DB[374]), .Z(n3154) );
  AND U4695 ( .A(n810), .B(n3155), .Z(n3153) );
  XOR U4696 ( .A(n3156), .B(n3157), .Z(n3155) );
  XOR U4697 ( .A(DB[374]), .B(DB[367]), .Z(n3157) );
  AND U4698 ( .A(n814), .B(n3158), .Z(n3156) );
  XOR U4699 ( .A(n3159), .B(n3160), .Z(n3158) );
  XOR U4700 ( .A(DB[367]), .B(DB[360]), .Z(n3160) );
  AND U4701 ( .A(n818), .B(n3161), .Z(n3159) );
  XOR U4702 ( .A(n3162), .B(n3163), .Z(n3161) );
  XOR U4703 ( .A(DB[360]), .B(DB[353]), .Z(n3163) );
  AND U4704 ( .A(n822), .B(n3164), .Z(n3162) );
  XOR U4705 ( .A(n3165), .B(n3166), .Z(n3164) );
  XOR U4706 ( .A(DB[353]), .B(DB[346]), .Z(n3166) );
  AND U4707 ( .A(n826), .B(n3167), .Z(n3165) );
  XOR U4708 ( .A(n3168), .B(n3169), .Z(n3167) );
  XOR U4709 ( .A(DB[346]), .B(DB[339]), .Z(n3169) );
  AND U4710 ( .A(n830), .B(n3170), .Z(n3168) );
  XOR U4711 ( .A(n3171), .B(n3172), .Z(n3170) );
  XOR U4712 ( .A(DB[339]), .B(DB[332]), .Z(n3172) );
  AND U4713 ( .A(n834), .B(n3173), .Z(n3171) );
  XOR U4714 ( .A(n3174), .B(n3175), .Z(n3173) );
  XOR U4715 ( .A(DB[332]), .B(DB[325]), .Z(n3175) );
  AND U4716 ( .A(n838), .B(n3176), .Z(n3174) );
  XOR U4717 ( .A(n3177), .B(n3178), .Z(n3176) );
  XOR U4718 ( .A(DB[325]), .B(DB[318]), .Z(n3178) );
  AND U4719 ( .A(n842), .B(n3179), .Z(n3177) );
  XOR U4720 ( .A(n3180), .B(n3181), .Z(n3179) );
  XOR U4721 ( .A(DB[318]), .B(DB[311]), .Z(n3181) );
  AND U4722 ( .A(n846), .B(n3182), .Z(n3180) );
  XOR U4723 ( .A(n3183), .B(n3184), .Z(n3182) );
  XOR U4724 ( .A(DB[311]), .B(DB[304]), .Z(n3184) );
  AND U4725 ( .A(n850), .B(n3185), .Z(n3183) );
  XOR U4726 ( .A(n3186), .B(n3187), .Z(n3185) );
  XOR U4727 ( .A(DB[304]), .B(DB[297]), .Z(n3187) );
  AND U4728 ( .A(n854), .B(n3188), .Z(n3186) );
  XOR U4729 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U4730 ( .A(DB[297]), .B(DB[290]), .Z(n3190) );
  AND U4731 ( .A(n858), .B(n3191), .Z(n3189) );
  XOR U4732 ( .A(n3192), .B(n3193), .Z(n3191) );
  XOR U4733 ( .A(DB[290]), .B(DB[283]), .Z(n3193) );
  AND U4734 ( .A(n862), .B(n3194), .Z(n3192) );
  XOR U4735 ( .A(n3195), .B(n3196), .Z(n3194) );
  XOR U4736 ( .A(DB[283]), .B(DB[276]), .Z(n3196) );
  AND U4737 ( .A(n866), .B(n3197), .Z(n3195) );
  XOR U4738 ( .A(n3198), .B(n3199), .Z(n3197) );
  XOR U4739 ( .A(DB[276]), .B(DB[269]), .Z(n3199) );
  AND U4740 ( .A(n870), .B(n3200), .Z(n3198) );
  XOR U4741 ( .A(n3201), .B(n3202), .Z(n3200) );
  XOR U4742 ( .A(DB[269]), .B(DB[262]), .Z(n3202) );
  AND U4743 ( .A(n874), .B(n3203), .Z(n3201) );
  XOR U4744 ( .A(n3204), .B(n3205), .Z(n3203) );
  XOR U4745 ( .A(DB[262]), .B(DB[255]), .Z(n3205) );
  AND U4746 ( .A(n878), .B(n3206), .Z(n3204) );
  XOR U4747 ( .A(n3207), .B(n3208), .Z(n3206) );
  XOR U4748 ( .A(DB[255]), .B(DB[248]), .Z(n3208) );
  AND U4749 ( .A(n882), .B(n3209), .Z(n3207) );
  XOR U4750 ( .A(n3210), .B(n3211), .Z(n3209) );
  XOR U4751 ( .A(DB[248]), .B(DB[241]), .Z(n3211) );
  AND U4752 ( .A(n886), .B(n3212), .Z(n3210) );
  XOR U4753 ( .A(n3213), .B(n3214), .Z(n3212) );
  XOR U4754 ( .A(DB[241]), .B(DB[234]), .Z(n3214) );
  AND U4755 ( .A(n890), .B(n3215), .Z(n3213) );
  XOR U4756 ( .A(n3216), .B(n3217), .Z(n3215) );
  XOR U4757 ( .A(DB[234]), .B(DB[227]), .Z(n3217) );
  AND U4758 ( .A(n894), .B(n3218), .Z(n3216) );
  XOR U4759 ( .A(n3219), .B(n3220), .Z(n3218) );
  XOR U4760 ( .A(DB[227]), .B(DB[220]), .Z(n3220) );
  AND U4761 ( .A(n898), .B(n3221), .Z(n3219) );
  XOR U4762 ( .A(n3222), .B(n3223), .Z(n3221) );
  XOR U4763 ( .A(DB[220]), .B(DB[213]), .Z(n3223) );
  AND U4764 ( .A(n902), .B(n3224), .Z(n3222) );
  XOR U4765 ( .A(n3225), .B(n3226), .Z(n3224) );
  XOR U4766 ( .A(DB[213]), .B(DB[206]), .Z(n3226) );
  AND U4767 ( .A(n906), .B(n3227), .Z(n3225) );
  XOR U4768 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR U4769 ( .A(DB[206]), .B(DB[199]), .Z(n3229) );
  AND U4770 ( .A(n910), .B(n3230), .Z(n3228) );
  XOR U4771 ( .A(n3231), .B(n3232), .Z(n3230) );
  XOR U4772 ( .A(DB[199]), .B(DB[192]), .Z(n3232) );
  AND U4773 ( .A(n914), .B(n3233), .Z(n3231) );
  XOR U4774 ( .A(n3234), .B(n3235), .Z(n3233) );
  XOR U4775 ( .A(DB[192]), .B(DB[185]), .Z(n3235) );
  AND U4776 ( .A(n918), .B(n3236), .Z(n3234) );
  XOR U4777 ( .A(n3237), .B(n3238), .Z(n3236) );
  XOR U4778 ( .A(DB[185]), .B(DB[178]), .Z(n3238) );
  AND U4779 ( .A(n922), .B(n3239), .Z(n3237) );
  XOR U4780 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U4781 ( .A(DB[178]), .B(DB[171]), .Z(n3241) );
  AND U4782 ( .A(n926), .B(n3242), .Z(n3240) );
  XOR U4783 ( .A(n3243), .B(n3244), .Z(n3242) );
  XOR U4784 ( .A(DB[171]), .B(DB[164]), .Z(n3244) );
  AND U4785 ( .A(n930), .B(n3245), .Z(n3243) );
  XOR U4786 ( .A(n3246), .B(n3247), .Z(n3245) );
  XOR U4787 ( .A(DB[164]), .B(DB[157]), .Z(n3247) );
  AND U4788 ( .A(n934), .B(n3248), .Z(n3246) );
  XOR U4789 ( .A(n3249), .B(n3250), .Z(n3248) );
  XOR U4790 ( .A(DB[157]), .B(DB[150]), .Z(n3250) );
  AND U4791 ( .A(n938), .B(n3251), .Z(n3249) );
  XOR U4792 ( .A(n3252), .B(n3253), .Z(n3251) );
  XOR U4793 ( .A(DB[150]), .B(DB[143]), .Z(n3253) );
  AND U4794 ( .A(n942), .B(n3254), .Z(n3252) );
  XOR U4795 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U4796 ( .A(DB[143]), .B(DB[136]), .Z(n3256) );
  AND U4797 ( .A(n946), .B(n3257), .Z(n3255) );
  XOR U4798 ( .A(n3258), .B(n3259), .Z(n3257) );
  XOR U4799 ( .A(DB[136]), .B(DB[129]), .Z(n3259) );
  AND U4800 ( .A(n950), .B(n3260), .Z(n3258) );
  XOR U4801 ( .A(n3261), .B(n3262), .Z(n3260) );
  XOR U4802 ( .A(DB[129]), .B(DB[122]), .Z(n3262) );
  AND U4803 ( .A(n954), .B(n3263), .Z(n3261) );
  XOR U4804 ( .A(n3264), .B(n3265), .Z(n3263) );
  XOR U4805 ( .A(DB[122]), .B(DB[115]), .Z(n3265) );
  AND U4806 ( .A(n958), .B(n3266), .Z(n3264) );
  XOR U4807 ( .A(n3267), .B(n3268), .Z(n3266) );
  XOR U4808 ( .A(DB[115]), .B(DB[108]), .Z(n3268) );
  AND U4809 ( .A(n962), .B(n3269), .Z(n3267) );
  XOR U4810 ( .A(n3270), .B(n3271), .Z(n3269) );
  XOR U4811 ( .A(DB[108]), .B(DB[101]), .Z(n3271) );
  AND U4812 ( .A(n966), .B(n3272), .Z(n3270) );
  XOR U4813 ( .A(n3273), .B(n3274), .Z(n3272) );
  XOR U4814 ( .A(DB[94]), .B(DB[101]), .Z(n3274) );
  AND U4815 ( .A(n970), .B(n3275), .Z(n3273) );
  XOR U4816 ( .A(n3276), .B(n3277), .Z(n3275) );
  XOR U4817 ( .A(DB[94]), .B(DB[87]), .Z(n3277) );
  AND U4818 ( .A(n974), .B(n3278), .Z(n3276) );
  XOR U4819 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR U4820 ( .A(DB[87]), .B(DB[80]), .Z(n3280) );
  AND U4821 ( .A(n978), .B(n3281), .Z(n3279) );
  XOR U4822 ( .A(n3282), .B(n3283), .Z(n3281) );
  XOR U4823 ( .A(DB[80]), .B(DB[73]), .Z(n3283) );
  AND U4824 ( .A(n982), .B(n3284), .Z(n3282) );
  XOR U4825 ( .A(n3285), .B(n3286), .Z(n3284) );
  XOR U4826 ( .A(DB[73]), .B(DB[66]), .Z(n3286) );
  AND U4827 ( .A(n986), .B(n3287), .Z(n3285) );
  XOR U4828 ( .A(n3288), .B(n3289), .Z(n3287) );
  XOR U4829 ( .A(DB[66]), .B(DB[59]), .Z(n3289) );
  AND U4830 ( .A(n990), .B(n3290), .Z(n3288) );
  XOR U4831 ( .A(n3291), .B(n3292), .Z(n3290) );
  XOR U4832 ( .A(DB[59]), .B(DB[52]), .Z(n3292) );
  AND U4833 ( .A(n994), .B(n3293), .Z(n3291) );
  XOR U4834 ( .A(n3294), .B(n3295), .Z(n3293) );
  XOR U4835 ( .A(DB[52]), .B(DB[45]), .Z(n3295) );
  AND U4836 ( .A(n998), .B(n3296), .Z(n3294) );
  XOR U4837 ( .A(n3297), .B(n3298), .Z(n3296) );
  XOR U4838 ( .A(DB[45]), .B(DB[38]), .Z(n3298) );
  AND U4839 ( .A(n1002), .B(n3299), .Z(n3297) );
  XOR U4840 ( .A(n3300), .B(n3301), .Z(n3299) );
  XOR U4841 ( .A(DB[38]), .B(DB[31]), .Z(n3301) );
  AND U4842 ( .A(n1006), .B(n3302), .Z(n3300) );
  XOR U4843 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR U4844 ( .A(DB[31]), .B(DB[24]), .Z(n3304) );
  AND U4845 ( .A(n1010), .B(n3305), .Z(n3303) );
  XOR U4846 ( .A(n3306), .B(n3307), .Z(n3305) );
  XOR U4847 ( .A(DB[24]), .B(DB[17]), .Z(n3307) );
  AND U4848 ( .A(n1014), .B(n3308), .Z(n3306) );
  XOR U4849 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR U4850 ( .A(DB[17]), .B(DB[10]), .Z(n3310) );
  AND U4851 ( .A(n1018), .B(n3311), .Z(n3309) );
  XOR U4852 ( .A(DB[3]), .B(DB[10]), .Z(n3311) );
  XOR U4853 ( .A(DB[1787]), .B(n3312), .Z(min_val_out[2]) );
  AND U4854 ( .A(n2), .B(n3313), .Z(n3312) );
  XOR U4855 ( .A(n3314), .B(n3315), .Z(n3313) );
  XOR U4856 ( .A(DB[1787]), .B(DB[1780]), .Z(n3315) );
  AND U4857 ( .A(n6), .B(n3316), .Z(n3314) );
  XOR U4858 ( .A(n3317), .B(n3318), .Z(n3316) );
  XOR U4859 ( .A(DB[1780]), .B(DB[1773]), .Z(n3318) );
  AND U4860 ( .A(n10), .B(n3319), .Z(n3317) );
  XOR U4861 ( .A(n3320), .B(n3321), .Z(n3319) );
  XOR U4862 ( .A(DB[1773]), .B(DB[1766]), .Z(n3321) );
  AND U4863 ( .A(n14), .B(n3322), .Z(n3320) );
  XOR U4864 ( .A(n3323), .B(n3324), .Z(n3322) );
  XOR U4865 ( .A(DB[1766]), .B(DB[1759]), .Z(n3324) );
  AND U4866 ( .A(n18), .B(n3325), .Z(n3323) );
  XOR U4867 ( .A(n3326), .B(n3327), .Z(n3325) );
  XOR U4868 ( .A(DB[1759]), .B(DB[1752]), .Z(n3327) );
  AND U4869 ( .A(n22), .B(n3328), .Z(n3326) );
  XOR U4870 ( .A(n3329), .B(n3330), .Z(n3328) );
  XOR U4871 ( .A(DB[1752]), .B(DB[1745]), .Z(n3330) );
  AND U4872 ( .A(n26), .B(n3331), .Z(n3329) );
  XOR U4873 ( .A(n3332), .B(n3333), .Z(n3331) );
  XOR U4874 ( .A(DB[1745]), .B(DB[1738]), .Z(n3333) );
  AND U4875 ( .A(n30), .B(n3334), .Z(n3332) );
  XOR U4876 ( .A(n3335), .B(n3336), .Z(n3334) );
  XOR U4877 ( .A(DB[1738]), .B(DB[1731]), .Z(n3336) );
  AND U4878 ( .A(n34), .B(n3337), .Z(n3335) );
  XOR U4879 ( .A(n3338), .B(n3339), .Z(n3337) );
  XOR U4880 ( .A(DB[1731]), .B(DB[1724]), .Z(n3339) );
  AND U4881 ( .A(n38), .B(n3340), .Z(n3338) );
  XOR U4882 ( .A(n3341), .B(n3342), .Z(n3340) );
  XOR U4883 ( .A(DB[1724]), .B(DB[1717]), .Z(n3342) );
  AND U4884 ( .A(n42), .B(n3343), .Z(n3341) );
  XOR U4885 ( .A(n3344), .B(n3345), .Z(n3343) );
  XOR U4886 ( .A(DB[1717]), .B(DB[1710]), .Z(n3345) );
  AND U4887 ( .A(n46), .B(n3346), .Z(n3344) );
  XOR U4888 ( .A(n3347), .B(n3348), .Z(n3346) );
  XOR U4889 ( .A(DB[1710]), .B(DB[1703]), .Z(n3348) );
  AND U4890 ( .A(n50), .B(n3349), .Z(n3347) );
  XOR U4891 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR U4892 ( .A(DB[1703]), .B(DB[1696]), .Z(n3351) );
  AND U4893 ( .A(n54), .B(n3352), .Z(n3350) );
  XOR U4894 ( .A(n3353), .B(n3354), .Z(n3352) );
  XOR U4895 ( .A(DB[1696]), .B(DB[1689]), .Z(n3354) );
  AND U4896 ( .A(n58), .B(n3355), .Z(n3353) );
  XOR U4897 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR U4898 ( .A(DB[1689]), .B(DB[1682]), .Z(n3357) );
  AND U4899 ( .A(n62), .B(n3358), .Z(n3356) );
  XOR U4900 ( .A(n3359), .B(n3360), .Z(n3358) );
  XOR U4901 ( .A(DB[1682]), .B(DB[1675]), .Z(n3360) );
  AND U4902 ( .A(n66), .B(n3361), .Z(n3359) );
  XOR U4903 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR U4904 ( .A(DB[1675]), .B(DB[1668]), .Z(n3363) );
  AND U4905 ( .A(n70), .B(n3364), .Z(n3362) );
  XOR U4906 ( .A(n3365), .B(n3366), .Z(n3364) );
  XOR U4907 ( .A(DB[1668]), .B(DB[1661]), .Z(n3366) );
  AND U4908 ( .A(n74), .B(n3367), .Z(n3365) );
  XOR U4909 ( .A(n3368), .B(n3369), .Z(n3367) );
  XOR U4910 ( .A(DB[1661]), .B(DB[1654]), .Z(n3369) );
  AND U4911 ( .A(n78), .B(n3370), .Z(n3368) );
  XOR U4912 ( .A(n3371), .B(n3372), .Z(n3370) );
  XOR U4913 ( .A(DB[1654]), .B(DB[1647]), .Z(n3372) );
  AND U4914 ( .A(n82), .B(n3373), .Z(n3371) );
  XOR U4915 ( .A(n3374), .B(n3375), .Z(n3373) );
  XOR U4916 ( .A(DB[1647]), .B(DB[1640]), .Z(n3375) );
  AND U4917 ( .A(n86), .B(n3376), .Z(n3374) );
  XOR U4918 ( .A(n3377), .B(n3378), .Z(n3376) );
  XOR U4919 ( .A(DB[1640]), .B(DB[1633]), .Z(n3378) );
  AND U4920 ( .A(n90), .B(n3379), .Z(n3377) );
  XOR U4921 ( .A(n3380), .B(n3381), .Z(n3379) );
  XOR U4922 ( .A(DB[1633]), .B(DB[1626]), .Z(n3381) );
  AND U4923 ( .A(n94), .B(n3382), .Z(n3380) );
  XOR U4924 ( .A(n3383), .B(n3384), .Z(n3382) );
  XOR U4925 ( .A(DB[1626]), .B(DB[1619]), .Z(n3384) );
  AND U4926 ( .A(n98), .B(n3385), .Z(n3383) );
  XOR U4927 ( .A(n3386), .B(n3387), .Z(n3385) );
  XOR U4928 ( .A(DB[1619]), .B(DB[1612]), .Z(n3387) );
  AND U4929 ( .A(n102), .B(n3388), .Z(n3386) );
  XOR U4930 ( .A(n3389), .B(n3390), .Z(n3388) );
  XOR U4931 ( .A(DB[1612]), .B(DB[1605]), .Z(n3390) );
  AND U4932 ( .A(n106), .B(n3391), .Z(n3389) );
  XOR U4933 ( .A(n3392), .B(n3393), .Z(n3391) );
  XOR U4934 ( .A(DB[1605]), .B(DB[1598]), .Z(n3393) );
  AND U4935 ( .A(n110), .B(n3394), .Z(n3392) );
  XOR U4936 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR U4937 ( .A(DB[1598]), .B(DB[1591]), .Z(n3396) );
  AND U4938 ( .A(n114), .B(n3397), .Z(n3395) );
  XOR U4939 ( .A(n3398), .B(n3399), .Z(n3397) );
  XOR U4940 ( .A(DB[1591]), .B(DB[1584]), .Z(n3399) );
  AND U4941 ( .A(n118), .B(n3400), .Z(n3398) );
  XOR U4942 ( .A(n3401), .B(n3402), .Z(n3400) );
  XOR U4943 ( .A(DB[1584]), .B(DB[1577]), .Z(n3402) );
  AND U4944 ( .A(n122), .B(n3403), .Z(n3401) );
  XOR U4945 ( .A(n3404), .B(n3405), .Z(n3403) );
  XOR U4946 ( .A(DB[1577]), .B(DB[1570]), .Z(n3405) );
  AND U4947 ( .A(n126), .B(n3406), .Z(n3404) );
  XOR U4948 ( .A(n3407), .B(n3408), .Z(n3406) );
  XOR U4949 ( .A(DB[1570]), .B(DB[1563]), .Z(n3408) );
  AND U4950 ( .A(n130), .B(n3409), .Z(n3407) );
  XOR U4951 ( .A(n3410), .B(n3411), .Z(n3409) );
  XOR U4952 ( .A(DB[1563]), .B(DB[1556]), .Z(n3411) );
  AND U4953 ( .A(n134), .B(n3412), .Z(n3410) );
  XOR U4954 ( .A(n3413), .B(n3414), .Z(n3412) );
  XOR U4955 ( .A(DB[1556]), .B(DB[1549]), .Z(n3414) );
  AND U4956 ( .A(n138), .B(n3415), .Z(n3413) );
  XOR U4957 ( .A(n3416), .B(n3417), .Z(n3415) );
  XOR U4958 ( .A(DB[1549]), .B(DB[1542]), .Z(n3417) );
  AND U4959 ( .A(n142), .B(n3418), .Z(n3416) );
  XOR U4960 ( .A(n3419), .B(n3420), .Z(n3418) );
  XOR U4961 ( .A(DB[1542]), .B(DB[1535]), .Z(n3420) );
  AND U4962 ( .A(n146), .B(n3421), .Z(n3419) );
  XOR U4963 ( .A(n3422), .B(n3423), .Z(n3421) );
  XOR U4964 ( .A(DB[1535]), .B(DB[1528]), .Z(n3423) );
  AND U4965 ( .A(n150), .B(n3424), .Z(n3422) );
  XOR U4966 ( .A(n3425), .B(n3426), .Z(n3424) );
  XOR U4967 ( .A(DB[1528]), .B(DB[1521]), .Z(n3426) );
  AND U4968 ( .A(n154), .B(n3427), .Z(n3425) );
  XOR U4969 ( .A(n3428), .B(n3429), .Z(n3427) );
  XOR U4970 ( .A(DB[1521]), .B(DB[1514]), .Z(n3429) );
  AND U4971 ( .A(n158), .B(n3430), .Z(n3428) );
  XOR U4972 ( .A(n3431), .B(n3432), .Z(n3430) );
  XOR U4973 ( .A(DB[1514]), .B(DB[1507]), .Z(n3432) );
  AND U4974 ( .A(n162), .B(n3433), .Z(n3431) );
  XOR U4975 ( .A(n3434), .B(n3435), .Z(n3433) );
  XOR U4976 ( .A(DB[1507]), .B(DB[1500]), .Z(n3435) );
  AND U4977 ( .A(n166), .B(n3436), .Z(n3434) );
  XOR U4978 ( .A(n3437), .B(n3438), .Z(n3436) );
  XOR U4979 ( .A(DB[1500]), .B(DB[1493]), .Z(n3438) );
  AND U4980 ( .A(n170), .B(n3439), .Z(n3437) );
  XOR U4981 ( .A(n3440), .B(n3441), .Z(n3439) );
  XOR U4982 ( .A(DB[1493]), .B(DB[1486]), .Z(n3441) );
  AND U4983 ( .A(n174), .B(n3442), .Z(n3440) );
  XOR U4984 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U4985 ( .A(DB[1486]), .B(DB[1479]), .Z(n3444) );
  AND U4986 ( .A(n178), .B(n3445), .Z(n3443) );
  XOR U4987 ( .A(n3446), .B(n3447), .Z(n3445) );
  XOR U4988 ( .A(DB[1479]), .B(DB[1472]), .Z(n3447) );
  AND U4989 ( .A(n182), .B(n3448), .Z(n3446) );
  XOR U4990 ( .A(n3449), .B(n3450), .Z(n3448) );
  XOR U4991 ( .A(DB[1472]), .B(DB[1465]), .Z(n3450) );
  AND U4992 ( .A(n186), .B(n3451), .Z(n3449) );
  XOR U4993 ( .A(n3452), .B(n3453), .Z(n3451) );
  XOR U4994 ( .A(DB[1465]), .B(DB[1458]), .Z(n3453) );
  AND U4995 ( .A(n190), .B(n3454), .Z(n3452) );
  XOR U4996 ( .A(n3455), .B(n3456), .Z(n3454) );
  XOR U4997 ( .A(DB[1458]), .B(DB[1451]), .Z(n3456) );
  AND U4998 ( .A(n194), .B(n3457), .Z(n3455) );
  XOR U4999 ( .A(n3458), .B(n3459), .Z(n3457) );
  XOR U5000 ( .A(DB[1451]), .B(DB[1444]), .Z(n3459) );
  AND U5001 ( .A(n198), .B(n3460), .Z(n3458) );
  XOR U5002 ( .A(n3461), .B(n3462), .Z(n3460) );
  XOR U5003 ( .A(DB[1444]), .B(DB[1437]), .Z(n3462) );
  AND U5004 ( .A(n202), .B(n3463), .Z(n3461) );
  XOR U5005 ( .A(n3464), .B(n3465), .Z(n3463) );
  XOR U5006 ( .A(DB[1437]), .B(DB[1430]), .Z(n3465) );
  AND U5007 ( .A(n206), .B(n3466), .Z(n3464) );
  XOR U5008 ( .A(n3467), .B(n3468), .Z(n3466) );
  XOR U5009 ( .A(DB[1430]), .B(DB[1423]), .Z(n3468) );
  AND U5010 ( .A(n210), .B(n3469), .Z(n3467) );
  XOR U5011 ( .A(n3470), .B(n3471), .Z(n3469) );
  XOR U5012 ( .A(DB[1423]), .B(DB[1416]), .Z(n3471) );
  AND U5013 ( .A(n214), .B(n3472), .Z(n3470) );
  XOR U5014 ( .A(n3473), .B(n3474), .Z(n3472) );
  XOR U5015 ( .A(DB[1416]), .B(DB[1409]), .Z(n3474) );
  AND U5016 ( .A(n218), .B(n3475), .Z(n3473) );
  XOR U5017 ( .A(n3476), .B(n3477), .Z(n3475) );
  XOR U5018 ( .A(DB[1409]), .B(DB[1402]), .Z(n3477) );
  AND U5019 ( .A(n222), .B(n3478), .Z(n3476) );
  XOR U5020 ( .A(n3479), .B(n3480), .Z(n3478) );
  XOR U5021 ( .A(DB[1402]), .B(DB[1395]), .Z(n3480) );
  AND U5022 ( .A(n226), .B(n3481), .Z(n3479) );
  XOR U5023 ( .A(n3482), .B(n3483), .Z(n3481) );
  XOR U5024 ( .A(DB[1395]), .B(DB[1388]), .Z(n3483) );
  AND U5025 ( .A(n230), .B(n3484), .Z(n3482) );
  XOR U5026 ( .A(n3485), .B(n3486), .Z(n3484) );
  XOR U5027 ( .A(DB[1388]), .B(DB[1381]), .Z(n3486) );
  AND U5028 ( .A(n234), .B(n3487), .Z(n3485) );
  XOR U5029 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR U5030 ( .A(DB[1381]), .B(DB[1374]), .Z(n3489) );
  AND U5031 ( .A(n238), .B(n3490), .Z(n3488) );
  XOR U5032 ( .A(n3491), .B(n3492), .Z(n3490) );
  XOR U5033 ( .A(DB[1374]), .B(DB[1367]), .Z(n3492) );
  AND U5034 ( .A(n242), .B(n3493), .Z(n3491) );
  XOR U5035 ( .A(n3494), .B(n3495), .Z(n3493) );
  XOR U5036 ( .A(DB[1367]), .B(DB[1360]), .Z(n3495) );
  AND U5037 ( .A(n246), .B(n3496), .Z(n3494) );
  XOR U5038 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR U5039 ( .A(DB[1360]), .B(DB[1353]), .Z(n3498) );
  AND U5040 ( .A(n250), .B(n3499), .Z(n3497) );
  XOR U5041 ( .A(n3500), .B(n3501), .Z(n3499) );
  XOR U5042 ( .A(DB[1353]), .B(DB[1346]), .Z(n3501) );
  AND U5043 ( .A(n254), .B(n3502), .Z(n3500) );
  XOR U5044 ( .A(n3503), .B(n3504), .Z(n3502) );
  XOR U5045 ( .A(DB[1346]), .B(DB[1339]), .Z(n3504) );
  AND U5046 ( .A(n258), .B(n3505), .Z(n3503) );
  XOR U5047 ( .A(n3506), .B(n3507), .Z(n3505) );
  XOR U5048 ( .A(DB[1339]), .B(DB[1332]), .Z(n3507) );
  AND U5049 ( .A(n262), .B(n3508), .Z(n3506) );
  XOR U5050 ( .A(n3509), .B(n3510), .Z(n3508) );
  XOR U5051 ( .A(DB[1332]), .B(DB[1325]), .Z(n3510) );
  AND U5052 ( .A(n266), .B(n3511), .Z(n3509) );
  XOR U5053 ( .A(n3512), .B(n3513), .Z(n3511) );
  XOR U5054 ( .A(DB[1325]), .B(DB[1318]), .Z(n3513) );
  AND U5055 ( .A(n270), .B(n3514), .Z(n3512) );
  XOR U5056 ( .A(n3515), .B(n3516), .Z(n3514) );
  XOR U5057 ( .A(DB[1318]), .B(DB[1311]), .Z(n3516) );
  AND U5058 ( .A(n274), .B(n3517), .Z(n3515) );
  XOR U5059 ( .A(n3518), .B(n3519), .Z(n3517) );
  XOR U5060 ( .A(DB[1311]), .B(DB[1304]), .Z(n3519) );
  AND U5061 ( .A(n278), .B(n3520), .Z(n3518) );
  XOR U5062 ( .A(n3521), .B(n3522), .Z(n3520) );
  XOR U5063 ( .A(DB[1304]), .B(DB[1297]), .Z(n3522) );
  AND U5064 ( .A(n282), .B(n3523), .Z(n3521) );
  XOR U5065 ( .A(n3524), .B(n3525), .Z(n3523) );
  XOR U5066 ( .A(DB[1297]), .B(DB[1290]), .Z(n3525) );
  AND U5067 ( .A(n286), .B(n3526), .Z(n3524) );
  XOR U5068 ( .A(n3527), .B(n3528), .Z(n3526) );
  XOR U5069 ( .A(DB[1290]), .B(DB[1283]), .Z(n3528) );
  AND U5070 ( .A(n290), .B(n3529), .Z(n3527) );
  XOR U5071 ( .A(n3530), .B(n3531), .Z(n3529) );
  XOR U5072 ( .A(DB[1283]), .B(DB[1276]), .Z(n3531) );
  AND U5073 ( .A(n294), .B(n3532), .Z(n3530) );
  XOR U5074 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR U5075 ( .A(DB[1276]), .B(DB[1269]), .Z(n3534) );
  AND U5076 ( .A(n298), .B(n3535), .Z(n3533) );
  XOR U5077 ( .A(n3536), .B(n3537), .Z(n3535) );
  XOR U5078 ( .A(DB[1269]), .B(DB[1262]), .Z(n3537) );
  AND U5079 ( .A(n302), .B(n3538), .Z(n3536) );
  XOR U5080 ( .A(n3539), .B(n3540), .Z(n3538) );
  XOR U5081 ( .A(DB[1262]), .B(DB[1255]), .Z(n3540) );
  AND U5082 ( .A(n306), .B(n3541), .Z(n3539) );
  XOR U5083 ( .A(n3542), .B(n3543), .Z(n3541) );
  XOR U5084 ( .A(DB[1255]), .B(DB[1248]), .Z(n3543) );
  AND U5085 ( .A(n310), .B(n3544), .Z(n3542) );
  XOR U5086 ( .A(n3545), .B(n3546), .Z(n3544) );
  XOR U5087 ( .A(DB[1248]), .B(DB[1241]), .Z(n3546) );
  AND U5088 ( .A(n314), .B(n3547), .Z(n3545) );
  XOR U5089 ( .A(n3548), .B(n3549), .Z(n3547) );
  XOR U5090 ( .A(DB[1241]), .B(DB[1234]), .Z(n3549) );
  AND U5091 ( .A(n318), .B(n3550), .Z(n3548) );
  XOR U5092 ( .A(n3551), .B(n3552), .Z(n3550) );
  XOR U5093 ( .A(DB[1234]), .B(DB[1227]), .Z(n3552) );
  AND U5094 ( .A(n322), .B(n3553), .Z(n3551) );
  XOR U5095 ( .A(n3554), .B(n3555), .Z(n3553) );
  XOR U5096 ( .A(DB[1227]), .B(DB[1220]), .Z(n3555) );
  AND U5097 ( .A(n326), .B(n3556), .Z(n3554) );
  XOR U5098 ( .A(n3557), .B(n3558), .Z(n3556) );
  XOR U5099 ( .A(DB[1220]), .B(DB[1213]), .Z(n3558) );
  AND U5100 ( .A(n330), .B(n3559), .Z(n3557) );
  XOR U5101 ( .A(n3560), .B(n3561), .Z(n3559) );
  XOR U5102 ( .A(DB[1213]), .B(DB[1206]), .Z(n3561) );
  AND U5103 ( .A(n334), .B(n3562), .Z(n3560) );
  XOR U5104 ( .A(n3563), .B(n3564), .Z(n3562) );
  XOR U5105 ( .A(DB[1206]), .B(DB[1199]), .Z(n3564) );
  AND U5106 ( .A(n338), .B(n3565), .Z(n3563) );
  XOR U5107 ( .A(n3566), .B(n3567), .Z(n3565) );
  XOR U5108 ( .A(DB[1199]), .B(DB[1192]), .Z(n3567) );
  AND U5109 ( .A(n342), .B(n3568), .Z(n3566) );
  XOR U5110 ( .A(n3569), .B(n3570), .Z(n3568) );
  XOR U5111 ( .A(DB[1192]), .B(DB[1185]), .Z(n3570) );
  AND U5112 ( .A(n346), .B(n3571), .Z(n3569) );
  XOR U5113 ( .A(n3572), .B(n3573), .Z(n3571) );
  XOR U5114 ( .A(DB[1185]), .B(DB[1178]), .Z(n3573) );
  AND U5115 ( .A(n350), .B(n3574), .Z(n3572) );
  XOR U5116 ( .A(n3575), .B(n3576), .Z(n3574) );
  XOR U5117 ( .A(DB[1178]), .B(DB[1171]), .Z(n3576) );
  AND U5118 ( .A(n354), .B(n3577), .Z(n3575) );
  XOR U5119 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U5120 ( .A(DB[1171]), .B(DB[1164]), .Z(n3579) );
  AND U5121 ( .A(n358), .B(n3580), .Z(n3578) );
  XOR U5122 ( .A(n3581), .B(n3582), .Z(n3580) );
  XOR U5123 ( .A(DB[1164]), .B(DB[1157]), .Z(n3582) );
  AND U5124 ( .A(n362), .B(n3583), .Z(n3581) );
  XOR U5125 ( .A(n3584), .B(n3585), .Z(n3583) );
  XOR U5126 ( .A(DB[1157]), .B(DB[1150]), .Z(n3585) );
  AND U5127 ( .A(n366), .B(n3586), .Z(n3584) );
  XOR U5128 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR U5129 ( .A(DB[1150]), .B(DB[1143]), .Z(n3588) );
  AND U5130 ( .A(n370), .B(n3589), .Z(n3587) );
  XOR U5131 ( .A(n3590), .B(n3591), .Z(n3589) );
  XOR U5132 ( .A(DB[1143]), .B(DB[1136]), .Z(n3591) );
  AND U5133 ( .A(n374), .B(n3592), .Z(n3590) );
  XOR U5134 ( .A(n3593), .B(n3594), .Z(n3592) );
  XOR U5135 ( .A(DB[1136]), .B(DB[1129]), .Z(n3594) );
  AND U5136 ( .A(n378), .B(n3595), .Z(n3593) );
  XOR U5137 ( .A(n3596), .B(n3597), .Z(n3595) );
  XOR U5138 ( .A(DB[1129]), .B(DB[1122]), .Z(n3597) );
  AND U5139 ( .A(n382), .B(n3598), .Z(n3596) );
  XOR U5140 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR U5141 ( .A(DB[1122]), .B(DB[1115]), .Z(n3600) );
  AND U5142 ( .A(n386), .B(n3601), .Z(n3599) );
  XOR U5143 ( .A(n3602), .B(n3603), .Z(n3601) );
  XOR U5144 ( .A(DB[1115]), .B(DB[1108]), .Z(n3603) );
  AND U5145 ( .A(n390), .B(n3604), .Z(n3602) );
  XOR U5146 ( .A(n3605), .B(n3606), .Z(n3604) );
  XOR U5147 ( .A(DB[1108]), .B(DB[1101]), .Z(n3606) );
  AND U5148 ( .A(n394), .B(n3607), .Z(n3605) );
  XOR U5149 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U5150 ( .A(DB[1101]), .B(DB[1094]), .Z(n3609) );
  AND U5151 ( .A(n398), .B(n3610), .Z(n3608) );
  XOR U5152 ( .A(n3611), .B(n3612), .Z(n3610) );
  XOR U5153 ( .A(DB[1094]), .B(DB[1087]), .Z(n3612) );
  AND U5154 ( .A(n402), .B(n3613), .Z(n3611) );
  XOR U5155 ( .A(n3614), .B(n3615), .Z(n3613) );
  XOR U5156 ( .A(DB[1087]), .B(DB[1080]), .Z(n3615) );
  AND U5157 ( .A(n406), .B(n3616), .Z(n3614) );
  XOR U5158 ( .A(n3617), .B(n3618), .Z(n3616) );
  XOR U5159 ( .A(DB[1080]), .B(DB[1073]), .Z(n3618) );
  AND U5160 ( .A(n410), .B(n3619), .Z(n3617) );
  XOR U5161 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U5162 ( .A(DB[1073]), .B(DB[1066]), .Z(n3621) );
  AND U5163 ( .A(n414), .B(n3622), .Z(n3620) );
  XOR U5164 ( .A(n3623), .B(n3624), .Z(n3622) );
  XOR U5165 ( .A(DB[1066]), .B(DB[1059]), .Z(n3624) );
  AND U5166 ( .A(n418), .B(n3625), .Z(n3623) );
  XOR U5167 ( .A(n3626), .B(n3627), .Z(n3625) );
  XOR U5168 ( .A(DB[1059]), .B(DB[1052]), .Z(n3627) );
  AND U5169 ( .A(n422), .B(n3628), .Z(n3626) );
  XOR U5170 ( .A(n3629), .B(n3630), .Z(n3628) );
  XOR U5171 ( .A(DB[1052]), .B(DB[1045]), .Z(n3630) );
  AND U5172 ( .A(n426), .B(n3631), .Z(n3629) );
  XOR U5173 ( .A(n3632), .B(n3633), .Z(n3631) );
  XOR U5174 ( .A(DB[1045]), .B(DB[1038]), .Z(n3633) );
  AND U5175 ( .A(n430), .B(n3634), .Z(n3632) );
  XOR U5176 ( .A(n3635), .B(n3636), .Z(n3634) );
  XOR U5177 ( .A(DB[1038]), .B(DB[1031]), .Z(n3636) );
  AND U5178 ( .A(n434), .B(n3637), .Z(n3635) );
  XOR U5179 ( .A(n3638), .B(n3639), .Z(n3637) );
  XOR U5180 ( .A(DB[1031]), .B(DB[1024]), .Z(n3639) );
  AND U5181 ( .A(n438), .B(n3640), .Z(n3638) );
  XOR U5182 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U5183 ( .A(DB[1024]), .B(DB[1017]), .Z(n3642) );
  AND U5184 ( .A(n442), .B(n3643), .Z(n3641) );
  XOR U5185 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U5186 ( .A(DB[1017]), .B(DB[1010]), .Z(n3645) );
  AND U5187 ( .A(n446), .B(n3646), .Z(n3644) );
  XOR U5188 ( .A(n3647), .B(n3648), .Z(n3646) );
  XOR U5189 ( .A(DB[1010]), .B(DB[1003]), .Z(n3648) );
  AND U5190 ( .A(n450), .B(n3649), .Z(n3647) );
  XOR U5191 ( .A(n3650), .B(n3651), .Z(n3649) );
  XOR U5192 ( .A(DB[996]), .B(DB[1003]), .Z(n3651) );
  AND U5193 ( .A(n454), .B(n3652), .Z(n3650) );
  XOR U5194 ( .A(n3653), .B(n3654), .Z(n3652) );
  XOR U5195 ( .A(DB[996]), .B(DB[989]), .Z(n3654) );
  AND U5196 ( .A(n458), .B(n3655), .Z(n3653) );
  XOR U5197 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR U5198 ( .A(DB[989]), .B(DB[982]), .Z(n3657) );
  AND U5199 ( .A(n462), .B(n3658), .Z(n3656) );
  XOR U5200 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U5201 ( .A(DB[982]), .B(DB[975]), .Z(n3660) );
  AND U5202 ( .A(n466), .B(n3661), .Z(n3659) );
  XOR U5203 ( .A(n3662), .B(n3663), .Z(n3661) );
  XOR U5204 ( .A(DB[975]), .B(DB[968]), .Z(n3663) );
  AND U5205 ( .A(n470), .B(n3664), .Z(n3662) );
  XOR U5206 ( .A(n3665), .B(n3666), .Z(n3664) );
  XOR U5207 ( .A(DB[968]), .B(DB[961]), .Z(n3666) );
  AND U5208 ( .A(n474), .B(n3667), .Z(n3665) );
  XOR U5209 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U5210 ( .A(DB[961]), .B(DB[954]), .Z(n3669) );
  AND U5211 ( .A(n478), .B(n3670), .Z(n3668) );
  XOR U5212 ( .A(n3671), .B(n3672), .Z(n3670) );
  XOR U5213 ( .A(DB[954]), .B(DB[947]), .Z(n3672) );
  AND U5214 ( .A(n482), .B(n3673), .Z(n3671) );
  XOR U5215 ( .A(n3674), .B(n3675), .Z(n3673) );
  XOR U5216 ( .A(DB[947]), .B(DB[940]), .Z(n3675) );
  AND U5217 ( .A(n486), .B(n3676), .Z(n3674) );
  XOR U5218 ( .A(n3677), .B(n3678), .Z(n3676) );
  XOR U5219 ( .A(DB[940]), .B(DB[933]), .Z(n3678) );
  AND U5220 ( .A(n490), .B(n3679), .Z(n3677) );
  XOR U5221 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR U5222 ( .A(DB[933]), .B(DB[926]), .Z(n3681) );
  AND U5223 ( .A(n494), .B(n3682), .Z(n3680) );
  XOR U5224 ( .A(n3683), .B(n3684), .Z(n3682) );
  XOR U5225 ( .A(DB[926]), .B(DB[919]), .Z(n3684) );
  AND U5226 ( .A(n498), .B(n3685), .Z(n3683) );
  XOR U5227 ( .A(n3686), .B(n3687), .Z(n3685) );
  XOR U5228 ( .A(DB[919]), .B(DB[912]), .Z(n3687) );
  AND U5229 ( .A(n502), .B(n3688), .Z(n3686) );
  XOR U5230 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U5231 ( .A(DB[912]), .B(DB[905]), .Z(n3690) );
  AND U5232 ( .A(n506), .B(n3691), .Z(n3689) );
  XOR U5233 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR U5234 ( .A(DB[905]), .B(DB[898]), .Z(n3693) );
  AND U5235 ( .A(n510), .B(n3694), .Z(n3692) );
  XOR U5236 ( .A(n3695), .B(n3696), .Z(n3694) );
  XOR U5237 ( .A(DB[898]), .B(DB[891]), .Z(n3696) );
  AND U5238 ( .A(n514), .B(n3697), .Z(n3695) );
  XOR U5239 ( .A(n3698), .B(n3699), .Z(n3697) );
  XOR U5240 ( .A(DB[891]), .B(DB[884]), .Z(n3699) );
  AND U5241 ( .A(n518), .B(n3700), .Z(n3698) );
  XOR U5242 ( .A(n3701), .B(n3702), .Z(n3700) );
  XOR U5243 ( .A(DB[884]), .B(DB[877]), .Z(n3702) );
  AND U5244 ( .A(n522), .B(n3703), .Z(n3701) );
  XOR U5245 ( .A(n3704), .B(n3705), .Z(n3703) );
  XOR U5246 ( .A(DB[877]), .B(DB[870]), .Z(n3705) );
  AND U5247 ( .A(n526), .B(n3706), .Z(n3704) );
  XOR U5248 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U5249 ( .A(DB[870]), .B(DB[863]), .Z(n3708) );
  AND U5250 ( .A(n530), .B(n3709), .Z(n3707) );
  XOR U5251 ( .A(n3710), .B(n3711), .Z(n3709) );
  XOR U5252 ( .A(DB[863]), .B(DB[856]), .Z(n3711) );
  AND U5253 ( .A(n534), .B(n3712), .Z(n3710) );
  XOR U5254 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U5255 ( .A(DB[856]), .B(DB[849]), .Z(n3714) );
  AND U5256 ( .A(n538), .B(n3715), .Z(n3713) );
  XOR U5257 ( .A(n3716), .B(n3717), .Z(n3715) );
  XOR U5258 ( .A(DB[849]), .B(DB[842]), .Z(n3717) );
  AND U5259 ( .A(n542), .B(n3718), .Z(n3716) );
  XOR U5260 ( .A(n3719), .B(n3720), .Z(n3718) );
  XOR U5261 ( .A(DB[842]), .B(DB[835]), .Z(n3720) );
  AND U5262 ( .A(n546), .B(n3721), .Z(n3719) );
  XOR U5263 ( .A(n3722), .B(n3723), .Z(n3721) );
  XOR U5264 ( .A(DB[835]), .B(DB[828]), .Z(n3723) );
  AND U5265 ( .A(n550), .B(n3724), .Z(n3722) );
  XOR U5266 ( .A(n3725), .B(n3726), .Z(n3724) );
  XOR U5267 ( .A(DB[828]), .B(DB[821]), .Z(n3726) );
  AND U5268 ( .A(n554), .B(n3727), .Z(n3725) );
  XOR U5269 ( .A(n3728), .B(n3729), .Z(n3727) );
  XOR U5270 ( .A(DB[821]), .B(DB[814]), .Z(n3729) );
  AND U5271 ( .A(n558), .B(n3730), .Z(n3728) );
  XOR U5272 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR U5273 ( .A(DB[814]), .B(DB[807]), .Z(n3732) );
  AND U5274 ( .A(n562), .B(n3733), .Z(n3731) );
  XOR U5275 ( .A(n3734), .B(n3735), .Z(n3733) );
  XOR U5276 ( .A(DB[807]), .B(DB[800]), .Z(n3735) );
  AND U5277 ( .A(n566), .B(n3736), .Z(n3734) );
  XOR U5278 ( .A(n3737), .B(n3738), .Z(n3736) );
  XOR U5279 ( .A(DB[800]), .B(DB[793]), .Z(n3738) );
  AND U5280 ( .A(n570), .B(n3739), .Z(n3737) );
  XOR U5281 ( .A(n3740), .B(n3741), .Z(n3739) );
  XOR U5282 ( .A(DB[793]), .B(DB[786]), .Z(n3741) );
  AND U5283 ( .A(n574), .B(n3742), .Z(n3740) );
  XOR U5284 ( .A(n3743), .B(n3744), .Z(n3742) );
  XOR U5285 ( .A(DB[786]), .B(DB[779]), .Z(n3744) );
  AND U5286 ( .A(n578), .B(n3745), .Z(n3743) );
  XOR U5287 ( .A(n3746), .B(n3747), .Z(n3745) );
  XOR U5288 ( .A(DB[779]), .B(DB[772]), .Z(n3747) );
  AND U5289 ( .A(n582), .B(n3748), .Z(n3746) );
  XOR U5290 ( .A(n3749), .B(n3750), .Z(n3748) );
  XOR U5291 ( .A(DB[772]), .B(DB[765]), .Z(n3750) );
  AND U5292 ( .A(n586), .B(n3751), .Z(n3749) );
  XOR U5293 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U5294 ( .A(DB[765]), .B(DB[758]), .Z(n3753) );
  AND U5295 ( .A(n590), .B(n3754), .Z(n3752) );
  XOR U5296 ( .A(n3755), .B(n3756), .Z(n3754) );
  XOR U5297 ( .A(DB[758]), .B(DB[751]), .Z(n3756) );
  AND U5298 ( .A(n594), .B(n3757), .Z(n3755) );
  XOR U5299 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR U5300 ( .A(DB[751]), .B(DB[744]), .Z(n3759) );
  AND U5301 ( .A(n598), .B(n3760), .Z(n3758) );
  XOR U5302 ( .A(n3761), .B(n3762), .Z(n3760) );
  XOR U5303 ( .A(DB[744]), .B(DB[737]), .Z(n3762) );
  AND U5304 ( .A(n602), .B(n3763), .Z(n3761) );
  XOR U5305 ( .A(n3764), .B(n3765), .Z(n3763) );
  XOR U5306 ( .A(DB[737]), .B(DB[730]), .Z(n3765) );
  AND U5307 ( .A(n606), .B(n3766), .Z(n3764) );
  XOR U5308 ( .A(n3767), .B(n3768), .Z(n3766) );
  XOR U5309 ( .A(DB[730]), .B(DB[723]), .Z(n3768) );
  AND U5310 ( .A(n610), .B(n3769), .Z(n3767) );
  XOR U5311 ( .A(n3770), .B(n3771), .Z(n3769) );
  XOR U5312 ( .A(DB[723]), .B(DB[716]), .Z(n3771) );
  AND U5313 ( .A(n614), .B(n3772), .Z(n3770) );
  XOR U5314 ( .A(n3773), .B(n3774), .Z(n3772) );
  XOR U5315 ( .A(DB[716]), .B(DB[709]), .Z(n3774) );
  AND U5316 ( .A(n618), .B(n3775), .Z(n3773) );
  XOR U5317 ( .A(n3776), .B(n3777), .Z(n3775) );
  XOR U5318 ( .A(DB[709]), .B(DB[702]), .Z(n3777) );
  AND U5319 ( .A(n622), .B(n3778), .Z(n3776) );
  XOR U5320 ( .A(n3779), .B(n3780), .Z(n3778) );
  XOR U5321 ( .A(DB[702]), .B(DB[695]), .Z(n3780) );
  AND U5322 ( .A(n626), .B(n3781), .Z(n3779) );
  XOR U5323 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U5324 ( .A(DB[695]), .B(DB[688]), .Z(n3783) );
  AND U5325 ( .A(n630), .B(n3784), .Z(n3782) );
  XOR U5326 ( .A(n3785), .B(n3786), .Z(n3784) );
  XOR U5327 ( .A(DB[688]), .B(DB[681]), .Z(n3786) );
  AND U5328 ( .A(n634), .B(n3787), .Z(n3785) );
  XOR U5329 ( .A(n3788), .B(n3789), .Z(n3787) );
  XOR U5330 ( .A(DB[681]), .B(DB[674]), .Z(n3789) );
  AND U5331 ( .A(n638), .B(n3790), .Z(n3788) );
  XOR U5332 ( .A(n3791), .B(n3792), .Z(n3790) );
  XOR U5333 ( .A(DB[674]), .B(DB[667]), .Z(n3792) );
  AND U5334 ( .A(n642), .B(n3793), .Z(n3791) );
  XOR U5335 ( .A(n3794), .B(n3795), .Z(n3793) );
  XOR U5336 ( .A(DB[667]), .B(DB[660]), .Z(n3795) );
  AND U5337 ( .A(n646), .B(n3796), .Z(n3794) );
  XOR U5338 ( .A(n3797), .B(n3798), .Z(n3796) );
  XOR U5339 ( .A(DB[660]), .B(DB[653]), .Z(n3798) );
  AND U5340 ( .A(n650), .B(n3799), .Z(n3797) );
  XOR U5341 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U5342 ( .A(DB[653]), .B(DB[646]), .Z(n3801) );
  AND U5343 ( .A(n654), .B(n3802), .Z(n3800) );
  XOR U5344 ( .A(n3803), .B(n3804), .Z(n3802) );
  XOR U5345 ( .A(DB[646]), .B(DB[639]), .Z(n3804) );
  AND U5346 ( .A(n658), .B(n3805), .Z(n3803) );
  XOR U5347 ( .A(n3806), .B(n3807), .Z(n3805) );
  XOR U5348 ( .A(DB[639]), .B(DB[632]), .Z(n3807) );
  AND U5349 ( .A(n662), .B(n3808), .Z(n3806) );
  XOR U5350 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U5351 ( .A(DB[632]), .B(DB[625]), .Z(n3810) );
  AND U5352 ( .A(n666), .B(n3811), .Z(n3809) );
  XOR U5353 ( .A(n3812), .B(n3813), .Z(n3811) );
  XOR U5354 ( .A(DB[625]), .B(DB[618]), .Z(n3813) );
  AND U5355 ( .A(n670), .B(n3814), .Z(n3812) );
  XOR U5356 ( .A(n3815), .B(n3816), .Z(n3814) );
  XOR U5357 ( .A(DB[618]), .B(DB[611]), .Z(n3816) );
  AND U5358 ( .A(n674), .B(n3817), .Z(n3815) );
  XOR U5359 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR U5360 ( .A(DB[611]), .B(DB[604]), .Z(n3819) );
  AND U5361 ( .A(n678), .B(n3820), .Z(n3818) );
  XOR U5362 ( .A(n3821), .B(n3822), .Z(n3820) );
  XOR U5363 ( .A(DB[604]), .B(DB[597]), .Z(n3822) );
  AND U5364 ( .A(n682), .B(n3823), .Z(n3821) );
  XOR U5365 ( .A(n3824), .B(n3825), .Z(n3823) );
  XOR U5366 ( .A(DB[597]), .B(DB[590]), .Z(n3825) );
  AND U5367 ( .A(n686), .B(n3826), .Z(n3824) );
  XOR U5368 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR U5369 ( .A(DB[590]), .B(DB[583]), .Z(n3828) );
  AND U5370 ( .A(n690), .B(n3829), .Z(n3827) );
  XOR U5371 ( .A(n3830), .B(n3831), .Z(n3829) );
  XOR U5372 ( .A(DB[583]), .B(DB[576]), .Z(n3831) );
  AND U5373 ( .A(n694), .B(n3832), .Z(n3830) );
  XOR U5374 ( .A(n3833), .B(n3834), .Z(n3832) );
  XOR U5375 ( .A(DB[576]), .B(DB[569]), .Z(n3834) );
  AND U5376 ( .A(n698), .B(n3835), .Z(n3833) );
  XOR U5377 ( .A(n3836), .B(n3837), .Z(n3835) );
  XOR U5378 ( .A(DB[569]), .B(DB[562]), .Z(n3837) );
  AND U5379 ( .A(n702), .B(n3838), .Z(n3836) );
  XOR U5380 ( .A(n3839), .B(n3840), .Z(n3838) );
  XOR U5381 ( .A(DB[562]), .B(DB[555]), .Z(n3840) );
  AND U5382 ( .A(n706), .B(n3841), .Z(n3839) );
  XOR U5383 ( .A(n3842), .B(n3843), .Z(n3841) );
  XOR U5384 ( .A(DB[555]), .B(DB[548]), .Z(n3843) );
  AND U5385 ( .A(n710), .B(n3844), .Z(n3842) );
  XOR U5386 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U5387 ( .A(DB[548]), .B(DB[541]), .Z(n3846) );
  AND U5388 ( .A(n714), .B(n3847), .Z(n3845) );
  XOR U5389 ( .A(n3848), .B(n3849), .Z(n3847) );
  XOR U5390 ( .A(DB[541]), .B(DB[534]), .Z(n3849) );
  AND U5391 ( .A(n718), .B(n3850), .Z(n3848) );
  XOR U5392 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR U5393 ( .A(DB[534]), .B(DB[527]), .Z(n3852) );
  AND U5394 ( .A(n722), .B(n3853), .Z(n3851) );
  XOR U5395 ( .A(n3854), .B(n3855), .Z(n3853) );
  XOR U5396 ( .A(DB[527]), .B(DB[520]), .Z(n3855) );
  AND U5397 ( .A(n726), .B(n3856), .Z(n3854) );
  XOR U5398 ( .A(n3857), .B(n3858), .Z(n3856) );
  XOR U5399 ( .A(DB[520]), .B(DB[513]), .Z(n3858) );
  AND U5400 ( .A(n730), .B(n3859), .Z(n3857) );
  XOR U5401 ( .A(n3860), .B(n3861), .Z(n3859) );
  XOR U5402 ( .A(DB[513]), .B(DB[506]), .Z(n3861) );
  AND U5403 ( .A(n734), .B(n3862), .Z(n3860) );
  XOR U5404 ( .A(n3863), .B(n3864), .Z(n3862) );
  XOR U5405 ( .A(DB[506]), .B(DB[499]), .Z(n3864) );
  AND U5406 ( .A(n738), .B(n3865), .Z(n3863) );
  XOR U5407 ( .A(n3866), .B(n3867), .Z(n3865) );
  XOR U5408 ( .A(DB[499]), .B(DB[492]), .Z(n3867) );
  AND U5409 ( .A(n742), .B(n3868), .Z(n3866) );
  XOR U5410 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U5411 ( .A(DB[492]), .B(DB[485]), .Z(n3870) );
  AND U5412 ( .A(n746), .B(n3871), .Z(n3869) );
  XOR U5413 ( .A(n3872), .B(n3873), .Z(n3871) );
  XOR U5414 ( .A(DB[485]), .B(DB[478]), .Z(n3873) );
  AND U5415 ( .A(n750), .B(n3874), .Z(n3872) );
  XOR U5416 ( .A(n3875), .B(n3876), .Z(n3874) );
  XOR U5417 ( .A(DB[478]), .B(DB[471]), .Z(n3876) );
  AND U5418 ( .A(n754), .B(n3877), .Z(n3875) );
  XOR U5419 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR U5420 ( .A(DB[471]), .B(DB[464]), .Z(n3879) );
  AND U5421 ( .A(n758), .B(n3880), .Z(n3878) );
  XOR U5422 ( .A(n3881), .B(n3882), .Z(n3880) );
  XOR U5423 ( .A(DB[464]), .B(DB[457]), .Z(n3882) );
  AND U5424 ( .A(n762), .B(n3883), .Z(n3881) );
  XOR U5425 ( .A(n3884), .B(n3885), .Z(n3883) );
  XOR U5426 ( .A(DB[457]), .B(DB[450]), .Z(n3885) );
  AND U5427 ( .A(n766), .B(n3886), .Z(n3884) );
  XOR U5428 ( .A(n3887), .B(n3888), .Z(n3886) );
  XOR U5429 ( .A(DB[450]), .B(DB[443]), .Z(n3888) );
  AND U5430 ( .A(n770), .B(n3889), .Z(n3887) );
  XOR U5431 ( .A(n3890), .B(n3891), .Z(n3889) );
  XOR U5432 ( .A(DB[443]), .B(DB[436]), .Z(n3891) );
  AND U5433 ( .A(n774), .B(n3892), .Z(n3890) );
  XOR U5434 ( .A(n3893), .B(n3894), .Z(n3892) );
  XOR U5435 ( .A(DB[436]), .B(DB[429]), .Z(n3894) );
  AND U5436 ( .A(n778), .B(n3895), .Z(n3893) );
  XOR U5437 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR U5438 ( .A(DB[429]), .B(DB[422]), .Z(n3897) );
  AND U5439 ( .A(n782), .B(n3898), .Z(n3896) );
  XOR U5440 ( .A(n3899), .B(n3900), .Z(n3898) );
  XOR U5441 ( .A(DB[422]), .B(DB[415]), .Z(n3900) );
  AND U5442 ( .A(n786), .B(n3901), .Z(n3899) );
  XOR U5443 ( .A(n3902), .B(n3903), .Z(n3901) );
  XOR U5444 ( .A(DB[415]), .B(DB[408]), .Z(n3903) );
  AND U5445 ( .A(n790), .B(n3904), .Z(n3902) );
  XOR U5446 ( .A(n3905), .B(n3906), .Z(n3904) );
  XOR U5447 ( .A(DB[408]), .B(DB[401]), .Z(n3906) );
  AND U5448 ( .A(n794), .B(n3907), .Z(n3905) );
  XOR U5449 ( .A(n3908), .B(n3909), .Z(n3907) );
  XOR U5450 ( .A(DB[401]), .B(DB[394]), .Z(n3909) );
  AND U5451 ( .A(n798), .B(n3910), .Z(n3908) );
  XOR U5452 ( .A(n3911), .B(n3912), .Z(n3910) );
  XOR U5453 ( .A(DB[394]), .B(DB[387]), .Z(n3912) );
  AND U5454 ( .A(n802), .B(n3913), .Z(n3911) );
  XOR U5455 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U5456 ( .A(DB[387]), .B(DB[380]), .Z(n3915) );
  AND U5457 ( .A(n806), .B(n3916), .Z(n3914) );
  XOR U5458 ( .A(n3917), .B(n3918), .Z(n3916) );
  XOR U5459 ( .A(DB[380]), .B(DB[373]), .Z(n3918) );
  AND U5460 ( .A(n810), .B(n3919), .Z(n3917) );
  XOR U5461 ( .A(n3920), .B(n3921), .Z(n3919) );
  XOR U5462 ( .A(DB[373]), .B(DB[366]), .Z(n3921) );
  AND U5463 ( .A(n814), .B(n3922), .Z(n3920) );
  XOR U5464 ( .A(n3923), .B(n3924), .Z(n3922) );
  XOR U5465 ( .A(DB[366]), .B(DB[359]), .Z(n3924) );
  AND U5466 ( .A(n818), .B(n3925), .Z(n3923) );
  XOR U5467 ( .A(n3926), .B(n3927), .Z(n3925) );
  XOR U5468 ( .A(DB[359]), .B(DB[352]), .Z(n3927) );
  AND U5469 ( .A(n822), .B(n3928), .Z(n3926) );
  XOR U5470 ( .A(n3929), .B(n3930), .Z(n3928) );
  XOR U5471 ( .A(DB[352]), .B(DB[345]), .Z(n3930) );
  AND U5472 ( .A(n826), .B(n3931), .Z(n3929) );
  XOR U5473 ( .A(n3932), .B(n3933), .Z(n3931) );
  XOR U5474 ( .A(DB[345]), .B(DB[338]), .Z(n3933) );
  AND U5475 ( .A(n830), .B(n3934), .Z(n3932) );
  XOR U5476 ( .A(n3935), .B(n3936), .Z(n3934) );
  XOR U5477 ( .A(DB[338]), .B(DB[331]), .Z(n3936) );
  AND U5478 ( .A(n834), .B(n3937), .Z(n3935) );
  XOR U5479 ( .A(n3938), .B(n3939), .Z(n3937) );
  XOR U5480 ( .A(DB[331]), .B(DB[324]), .Z(n3939) );
  AND U5481 ( .A(n838), .B(n3940), .Z(n3938) );
  XOR U5482 ( .A(n3941), .B(n3942), .Z(n3940) );
  XOR U5483 ( .A(DB[324]), .B(DB[317]), .Z(n3942) );
  AND U5484 ( .A(n842), .B(n3943), .Z(n3941) );
  XOR U5485 ( .A(n3944), .B(n3945), .Z(n3943) );
  XOR U5486 ( .A(DB[317]), .B(DB[310]), .Z(n3945) );
  AND U5487 ( .A(n846), .B(n3946), .Z(n3944) );
  XOR U5488 ( .A(n3947), .B(n3948), .Z(n3946) );
  XOR U5489 ( .A(DB[310]), .B(DB[303]), .Z(n3948) );
  AND U5490 ( .A(n850), .B(n3949), .Z(n3947) );
  XOR U5491 ( .A(n3950), .B(n3951), .Z(n3949) );
  XOR U5492 ( .A(DB[303]), .B(DB[296]), .Z(n3951) );
  AND U5493 ( .A(n854), .B(n3952), .Z(n3950) );
  XOR U5494 ( .A(n3953), .B(n3954), .Z(n3952) );
  XOR U5495 ( .A(DB[296]), .B(DB[289]), .Z(n3954) );
  AND U5496 ( .A(n858), .B(n3955), .Z(n3953) );
  XOR U5497 ( .A(n3956), .B(n3957), .Z(n3955) );
  XOR U5498 ( .A(DB[289]), .B(DB[282]), .Z(n3957) );
  AND U5499 ( .A(n862), .B(n3958), .Z(n3956) );
  XOR U5500 ( .A(n3959), .B(n3960), .Z(n3958) );
  XOR U5501 ( .A(DB[282]), .B(DB[275]), .Z(n3960) );
  AND U5502 ( .A(n866), .B(n3961), .Z(n3959) );
  XOR U5503 ( .A(n3962), .B(n3963), .Z(n3961) );
  XOR U5504 ( .A(DB[275]), .B(DB[268]), .Z(n3963) );
  AND U5505 ( .A(n870), .B(n3964), .Z(n3962) );
  XOR U5506 ( .A(n3965), .B(n3966), .Z(n3964) );
  XOR U5507 ( .A(DB[268]), .B(DB[261]), .Z(n3966) );
  AND U5508 ( .A(n874), .B(n3967), .Z(n3965) );
  XOR U5509 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U5510 ( .A(DB[261]), .B(DB[254]), .Z(n3969) );
  AND U5511 ( .A(n878), .B(n3970), .Z(n3968) );
  XOR U5512 ( .A(n3971), .B(n3972), .Z(n3970) );
  XOR U5513 ( .A(DB[254]), .B(DB[247]), .Z(n3972) );
  AND U5514 ( .A(n882), .B(n3973), .Z(n3971) );
  XOR U5515 ( .A(n3974), .B(n3975), .Z(n3973) );
  XOR U5516 ( .A(DB[247]), .B(DB[240]), .Z(n3975) );
  AND U5517 ( .A(n886), .B(n3976), .Z(n3974) );
  XOR U5518 ( .A(n3977), .B(n3978), .Z(n3976) );
  XOR U5519 ( .A(DB[240]), .B(DB[233]), .Z(n3978) );
  AND U5520 ( .A(n890), .B(n3979), .Z(n3977) );
  XOR U5521 ( .A(n3980), .B(n3981), .Z(n3979) );
  XOR U5522 ( .A(DB[233]), .B(DB[226]), .Z(n3981) );
  AND U5523 ( .A(n894), .B(n3982), .Z(n3980) );
  XOR U5524 ( .A(n3983), .B(n3984), .Z(n3982) );
  XOR U5525 ( .A(DB[226]), .B(DB[219]), .Z(n3984) );
  AND U5526 ( .A(n898), .B(n3985), .Z(n3983) );
  XOR U5527 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U5528 ( .A(DB[219]), .B(DB[212]), .Z(n3987) );
  AND U5529 ( .A(n902), .B(n3988), .Z(n3986) );
  XOR U5530 ( .A(n3989), .B(n3990), .Z(n3988) );
  XOR U5531 ( .A(DB[212]), .B(DB[205]), .Z(n3990) );
  AND U5532 ( .A(n906), .B(n3991), .Z(n3989) );
  XOR U5533 ( .A(n3992), .B(n3993), .Z(n3991) );
  XOR U5534 ( .A(DB[205]), .B(DB[198]), .Z(n3993) );
  AND U5535 ( .A(n910), .B(n3994), .Z(n3992) );
  XOR U5536 ( .A(n3995), .B(n3996), .Z(n3994) );
  XOR U5537 ( .A(DB[198]), .B(DB[191]), .Z(n3996) );
  AND U5538 ( .A(n914), .B(n3997), .Z(n3995) );
  XOR U5539 ( .A(n3998), .B(n3999), .Z(n3997) );
  XOR U5540 ( .A(DB[191]), .B(DB[184]), .Z(n3999) );
  AND U5541 ( .A(n918), .B(n4000), .Z(n3998) );
  XOR U5542 ( .A(n4001), .B(n4002), .Z(n4000) );
  XOR U5543 ( .A(DB[184]), .B(DB[177]), .Z(n4002) );
  AND U5544 ( .A(n922), .B(n4003), .Z(n4001) );
  XOR U5545 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U5546 ( .A(DB[177]), .B(DB[170]), .Z(n4005) );
  AND U5547 ( .A(n926), .B(n4006), .Z(n4004) );
  XOR U5548 ( .A(n4007), .B(n4008), .Z(n4006) );
  XOR U5549 ( .A(DB[170]), .B(DB[163]), .Z(n4008) );
  AND U5550 ( .A(n930), .B(n4009), .Z(n4007) );
  XOR U5551 ( .A(n4010), .B(n4011), .Z(n4009) );
  XOR U5552 ( .A(DB[163]), .B(DB[156]), .Z(n4011) );
  AND U5553 ( .A(n934), .B(n4012), .Z(n4010) );
  XOR U5554 ( .A(n4013), .B(n4014), .Z(n4012) );
  XOR U5555 ( .A(DB[156]), .B(DB[149]), .Z(n4014) );
  AND U5556 ( .A(n938), .B(n4015), .Z(n4013) );
  XOR U5557 ( .A(n4016), .B(n4017), .Z(n4015) );
  XOR U5558 ( .A(DB[149]), .B(DB[142]), .Z(n4017) );
  AND U5559 ( .A(n942), .B(n4018), .Z(n4016) );
  XOR U5560 ( .A(n4019), .B(n4020), .Z(n4018) );
  XOR U5561 ( .A(DB[142]), .B(DB[135]), .Z(n4020) );
  AND U5562 ( .A(n946), .B(n4021), .Z(n4019) );
  XOR U5563 ( .A(n4022), .B(n4023), .Z(n4021) );
  XOR U5564 ( .A(DB[135]), .B(DB[128]), .Z(n4023) );
  AND U5565 ( .A(n950), .B(n4024), .Z(n4022) );
  XOR U5566 ( .A(n4025), .B(n4026), .Z(n4024) );
  XOR U5567 ( .A(DB[128]), .B(DB[121]), .Z(n4026) );
  AND U5568 ( .A(n954), .B(n4027), .Z(n4025) );
  XOR U5569 ( .A(n4028), .B(n4029), .Z(n4027) );
  XOR U5570 ( .A(DB[121]), .B(DB[114]), .Z(n4029) );
  AND U5571 ( .A(n958), .B(n4030), .Z(n4028) );
  XOR U5572 ( .A(n4031), .B(n4032), .Z(n4030) );
  XOR U5573 ( .A(DB[114]), .B(DB[107]), .Z(n4032) );
  AND U5574 ( .A(n962), .B(n4033), .Z(n4031) );
  XOR U5575 ( .A(n4034), .B(n4035), .Z(n4033) );
  XOR U5576 ( .A(DB[107]), .B(DB[100]), .Z(n4035) );
  AND U5577 ( .A(n966), .B(n4036), .Z(n4034) );
  XOR U5578 ( .A(n4037), .B(n4038), .Z(n4036) );
  XOR U5579 ( .A(DB[93]), .B(DB[100]), .Z(n4038) );
  AND U5580 ( .A(n970), .B(n4039), .Z(n4037) );
  XOR U5581 ( .A(n4040), .B(n4041), .Z(n4039) );
  XOR U5582 ( .A(DB[93]), .B(DB[86]), .Z(n4041) );
  AND U5583 ( .A(n974), .B(n4042), .Z(n4040) );
  XOR U5584 ( .A(n4043), .B(n4044), .Z(n4042) );
  XOR U5585 ( .A(DB[86]), .B(DB[79]), .Z(n4044) );
  AND U5586 ( .A(n978), .B(n4045), .Z(n4043) );
  XOR U5587 ( .A(n4046), .B(n4047), .Z(n4045) );
  XOR U5588 ( .A(DB[79]), .B(DB[72]), .Z(n4047) );
  AND U5589 ( .A(n982), .B(n4048), .Z(n4046) );
  XOR U5590 ( .A(n4049), .B(n4050), .Z(n4048) );
  XOR U5591 ( .A(DB[72]), .B(DB[65]), .Z(n4050) );
  AND U5592 ( .A(n986), .B(n4051), .Z(n4049) );
  XOR U5593 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U5594 ( .A(DB[65]), .B(DB[58]), .Z(n4053) );
  AND U5595 ( .A(n990), .B(n4054), .Z(n4052) );
  XOR U5596 ( .A(n4055), .B(n4056), .Z(n4054) );
  XOR U5597 ( .A(DB[58]), .B(DB[51]), .Z(n4056) );
  AND U5598 ( .A(n994), .B(n4057), .Z(n4055) );
  XOR U5599 ( .A(n4058), .B(n4059), .Z(n4057) );
  XOR U5600 ( .A(DB[51]), .B(DB[44]), .Z(n4059) );
  AND U5601 ( .A(n998), .B(n4060), .Z(n4058) );
  XOR U5602 ( .A(n4061), .B(n4062), .Z(n4060) );
  XOR U5603 ( .A(DB[44]), .B(DB[37]), .Z(n4062) );
  AND U5604 ( .A(n1002), .B(n4063), .Z(n4061) );
  XOR U5605 ( .A(n4064), .B(n4065), .Z(n4063) );
  XOR U5606 ( .A(DB[37]), .B(DB[30]), .Z(n4065) );
  AND U5607 ( .A(n1006), .B(n4066), .Z(n4064) );
  XOR U5608 ( .A(n4067), .B(n4068), .Z(n4066) );
  XOR U5609 ( .A(DB[30]), .B(DB[23]), .Z(n4068) );
  AND U5610 ( .A(n1010), .B(n4069), .Z(n4067) );
  XOR U5611 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR U5612 ( .A(DB[23]), .B(DB[16]), .Z(n4071) );
  AND U5613 ( .A(n1014), .B(n4072), .Z(n4070) );
  XOR U5614 ( .A(n4073), .B(n4074), .Z(n4072) );
  XOR U5615 ( .A(DB[9]), .B(DB[16]), .Z(n4074) );
  AND U5616 ( .A(n1018), .B(n4075), .Z(n4073) );
  XOR U5617 ( .A(DB[9]), .B(DB[2]), .Z(n4075) );
  XOR U5618 ( .A(DB[1786]), .B(n4076), .Z(min_val_out[1]) );
  AND U5619 ( .A(n2), .B(n4077), .Z(n4076) );
  XOR U5620 ( .A(n4078), .B(n4079), .Z(n4077) );
  XOR U5621 ( .A(DB[1786]), .B(DB[1779]), .Z(n4079) );
  AND U5622 ( .A(n6), .B(n4080), .Z(n4078) );
  XOR U5623 ( .A(n4081), .B(n4082), .Z(n4080) );
  XOR U5624 ( .A(DB[1779]), .B(DB[1772]), .Z(n4082) );
  AND U5625 ( .A(n10), .B(n4083), .Z(n4081) );
  XOR U5626 ( .A(n4084), .B(n4085), .Z(n4083) );
  XOR U5627 ( .A(DB[1772]), .B(DB[1765]), .Z(n4085) );
  AND U5628 ( .A(n14), .B(n4086), .Z(n4084) );
  XOR U5629 ( .A(n4087), .B(n4088), .Z(n4086) );
  XOR U5630 ( .A(DB[1765]), .B(DB[1758]), .Z(n4088) );
  AND U5631 ( .A(n18), .B(n4089), .Z(n4087) );
  XOR U5632 ( .A(n4090), .B(n4091), .Z(n4089) );
  XOR U5633 ( .A(DB[1758]), .B(DB[1751]), .Z(n4091) );
  AND U5634 ( .A(n22), .B(n4092), .Z(n4090) );
  XOR U5635 ( .A(n4093), .B(n4094), .Z(n4092) );
  XOR U5636 ( .A(DB[1751]), .B(DB[1744]), .Z(n4094) );
  AND U5637 ( .A(n26), .B(n4095), .Z(n4093) );
  XOR U5638 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U5639 ( .A(DB[1744]), .B(DB[1737]), .Z(n4097) );
  AND U5640 ( .A(n30), .B(n4098), .Z(n4096) );
  XOR U5641 ( .A(n4099), .B(n4100), .Z(n4098) );
  XOR U5642 ( .A(DB[1737]), .B(DB[1730]), .Z(n4100) );
  AND U5643 ( .A(n34), .B(n4101), .Z(n4099) );
  XOR U5644 ( .A(n4102), .B(n4103), .Z(n4101) );
  XOR U5645 ( .A(DB[1730]), .B(DB[1723]), .Z(n4103) );
  AND U5646 ( .A(n38), .B(n4104), .Z(n4102) );
  XOR U5647 ( .A(n4105), .B(n4106), .Z(n4104) );
  XOR U5648 ( .A(DB[1723]), .B(DB[1716]), .Z(n4106) );
  AND U5649 ( .A(n42), .B(n4107), .Z(n4105) );
  XOR U5650 ( .A(n4108), .B(n4109), .Z(n4107) );
  XOR U5651 ( .A(DB[1716]), .B(DB[1709]), .Z(n4109) );
  AND U5652 ( .A(n46), .B(n4110), .Z(n4108) );
  XOR U5653 ( .A(n4111), .B(n4112), .Z(n4110) );
  XOR U5654 ( .A(DB[1709]), .B(DB[1702]), .Z(n4112) );
  AND U5655 ( .A(n50), .B(n4113), .Z(n4111) );
  XOR U5656 ( .A(n4114), .B(n4115), .Z(n4113) );
  XOR U5657 ( .A(DB[1702]), .B(DB[1695]), .Z(n4115) );
  AND U5658 ( .A(n54), .B(n4116), .Z(n4114) );
  XOR U5659 ( .A(n4117), .B(n4118), .Z(n4116) );
  XOR U5660 ( .A(DB[1695]), .B(DB[1688]), .Z(n4118) );
  AND U5661 ( .A(n58), .B(n4119), .Z(n4117) );
  XOR U5662 ( .A(n4120), .B(n4121), .Z(n4119) );
  XOR U5663 ( .A(DB[1688]), .B(DB[1681]), .Z(n4121) );
  AND U5664 ( .A(n62), .B(n4122), .Z(n4120) );
  XOR U5665 ( .A(n4123), .B(n4124), .Z(n4122) );
  XOR U5666 ( .A(DB[1681]), .B(DB[1674]), .Z(n4124) );
  AND U5667 ( .A(n66), .B(n4125), .Z(n4123) );
  XOR U5668 ( .A(n4126), .B(n4127), .Z(n4125) );
  XOR U5669 ( .A(DB[1674]), .B(DB[1667]), .Z(n4127) );
  AND U5670 ( .A(n70), .B(n4128), .Z(n4126) );
  XOR U5671 ( .A(n4129), .B(n4130), .Z(n4128) );
  XOR U5672 ( .A(DB[1667]), .B(DB[1660]), .Z(n4130) );
  AND U5673 ( .A(n74), .B(n4131), .Z(n4129) );
  XOR U5674 ( .A(n4132), .B(n4133), .Z(n4131) );
  XOR U5675 ( .A(DB[1660]), .B(DB[1653]), .Z(n4133) );
  AND U5676 ( .A(n78), .B(n4134), .Z(n4132) );
  XOR U5677 ( .A(n4135), .B(n4136), .Z(n4134) );
  XOR U5678 ( .A(DB[1653]), .B(DB[1646]), .Z(n4136) );
  AND U5679 ( .A(n82), .B(n4137), .Z(n4135) );
  XOR U5680 ( .A(n4138), .B(n4139), .Z(n4137) );
  XOR U5681 ( .A(DB[1646]), .B(DB[1639]), .Z(n4139) );
  AND U5682 ( .A(n86), .B(n4140), .Z(n4138) );
  XOR U5683 ( .A(n4141), .B(n4142), .Z(n4140) );
  XOR U5684 ( .A(DB[1639]), .B(DB[1632]), .Z(n4142) );
  AND U5685 ( .A(n90), .B(n4143), .Z(n4141) );
  XOR U5686 ( .A(n4144), .B(n4145), .Z(n4143) );
  XOR U5687 ( .A(DB[1632]), .B(DB[1625]), .Z(n4145) );
  AND U5688 ( .A(n94), .B(n4146), .Z(n4144) );
  XOR U5689 ( .A(n4147), .B(n4148), .Z(n4146) );
  XOR U5690 ( .A(DB[1625]), .B(DB[1618]), .Z(n4148) );
  AND U5691 ( .A(n98), .B(n4149), .Z(n4147) );
  XOR U5692 ( .A(n4150), .B(n4151), .Z(n4149) );
  XOR U5693 ( .A(DB[1618]), .B(DB[1611]), .Z(n4151) );
  AND U5694 ( .A(n102), .B(n4152), .Z(n4150) );
  XOR U5695 ( .A(n4153), .B(n4154), .Z(n4152) );
  XOR U5696 ( .A(DB[1611]), .B(DB[1604]), .Z(n4154) );
  AND U5697 ( .A(n106), .B(n4155), .Z(n4153) );
  XOR U5698 ( .A(n4156), .B(n4157), .Z(n4155) );
  XOR U5699 ( .A(DB[1604]), .B(DB[1597]), .Z(n4157) );
  AND U5700 ( .A(n110), .B(n4158), .Z(n4156) );
  XOR U5701 ( .A(n4159), .B(n4160), .Z(n4158) );
  XOR U5702 ( .A(DB[1597]), .B(DB[1590]), .Z(n4160) );
  AND U5703 ( .A(n114), .B(n4161), .Z(n4159) );
  XOR U5704 ( .A(n4162), .B(n4163), .Z(n4161) );
  XOR U5705 ( .A(DB[1590]), .B(DB[1583]), .Z(n4163) );
  AND U5706 ( .A(n118), .B(n4164), .Z(n4162) );
  XOR U5707 ( .A(n4165), .B(n4166), .Z(n4164) );
  XOR U5708 ( .A(DB[1583]), .B(DB[1576]), .Z(n4166) );
  AND U5709 ( .A(n122), .B(n4167), .Z(n4165) );
  XOR U5710 ( .A(n4168), .B(n4169), .Z(n4167) );
  XOR U5711 ( .A(DB[1576]), .B(DB[1569]), .Z(n4169) );
  AND U5712 ( .A(n126), .B(n4170), .Z(n4168) );
  XOR U5713 ( .A(n4171), .B(n4172), .Z(n4170) );
  XOR U5714 ( .A(DB[1569]), .B(DB[1562]), .Z(n4172) );
  AND U5715 ( .A(n130), .B(n4173), .Z(n4171) );
  XOR U5716 ( .A(n4174), .B(n4175), .Z(n4173) );
  XOR U5717 ( .A(DB[1562]), .B(DB[1555]), .Z(n4175) );
  AND U5718 ( .A(n134), .B(n4176), .Z(n4174) );
  XOR U5719 ( .A(n4177), .B(n4178), .Z(n4176) );
  XOR U5720 ( .A(DB[1555]), .B(DB[1548]), .Z(n4178) );
  AND U5721 ( .A(n138), .B(n4179), .Z(n4177) );
  XOR U5722 ( .A(n4180), .B(n4181), .Z(n4179) );
  XOR U5723 ( .A(DB[1548]), .B(DB[1541]), .Z(n4181) );
  AND U5724 ( .A(n142), .B(n4182), .Z(n4180) );
  XOR U5725 ( .A(n4183), .B(n4184), .Z(n4182) );
  XOR U5726 ( .A(DB[1541]), .B(DB[1534]), .Z(n4184) );
  AND U5727 ( .A(n146), .B(n4185), .Z(n4183) );
  XOR U5728 ( .A(n4186), .B(n4187), .Z(n4185) );
  XOR U5729 ( .A(DB[1534]), .B(DB[1527]), .Z(n4187) );
  AND U5730 ( .A(n150), .B(n4188), .Z(n4186) );
  XOR U5731 ( .A(n4189), .B(n4190), .Z(n4188) );
  XOR U5732 ( .A(DB[1527]), .B(DB[1520]), .Z(n4190) );
  AND U5733 ( .A(n154), .B(n4191), .Z(n4189) );
  XOR U5734 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR U5735 ( .A(DB[1520]), .B(DB[1513]), .Z(n4193) );
  AND U5736 ( .A(n158), .B(n4194), .Z(n4192) );
  XOR U5737 ( .A(n4195), .B(n4196), .Z(n4194) );
  XOR U5738 ( .A(DB[1513]), .B(DB[1506]), .Z(n4196) );
  AND U5739 ( .A(n162), .B(n4197), .Z(n4195) );
  XOR U5740 ( .A(n4198), .B(n4199), .Z(n4197) );
  XOR U5741 ( .A(DB[1506]), .B(DB[1499]), .Z(n4199) );
  AND U5742 ( .A(n166), .B(n4200), .Z(n4198) );
  XOR U5743 ( .A(n4201), .B(n4202), .Z(n4200) );
  XOR U5744 ( .A(DB[1499]), .B(DB[1492]), .Z(n4202) );
  AND U5745 ( .A(n170), .B(n4203), .Z(n4201) );
  XOR U5746 ( .A(n4204), .B(n4205), .Z(n4203) );
  XOR U5747 ( .A(DB[1492]), .B(DB[1485]), .Z(n4205) );
  AND U5748 ( .A(n174), .B(n4206), .Z(n4204) );
  XOR U5749 ( .A(n4207), .B(n4208), .Z(n4206) );
  XOR U5750 ( .A(DB[1485]), .B(DB[1478]), .Z(n4208) );
  AND U5751 ( .A(n178), .B(n4209), .Z(n4207) );
  XOR U5752 ( .A(n4210), .B(n4211), .Z(n4209) );
  XOR U5753 ( .A(DB[1478]), .B(DB[1471]), .Z(n4211) );
  AND U5754 ( .A(n182), .B(n4212), .Z(n4210) );
  XOR U5755 ( .A(n4213), .B(n4214), .Z(n4212) );
  XOR U5756 ( .A(DB[1471]), .B(DB[1464]), .Z(n4214) );
  AND U5757 ( .A(n186), .B(n4215), .Z(n4213) );
  XOR U5758 ( .A(n4216), .B(n4217), .Z(n4215) );
  XOR U5759 ( .A(DB[1464]), .B(DB[1457]), .Z(n4217) );
  AND U5760 ( .A(n190), .B(n4218), .Z(n4216) );
  XOR U5761 ( .A(n4219), .B(n4220), .Z(n4218) );
  XOR U5762 ( .A(DB[1457]), .B(DB[1450]), .Z(n4220) );
  AND U5763 ( .A(n194), .B(n4221), .Z(n4219) );
  XOR U5764 ( .A(n4222), .B(n4223), .Z(n4221) );
  XOR U5765 ( .A(DB[1450]), .B(DB[1443]), .Z(n4223) );
  AND U5766 ( .A(n198), .B(n4224), .Z(n4222) );
  XOR U5767 ( .A(n4225), .B(n4226), .Z(n4224) );
  XOR U5768 ( .A(DB[1443]), .B(DB[1436]), .Z(n4226) );
  AND U5769 ( .A(n202), .B(n4227), .Z(n4225) );
  XOR U5770 ( .A(n4228), .B(n4229), .Z(n4227) );
  XOR U5771 ( .A(DB[1436]), .B(DB[1429]), .Z(n4229) );
  AND U5772 ( .A(n206), .B(n4230), .Z(n4228) );
  XOR U5773 ( .A(n4231), .B(n4232), .Z(n4230) );
  XOR U5774 ( .A(DB[1429]), .B(DB[1422]), .Z(n4232) );
  AND U5775 ( .A(n210), .B(n4233), .Z(n4231) );
  XOR U5776 ( .A(n4234), .B(n4235), .Z(n4233) );
  XOR U5777 ( .A(DB[1422]), .B(DB[1415]), .Z(n4235) );
  AND U5778 ( .A(n214), .B(n4236), .Z(n4234) );
  XOR U5779 ( .A(n4237), .B(n4238), .Z(n4236) );
  XOR U5780 ( .A(DB[1415]), .B(DB[1408]), .Z(n4238) );
  AND U5781 ( .A(n218), .B(n4239), .Z(n4237) );
  XOR U5782 ( .A(n4240), .B(n4241), .Z(n4239) );
  XOR U5783 ( .A(DB[1408]), .B(DB[1401]), .Z(n4241) );
  AND U5784 ( .A(n222), .B(n4242), .Z(n4240) );
  XOR U5785 ( .A(n4243), .B(n4244), .Z(n4242) );
  XOR U5786 ( .A(DB[1401]), .B(DB[1394]), .Z(n4244) );
  AND U5787 ( .A(n226), .B(n4245), .Z(n4243) );
  XOR U5788 ( .A(n4246), .B(n4247), .Z(n4245) );
  XOR U5789 ( .A(DB[1394]), .B(DB[1387]), .Z(n4247) );
  AND U5790 ( .A(n230), .B(n4248), .Z(n4246) );
  XOR U5791 ( .A(n4249), .B(n4250), .Z(n4248) );
  XOR U5792 ( .A(DB[1387]), .B(DB[1380]), .Z(n4250) );
  AND U5793 ( .A(n234), .B(n4251), .Z(n4249) );
  XOR U5794 ( .A(n4252), .B(n4253), .Z(n4251) );
  XOR U5795 ( .A(DB[1380]), .B(DB[1373]), .Z(n4253) );
  AND U5796 ( .A(n238), .B(n4254), .Z(n4252) );
  XOR U5797 ( .A(n4255), .B(n4256), .Z(n4254) );
  XOR U5798 ( .A(DB[1373]), .B(DB[1366]), .Z(n4256) );
  AND U5799 ( .A(n242), .B(n4257), .Z(n4255) );
  XOR U5800 ( .A(n4258), .B(n4259), .Z(n4257) );
  XOR U5801 ( .A(DB[1366]), .B(DB[1359]), .Z(n4259) );
  AND U5802 ( .A(n246), .B(n4260), .Z(n4258) );
  XOR U5803 ( .A(n4261), .B(n4262), .Z(n4260) );
  XOR U5804 ( .A(DB[1359]), .B(DB[1352]), .Z(n4262) );
  AND U5805 ( .A(n250), .B(n4263), .Z(n4261) );
  XOR U5806 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U5807 ( .A(DB[1352]), .B(DB[1345]), .Z(n4265) );
  AND U5808 ( .A(n254), .B(n4266), .Z(n4264) );
  XOR U5809 ( .A(n4267), .B(n4268), .Z(n4266) );
  XOR U5810 ( .A(DB[1345]), .B(DB[1338]), .Z(n4268) );
  AND U5811 ( .A(n258), .B(n4269), .Z(n4267) );
  XOR U5812 ( .A(n4270), .B(n4271), .Z(n4269) );
  XOR U5813 ( .A(DB[1338]), .B(DB[1331]), .Z(n4271) );
  AND U5814 ( .A(n262), .B(n4272), .Z(n4270) );
  XOR U5815 ( .A(n4273), .B(n4274), .Z(n4272) );
  XOR U5816 ( .A(DB[1331]), .B(DB[1324]), .Z(n4274) );
  AND U5817 ( .A(n266), .B(n4275), .Z(n4273) );
  XOR U5818 ( .A(n4276), .B(n4277), .Z(n4275) );
  XOR U5819 ( .A(DB[1324]), .B(DB[1317]), .Z(n4277) );
  AND U5820 ( .A(n270), .B(n4278), .Z(n4276) );
  XOR U5821 ( .A(n4279), .B(n4280), .Z(n4278) );
  XOR U5822 ( .A(DB[1317]), .B(DB[1310]), .Z(n4280) );
  AND U5823 ( .A(n274), .B(n4281), .Z(n4279) );
  XOR U5824 ( .A(n4282), .B(n4283), .Z(n4281) );
  XOR U5825 ( .A(DB[1310]), .B(DB[1303]), .Z(n4283) );
  AND U5826 ( .A(n278), .B(n4284), .Z(n4282) );
  XOR U5827 ( .A(n4285), .B(n4286), .Z(n4284) );
  XOR U5828 ( .A(DB[1303]), .B(DB[1296]), .Z(n4286) );
  AND U5829 ( .A(n282), .B(n4287), .Z(n4285) );
  XOR U5830 ( .A(n4288), .B(n4289), .Z(n4287) );
  XOR U5831 ( .A(DB[1296]), .B(DB[1289]), .Z(n4289) );
  AND U5832 ( .A(n286), .B(n4290), .Z(n4288) );
  XOR U5833 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR U5834 ( .A(DB[1289]), .B(DB[1282]), .Z(n4292) );
  AND U5835 ( .A(n290), .B(n4293), .Z(n4291) );
  XOR U5836 ( .A(n4294), .B(n4295), .Z(n4293) );
  XOR U5837 ( .A(DB[1282]), .B(DB[1275]), .Z(n4295) );
  AND U5838 ( .A(n294), .B(n4296), .Z(n4294) );
  XOR U5839 ( .A(n4297), .B(n4298), .Z(n4296) );
  XOR U5840 ( .A(DB[1275]), .B(DB[1268]), .Z(n4298) );
  AND U5841 ( .A(n298), .B(n4299), .Z(n4297) );
  XOR U5842 ( .A(n4300), .B(n4301), .Z(n4299) );
  XOR U5843 ( .A(DB[1268]), .B(DB[1261]), .Z(n4301) );
  AND U5844 ( .A(n302), .B(n4302), .Z(n4300) );
  XOR U5845 ( .A(n4303), .B(n4304), .Z(n4302) );
  XOR U5846 ( .A(DB[1261]), .B(DB[1254]), .Z(n4304) );
  AND U5847 ( .A(n306), .B(n4305), .Z(n4303) );
  XOR U5848 ( .A(n4306), .B(n4307), .Z(n4305) );
  XOR U5849 ( .A(DB[1254]), .B(DB[1247]), .Z(n4307) );
  AND U5850 ( .A(n310), .B(n4308), .Z(n4306) );
  XOR U5851 ( .A(n4309), .B(n4310), .Z(n4308) );
  XOR U5852 ( .A(DB[1247]), .B(DB[1240]), .Z(n4310) );
  AND U5853 ( .A(n314), .B(n4311), .Z(n4309) );
  XOR U5854 ( .A(n4312), .B(n4313), .Z(n4311) );
  XOR U5855 ( .A(DB[1240]), .B(DB[1233]), .Z(n4313) );
  AND U5856 ( .A(n318), .B(n4314), .Z(n4312) );
  XOR U5857 ( .A(n4315), .B(n4316), .Z(n4314) );
  XOR U5858 ( .A(DB[1233]), .B(DB[1226]), .Z(n4316) );
  AND U5859 ( .A(n322), .B(n4317), .Z(n4315) );
  XOR U5860 ( .A(n4318), .B(n4319), .Z(n4317) );
  XOR U5861 ( .A(DB[1226]), .B(DB[1219]), .Z(n4319) );
  AND U5862 ( .A(n326), .B(n4320), .Z(n4318) );
  XOR U5863 ( .A(n4321), .B(n4322), .Z(n4320) );
  XOR U5864 ( .A(DB[1219]), .B(DB[1212]), .Z(n4322) );
  AND U5865 ( .A(n330), .B(n4323), .Z(n4321) );
  XOR U5866 ( .A(n4324), .B(n4325), .Z(n4323) );
  XOR U5867 ( .A(DB[1212]), .B(DB[1205]), .Z(n4325) );
  AND U5868 ( .A(n334), .B(n4326), .Z(n4324) );
  XOR U5869 ( .A(n4327), .B(n4328), .Z(n4326) );
  XOR U5870 ( .A(DB[1205]), .B(DB[1198]), .Z(n4328) );
  AND U5871 ( .A(n338), .B(n4329), .Z(n4327) );
  XOR U5872 ( .A(n4330), .B(n4331), .Z(n4329) );
  XOR U5873 ( .A(DB[1198]), .B(DB[1191]), .Z(n4331) );
  AND U5874 ( .A(n342), .B(n4332), .Z(n4330) );
  XOR U5875 ( .A(n4333), .B(n4334), .Z(n4332) );
  XOR U5876 ( .A(DB[1191]), .B(DB[1184]), .Z(n4334) );
  AND U5877 ( .A(n346), .B(n4335), .Z(n4333) );
  XOR U5878 ( .A(n4336), .B(n4337), .Z(n4335) );
  XOR U5879 ( .A(DB[1184]), .B(DB[1177]), .Z(n4337) );
  AND U5880 ( .A(n350), .B(n4338), .Z(n4336) );
  XOR U5881 ( .A(n4339), .B(n4340), .Z(n4338) );
  XOR U5882 ( .A(DB[1177]), .B(DB[1170]), .Z(n4340) );
  AND U5883 ( .A(n354), .B(n4341), .Z(n4339) );
  XOR U5884 ( .A(n4342), .B(n4343), .Z(n4341) );
  XOR U5885 ( .A(DB[1170]), .B(DB[1163]), .Z(n4343) );
  AND U5886 ( .A(n358), .B(n4344), .Z(n4342) );
  XOR U5887 ( .A(n4345), .B(n4346), .Z(n4344) );
  XOR U5888 ( .A(DB[1163]), .B(DB[1156]), .Z(n4346) );
  AND U5889 ( .A(n362), .B(n4347), .Z(n4345) );
  XOR U5890 ( .A(n4348), .B(n4349), .Z(n4347) );
  XOR U5891 ( .A(DB[1156]), .B(DB[1149]), .Z(n4349) );
  AND U5892 ( .A(n366), .B(n4350), .Z(n4348) );
  XOR U5893 ( .A(n4351), .B(n4352), .Z(n4350) );
  XOR U5894 ( .A(DB[1149]), .B(DB[1142]), .Z(n4352) );
  AND U5895 ( .A(n370), .B(n4353), .Z(n4351) );
  XOR U5896 ( .A(n4354), .B(n4355), .Z(n4353) );
  XOR U5897 ( .A(DB[1142]), .B(DB[1135]), .Z(n4355) );
  AND U5898 ( .A(n374), .B(n4356), .Z(n4354) );
  XOR U5899 ( .A(n4357), .B(n4358), .Z(n4356) );
  XOR U5900 ( .A(DB[1135]), .B(DB[1128]), .Z(n4358) );
  AND U5901 ( .A(n378), .B(n4359), .Z(n4357) );
  XOR U5902 ( .A(n4360), .B(n4361), .Z(n4359) );
  XOR U5903 ( .A(DB[1128]), .B(DB[1121]), .Z(n4361) );
  AND U5904 ( .A(n382), .B(n4362), .Z(n4360) );
  XOR U5905 ( .A(n4363), .B(n4364), .Z(n4362) );
  XOR U5906 ( .A(DB[1121]), .B(DB[1114]), .Z(n4364) );
  AND U5907 ( .A(n386), .B(n4365), .Z(n4363) );
  XOR U5908 ( .A(n4366), .B(n4367), .Z(n4365) );
  XOR U5909 ( .A(DB[1114]), .B(DB[1107]), .Z(n4367) );
  AND U5910 ( .A(n390), .B(n4368), .Z(n4366) );
  XOR U5911 ( .A(n4369), .B(n4370), .Z(n4368) );
  XOR U5912 ( .A(DB[1107]), .B(DB[1100]), .Z(n4370) );
  AND U5913 ( .A(n394), .B(n4371), .Z(n4369) );
  XOR U5914 ( .A(n4372), .B(n4373), .Z(n4371) );
  XOR U5915 ( .A(DB[1100]), .B(DB[1093]), .Z(n4373) );
  AND U5916 ( .A(n398), .B(n4374), .Z(n4372) );
  XOR U5917 ( .A(n4375), .B(n4376), .Z(n4374) );
  XOR U5918 ( .A(DB[1093]), .B(DB[1086]), .Z(n4376) );
  AND U5919 ( .A(n402), .B(n4377), .Z(n4375) );
  XOR U5920 ( .A(n4378), .B(n4379), .Z(n4377) );
  XOR U5921 ( .A(DB[1086]), .B(DB[1079]), .Z(n4379) );
  AND U5922 ( .A(n406), .B(n4380), .Z(n4378) );
  XOR U5923 ( .A(n4381), .B(n4382), .Z(n4380) );
  XOR U5924 ( .A(DB[1079]), .B(DB[1072]), .Z(n4382) );
  AND U5925 ( .A(n410), .B(n4383), .Z(n4381) );
  XOR U5926 ( .A(n4384), .B(n4385), .Z(n4383) );
  XOR U5927 ( .A(DB[1072]), .B(DB[1065]), .Z(n4385) );
  AND U5928 ( .A(n414), .B(n4386), .Z(n4384) );
  XOR U5929 ( .A(n4387), .B(n4388), .Z(n4386) );
  XOR U5930 ( .A(DB[1065]), .B(DB[1058]), .Z(n4388) );
  AND U5931 ( .A(n418), .B(n4389), .Z(n4387) );
  XOR U5932 ( .A(n4390), .B(n4391), .Z(n4389) );
  XOR U5933 ( .A(DB[1058]), .B(DB[1051]), .Z(n4391) );
  AND U5934 ( .A(n422), .B(n4392), .Z(n4390) );
  XOR U5935 ( .A(n4393), .B(n4394), .Z(n4392) );
  XOR U5936 ( .A(DB[1051]), .B(DB[1044]), .Z(n4394) );
  AND U5937 ( .A(n426), .B(n4395), .Z(n4393) );
  XOR U5938 ( .A(n4396), .B(n4397), .Z(n4395) );
  XOR U5939 ( .A(DB[1044]), .B(DB[1037]), .Z(n4397) );
  AND U5940 ( .A(n430), .B(n4398), .Z(n4396) );
  XOR U5941 ( .A(n4399), .B(n4400), .Z(n4398) );
  XOR U5942 ( .A(DB[1037]), .B(DB[1030]), .Z(n4400) );
  AND U5943 ( .A(n434), .B(n4401), .Z(n4399) );
  XOR U5944 ( .A(n4402), .B(n4403), .Z(n4401) );
  XOR U5945 ( .A(DB[1030]), .B(DB[1023]), .Z(n4403) );
  AND U5946 ( .A(n438), .B(n4404), .Z(n4402) );
  XOR U5947 ( .A(n4405), .B(n4406), .Z(n4404) );
  XOR U5948 ( .A(DB[1023]), .B(DB[1016]), .Z(n4406) );
  AND U5949 ( .A(n442), .B(n4407), .Z(n4405) );
  XOR U5950 ( .A(n4408), .B(n4409), .Z(n4407) );
  XOR U5951 ( .A(DB[1016]), .B(DB[1009]), .Z(n4409) );
  AND U5952 ( .A(n446), .B(n4410), .Z(n4408) );
  XOR U5953 ( .A(n4411), .B(n4412), .Z(n4410) );
  XOR U5954 ( .A(DB[1009]), .B(DB[1002]), .Z(n4412) );
  AND U5955 ( .A(n450), .B(n4413), .Z(n4411) );
  XOR U5956 ( .A(n4414), .B(n4415), .Z(n4413) );
  XOR U5957 ( .A(DB[995]), .B(DB[1002]), .Z(n4415) );
  AND U5958 ( .A(n454), .B(n4416), .Z(n4414) );
  XOR U5959 ( .A(n4417), .B(n4418), .Z(n4416) );
  XOR U5960 ( .A(DB[995]), .B(DB[988]), .Z(n4418) );
  AND U5961 ( .A(n458), .B(n4419), .Z(n4417) );
  XOR U5962 ( .A(n4420), .B(n4421), .Z(n4419) );
  XOR U5963 ( .A(DB[988]), .B(DB[981]), .Z(n4421) );
  AND U5964 ( .A(n462), .B(n4422), .Z(n4420) );
  XOR U5965 ( .A(n4423), .B(n4424), .Z(n4422) );
  XOR U5966 ( .A(DB[981]), .B(DB[974]), .Z(n4424) );
  AND U5967 ( .A(n466), .B(n4425), .Z(n4423) );
  XOR U5968 ( .A(n4426), .B(n4427), .Z(n4425) );
  XOR U5969 ( .A(DB[974]), .B(DB[967]), .Z(n4427) );
  AND U5970 ( .A(n470), .B(n4428), .Z(n4426) );
  XOR U5971 ( .A(n4429), .B(n4430), .Z(n4428) );
  XOR U5972 ( .A(DB[967]), .B(DB[960]), .Z(n4430) );
  AND U5973 ( .A(n474), .B(n4431), .Z(n4429) );
  XOR U5974 ( .A(n4432), .B(n4433), .Z(n4431) );
  XOR U5975 ( .A(DB[960]), .B(DB[953]), .Z(n4433) );
  AND U5976 ( .A(n478), .B(n4434), .Z(n4432) );
  XOR U5977 ( .A(n4435), .B(n4436), .Z(n4434) );
  XOR U5978 ( .A(DB[953]), .B(DB[946]), .Z(n4436) );
  AND U5979 ( .A(n482), .B(n4437), .Z(n4435) );
  XOR U5980 ( .A(n4438), .B(n4439), .Z(n4437) );
  XOR U5981 ( .A(DB[946]), .B(DB[939]), .Z(n4439) );
  AND U5982 ( .A(n486), .B(n4440), .Z(n4438) );
  XOR U5983 ( .A(n4441), .B(n4442), .Z(n4440) );
  XOR U5984 ( .A(DB[939]), .B(DB[932]), .Z(n4442) );
  AND U5985 ( .A(n490), .B(n4443), .Z(n4441) );
  XOR U5986 ( .A(n4444), .B(n4445), .Z(n4443) );
  XOR U5987 ( .A(DB[932]), .B(DB[925]), .Z(n4445) );
  AND U5988 ( .A(n494), .B(n4446), .Z(n4444) );
  XOR U5989 ( .A(n4447), .B(n4448), .Z(n4446) );
  XOR U5990 ( .A(DB[925]), .B(DB[918]), .Z(n4448) );
  AND U5991 ( .A(n498), .B(n4449), .Z(n4447) );
  XOR U5992 ( .A(n4450), .B(n4451), .Z(n4449) );
  XOR U5993 ( .A(DB[918]), .B(DB[911]), .Z(n4451) );
  AND U5994 ( .A(n502), .B(n4452), .Z(n4450) );
  XOR U5995 ( .A(n4453), .B(n4454), .Z(n4452) );
  XOR U5996 ( .A(DB[911]), .B(DB[904]), .Z(n4454) );
  AND U5997 ( .A(n506), .B(n4455), .Z(n4453) );
  XOR U5998 ( .A(n4456), .B(n4457), .Z(n4455) );
  XOR U5999 ( .A(DB[904]), .B(DB[897]), .Z(n4457) );
  AND U6000 ( .A(n510), .B(n4458), .Z(n4456) );
  XOR U6001 ( .A(n4459), .B(n4460), .Z(n4458) );
  XOR U6002 ( .A(DB[897]), .B(DB[890]), .Z(n4460) );
  AND U6003 ( .A(n514), .B(n4461), .Z(n4459) );
  XOR U6004 ( .A(n4462), .B(n4463), .Z(n4461) );
  XOR U6005 ( .A(DB[890]), .B(DB[883]), .Z(n4463) );
  AND U6006 ( .A(n518), .B(n4464), .Z(n4462) );
  XOR U6007 ( .A(n4465), .B(n4466), .Z(n4464) );
  XOR U6008 ( .A(DB[883]), .B(DB[876]), .Z(n4466) );
  AND U6009 ( .A(n522), .B(n4467), .Z(n4465) );
  XOR U6010 ( .A(n4468), .B(n4469), .Z(n4467) );
  XOR U6011 ( .A(DB[876]), .B(DB[869]), .Z(n4469) );
  AND U6012 ( .A(n526), .B(n4470), .Z(n4468) );
  XOR U6013 ( .A(n4471), .B(n4472), .Z(n4470) );
  XOR U6014 ( .A(DB[869]), .B(DB[862]), .Z(n4472) );
  AND U6015 ( .A(n530), .B(n4473), .Z(n4471) );
  XOR U6016 ( .A(n4474), .B(n4475), .Z(n4473) );
  XOR U6017 ( .A(DB[862]), .B(DB[855]), .Z(n4475) );
  AND U6018 ( .A(n534), .B(n4476), .Z(n4474) );
  XOR U6019 ( .A(n4477), .B(n4478), .Z(n4476) );
  XOR U6020 ( .A(DB[855]), .B(DB[848]), .Z(n4478) );
  AND U6021 ( .A(n538), .B(n4479), .Z(n4477) );
  XOR U6022 ( .A(n4480), .B(n4481), .Z(n4479) );
  XOR U6023 ( .A(DB[848]), .B(DB[841]), .Z(n4481) );
  AND U6024 ( .A(n542), .B(n4482), .Z(n4480) );
  XOR U6025 ( .A(n4483), .B(n4484), .Z(n4482) );
  XOR U6026 ( .A(DB[841]), .B(DB[834]), .Z(n4484) );
  AND U6027 ( .A(n546), .B(n4485), .Z(n4483) );
  XOR U6028 ( .A(n4486), .B(n4487), .Z(n4485) );
  XOR U6029 ( .A(DB[834]), .B(DB[827]), .Z(n4487) );
  AND U6030 ( .A(n550), .B(n4488), .Z(n4486) );
  XOR U6031 ( .A(n4489), .B(n4490), .Z(n4488) );
  XOR U6032 ( .A(DB[827]), .B(DB[820]), .Z(n4490) );
  AND U6033 ( .A(n554), .B(n4491), .Z(n4489) );
  XOR U6034 ( .A(n4492), .B(n4493), .Z(n4491) );
  XOR U6035 ( .A(DB[820]), .B(DB[813]), .Z(n4493) );
  AND U6036 ( .A(n558), .B(n4494), .Z(n4492) );
  XOR U6037 ( .A(n4495), .B(n4496), .Z(n4494) );
  XOR U6038 ( .A(DB[813]), .B(DB[806]), .Z(n4496) );
  AND U6039 ( .A(n562), .B(n4497), .Z(n4495) );
  XOR U6040 ( .A(n4498), .B(n4499), .Z(n4497) );
  XOR U6041 ( .A(DB[806]), .B(DB[799]), .Z(n4499) );
  AND U6042 ( .A(n566), .B(n4500), .Z(n4498) );
  XOR U6043 ( .A(n4501), .B(n4502), .Z(n4500) );
  XOR U6044 ( .A(DB[799]), .B(DB[792]), .Z(n4502) );
  AND U6045 ( .A(n570), .B(n4503), .Z(n4501) );
  XOR U6046 ( .A(n4504), .B(n4505), .Z(n4503) );
  XOR U6047 ( .A(DB[792]), .B(DB[785]), .Z(n4505) );
  AND U6048 ( .A(n574), .B(n4506), .Z(n4504) );
  XOR U6049 ( .A(n4507), .B(n4508), .Z(n4506) );
  XOR U6050 ( .A(DB[785]), .B(DB[778]), .Z(n4508) );
  AND U6051 ( .A(n578), .B(n4509), .Z(n4507) );
  XOR U6052 ( .A(n4510), .B(n4511), .Z(n4509) );
  XOR U6053 ( .A(DB[778]), .B(DB[771]), .Z(n4511) );
  AND U6054 ( .A(n582), .B(n4512), .Z(n4510) );
  XOR U6055 ( .A(n4513), .B(n4514), .Z(n4512) );
  XOR U6056 ( .A(DB[771]), .B(DB[764]), .Z(n4514) );
  AND U6057 ( .A(n586), .B(n4515), .Z(n4513) );
  XOR U6058 ( .A(n4516), .B(n4517), .Z(n4515) );
  XOR U6059 ( .A(DB[764]), .B(DB[757]), .Z(n4517) );
  AND U6060 ( .A(n590), .B(n4518), .Z(n4516) );
  XOR U6061 ( .A(n4519), .B(n4520), .Z(n4518) );
  XOR U6062 ( .A(DB[757]), .B(DB[750]), .Z(n4520) );
  AND U6063 ( .A(n594), .B(n4521), .Z(n4519) );
  XOR U6064 ( .A(n4522), .B(n4523), .Z(n4521) );
  XOR U6065 ( .A(DB[750]), .B(DB[743]), .Z(n4523) );
  AND U6066 ( .A(n598), .B(n4524), .Z(n4522) );
  XOR U6067 ( .A(n4525), .B(n4526), .Z(n4524) );
  XOR U6068 ( .A(DB[743]), .B(DB[736]), .Z(n4526) );
  AND U6069 ( .A(n602), .B(n4527), .Z(n4525) );
  XOR U6070 ( .A(n4528), .B(n4529), .Z(n4527) );
  XOR U6071 ( .A(DB[736]), .B(DB[729]), .Z(n4529) );
  AND U6072 ( .A(n606), .B(n4530), .Z(n4528) );
  XOR U6073 ( .A(n4531), .B(n4532), .Z(n4530) );
  XOR U6074 ( .A(DB[729]), .B(DB[722]), .Z(n4532) );
  AND U6075 ( .A(n610), .B(n4533), .Z(n4531) );
  XOR U6076 ( .A(n4534), .B(n4535), .Z(n4533) );
  XOR U6077 ( .A(DB[722]), .B(DB[715]), .Z(n4535) );
  AND U6078 ( .A(n614), .B(n4536), .Z(n4534) );
  XOR U6079 ( .A(n4537), .B(n4538), .Z(n4536) );
  XOR U6080 ( .A(DB[715]), .B(DB[708]), .Z(n4538) );
  AND U6081 ( .A(n618), .B(n4539), .Z(n4537) );
  XOR U6082 ( .A(n4540), .B(n4541), .Z(n4539) );
  XOR U6083 ( .A(DB[708]), .B(DB[701]), .Z(n4541) );
  AND U6084 ( .A(n622), .B(n4542), .Z(n4540) );
  XOR U6085 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U6086 ( .A(DB[701]), .B(DB[694]), .Z(n4544) );
  AND U6087 ( .A(n626), .B(n4545), .Z(n4543) );
  XOR U6088 ( .A(n4546), .B(n4547), .Z(n4545) );
  XOR U6089 ( .A(DB[694]), .B(DB[687]), .Z(n4547) );
  AND U6090 ( .A(n630), .B(n4548), .Z(n4546) );
  XOR U6091 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U6092 ( .A(DB[687]), .B(DB[680]), .Z(n4550) );
  AND U6093 ( .A(n634), .B(n4551), .Z(n4549) );
  XOR U6094 ( .A(n4552), .B(n4553), .Z(n4551) );
  XOR U6095 ( .A(DB[680]), .B(DB[673]), .Z(n4553) );
  AND U6096 ( .A(n638), .B(n4554), .Z(n4552) );
  XOR U6097 ( .A(n4555), .B(n4556), .Z(n4554) );
  XOR U6098 ( .A(DB[673]), .B(DB[666]), .Z(n4556) );
  AND U6099 ( .A(n642), .B(n4557), .Z(n4555) );
  XOR U6100 ( .A(n4558), .B(n4559), .Z(n4557) );
  XOR U6101 ( .A(DB[666]), .B(DB[659]), .Z(n4559) );
  AND U6102 ( .A(n646), .B(n4560), .Z(n4558) );
  XOR U6103 ( .A(n4561), .B(n4562), .Z(n4560) );
  XOR U6104 ( .A(DB[659]), .B(DB[652]), .Z(n4562) );
  AND U6105 ( .A(n650), .B(n4563), .Z(n4561) );
  XOR U6106 ( .A(n4564), .B(n4565), .Z(n4563) );
  XOR U6107 ( .A(DB[652]), .B(DB[645]), .Z(n4565) );
  AND U6108 ( .A(n654), .B(n4566), .Z(n4564) );
  XOR U6109 ( .A(n4567), .B(n4568), .Z(n4566) );
  XOR U6110 ( .A(DB[645]), .B(DB[638]), .Z(n4568) );
  AND U6111 ( .A(n658), .B(n4569), .Z(n4567) );
  XOR U6112 ( .A(n4570), .B(n4571), .Z(n4569) );
  XOR U6113 ( .A(DB[638]), .B(DB[631]), .Z(n4571) );
  AND U6114 ( .A(n662), .B(n4572), .Z(n4570) );
  XOR U6115 ( .A(n4573), .B(n4574), .Z(n4572) );
  XOR U6116 ( .A(DB[631]), .B(DB[624]), .Z(n4574) );
  AND U6117 ( .A(n666), .B(n4575), .Z(n4573) );
  XOR U6118 ( .A(n4576), .B(n4577), .Z(n4575) );
  XOR U6119 ( .A(DB[624]), .B(DB[617]), .Z(n4577) );
  AND U6120 ( .A(n670), .B(n4578), .Z(n4576) );
  XOR U6121 ( .A(n4579), .B(n4580), .Z(n4578) );
  XOR U6122 ( .A(DB[617]), .B(DB[610]), .Z(n4580) );
  AND U6123 ( .A(n674), .B(n4581), .Z(n4579) );
  XOR U6124 ( .A(n4582), .B(n4583), .Z(n4581) );
  XOR U6125 ( .A(DB[610]), .B(DB[603]), .Z(n4583) );
  AND U6126 ( .A(n678), .B(n4584), .Z(n4582) );
  XOR U6127 ( .A(n4585), .B(n4586), .Z(n4584) );
  XOR U6128 ( .A(DB[603]), .B(DB[596]), .Z(n4586) );
  AND U6129 ( .A(n682), .B(n4587), .Z(n4585) );
  XOR U6130 ( .A(n4588), .B(n4589), .Z(n4587) );
  XOR U6131 ( .A(DB[596]), .B(DB[589]), .Z(n4589) );
  AND U6132 ( .A(n686), .B(n4590), .Z(n4588) );
  XOR U6133 ( .A(n4591), .B(n4592), .Z(n4590) );
  XOR U6134 ( .A(DB[589]), .B(DB[582]), .Z(n4592) );
  AND U6135 ( .A(n690), .B(n4593), .Z(n4591) );
  XOR U6136 ( .A(n4594), .B(n4595), .Z(n4593) );
  XOR U6137 ( .A(DB[582]), .B(DB[575]), .Z(n4595) );
  AND U6138 ( .A(n694), .B(n4596), .Z(n4594) );
  XOR U6139 ( .A(n4597), .B(n4598), .Z(n4596) );
  XOR U6140 ( .A(DB[575]), .B(DB[568]), .Z(n4598) );
  AND U6141 ( .A(n698), .B(n4599), .Z(n4597) );
  XOR U6142 ( .A(n4600), .B(n4601), .Z(n4599) );
  XOR U6143 ( .A(DB[568]), .B(DB[561]), .Z(n4601) );
  AND U6144 ( .A(n702), .B(n4602), .Z(n4600) );
  XOR U6145 ( .A(n4603), .B(n4604), .Z(n4602) );
  XOR U6146 ( .A(DB[561]), .B(DB[554]), .Z(n4604) );
  AND U6147 ( .A(n706), .B(n4605), .Z(n4603) );
  XOR U6148 ( .A(n4606), .B(n4607), .Z(n4605) );
  XOR U6149 ( .A(DB[554]), .B(DB[547]), .Z(n4607) );
  AND U6150 ( .A(n710), .B(n4608), .Z(n4606) );
  XOR U6151 ( .A(n4609), .B(n4610), .Z(n4608) );
  XOR U6152 ( .A(DB[547]), .B(DB[540]), .Z(n4610) );
  AND U6153 ( .A(n714), .B(n4611), .Z(n4609) );
  XOR U6154 ( .A(n4612), .B(n4613), .Z(n4611) );
  XOR U6155 ( .A(DB[540]), .B(DB[533]), .Z(n4613) );
  AND U6156 ( .A(n718), .B(n4614), .Z(n4612) );
  XOR U6157 ( .A(n4615), .B(n4616), .Z(n4614) );
  XOR U6158 ( .A(DB[533]), .B(DB[526]), .Z(n4616) );
  AND U6159 ( .A(n722), .B(n4617), .Z(n4615) );
  XOR U6160 ( .A(n4618), .B(n4619), .Z(n4617) );
  XOR U6161 ( .A(DB[526]), .B(DB[519]), .Z(n4619) );
  AND U6162 ( .A(n726), .B(n4620), .Z(n4618) );
  XOR U6163 ( .A(n4621), .B(n4622), .Z(n4620) );
  XOR U6164 ( .A(DB[519]), .B(DB[512]), .Z(n4622) );
  AND U6165 ( .A(n730), .B(n4623), .Z(n4621) );
  XOR U6166 ( .A(n4624), .B(n4625), .Z(n4623) );
  XOR U6167 ( .A(DB[512]), .B(DB[505]), .Z(n4625) );
  AND U6168 ( .A(n734), .B(n4626), .Z(n4624) );
  XOR U6169 ( .A(n4627), .B(n4628), .Z(n4626) );
  XOR U6170 ( .A(DB[505]), .B(DB[498]), .Z(n4628) );
  AND U6171 ( .A(n738), .B(n4629), .Z(n4627) );
  XOR U6172 ( .A(n4630), .B(n4631), .Z(n4629) );
  XOR U6173 ( .A(DB[498]), .B(DB[491]), .Z(n4631) );
  AND U6174 ( .A(n742), .B(n4632), .Z(n4630) );
  XOR U6175 ( .A(n4633), .B(n4634), .Z(n4632) );
  XOR U6176 ( .A(DB[491]), .B(DB[484]), .Z(n4634) );
  AND U6177 ( .A(n746), .B(n4635), .Z(n4633) );
  XOR U6178 ( .A(n4636), .B(n4637), .Z(n4635) );
  XOR U6179 ( .A(DB[484]), .B(DB[477]), .Z(n4637) );
  AND U6180 ( .A(n750), .B(n4638), .Z(n4636) );
  XOR U6181 ( .A(n4639), .B(n4640), .Z(n4638) );
  XOR U6182 ( .A(DB[477]), .B(DB[470]), .Z(n4640) );
  AND U6183 ( .A(n754), .B(n4641), .Z(n4639) );
  XOR U6184 ( .A(n4642), .B(n4643), .Z(n4641) );
  XOR U6185 ( .A(DB[470]), .B(DB[463]), .Z(n4643) );
  AND U6186 ( .A(n758), .B(n4644), .Z(n4642) );
  XOR U6187 ( .A(n4645), .B(n4646), .Z(n4644) );
  XOR U6188 ( .A(DB[463]), .B(DB[456]), .Z(n4646) );
  AND U6189 ( .A(n762), .B(n4647), .Z(n4645) );
  XOR U6190 ( .A(n4648), .B(n4649), .Z(n4647) );
  XOR U6191 ( .A(DB[456]), .B(DB[449]), .Z(n4649) );
  AND U6192 ( .A(n766), .B(n4650), .Z(n4648) );
  XOR U6193 ( .A(n4651), .B(n4652), .Z(n4650) );
  XOR U6194 ( .A(DB[449]), .B(DB[442]), .Z(n4652) );
  AND U6195 ( .A(n770), .B(n4653), .Z(n4651) );
  XOR U6196 ( .A(n4654), .B(n4655), .Z(n4653) );
  XOR U6197 ( .A(DB[442]), .B(DB[435]), .Z(n4655) );
  AND U6198 ( .A(n774), .B(n4656), .Z(n4654) );
  XOR U6199 ( .A(n4657), .B(n4658), .Z(n4656) );
  XOR U6200 ( .A(DB[435]), .B(DB[428]), .Z(n4658) );
  AND U6201 ( .A(n778), .B(n4659), .Z(n4657) );
  XOR U6202 ( .A(n4660), .B(n4661), .Z(n4659) );
  XOR U6203 ( .A(DB[428]), .B(DB[421]), .Z(n4661) );
  AND U6204 ( .A(n782), .B(n4662), .Z(n4660) );
  XOR U6205 ( .A(n4663), .B(n4664), .Z(n4662) );
  XOR U6206 ( .A(DB[421]), .B(DB[414]), .Z(n4664) );
  AND U6207 ( .A(n786), .B(n4665), .Z(n4663) );
  XOR U6208 ( .A(n4666), .B(n4667), .Z(n4665) );
  XOR U6209 ( .A(DB[414]), .B(DB[407]), .Z(n4667) );
  AND U6210 ( .A(n790), .B(n4668), .Z(n4666) );
  XOR U6211 ( .A(n4669), .B(n4670), .Z(n4668) );
  XOR U6212 ( .A(DB[407]), .B(DB[400]), .Z(n4670) );
  AND U6213 ( .A(n794), .B(n4671), .Z(n4669) );
  XOR U6214 ( .A(n4672), .B(n4673), .Z(n4671) );
  XOR U6215 ( .A(DB[400]), .B(DB[393]), .Z(n4673) );
  AND U6216 ( .A(n798), .B(n4674), .Z(n4672) );
  XOR U6217 ( .A(n4675), .B(n4676), .Z(n4674) );
  XOR U6218 ( .A(DB[393]), .B(DB[386]), .Z(n4676) );
  AND U6219 ( .A(n802), .B(n4677), .Z(n4675) );
  XOR U6220 ( .A(n4678), .B(n4679), .Z(n4677) );
  XOR U6221 ( .A(DB[386]), .B(DB[379]), .Z(n4679) );
  AND U6222 ( .A(n806), .B(n4680), .Z(n4678) );
  XOR U6223 ( .A(n4681), .B(n4682), .Z(n4680) );
  XOR U6224 ( .A(DB[379]), .B(DB[372]), .Z(n4682) );
  AND U6225 ( .A(n810), .B(n4683), .Z(n4681) );
  XOR U6226 ( .A(n4684), .B(n4685), .Z(n4683) );
  XOR U6227 ( .A(DB[372]), .B(DB[365]), .Z(n4685) );
  AND U6228 ( .A(n814), .B(n4686), .Z(n4684) );
  XOR U6229 ( .A(n4687), .B(n4688), .Z(n4686) );
  XOR U6230 ( .A(DB[365]), .B(DB[358]), .Z(n4688) );
  AND U6231 ( .A(n818), .B(n4689), .Z(n4687) );
  XOR U6232 ( .A(n4690), .B(n4691), .Z(n4689) );
  XOR U6233 ( .A(DB[358]), .B(DB[351]), .Z(n4691) );
  AND U6234 ( .A(n822), .B(n4692), .Z(n4690) );
  XOR U6235 ( .A(n4693), .B(n4694), .Z(n4692) );
  XOR U6236 ( .A(DB[351]), .B(DB[344]), .Z(n4694) );
  AND U6237 ( .A(n826), .B(n4695), .Z(n4693) );
  XOR U6238 ( .A(n4696), .B(n4697), .Z(n4695) );
  XOR U6239 ( .A(DB[344]), .B(DB[337]), .Z(n4697) );
  AND U6240 ( .A(n830), .B(n4698), .Z(n4696) );
  XOR U6241 ( .A(n4699), .B(n4700), .Z(n4698) );
  XOR U6242 ( .A(DB[337]), .B(DB[330]), .Z(n4700) );
  AND U6243 ( .A(n834), .B(n4701), .Z(n4699) );
  XOR U6244 ( .A(n4702), .B(n4703), .Z(n4701) );
  XOR U6245 ( .A(DB[330]), .B(DB[323]), .Z(n4703) );
  AND U6246 ( .A(n838), .B(n4704), .Z(n4702) );
  XOR U6247 ( .A(n4705), .B(n4706), .Z(n4704) );
  XOR U6248 ( .A(DB[323]), .B(DB[316]), .Z(n4706) );
  AND U6249 ( .A(n842), .B(n4707), .Z(n4705) );
  XOR U6250 ( .A(n4708), .B(n4709), .Z(n4707) );
  XOR U6251 ( .A(DB[316]), .B(DB[309]), .Z(n4709) );
  AND U6252 ( .A(n846), .B(n4710), .Z(n4708) );
  XOR U6253 ( .A(n4711), .B(n4712), .Z(n4710) );
  XOR U6254 ( .A(DB[309]), .B(DB[302]), .Z(n4712) );
  AND U6255 ( .A(n850), .B(n4713), .Z(n4711) );
  XOR U6256 ( .A(n4714), .B(n4715), .Z(n4713) );
  XOR U6257 ( .A(DB[302]), .B(DB[295]), .Z(n4715) );
  AND U6258 ( .A(n854), .B(n4716), .Z(n4714) );
  XOR U6259 ( .A(n4717), .B(n4718), .Z(n4716) );
  XOR U6260 ( .A(DB[295]), .B(DB[288]), .Z(n4718) );
  AND U6261 ( .A(n858), .B(n4719), .Z(n4717) );
  XOR U6262 ( .A(n4720), .B(n4721), .Z(n4719) );
  XOR U6263 ( .A(DB[288]), .B(DB[281]), .Z(n4721) );
  AND U6264 ( .A(n862), .B(n4722), .Z(n4720) );
  XOR U6265 ( .A(n4723), .B(n4724), .Z(n4722) );
  XOR U6266 ( .A(DB[281]), .B(DB[274]), .Z(n4724) );
  AND U6267 ( .A(n866), .B(n4725), .Z(n4723) );
  XOR U6268 ( .A(n4726), .B(n4727), .Z(n4725) );
  XOR U6269 ( .A(DB[274]), .B(DB[267]), .Z(n4727) );
  AND U6270 ( .A(n870), .B(n4728), .Z(n4726) );
  XOR U6271 ( .A(n4729), .B(n4730), .Z(n4728) );
  XOR U6272 ( .A(DB[267]), .B(DB[260]), .Z(n4730) );
  AND U6273 ( .A(n874), .B(n4731), .Z(n4729) );
  XOR U6274 ( .A(n4732), .B(n4733), .Z(n4731) );
  XOR U6275 ( .A(DB[260]), .B(DB[253]), .Z(n4733) );
  AND U6276 ( .A(n878), .B(n4734), .Z(n4732) );
  XOR U6277 ( .A(n4735), .B(n4736), .Z(n4734) );
  XOR U6278 ( .A(DB[253]), .B(DB[246]), .Z(n4736) );
  AND U6279 ( .A(n882), .B(n4737), .Z(n4735) );
  XOR U6280 ( .A(n4738), .B(n4739), .Z(n4737) );
  XOR U6281 ( .A(DB[246]), .B(DB[239]), .Z(n4739) );
  AND U6282 ( .A(n886), .B(n4740), .Z(n4738) );
  XOR U6283 ( .A(n4741), .B(n4742), .Z(n4740) );
  XOR U6284 ( .A(DB[239]), .B(DB[232]), .Z(n4742) );
  AND U6285 ( .A(n890), .B(n4743), .Z(n4741) );
  XOR U6286 ( .A(n4744), .B(n4745), .Z(n4743) );
  XOR U6287 ( .A(DB[232]), .B(DB[225]), .Z(n4745) );
  AND U6288 ( .A(n894), .B(n4746), .Z(n4744) );
  XOR U6289 ( .A(n4747), .B(n4748), .Z(n4746) );
  XOR U6290 ( .A(DB[225]), .B(DB[218]), .Z(n4748) );
  AND U6291 ( .A(n898), .B(n4749), .Z(n4747) );
  XOR U6292 ( .A(n4750), .B(n4751), .Z(n4749) );
  XOR U6293 ( .A(DB[218]), .B(DB[211]), .Z(n4751) );
  AND U6294 ( .A(n902), .B(n4752), .Z(n4750) );
  XOR U6295 ( .A(n4753), .B(n4754), .Z(n4752) );
  XOR U6296 ( .A(DB[211]), .B(DB[204]), .Z(n4754) );
  AND U6297 ( .A(n906), .B(n4755), .Z(n4753) );
  XOR U6298 ( .A(n4756), .B(n4757), .Z(n4755) );
  XOR U6299 ( .A(DB[204]), .B(DB[197]), .Z(n4757) );
  AND U6300 ( .A(n910), .B(n4758), .Z(n4756) );
  XOR U6301 ( .A(n4759), .B(n4760), .Z(n4758) );
  XOR U6302 ( .A(DB[197]), .B(DB[190]), .Z(n4760) );
  AND U6303 ( .A(n914), .B(n4761), .Z(n4759) );
  XOR U6304 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U6305 ( .A(DB[190]), .B(DB[183]), .Z(n4763) );
  AND U6306 ( .A(n918), .B(n4764), .Z(n4762) );
  XOR U6307 ( .A(n4765), .B(n4766), .Z(n4764) );
  XOR U6308 ( .A(DB[183]), .B(DB[176]), .Z(n4766) );
  AND U6309 ( .A(n922), .B(n4767), .Z(n4765) );
  XOR U6310 ( .A(n4768), .B(n4769), .Z(n4767) );
  XOR U6311 ( .A(DB[176]), .B(DB[169]), .Z(n4769) );
  AND U6312 ( .A(n926), .B(n4770), .Z(n4768) );
  XOR U6313 ( .A(n4771), .B(n4772), .Z(n4770) );
  XOR U6314 ( .A(DB[169]), .B(DB[162]), .Z(n4772) );
  AND U6315 ( .A(n930), .B(n4773), .Z(n4771) );
  XOR U6316 ( .A(n4774), .B(n4775), .Z(n4773) );
  XOR U6317 ( .A(DB[162]), .B(DB[155]), .Z(n4775) );
  AND U6318 ( .A(n934), .B(n4776), .Z(n4774) );
  XOR U6319 ( .A(n4777), .B(n4778), .Z(n4776) );
  XOR U6320 ( .A(DB[155]), .B(DB[148]), .Z(n4778) );
  AND U6321 ( .A(n938), .B(n4779), .Z(n4777) );
  XOR U6322 ( .A(n4780), .B(n4781), .Z(n4779) );
  XOR U6323 ( .A(DB[148]), .B(DB[141]), .Z(n4781) );
  AND U6324 ( .A(n942), .B(n4782), .Z(n4780) );
  XOR U6325 ( .A(n4783), .B(n4784), .Z(n4782) );
  XOR U6326 ( .A(DB[141]), .B(DB[134]), .Z(n4784) );
  AND U6327 ( .A(n946), .B(n4785), .Z(n4783) );
  XOR U6328 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U6329 ( .A(DB[134]), .B(DB[127]), .Z(n4787) );
  AND U6330 ( .A(n950), .B(n4788), .Z(n4786) );
  XOR U6331 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U6332 ( .A(DB[127]), .B(DB[120]), .Z(n4790) );
  AND U6333 ( .A(n954), .B(n4791), .Z(n4789) );
  XOR U6334 ( .A(n4792), .B(n4793), .Z(n4791) );
  XOR U6335 ( .A(DB[120]), .B(DB[113]), .Z(n4793) );
  AND U6336 ( .A(n958), .B(n4794), .Z(n4792) );
  XOR U6337 ( .A(n4795), .B(n4796), .Z(n4794) );
  XOR U6338 ( .A(DB[113]), .B(DB[106]), .Z(n4796) );
  AND U6339 ( .A(n962), .B(n4797), .Z(n4795) );
  XOR U6340 ( .A(n4798), .B(n4799), .Z(n4797) );
  XOR U6341 ( .A(DB[99]), .B(DB[106]), .Z(n4799) );
  AND U6342 ( .A(n966), .B(n4800), .Z(n4798) );
  XOR U6343 ( .A(n4801), .B(n4802), .Z(n4800) );
  XOR U6344 ( .A(DB[99]), .B(DB[92]), .Z(n4802) );
  AND U6345 ( .A(n970), .B(n4803), .Z(n4801) );
  XOR U6346 ( .A(n4804), .B(n4805), .Z(n4803) );
  XOR U6347 ( .A(DB[92]), .B(DB[85]), .Z(n4805) );
  AND U6348 ( .A(n974), .B(n4806), .Z(n4804) );
  XOR U6349 ( .A(n4807), .B(n4808), .Z(n4806) );
  XOR U6350 ( .A(DB[85]), .B(DB[78]), .Z(n4808) );
  AND U6351 ( .A(n978), .B(n4809), .Z(n4807) );
  XOR U6352 ( .A(n4810), .B(n4811), .Z(n4809) );
  XOR U6353 ( .A(DB[78]), .B(DB[71]), .Z(n4811) );
  AND U6354 ( .A(n982), .B(n4812), .Z(n4810) );
  XOR U6355 ( .A(n4813), .B(n4814), .Z(n4812) );
  XOR U6356 ( .A(DB[71]), .B(DB[64]), .Z(n4814) );
  AND U6357 ( .A(n986), .B(n4815), .Z(n4813) );
  XOR U6358 ( .A(n4816), .B(n4817), .Z(n4815) );
  XOR U6359 ( .A(DB[64]), .B(DB[57]), .Z(n4817) );
  AND U6360 ( .A(n990), .B(n4818), .Z(n4816) );
  XOR U6361 ( .A(n4819), .B(n4820), .Z(n4818) );
  XOR U6362 ( .A(DB[57]), .B(DB[50]), .Z(n4820) );
  AND U6363 ( .A(n994), .B(n4821), .Z(n4819) );
  XOR U6364 ( .A(n4822), .B(n4823), .Z(n4821) );
  XOR U6365 ( .A(DB[50]), .B(DB[43]), .Z(n4823) );
  AND U6366 ( .A(n998), .B(n4824), .Z(n4822) );
  XOR U6367 ( .A(n4825), .B(n4826), .Z(n4824) );
  XOR U6368 ( .A(DB[43]), .B(DB[36]), .Z(n4826) );
  AND U6369 ( .A(n1002), .B(n4827), .Z(n4825) );
  XOR U6370 ( .A(n4828), .B(n4829), .Z(n4827) );
  XOR U6371 ( .A(DB[36]), .B(DB[29]), .Z(n4829) );
  AND U6372 ( .A(n1006), .B(n4830), .Z(n4828) );
  XOR U6373 ( .A(n4831), .B(n4832), .Z(n4830) );
  XOR U6374 ( .A(DB[29]), .B(DB[22]), .Z(n4832) );
  AND U6375 ( .A(n1010), .B(n4833), .Z(n4831) );
  XOR U6376 ( .A(n4834), .B(n4835), .Z(n4833) );
  XOR U6377 ( .A(DB[22]), .B(DB[15]), .Z(n4835) );
  AND U6378 ( .A(n1014), .B(n4836), .Z(n4834) );
  XOR U6379 ( .A(n4837), .B(n4838), .Z(n4836) );
  XOR U6380 ( .A(DB[8]), .B(DB[15]), .Z(n4838) );
  AND U6381 ( .A(n1018), .B(n4839), .Z(n4837) );
  XOR U6382 ( .A(DB[8]), .B(DB[1]), .Z(n4839) );
  XOR U6383 ( .A(DB[1785]), .B(n4840), .Z(min_val_out[0]) );
  AND U6384 ( .A(n2), .B(n4841), .Z(n4840) );
  XOR U6385 ( .A(n4842), .B(n4843), .Z(n4841) );
  XOR U6386 ( .A(DB[1785]), .B(DB[1778]), .Z(n4843) );
  AND U6387 ( .A(n6), .B(n4844), .Z(n4842) );
  XOR U6388 ( .A(n4845), .B(n4846), .Z(n4844) );
  XOR U6389 ( .A(DB[1778]), .B(DB[1771]), .Z(n4846) );
  AND U6390 ( .A(n10), .B(n4847), .Z(n4845) );
  XOR U6391 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U6392 ( .A(DB[1771]), .B(DB[1764]), .Z(n4849) );
  AND U6393 ( .A(n14), .B(n4850), .Z(n4848) );
  XOR U6394 ( .A(n4851), .B(n4852), .Z(n4850) );
  XOR U6395 ( .A(DB[1764]), .B(DB[1757]), .Z(n4852) );
  AND U6396 ( .A(n18), .B(n4853), .Z(n4851) );
  XOR U6397 ( .A(n4854), .B(n4855), .Z(n4853) );
  XOR U6398 ( .A(DB[1757]), .B(DB[1750]), .Z(n4855) );
  AND U6399 ( .A(n22), .B(n4856), .Z(n4854) );
  XOR U6400 ( .A(n4857), .B(n4858), .Z(n4856) );
  XOR U6401 ( .A(DB[1750]), .B(DB[1743]), .Z(n4858) );
  AND U6402 ( .A(n26), .B(n4859), .Z(n4857) );
  XOR U6403 ( .A(n4860), .B(n4861), .Z(n4859) );
  XOR U6404 ( .A(DB[1743]), .B(DB[1736]), .Z(n4861) );
  AND U6405 ( .A(n30), .B(n4862), .Z(n4860) );
  XOR U6406 ( .A(n4863), .B(n4864), .Z(n4862) );
  XOR U6407 ( .A(DB[1736]), .B(DB[1729]), .Z(n4864) );
  AND U6408 ( .A(n34), .B(n4865), .Z(n4863) );
  XOR U6409 ( .A(n4866), .B(n4867), .Z(n4865) );
  XOR U6410 ( .A(DB[1729]), .B(DB[1722]), .Z(n4867) );
  AND U6411 ( .A(n38), .B(n4868), .Z(n4866) );
  XOR U6412 ( .A(n4869), .B(n4870), .Z(n4868) );
  XOR U6413 ( .A(DB[1722]), .B(DB[1715]), .Z(n4870) );
  AND U6414 ( .A(n42), .B(n4871), .Z(n4869) );
  XOR U6415 ( .A(n4872), .B(n4873), .Z(n4871) );
  XOR U6416 ( .A(DB[1715]), .B(DB[1708]), .Z(n4873) );
  AND U6417 ( .A(n46), .B(n4874), .Z(n4872) );
  XOR U6418 ( .A(n4875), .B(n4876), .Z(n4874) );
  XOR U6419 ( .A(DB[1708]), .B(DB[1701]), .Z(n4876) );
  AND U6420 ( .A(n50), .B(n4877), .Z(n4875) );
  XOR U6421 ( .A(n4878), .B(n4879), .Z(n4877) );
  XOR U6422 ( .A(DB[1701]), .B(DB[1694]), .Z(n4879) );
  AND U6423 ( .A(n54), .B(n4880), .Z(n4878) );
  XOR U6424 ( .A(n4881), .B(n4882), .Z(n4880) );
  XOR U6425 ( .A(DB[1694]), .B(DB[1687]), .Z(n4882) );
  AND U6426 ( .A(n58), .B(n4883), .Z(n4881) );
  XOR U6427 ( .A(n4884), .B(n4885), .Z(n4883) );
  XOR U6428 ( .A(DB[1687]), .B(DB[1680]), .Z(n4885) );
  AND U6429 ( .A(n62), .B(n4886), .Z(n4884) );
  XOR U6430 ( .A(n4887), .B(n4888), .Z(n4886) );
  XOR U6431 ( .A(DB[1680]), .B(DB[1673]), .Z(n4888) );
  AND U6432 ( .A(n66), .B(n4889), .Z(n4887) );
  XOR U6433 ( .A(n4890), .B(n4891), .Z(n4889) );
  XOR U6434 ( .A(DB[1673]), .B(DB[1666]), .Z(n4891) );
  AND U6435 ( .A(n70), .B(n4892), .Z(n4890) );
  XOR U6436 ( .A(n4893), .B(n4894), .Z(n4892) );
  XOR U6437 ( .A(DB[1666]), .B(DB[1659]), .Z(n4894) );
  AND U6438 ( .A(n74), .B(n4895), .Z(n4893) );
  XOR U6439 ( .A(n4896), .B(n4897), .Z(n4895) );
  XOR U6440 ( .A(DB[1659]), .B(DB[1652]), .Z(n4897) );
  AND U6441 ( .A(n78), .B(n4898), .Z(n4896) );
  XOR U6442 ( .A(n4899), .B(n4900), .Z(n4898) );
  XOR U6443 ( .A(DB[1652]), .B(DB[1645]), .Z(n4900) );
  AND U6444 ( .A(n82), .B(n4901), .Z(n4899) );
  XOR U6445 ( .A(n4902), .B(n4903), .Z(n4901) );
  XOR U6446 ( .A(DB[1645]), .B(DB[1638]), .Z(n4903) );
  AND U6447 ( .A(n86), .B(n4904), .Z(n4902) );
  XOR U6448 ( .A(n4905), .B(n4906), .Z(n4904) );
  XOR U6449 ( .A(DB[1638]), .B(DB[1631]), .Z(n4906) );
  AND U6450 ( .A(n90), .B(n4907), .Z(n4905) );
  XOR U6451 ( .A(n4908), .B(n4909), .Z(n4907) );
  XOR U6452 ( .A(DB[1631]), .B(DB[1624]), .Z(n4909) );
  AND U6453 ( .A(n94), .B(n4910), .Z(n4908) );
  XOR U6454 ( .A(n4911), .B(n4912), .Z(n4910) );
  XOR U6455 ( .A(DB[1624]), .B(DB[1617]), .Z(n4912) );
  AND U6456 ( .A(n98), .B(n4913), .Z(n4911) );
  XOR U6457 ( .A(n4914), .B(n4915), .Z(n4913) );
  XOR U6458 ( .A(DB[1617]), .B(DB[1610]), .Z(n4915) );
  AND U6459 ( .A(n102), .B(n4916), .Z(n4914) );
  XOR U6460 ( .A(n4917), .B(n4918), .Z(n4916) );
  XOR U6461 ( .A(DB[1610]), .B(DB[1603]), .Z(n4918) );
  AND U6462 ( .A(n106), .B(n4919), .Z(n4917) );
  XOR U6463 ( .A(n4920), .B(n4921), .Z(n4919) );
  XOR U6464 ( .A(DB[1603]), .B(DB[1596]), .Z(n4921) );
  AND U6465 ( .A(n110), .B(n4922), .Z(n4920) );
  XOR U6466 ( .A(n4923), .B(n4924), .Z(n4922) );
  XOR U6467 ( .A(DB[1596]), .B(DB[1589]), .Z(n4924) );
  AND U6468 ( .A(n114), .B(n4925), .Z(n4923) );
  XOR U6469 ( .A(n4926), .B(n4927), .Z(n4925) );
  XOR U6470 ( .A(DB[1589]), .B(DB[1582]), .Z(n4927) );
  AND U6471 ( .A(n118), .B(n4928), .Z(n4926) );
  XOR U6472 ( .A(n4929), .B(n4930), .Z(n4928) );
  XOR U6473 ( .A(DB[1582]), .B(DB[1575]), .Z(n4930) );
  AND U6474 ( .A(n122), .B(n4931), .Z(n4929) );
  XOR U6475 ( .A(n4932), .B(n4933), .Z(n4931) );
  XOR U6476 ( .A(DB[1575]), .B(DB[1568]), .Z(n4933) );
  AND U6477 ( .A(n126), .B(n4934), .Z(n4932) );
  XOR U6478 ( .A(n4935), .B(n4936), .Z(n4934) );
  XOR U6479 ( .A(DB[1568]), .B(DB[1561]), .Z(n4936) );
  AND U6480 ( .A(n130), .B(n4937), .Z(n4935) );
  XOR U6481 ( .A(n4938), .B(n4939), .Z(n4937) );
  XOR U6482 ( .A(DB[1561]), .B(DB[1554]), .Z(n4939) );
  AND U6483 ( .A(n134), .B(n4940), .Z(n4938) );
  XOR U6484 ( .A(n4941), .B(n4942), .Z(n4940) );
  XOR U6485 ( .A(DB[1554]), .B(DB[1547]), .Z(n4942) );
  AND U6486 ( .A(n138), .B(n4943), .Z(n4941) );
  XOR U6487 ( .A(n4944), .B(n4945), .Z(n4943) );
  XOR U6488 ( .A(DB[1547]), .B(DB[1540]), .Z(n4945) );
  AND U6489 ( .A(n142), .B(n4946), .Z(n4944) );
  XOR U6490 ( .A(n4947), .B(n4948), .Z(n4946) );
  XOR U6491 ( .A(DB[1540]), .B(DB[1533]), .Z(n4948) );
  AND U6492 ( .A(n146), .B(n4949), .Z(n4947) );
  XOR U6493 ( .A(n4950), .B(n4951), .Z(n4949) );
  XOR U6494 ( .A(DB[1533]), .B(DB[1526]), .Z(n4951) );
  AND U6495 ( .A(n150), .B(n4952), .Z(n4950) );
  XOR U6496 ( .A(n4953), .B(n4954), .Z(n4952) );
  XOR U6497 ( .A(DB[1526]), .B(DB[1519]), .Z(n4954) );
  AND U6498 ( .A(n154), .B(n4955), .Z(n4953) );
  XOR U6499 ( .A(n4956), .B(n4957), .Z(n4955) );
  XOR U6500 ( .A(DB[1519]), .B(DB[1512]), .Z(n4957) );
  AND U6501 ( .A(n158), .B(n4958), .Z(n4956) );
  XOR U6502 ( .A(n4959), .B(n4960), .Z(n4958) );
  XOR U6503 ( .A(DB[1512]), .B(DB[1505]), .Z(n4960) );
  AND U6504 ( .A(n162), .B(n4961), .Z(n4959) );
  XOR U6505 ( .A(n4962), .B(n4963), .Z(n4961) );
  XOR U6506 ( .A(DB[1505]), .B(DB[1498]), .Z(n4963) );
  AND U6507 ( .A(n166), .B(n4964), .Z(n4962) );
  XOR U6508 ( .A(n4965), .B(n4966), .Z(n4964) );
  XOR U6509 ( .A(DB[1498]), .B(DB[1491]), .Z(n4966) );
  AND U6510 ( .A(n170), .B(n4967), .Z(n4965) );
  XOR U6511 ( .A(n4968), .B(n4969), .Z(n4967) );
  XOR U6512 ( .A(DB[1491]), .B(DB[1484]), .Z(n4969) );
  AND U6513 ( .A(n174), .B(n4970), .Z(n4968) );
  XOR U6514 ( .A(n4971), .B(n4972), .Z(n4970) );
  XOR U6515 ( .A(DB[1484]), .B(DB[1477]), .Z(n4972) );
  AND U6516 ( .A(n178), .B(n4973), .Z(n4971) );
  XOR U6517 ( .A(n4974), .B(n4975), .Z(n4973) );
  XOR U6518 ( .A(DB[1477]), .B(DB[1470]), .Z(n4975) );
  AND U6519 ( .A(n182), .B(n4976), .Z(n4974) );
  XOR U6520 ( .A(n4977), .B(n4978), .Z(n4976) );
  XOR U6521 ( .A(DB[1470]), .B(DB[1463]), .Z(n4978) );
  AND U6522 ( .A(n186), .B(n4979), .Z(n4977) );
  XOR U6523 ( .A(n4980), .B(n4981), .Z(n4979) );
  XOR U6524 ( .A(DB[1463]), .B(DB[1456]), .Z(n4981) );
  AND U6525 ( .A(n190), .B(n4982), .Z(n4980) );
  XOR U6526 ( .A(n4983), .B(n4984), .Z(n4982) );
  XOR U6527 ( .A(DB[1456]), .B(DB[1449]), .Z(n4984) );
  AND U6528 ( .A(n194), .B(n4985), .Z(n4983) );
  XOR U6529 ( .A(n4986), .B(n4987), .Z(n4985) );
  XOR U6530 ( .A(DB[1449]), .B(DB[1442]), .Z(n4987) );
  AND U6531 ( .A(n198), .B(n4988), .Z(n4986) );
  XOR U6532 ( .A(n4989), .B(n4990), .Z(n4988) );
  XOR U6533 ( .A(DB[1442]), .B(DB[1435]), .Z(n4990) );
  AND U6534 ( .A(n202), .B(n4991), .Z(n4989) );
  XOR U6535 ( .A(n4992), .B(n4993), .Z(n4991) );
  XOR U6536 ( .A(DB[1435]), .B(DB[1428]), .Z(n4993) );
  AND U6537 ( .A(n206), .B(n4994), .Z(n4992) );
  XOR U6538 ( .A(n4995), .B(n4996), .Z(n4994) );
  XOR U6539 ( .A(DB[1428]), .B(DB[1421]), .Z(n4996) );
  AND U6540 ( .A(n210), .B(n4997), .Z(n4995) );
  XOR U6541 ( .A(n4998), .B(n4999), .Z(n4997) );
  XOR U6542 ( .A(DB[1421]), .B(DB[1414]), .Z(n4999) );
  AND U6543 ( .A(n214), .B(n5000), .Z(n4998) );
  XOR U6544 ( .A(n5001), .B(n5002), .Z(n5000) );
  XOR U6545 ( .A(DB[1414]), .B(DB[1407]), .Z(n5002) );
  AND U6546 ( .A(n218), .B(n5003), .Z(n5001) );
  XOR U6547 ( .A(n5004), .B(n5005), .Z(n5003) );
  XOR U6548 ( .A(DB[1407]), .B(DB[1400]), .Z(n5005) );
  AND U6549 ( .A(n222), .B(n5006), .Z(n5004) );
  XOR U6550 ( .A(n5007), .B(n5008), .Z(n5006) );
  XOR U6551 ( .A(DB[1400]), .B(DB[1393]), .Z(n5008) );
  AND U6552 ( .A(n226), .B(n5009), .Z(n5007) );
  XOR U6553 ( .A(n5010), .B(n5011), .Z(n5009) );
  XOR U6554 ( .A(DB[1393]), .B(DB[1386]), .Z(n5011) );
  AND U6555 ( .A(n230), .B(n5012), .Z(n5010) );
  XOR U6556 ( .A(n5013), .B(n5014), .Z(n5012) );
  XOR U6557 ( .A(DB[1386]), .B(DB[1379]), .Z(n5014) );
  AND U6558 ( .A(n234), .B(n5015), .Z(n5013) );
  XOR U6559 ( .A(n5016), .B(n5017), .Z(n5015) );
  XOR U6560 ( .A(DB[1379]), .B(DB[1372]), .Z(n5017) );
  AND U6561 ( .A(n238), .B(n5018), .Z(n5016) );
  XOR U6562 ( .A(n5019), .B(n5020), .Z(n5018) );
  XOR U6563 ( .A(DB[1372]), .B(DB[1365]), .Z(n5020) );
  AND U6564 ( .A(n242), .B(n5021), .Z(n5019) );
  XOR U6565 ( .A(n5022), .B(n5023), .Z(n5021) );
  XOR U6566 ( .A(DB[1365]), .B(DB[1358]), .Z(n5023) );
  AND U6567 ( .A(n246), .B(n5024), .Z(n5022) );
  XOR U6568 ( .A(n5025), .B(n5026), .Z(n5024) );
  XOR U6569 ( .A(DB[1358]), .B(DB[1351]), .Z(n5026) );
  AND U6570 ( .A(n250), .B(n5027), .Z(n5025) );
  XOR U6571 ( .A(n5028), .B(n5029), .Z(n5027) );
  XOR U6572 ( .A(DB[1351]), .B(DB[1344]), .Z(n5029) );
  AND U6573 ( .A(n254), .B(n5030), .Z(n5028) );
  XOR U6574 ( .A(n5031), .B(n5032), .Z(n5030) );
  XOR U6575 ( .A(DB[1344]), .B(DB[1337]), .Z(n5032) );
  AND U6576 ( .A(n258), .B(n5033), .Z(n5031) );
  XOR U6577 ( .A(n5034), .B(n5035), .Z(n5033) );
  XOR U6578 ( .A(DB[1337]), .B(DB[1330]), .Z(n5035) );
  AND U6579 ( .A(n262), .B(n5036), .Z(n5034) );
  XOR U6580 ( .A(n5037), .B(n5038), .Z(n5036) );
  XOR U6581 ( .A(DB[1330]), .B(DB[1323]), .Z(n5038) );
  AND U6582 ( .A(n266), .B(n5039), .Z(n5037) );
  XOR U6583 ( .A(n5040), .B(n5041), .Z(n5039) );
  XOR U6584 ( .A(DB[1323]), .B(DB[1316]), .Z(n5041) );
  AND U6585 ( .A(n270), .B(n5042), .Z(n5040) );
  XOR U6586 ( .A(n5043), .B(n5044), .Z(n5042) );
  XOR U6587 ( .A(DB[1316]), .B(DB[1309]), .Z(n5044) );
  AND U6588 ( .A(n274), .B(n5045), .Z(n5043) );
  XOR U6589 ( .A(n5046), .B(n5047), .Z(n5045) );
  XOR U6590 ( .A(DB[1309]), .B(DB[1302]), .Z(n5047) );
  AND U6591 ( .A(n278), .B(n5048), .Z(n5046) );
  XOR U6592 ( .A(n5049), .B(n5050), .Z(n5048) );
  XOR U6593 ( .A(DB[1302]), .B(DB[1295]), .Z(n5050) );
  AND U6594 ( .A(n282), .B(n5051), .Z(n5049) );
  XOR U6595 ( .A(n5052), .B(n5053), .Z(n5051) );
  XOR U6596 ( .A(DB[1295]), .B(DB[1288]), .Z(n5053) );
  AND U6597 ( .A(n286), .B(n5054), .Z(n5052) );
  XOR U6598 ( .A(n5055), .B(n5056), .Z(n5054) );
  XOR U6599 ( .A(DB[1288]), .B(DB[1281]), .Z(n5056) );
  AND U6600 ( .A(n290), .B(n5057), .Z(n5055) );
  XOR U6601 ( .A(n5058), .B(n5059), .Z(n5057) );
  XOR U6602 ( .A(DB[1281]), .B(DB[1274]), .Z(n5059) );
  AND U6603 ( .A(n294), .B(n5060), .Z(n5058) );
  XOR U6604 ( .A(n5061), .B(n5062), .Z(n5060) );
  XOR U6605 ( .A(DB[1274]), .B(DB[1267]), .Z(n5062) );
  AND U6606 ( .A(n298), .B(n5063), .Z(n5061) );
  XOR U6607 ( .A(n5064), .B(n5065), .Z(n5063) );
  XOR U6608 ( .A(DB[1267]), .B(DB[1260]), .Z(n5065) );
  AND U6609 ( .A(n302), .B(n5066), .Z(n5064) );
  XOR U6610 ( .A(n5067), .B(n5068), .Z(n5066) );
  XOR U6611 ( .A(DB[1260]), .B(DB[1253]), .Z(n5068) );
  AND U6612 ( .A(n306), .B(n5069), .Z(n5067) );
  XOR U6613 ( .A(n5070), .B(n5071), .Z(n5069) );
  XOR U6614 ( .A(DB[1253]), .B(DB[1246]), .Z(n5071) );
  AND U6615 ( .A(n310), .B(n5072), .Z(n5070) );
  XOR U6616 ( .A(n5073), .B(n5074), .Z(n5072) );
  XOR U6617 ( .A(DB[1246]), .B(DB[1239]), .Z(n5074) );
  AND U6618 ( .A(n314), .B(n5075), .Z(n5073) );
  XOR U6619 ( .A(n5076), .B(n5077), .Z(n5075) );
  XOR U6620 ( .A(DB[1239]), .B(DB[1232]), .Z(n5077) );
  AND U6621 ( .A(n318), .B(n5078), .Z(n5076) );
  XOR U6622 ( .A(n5079), .B(n5080), .Z(n5078) );
  XOR U6623 ( .A(DB[1232]), .B(DB[1225]), .Z(n5080) );
  AND U6624 ( .A(n322), .B(n5081), .Z(n5079) );
  XOR U6625 ( .A(n5082), .B(n5083), .Z(n5081) );
  XOR U6626 ( .A(DB[1225]), .B(DB[1218]), .Z(n5083) );
  AND U6627 ( .A(n326), .B(n5084), .Z(n5082) );
  XOR U6628 ( .A(n5085), .B(n5086), .Z(n5084) );
  XOR U6629 ( .A(DB[1218]), .B(DB[1211]), .Z(n5086) );
  AND U6630 ( .A(n330), .B(n5087), .Z(n5085) );
  XOR U6631 ( .A(n5088), .B(n5089), .Z(n5087) );
  XOR U6632 ( .A(DB[1211]), .B(DB[1204]), .Z(n5089) );
  AND U6633 ( .A(n334), .B(n5090), .Z(n5088) );
  XOR U6634 ( .A(n5091), .B(n5092), .Z(n5090) );
  XOR U6635 ( .A(DB[1204]), .B(DB[1197]), .Z(n5092) );
  AND U6636 ( .A(n338), .B(n5093), .Z(n5091) );
  XOR U6637 ( .A(n5094), .B(n5095), .Z(n5093) );
  XOR U6638 ( .A(DB[1197]), .B(DB[1190]), .Z(n5095) );
  AND U6639 ( .A(n342), .B(n5096), .Z(n5094) );
  XOR U6640 ( .A(n5097), .B(n5098), .Z(n5096) );
  XOR U6641 ( .A(DB[1190]), .B(DB[1183]), .Z(n5098) );
  AND U6642 ( .A(n346), .B(n5099), .Z(n5097) );
  XOR U6643 ( .A(n5100), .B(n5101), .Z(n5099) );
  XOR U6644 ( .A(DB[1183]), .B(DB[1176]), .Z(n5101) );
  AND U6645 ( .A(n350), .B(n5102), .Z(n5100) );
  XOR U6646 ( .A(n5103), .B(n5104), .Z(n5102) );
  XOR U6647 ( .A(DB[1176]), .B(DB[1169]), .Z(n5104) );
  AND U6648 ( .A(n354), .B(n5105), .Z(n5103) );
  XOR U6649 ( .A(n5106), .B(n5107), .Z(n5105) );
  XOR U6650 ( .A(DB[1169]), .B(DB[1162]), .Z(n5107) );
  AND U6651 ( .A(n358), .B(n5108), .Z(n5106) );
  XOR U6652 ( .A(n5109), .B(n5110), .Z(n5108) );
  XOR U6653 ( .A(DB[1162]), .B(DB[1155]), .Z(n5110) );
  AND U6654 ( .A(n362), .B(n5111), .Z(n5109) );
  XOR U6655 ( .A(n5112), .B(n5113), .Z(n5111) );
  XOR U6656 ( .A(DB[1155]), .B(DB[1148]), .Z(n5113) );
  AND U6657 ( .A(n366), .B(n5114), .Z(n5112) );
  XOR U6658 ( .A(n5115), .B(n5116), .Z(n5114) );
  XOR U6659 ( .A(DB[1148]), .B(DB[1141]), .Z(n5116) );
  AND U6660 ( .A(n370), .B(n5117), .Z(n5115) );
  XOR U6661 ( .A(n5118), .B(n5119), .Z(n5117) );
  XOR U6662 ( .A(DB[1141]), .B(DB[1134]), .Z(n5119) );
  AND U6663 ( .A(n374), .B(n5120), .Z(n5118) );
  XOR U6664 ( .A(n5121), .B(n5122), .Z(n5120) );
  XOR U6665 ( .A(DB[1134]), .B(DB[1127]), .Z(n5122) );
  AND U6666 ( .A(n378), .B(n5123), .Z(n5121) );
  XOR U6667 ( .A(n5124), .B(n5125), .Z(n5123) );
  XOR U6668 ( .A(DB[1127]), .B(DB[1120]), .Z(n5125) );
  AND U6669 ( .A(n382), .B(n5126), .Z(n5124) );
  XOR U6670 ( .A(n5127), .B(n5128), .Z(n5126) );
  XOR U6671 ( .A(DB[1120]), .B(DB[1113]), .Z(n5128) );
  AND U6672 ( .A(n386), .B(n5129), .Z(n5127) );
  XOR U6673 ( .A(n5130), .B(n5131), .Z(n5129) );
  XOR U6674 ( .A(DB[1113]), .B(DB[1106]), .Z(n5131) );
  AND U6675 ( .A(n390), .B(n5132), .Z(n5130) );
  XOR U6676 ( .A(n5133), .B(n5134), .Z(n5132) );
  XOR U6677 ( .A(DB[1106]), .B(DB[1099]), .Z(n5134) );
  AND U6678 ( .A(n394), .B(n5135), .Z(n5133) );
  XOR U6679 ( .A(n5136), .B(n5137), .Z(n5135) );
  XOR U6680 ( .A(DB[1099]), .B(DB[1092]), .Z(n5137) );
  AND U6681 ( .A(n398), .B(n5138), .Z(n5136) );
  XOR U6682 ( .A(n5139), .B(n5140), .Z(n5138) );
  XOR U6683 ( .A(DB[1092]), .B(DB[1085]), .Z(n5140) );
  AND U6684 ( .A(n402), .B(n5141), .Z(n5139) );
  XOR U6685 ( .A(n5142), .B(n5143), .Z(n5141) );
  XOR U6686 ( .A(DB[1085]), .B(DB[1078]), .Z(n5143) );
  AND U6687 ( .A(n406), .B(n5144), .Z(n5142) );
  XOR U6688 ( .A(n5145), .B(n5146), .Z(n5144) );
  XOR U6689 ( .A(DB[1078]), .B(DB[1071]), .Z(n5146) );
  AND U6690 ( .A(n410), .B(n5147), .Z(n5145) );
  XOR U6691 ( .A(n5148), .B(n5149), .Z(n5147) );
  XOR U6692 ( .A(DB[1071]), .B(DB[1064]), .Z(n5149) );
  AND U6693 ( .A(n414), .B(n5150), .Z(n5148) );
  XOR U6694 ( .A(n5151), .B(n5152), .Z(n5150) );
  XOR U6695 ( .A(DB[1064]), .B(DB[1057]), .Z(n5152) );
  AND U6696 ( .A(n418), .B(n5153), .Z(n5151) );
  XOR U6697 ( .A(n5154), .B(n5155), .Z(n5153) );
  XOR U6698 ( .A(DB[1057]), .B(DB[1050]), .Z(n5155) );
  AND U6699 ( .A(n422), .B(n5156), .Z(n5154) );
  XOR U6700 ( .A(n5157), .B(n5158), .Z(n5156) );
  XOR U6701 ( .A(DB[1050]), .B(DB[1043]), .Z(n5158) );
  AND U6702 ( .A(n426), .B(n5159), .Z(n5157) );
  XOR U6703 ( .A(n5160), .B(n5161), .Z(n5159) );
  XOR U6704 ( .A(DB[1043]), .B(DB[1036]), .Z(n5161) );
  AND U6705 ( .A(n430), .B(n5162), .Z(n5160) );
  XOR U6706 ( .A(n5163), .B(n5164), .Z(n5162) );
  XOR U6707 ( .A(DB[1036]), .B(DB[1029]), .Z(n5164) );
  AND U6708 ( .A(n434), .B(n5165), .Z(n5163) );
  XOR U6709 ( .A(n5166), .B(n5167), .Z(n5165) );
  XOR U6710 ( .A(DB[1029]), .B(DB[1022]), .Z(n5167) );
  AND U6711 ( .A(n438), .B(n5168), .Z(n5166) );
  XOR U6712 ( .A(n5169), .B(n5170), .Z(n5168) );
  XOR U6713 ( .A(DB[1022]), .B(DB[1015]), .Z(n5170) );
  AND U6714 ( .A(n442), .B(n5171), .Z(n5169) );
  XOR U6715 ( .A(n5172), .B(n5173), .Z(n5171) );
  XOR U6716 ( .A(DB[1015]), .B(DB[1008]), .Z(n5173) );
  AND U6717 ( .A(n446), .B(n5174), .Z(n5172) );
  XOR U6718 ( .A(n5175), .B(n5176), .Z(n5174) );
  XOR U6719 ( .A(DB[1008]), .B(DB[1001]), .Z(n5176) );
  AND U6720 ( .A(n450), .B(n5177), .Z(n5175) );
  XOR U6721 ( .A(n5178), .B(n5179), .Z(n5177) );
  XOR U6722 ( .A(DB[994]), .B(DB[1001]), .Z(n5179) );
  AND U6723 ( .A(n454), .B(n5180), .Z(n5178) );
  XOR U6724 ( .A(n5181), .B(n5182), .Z(n5180) );
  XOR U6725 ( .A(DB[994]), .B(DB[987]), .Z(n5182) );
  AND U6726 ( .A(n458), .B(n5183), .Z(n5181) );
  XOR U6727 ( .A(n5184), .B(n5185), .Z(n5183) );
  XOR U6728 ( .A(DB[987]), .B(DB[980]), .Z(n5185) );
  AND U6729 ( .A(n462), .B(n5186), .Z(n5184) );
  XOR U6730 ( .A(n5187), .B(n5188), .Z(n5186) );
  XOR U6731 ( .A(DB[980]), .B(DB[973]), .Z(n5188) );
  AND U6732 ( .A(n466), .B(n5189), .Z(n5187) );
  XOR U6733 ( .A(n5190), .B(n5191), .Z(n5189) );
  XOR U6734 ( .A(DB[973]), .B(DB[966]), .Z(n5191) );
  AND U6735 ( .A(n470), .B(n5192), .Z(n5190) );
  XOR U6736 ( .A(n5193), .B(n5194), .Z(n5192) );
  XOR U6737 ( .A(DB[966]), .B(DB[959]), .Z(n5194) );
  AND U6738 ( .A(n474), .B(n5195), .Z(n5193) );
  XOR U6739 ( .A(n5196), .B(n5197), .Z(n5195) );
  XOR U6740 ( .A(DB[959]), .B(DB[952]), .Z(n5197) );
  AND U6741 ( .A(n478), .B(n5198), .Z(n5196) );
  XOR U6742 ( .A(n5199), .B(n5200), .Z(n5198) );
  XOR U6743 ( .A(DB[952]), .B(DB[945]), .Z(n5200) );
  AND U6744 ( .A(n482), .B(n5201), .Z(n5199) );
  XOR U6745 ( .A(n5202), .B(n5203), .Z(n5201) );
  XOR U6746 ( .A(DB[945]), .B(DB[938]), .Z(n5203) );
  AND U6747 ( .A(n486), .B(n5204), .Z(n5202) );
  XOR U6748 ( .A(n5205), .B(n5206), .Z(n5204) );
  XOR U6749 ( .A(DB[938]), .B(DB[931]), .Z(n5206) );
  AND U6750 ( .A(n490), .B(n5207), .Z(n5205) );
  XOR U6751 ( .A(n5208), .B(n5209), .Z(n5207) );
  XOR U6752 ( .A(DB[931]), .B(DB[924]), .Z(n5209) );
  AND U6753 ( .A(n494), .B(n5210), .Z(n5208) );
  XOR U6754 ( .A(n5211), .B(n5212), .Z(n5210) );
  XOR U6755 ( .A(DB[924]), .B(DB[917]), .Z(n5212) );
  AND U6756 ( .A(n498), .B(n5213), .Z(n5211) );
  XOR U6757 ( .A(n5214), .B(n5215), .Z(n5213) );
  XOR U6758 ( .A(DB[917]), .B(DB[910]), .Z(n5215) );
  AND U6759 ( .A(n502), .B(n5216), .Z(n5214) );
  XOR U6760 ( .A(n5217), .B(n5218), .Z(n5216) );
  XOR U6761 ( .A(DB[910]), .B(DB[903]), .Z(n5218) );
  AND U6762 ( .A(n506), .B(n5219), .Z(n5217) );
  XOR U6763 ( .A(n5220), .B(n5221), .Z(n5219) );
  XOR U6764 ( .A(DB[903]), .B(DB[896]), .Z(n5221) );
  AND U6765 ( .A(n510), .B(n5222), .Z(n5220) );
  XOR U6766 ( .A(n5223), .B(n5224), .Z(n5222) );
  XOR U6767 ( .A(DB[896]), .B(DB[889]), .Z(n5224) );
  AND U6768 ( .A(n514), .B(n5225), .Z(n5223) );
  XOR U6769 ( .A(n5226), .B(n5227), .Z(n5225) );
  XOR U6770 ( .A(DB[889]), .B(DB[882]), .Z(n5227) );
  AND U6771 ( .A(n518), .B(n5228), .Z(n5226) );
  XOR U6772 ( .A(n5229), .B(n5230), .Z(n5228) );
  XOR U6773 ( .A(DB[882]), .B(DB[875]), .Z(n5230) );
  AND U6774 ( .A(n522), .B(n5231), .Z(n5229) );
  XOR U6775 ( .A(n5232), .B(n5233), .Z(n5231) );
  XOR U6776 ( .A(DB[875]), .B(DB[868]), .Z(n5233) );
  AND U6777 ( .A(n526), .B(n5234), .Z(n5232) );
  XOR U6778 ( .A(n5235), .B(n5236), .Z(n5234) );
  XOR U6779 ( .A(DB[868]), .B(DB[861]), .Z(n5236) );
  AND U6780 ( .A(n530), .B(n5237), .Z(n5235) );
  XOR U6781 ( .A(n5238), .B(n5239), .Z(n5237) );
  XOR U6782 ( .A(DB[861]), .B(DB[854]), .Z(n5239) );
  AND U6783 ( .A(n534), .B(n5240), .Z(n5238) );
  XOR U6784 ( .A(n5241), .B(n5242), .Z(n5240) );
  XOR U6785 ( .A(DB[854]), .B(DB[847]), .Z(n5242) );
  AND U6786 ( .A(n538), .B(n5243), .Z(n5241) );
  XOR U6787 ( .A(n5244), .B(n5245), .Z(n5243) );
  XOR U6788 ( .A(DB[847]), .B(DB[840]), .Z(n5245) );
  AND U6789 ( .A(n542), .B(n5246), .Z(n5244) );
  XOR U6790 ( .A(n5247), .B(n5248), .Z(n5246) );
  XOR U6791 ( .A(DB[840]), .B(DB[833]), .Z(n5248) );
  AND U6792 ( .A(n546), .B(n5249), .Z(n5247) );
  XOR U6793 ( .A(n5250), .B(n5251), .Z(n5249) );
  XOR U6794 ( .A(DB[833]), .B(DB[826]), .Z(n5251) );
  AND U6795 ( .A(n550), .B(n5252), .Z(n5250) );
  XOR U6796 ( .A(n5253), .B(n5254), .Z(n5252) );
  XOR U6797 ( .A(DB[826]), .B(DB[819]), .Z(n5254) );
  AND U6798 ( .A(n554), .B(n5255), .Z(n5253) );
  XOR U6799 ( .A(n5256), .B(n5257), .Z(n5255) );
  XOR U6800 ( .A(DB[819]), .B(DB[812]), .Z(n5257) );
  AND U6801 ( .A(n558), .B(n5258), .Z(n5256) );
  XOR U6802 ( .A(n5259), .B(n5260), .Z(n5258) );
  XOR U6803 ( .A(DB[812]), .B(DB[805]), .Z(n5260) );
  AND U6804 ( .A(n562), .B(n5261), .Z(n5259) );
  XOR U6805 ( .A(n5262), .B(n5263), .Z(n5261) );
  XOR U6806 ( .A(DB[805]), .B(DB[798]), .Z(n5263) );
  AND U6807 ( .A(n566), .B(n5264), .Z(n5262) );
  XOR U6808 ( .A(n5265), .B(n5266), .Z(n5264) );
  XOR U6809 ( .A(DB[798]), .B(DB[791]), .Z(n5266) );
  AND U6810 ( .A(n570), .B(n5267), .Z(n5265) );
  XOR U6811 ( .A(n5268), .B(n5269), .Z(n5267) );
  XOR U6812 ( .A(DB[791]), .B(DB[784]), .Z(n5269) );
  AND U6813 ( .A(n574), .B(n5270), .Z(n5268) );
  XOR U6814 ( .A(n5271), .B(n5272), .Z(n5270) );
  XOR U6815 ( .A(DB[784]), .B(DB[777]), .Z(n5272) );
  AND U6816 ( .A(n578), .B(n5273), .Z(n5271) );
  XOR U6817 ( .A(n5274), .B(n5275), .Z(n5273) );
  XOR U6818 ( .A(DB[777]), .B(DB[770]), .Z(n5275) );
  AND U6819 ( .A(n582), .B(n5276), .Z(n5274) );
  XOR U6820 ( .A(n5277), .B(n5278), .Z(n5276) );
  XOR U6821 ( .A(DB[770]), .B(DB[763]), .Z(n5278) );
  AND U6822 ( .A(n586), .B(n5279), .Z(n5277) );
  XOR U6823 ( .A(n5280), .B(n5281), .Z(n5279) );
  XOR U6824 ( .A(DB[763]), .B(DB[756]), .Z(n5281) );
  AND U6825 ( .A(n590), .B(n5282), .Z(n5280) );
  XOR U6826 ( .A(n5283), .B(n5284), .Z(n5282) );
  XOR U6827 ( .A(DB[756]), .B(DB[749]), .Z(n5284) );
  AND U6828 ( .A(n594), .B(n5285), .Z(n5283) );
  XOR U6829 ( .A(n5286), .B(n5287), .Z(n5285) );
  XOR U6830 ( .A(DB[749]), .B(DB[742]), .Z(n5287) );
  AND U6831 ( .A(n598), .B(n5288), .Z(n5286) );
  XOR U6832 ( .A(n5289), .B(n5290), .Z(n5288) );
  XOR U6833 ( .A(DB[742]), .B(DB[735]), .Z(n5290) );
  AND U6834 ( .A(n602), .B(n5291), .Z(n5289) );
  XOR U6835 ( .A(n5292), .B(n5293), .Z(n5291) );
  XOR U6836 ( .A(DB[735]), .B(DB[728]), .Z(n5293) );
  AND U6837 ( .A(n606), .B(n5294), .Z(n5292) );
  XOR U6838 ( .A(n5295), .B(n5296), .Z(n5294) );
  XOR U6839 ( .A(DB[728]), .B(DB[721]), .Z(n5296) );
  AND U6840 ( .A(n610), .B(n5297), .Z(n5295) );
  XOR U6841 ( .A(n5298), .B(n5299), .Z(n5297) );
  XOR U6842 ( .A(DB[721]), .B(DB[714]), .Z(n5299) );
  AND U6843 ( .A(n614), .B(n5300), .Z(n5298) );
  XOR U6844 ( .A(n5301), .B(n5302), .Z(n5300) );
  XOR U6845 ( .A(DB[714]), .B(DB[707]), .Z(n5302) );
  AND U6846 ( .A(n618), .B(n5303), .Z(n5301) );
  XOR U6847 ( .A(n5304), .B(n5305), .Z(n5303) );
  XOR U6848 ( .A(DB[707]), .B(DB[700]), .Z(n5305) );
  AND U6849 ( .A(n622), .B(n5306), .Z(n5304) );
  XOR U6850 ( .A(n5307), .B(n5308), .Z(n5306) );
  XOR U6851 ( .A(DB[700]), .B(DB[693]), .Z(n5308) );
  AND U6852 ( .A(n626), .B(n5309), .Z(n5307) );
  XOR U6853 ( .A(n5310), .B(n5311), .Z(n5309) );
  XOR U6854 ( .A(DB[693]), .B(DB[686]), .Z(n5311) );
  AND U6855 ( .A(n630), .B(n5312), .Z(n5310) );
  XOR U6856 ( .A(n5313), .B(n5314), .Z(n5312) );
  XOR U6857 ( .A(DB[686]), .B(DB[679]), .Z(n5314) );
  AND U6858 ( .A(n634), .B(n5315), .Z(n5313) );
  XOR U6859 ( .A(n5316), .B(n5317), .Z(n5315) );
  XOR U6860 ( .A(DB[679]), .B(DB[672]), .Z(n5317) );
  AND U6861 ( .A(n638), .B(n5318), .Z(n5316) );
  XOR U6862 ( .A(n5319), .B(n5320), .Z(n5318) );
  XOR U6863 ( .A(DB[672]), .B(DB[665]), .Z(n5320) );
  AND U6864 ( .A(n642), .B(n5321), .Z(n5319) );
  XOR U6865 ( .A(n5322), .B(n5323), .Z(n5321) );
  XOR U6866 ( .A(DB[665]), .B(DB[658]), .Z(n5323) );
  AND U6867 ( .A(n646), .B(n5324), .Z(n5322) );
  XOR U6868 ( .A(n5325), .B(n5326), .Z(n5324) );
  XOR U6869 ( .A(DB[658]), .B(DB[651]), .Z(n5326) );
  AND U6870 ( .A(n650), .B(n5327), .Z(n5325) );
  XOR U6871 ( .A(n5328), .B(n5329), .Z(n5327) );
  XOR U6872 ( .A(DB[651]), .B(DB[644]), .Z(n5329) );
  AND U6873 ( .A(n654), .B(n5330), .Z(n5328) );
  XOR U6874 ( .A(n5331), .B(n5332), .Z(n5330) );
  XOR U6875 ( .A(DB[644]), .B(DB[637]), .Z(n5332) );
  AND U6876 ( .A(n658), .B(n5333), .Z(n5331) );
  XOR U6877 ( .A(n5334), .B(n5335), .Z(n5333) );
  XOR U6878 ( .A(DB[637]), .B(DB[630]), .Z(n5335) );
  AND U6879 ( .A(n662), .B(n5336), .Z(n5334) );
  XOR U6880 ( .A(n5337), .B(n5338), .Z(n5336) );
  XOR U6881 ( .A(DB[630]), .B(DB[623]), .Z(n5338) );
  AND U6882 ( .A(n666), .B(n5339), .Z(n5337) );
  XOR U6883 ( .A(n5340), .B(n5341), .Z(n5339) );
  XOR U6884 ( .A(DB[623]), .B(DB[616]), .Z(n5341) );
  AND U6885 ( .A(n670), .B(n5342), .Z(n5340) );
  XOR U6886 ( .A(n5343), .B(n5344), .Z(n5342) );
  XOR U6887 ( .A(DB[616]), .B(DB[609]), .Z(n5344) );
  AND U6888 ( .A(n674), .B(n5345), .Z(n5343) );
  XOR U6889 ( .A(n5346), .B(n5347), .Z(n5345) );
  XOR U6890 ( .A(DB[609]), .B(DB[602]), .Z(n5347) );
  AND U6891 ( .A(n678), .B(n5348), .Z(n5346) );
  XOR U6892 ( .A(n5349), .B(n5350), .Z(n5348) );
  XOR U6893 ( .A(DB[602]), .B(DB[595]), .Z(n5350) );
  AND U6894 ( .A(n682), .B(n5351), .Z(n5349) );
  XOR U6895 ( .A(n5352), .B(n5353), .Z(n5351) );
  XOR U6896 ( .A(DB[595]), .B(DB[588]), .Z(n5353) );
  AND U6897 ( .A(n686), .B(n5354), .Z(n5352) );
  XOR U6898 ( .A(n5355), .B(n5356), .Z(n5354) );
  XOR U6899 ( .A(DB[588]), .B(DB[581]), .Z(n5356) );
  AND U6900 ( .A(n690), .B(n5357), .Z(n5355) );
  XOR U6901 ( .A(n5358), .B(n5359), .Z(n5357) );
  XOR U6902 ( .A(DB[581]), .B(DB[574]), .Z(n5359) );
  AND U6903 ( .A(n694), .B(n5360), .Z(n5358) );
  XOR U6904 ( .A(n5361), .B(n5362), .Z(n5360) );
  XOR U6905 ( .A(DB[574]), .B(DB[567]), .Z(n5362) );
  AND U6906 ( .A(n698), .B(n5363), .Z(n5361) );
  XOR U6907 ( .A(n5364), .B(n5365), .Z(n5363) );
  XOR U6908 ( .A(DB[567]), .B(DB[560]), .Z(n5365) );
  AND U6909 ( .A(n702), .B(n5366), .Z(n5364) );
  XOR U6910 ( .A(n5367), .B(n5368), .Z(n5366) );
  XOR U6911 ( .A(DB[560]), .B(DB[553]), .Z(n5368) );
  AND U6912 ( .A(n706), .B(n5369), .Z(n5367) );
  XOR U6913 ( .A(n5370), .B(n5371), .Z(n5369) );
  XOR U6914 ( .A(DB[553]), .B(DB[546]), .Z(n5371) );
  AND U6915 ( .A(n710), .B(n5372), .Z(n5370) );
  XOR U6916 ( .A(n5373), .B(n5374), .Z(n5372) );
  XOR U6917 ( .A(DB[546]), .B(DB[539]), .Z(n5374) );
  AND U6918 ( .A(n714), .B(n5375), .Z(n5373) );
  XOR U6919 ( .A(n5376), .B(n5377), .Z(n5375) );
  XOR U6920 ( .A(DB[539]), .B(DB[532]), .Z(n5377) );
  AND U6921 ( .A(n718), .B(n5378), .Z(n5376) );
  XOR U6922 ( .A(n5379), .B(n5380), .Z(n5378) );
  XOR U6923 ( .A(DB[532]), .B(DB[525]), .Z(n5380) );
  AND U6924 ( .A(n722), .B(n5381), .Z(n5379) );
  XOR U6925 ( .A(n5382), .B(n5383), .Z(n5381) );
  XOR U6926 ( .A(DB[525]), .B(DB[518]), .Z(n5383) );
  AND U6927 ( .A(n726), .B(n5384), .Z(n5382) );
  XOR U6928 ( .A(n5385), .B(n5386), .Z(n5384) );
  XOR U6929 ( .A(DB[518]), .B(DB[511]), .Z(n5386) );
  AND U6930 ( .A(n730), .B(n5387), .Z(n5385) );
  XOR U6931 ( .A(n5388), .B(n5389), .Z(n5387) );
  XOR U6932 ( .A(DB[511]), .B(DB[504]), .Z(n5389) );
  AND U6933 ( .A(n734), .B(n5390), .Z(n5388) );
  XOR U6934 ( .A(n5391), .B(n5392), .Z(n5390) );
  XOR U6935 ( .A(DB[504]), .B(DB[497]), .Z(n5392) );
  AND U6936 ( .A(n738), .B(n5393), .Z(n5391) );
  XOR U6937 ( .A(n5394), .B(n5395), .Z(n5393) );
  XOR U6938 ( .A(DB[497]), .B(DB[490]), .Z(n5395) );
  AND U6939 ( .A(n742), .B(n5396), .Z(n5394) );
  XOR U6940 ( .A(n5397), .B(n5398), .Z(n5396) );
  XOR U6941 ( .A(DB[490]), .B(DB[483]), .Z(n5398) );
  AND U6942 ( .A(n746), .B(n5399), .Z(n5397) );
  XOR U6943 ( .A(n5400), .B(n5401), .Z(n5399) );
  XOR U6944 ( .A(DB[483]), .B(DB[476]), .Z(n5401) );
  AND U6945 ( .A(n750), .B(n5402), .Z(n5400) );
  XOR U6946 ( .A(n5403), .B(n5404), .Z(n5402) );
  XOR U6947 ( .A(DB[476]), .B(DB[469]), .Z(n5404) );
  AND U6948 ( .A(n754), .B(n5405), .Z(n5403) );
  XOR U6949 ( .A(n5406), .B(n5407), .Z(n5405) );
  XOR U6950 ( .A(DB[469]), .B(DB[462]), .Z(n5407) );
  AND U6951 ( .A(n758), .B(n5408), .Z(n5406) );
  XOR U6952 ( .A(n5409), .B(n5410), .Z(n5408) );
  XOR U6953 ( .A(DB[462]), .B(DB[455]), .Z(n5410) );
  AND U6954 ( .A(n762), .B(n5411), .Z(n5409) );
  XOR U6955 ( .A(n5412), .B(n5413), .Z(n5411) );
  XOR U6956 ( .A(DB[455]), .B(DB[448]), .Z(n5413) );
  AND U6957 ( .A(n766), .B(n5414), .Z(n5412) );
  XOR U6958 ( .A(n5415), .B(n5416), .Z(n5414) );
  XOR U6959 ( .A(DB[448]), .B(DB[441]), .Z(n5416) );
  AND U6960 ( .A(n770), .B(n5417), .Z(n5415) );
  XOR U6961 ( .A(n5418), .B(n5419), .Z(n5417) );
  XOR U6962 ( .A(DB[441]), .B(DB[434]), .Z(n5419) );
  AND U6963 ( .A(n774), .B(n5420), .Z(n5418) );
  XOR U6964 ( .A(n5421), .B(n5422), .Z(n5420) );
  XOR U6965 ( .A(DB[434]), .B(DB[427]), .Z(n5422) );
  AND U6966 ( .A(n778), .B(n5423), .Z(n5421) );
  XOR U6967 ( .A(n5424), .B(n5425), .Z(n5423) );
  XOR U6968 ( .A(DB[427]), .B(DB[420]), .Z(n5425) );
  AND U6969 ( .A(n782), .B(n5426), .Z(n5424) );
  XOR U6970 ( .A(n5427), .B(n5428), .Z(n5426) );
  XOR U6971 ( .A(DB[420]), .B(DB[413]), .Z(n5428) );
  AND U6972 ( .A(n786), .B(n5429), .Z(n5427) );
  XOR U6973 ( .A(n5430), .B(n5431), .Z(n5429) );
  XOR U6974 ( .A(DB[413]), .B(DB[406]), .Z(n5431) );
  AND U6975 ( .A(n790), .B(n5432), .Z(n5430) );
  XOR U6976 ( .A(n5433), .B(n5434), .Z(n5432) );
  XOR U6977 ( .A(DB[406]), .B(DB[399]), .Z(n5434) );
  AND U6978 ( .A(n794), .B(n5435), .Z(n5433) );
  XOR U6979 ( .A(n5436), .B(n5437), .Z(n5435) );
  XOR U6980 ( .A(DB[399]), .B(DB[392]), .Z(n5437) );
  AND U6981 ( .A(n798), .B(n5438), .Z(n5436) );
  XOR U6982 ( .A(n5439), .B(n5440), .Z(n5438) );
  XOR U6983 ( .A(DB[392]), .B(DB[385]), .Z(n5440) );
  AND U6984 ( .A(n802), .B(n5441), .Z(n5439) );
  XOR U6985 ( .A(n5442), .B(n5443), .Z(n5441) );
  XOR U6986 ( .A(DB[385]), .B(DB[378]), .Z(n5443) );
  AND U6987 ( .A(n806), .B(n5444), .Z(n5442) );
  XOR U6988 ( .A(n5445), .B(n5446), .Z(n5444) );
  XOR U6989 ( .A(DB[378]), .B(DB[371]), .Z(n5446) );
  AND U6990 ( .A(n810), .B(n5447), .Z(n5445) );
  XOR U6991 ( .A(n5448), .B(n5449), .Z(n5447) );
  XOR U6992 ( .A(DB[371]), .B(DB[364]), .Z(n5449) );
  AND U6993 ( .A(n814), .B(n5450), .Z(n5448) );
  XOR U6994 ( .A(n5451), .B(n5452), .Z(n5450) );
  XOR U6995 ( .A(DB[364]), .B(DB[357]), .Z(n5452) );
  AND U6996 ( .A(n818), .B(n5453), .Z(n5451) );
  XOR U6997 ( .A(n5454), .B(n5455), .Z(n5453) );
  XOR U6998 ( .A(DB[357]), .B(DB[350]), .Z(n5455) );
  AND U6999 ( .A(n822), .B(n5456), .Z(n5454) );
  XOR U7000 ( .A(n5457), .B(n5458), .Z(n5456) );
  XOR U7001 ( .A(DB[350]), .B(DB[343]), .Z(n5458) );
  AND U7002 ( .A(n826), .B(n5459), .Z(n5457) );
  XOR U7003 ( .A(n5460), .B(n5461), .Z(n5459) );
  XOR U7004 ( .A(DB[343]), .B(DB[336]), .Z(n5461) );
  AND U7005 ( .A(n830), .B(n5462), .Z(n5460) );
  XOR U7006 ( .A(n5463), .B(n5464), .Z(n5462) );
  XOR U7007 ( .A(DB[336]), .B(DB[329]), .Z(n5464) );
  AND U7008 ( .A(n834), .B(n5465), .Z(n5463) );
  XOR U7009 ( .A(n5466), .B(n5467), .Z(n5465) );
  XOR U7010 ( .A(DB[329]), .B(DB[322]), .Z(n5467) );
  AND U7011 ( .A(n838), .B(n5468), .Z(n5466) );
  XOR U7012 ( .A(n5469), .B(n5470), .Z(n5468) );
  XOR U7013 ( .A(DB[322]), .B(DB[315]), .Z(n5470) );
  AND U7014 ( .A(n842), .B(n5471), .Z(n5469) );
  XOR U7015 ( .A(n5472), .B(n5473), .Z(n5471) );
  XOR U7016 ( .A(DB[315]), .B(DB[308]), .Z(n5473) );
  AND U7017 ( .A(n846), .B(n5474), .Z(n5472) );
  XOR U7018 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U7019 ( .A(DB[308]), .B(DB[301]), .Z(n5476) );
  AND U7020 ( .A(n850), .B(n5477), .Z(n5475) );
  XOR U7021 ( .A(n5478), .B(n5479), .Z(n5477) );
  XOR U7022 ( .A(DB[301]), .B(DB[294]), .Z(n5479) );
  AND U7023 ( .A(n854), .B(n5480), .Z(n5478) );
  XOR U7024 ( .A(n5481), .B(n5482), .Z(n5480) );
  XOR U7025 ( .A(DB[294]), .B(DB[287]), .Z(n5482) );
  AND U7026 ( .A(n858), .B(n5483), .Z(n5481) );
  XOR U7027 ( .A(n5484), .B(n5485), .Z(n5483) );
  XOR U7028 ( .A(DB[287]), .B(DB[280]), .Z(n5485) );
  AND U7029 ( .A(n862), .B(n5486), .Z(n5484) );
  XOR U7030 ( .A(n5487), .B(n5488), .Z(n5486) );
  XOR U7031 ( .A(DB[280]), .B(DB[273]), .Z(n5488) );
  AND U7032 ( .A(n866), .B(n5489), .Z(n5487) );
  XOR U7033 ( .A(n5490), .B(n5491), .Z(n5489) );
  XOR U7034 ( .A(DB[273]), .B(DB[266]), .Z(n5491) );
  AND U7035 ( .A(n870), .B(n5492), .Z(n5490) );
  XOR U7036 ( .A(n5493), .B(n5494), .Z(n5492) );
  XOR U7037 ( .A(DB[266]), .B(DB[259]), .Z(n5494) );
  AND U7038 ( .A(n874), .B(n5495), .Z(n5493) );
  XOR U7039 ( .A(n5496), .B(n5497), .Z(n5495) );
  XOR U7040 ( .A(DB[259]), .B(DB[252]), .Z(n5497) );
  AND U7041 ( .A(n878), .B(n5498), .Z(n5496) );
  XOR U7042 ( .A(n5499), .B(n5500), .Z(n5498) );
  XOR U7043 ( .A(DB[252]), .B(DB[245]), .Z(n5500) );
  AND U7044 ( .A(n882), .B(n5501), .Z(n5499) );
  XOR U7045 ( .A(n5502), .B(n5503), .Z(n5501) );
  XOR U7046 ( .A(DB[245]), .B(DB[238]), .Z(n5503) );
  AND U7047 ( .A(n886), .B(n5504), .Z(n5502) );
  XOR U7048 ( .A(n5505), .B(n5506), .Z(n5504) );
  XOR U7049 ( .A(DB[238]), .B(DB[231]), .Z(n5506) );
  AND U7050 ( .A(n890), .B(n5507), .Z(n5505) );
  XOR U7051 ( .A(n5508), .B(n5509), .Z(n5507) );
  XOR U7052 ( .A(DB[231]), .B(DB[224]), .Z(n5509) );
  AND U7053 ( .A(n894), .B(n5510), .Z(n5508) );
  XOR U7054 ( .A(n5511), .B(n5512), .Z(n5510) );
  XOR U7055 ( .A(DB[224]), .B(DB[217]), .Z(n5512) );
  AND U7056 ( .A(n898), .B(n5513), .Z(n5511) );
  XOR U7057 ( .A(n5514), .B(n5515), .Z(n5513) );
  XOR U7058 ( .A(DB[217]), .B(DB[210]), .Z(n5515) );
  AND U7059 ( .A(n902), .B(n5516), .Z(n5514) );
  XOR U7060 ( .A(n5517), .B(n5518), .Z(n5516) );
  XOR U7061 ( .A(DB[210]), .B(DB[203]), .Z(n5518) );
  AND U7062 ( .A(n906), .B(n5519), .Z(n5517) );
  XOR U7063 ( .A(n5520), .B(n5521), .Z(n5519) );
  XOR U7064 ( .A(DB[203]), .B(DB[196]), .Z(n5521) );
  AND U7065 ( .A(n910), .B(n5522), .Z(n5520) );
  XOR U7066 ( .A(n5523), .B(n5524), .Z(n5522) );
  XOR U7067 ( .A(DB[196]), .B(DB[189]), .Z(n5524) );
  AND U7068 ( .A(n914), .B(n5525), .Z(n5523) );
  XOR U7069 ( .A(n5526), .B(n5527), .Z(n5525) );
  XOR U7070 ( .A(DB[189]), .B(DB[182]), .Z(n5527) );
  AND U7071 ( .A(n918), .B(n5528), .Z(n5526) );
  XOR U7072 ( .A(n5529), .B(n5530), .Z(n5528) );
  XOR U7073 ( .A(DB[182]), .B(DB[175]), .Z(n5530) );
  AND U7074 ( .A(n922), .B(n5531), .Z(n5529) );
  XOR U7075 ( .A(n5532), .B(n5533), .Z(n5531) );
  XOR U7076 ( .A(DB[175]), .B(DB[168]), .Z(n5533) );
  AND U7077 ( .A(n926), .B(n5534), .Z(n5532) );
  XOR U7078 ( .A(n5535), .B(n5536), .Z(n5534) );
  XOR U7079 ( .A(DB[168]), .B(DB[161]), .Z(n5536) );
  AND U7080 ( .A(n930), .B(n5537), .Z(n5535) );
  XOR U7081 ( .A(n5538), .B(n5539), .Z(n5537) );
  XOR U7082 ( .A(DB[161]), .B(DB[154]), .Z(n5539) );
  AND U7083 ( .A(n934), .B(n5540), .Z(n5538) );
  XOR U7084 ( .A(n5541), .B(n5542), .Z(n5540) );
  XOR U7085 ( .A(DB[154]), .B(DB[147]), .Z(n5542) );
  AND U7086 ( .A(n938), .B(n5543), .Z(n5541) );
  XOR U7087 ( .A(n5544), .B(n5545), .Z(n5543) );
  XOR U7088 ( .A(DB[147]), .B(DB[140]), .Z(n5545) );
  AND U7089 ( .A(n942), .B(n5546), .Z(n5544) );
  XOR U7090 ( .A(n5547), .B(n5548), .Z(n5546) );
  XOR U7091 ( .A(DB[140]), .B(DB[133]), .Z(n5548) );
  AND U7092 ( .A(n946), .B(n5549), .Z(n5547) );
  XOR U7093 ( .A(n5550), .B(n5551), .Z(n5549) );
  XOR U7094 ( .A(DB[133]), .B(DB[126]), .Z(n5551) );
  AND U7095 ( .A(n950), .B(n5552), .Z(n5550) );
  XOR U7096 ( .A(n5553), .B(n5554), .Z(n5552) );
  XOR U7097 ( .A(DB[126]), .B(DB[119]), .Z(n5554) );
  AND U7098 ( .A(n954), .B(n5555), .Z(n5553) );
  XOR U7099 ( .A(n5556), .B(n5557), .Z(n5555) );
  XOR U7100 ( .A(DB[119]), .B(DB[112]), .Z(n5557) );
  AND U7101 ( .A(n958), .B(n5558), .Z(n5556) );
  XOR U7102 ( .A(n5559), .B(n5560), .Z(n5558) );
  XOR U7103 ( .A(DB[112]), .B(DB[105]), .Z(n5560) );
  AND U7104 ( .A(n962), .B(n5561), .Z(n5559) );
  XOR U7105 ( .A(n5562), .B(n5563), .Z(n5561) );
  XOR U7106 ( .A(DB[98]), .B(DB[105]), .Z(n5563) );
  AND U7107 ( .A(n966), .B(n5564), .Z(n5562) );
  XOR U7108 ( .A(n5565), .B(n5566), .Z(n5564) );
  XOR U7109 ( .A(DB[98]), .B(DB[91]), .Z(n5566) );
  AND U7110 ( .A(n970), .B(n5567), .Z(n5565) );
  XOR U7111 ( .A(n5568), .B(n5569), .Z(n5567) );
  XOR U7112 ( .A(DB[91]), .B(DB[84]), .Z(n5569) );
  AND U7113 ( .A(n974), .B(n5570), .Z(n5568) );
  XOR U7114 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U7115 ( .A(DB[84]), .B(DB[77]), .Z(n5572) );
  AND U7116 ( .A(n978), .B(n5573), .Z(n5571) );
  XOR U7117 ( .A(n5574), .B(n5575), .Z(n5573) );
  XOR U7118 ( .A(DB[77]), .B(DB[70]), .Z(n5575) );
  AND U7119 ( .A(n982), .B(n5576), .Z(n5574) );
  XOR U7120 ( .A(n5577), .B(n5578), .Z(n5576) );
  XOR U7121 ( .A(DB[70]), .B(DB[63]), .Z(n5578) );
  AND U7122 ( .A(n986), .B(n5579), .Z(n5577) );
  XOR U7123 ( .A(n5580), .B(n5581), .Z(n5579) );
  XOR U7124 ( .A(DB[63]), .B(DB[56]), .Z(n5581) );
  AND U7125 ( .A(n990), .B(n5582), .Z(n5580) );
  XOR U7126 ( .A(n5583), .B(n5584), .Z(n5582) );
  XOR U7127 ( .A(DB[56]), .B(DB[49]), .Z(n5584) );
  AND U7128 ( .A(n994), .B(n5585), .Z(n5583) );
  XOR U7129 ( .A(n5586), .B(n5587), .Z(n5585) );
  XOR U7130 ( .A(DB[49]), .B(DB[42]), .Z(n5587) );
  AND U7131 ( .A(n998), .B(n5588), .Z(n5586) );
  XOR U7132 ( .A(n5589), .B(n5590), .Z(n5588) );
  XOR U7133 ( .A(DB[42]), .B(DB[35]), .Z(n5590) );
  AND U7134 ( .A(n1002), .B(n5591), .Z(n5589) );
  XOR U7135 ( .A(n5592), .B(n5593), .Z(n5591) );
  XOR U7136 ( .A(DB[35]), .B(DB[28]), .Z(n5593) );
  AND U7137 ( .A(n1006), .B(n5594), .Z(n5592) );
  XOR U7138 ( .A(n5595), .B(n5596), .Z(n5594) );
  XOR U7139 ( .A(DB[28]), .B(DB[21]), .Z(n5596) );
  AND U7140 ( .A(n1010), .B(n5597), .Z(n5595) );
  XOR U7141 ( .A(n5598), .B(n5599), .Z(n5597) );
  XOR U7142 ( .A(DB[21]), .B(DB[14]), .Z(n5599) );
  AND U7143 ( .A(n1014), .B(n5600), .Z(n5598) );
  XOR U7144 ( .A(n5601), .B(n5602), .Z(n5600) );
  XOR U7145 ( .A(DB[7]), .B(DB[14]), .Z(n5602) );
  AND U7146 ( .A(n1018), .B(n5603), .Z(n5601) );
  XOR U7147 ( .A(DB[7]), .B(DB[0]), .Z(n5603) );
  XOR U7148 ( .A(n5604), .B(n5605), .Z(n2) );
  AND U7149 ( .A(n5606), .B(n5607), .Z(n5604) );
  XNOR U7150 ( .A(n5605), .B(n5608), .Z(n5607) );
  XOR U7151 ( .A(n5609), .B(n5610), .Z(n5608) );
  AND U7152 ( .A(n5611), .B(n5612), .Z(n5609) );
  XNOR U7153 ( .A(n5613), .B(n5614), .Z(n5612) );
  XNOR U7154 ( .A(n5605), .B(n5615), .Z(n5606) );
  XNOR U7155 ( .A(n5616), .B(n5617), .Z(n5615) );
  AND U7156 ( .A(n6), .B(n5618), .Z(n5616) );
  XOR U7157 ( .A(n5619), .B(n5617), .Z(n5618) );
  XNOR U7158 ( .A(n5620), .B(n5621), .Z(n5605) );
  NAND U7159 ( .A(n5622), .B(n5623), .Z(n5621) );
  XOR U7160 ( .A(n5611), .B(n5624), .Z(n5623) );
  XNOR U7161 ( .A(n5620), .B(n5613), .Z(n5624) );
  XOR U7162 ( .A(n5625), .B(n5626), .Z(n5613) );
  ANDN U7163 ( .B(n5627), .A(n5628), .Z(n5625) );
  XNOR U7164 ( .A(n5626), .B(n5629), .Z(n5627) );
  XNOR U7165 ( .A(n5610), .B(n5630), .Z(n5611) );
  XNOR U7166 ( .A(n5631), .B(n5632), .Z(n5630) );
  ANDN U7167 ( .B(n5633), .A(n5634), .Z(n5631) );
  XNOR U7168 ( .A(n5635), .B(n5636), .Z(n5633) );
  IV U7169 ( .A(n5632), .Z(n5636) );
  IV U7170 ( .A(n5614), .Z(n5610) );
  XNOR U7171 ( .A(n5637), .B(n5638), .Z(n5614) );
  AND U7172 ( .A(n5639), .B(n5640), .Z(n5637) );
  XNOR U7173 ( .A(n5638), .B(n5641), .Z(n5640) );
  XOR U7174 ( .A(n5642), .B(n5643), .Z(n5622) );
  XNOR U7175 ( .A(n5620), .B(n5644), .Z(n5643) );
  NAND U7176 ( .A(n5645), .B(n6), .Z(n5644) );
  XOR U7177 ( .A(n5646), .B(n5642), .Z(n5645) );
  NAND U7178 ( .A(n5647), .B(n5648), .Z(n5620) );
  XNOR U7179 ( .A(n5639), .B(n5641), .Z(n5648) );
  XOR U7180 ( .A(n5649), .B(n5629), .Z(n5641) );
  XNOR U7181 ( .A(q[6]), .B(DB[1791]), .Z(n5629) );
  IV U7182 ( .A(n5628), .Z(n5649) );
  XOR U7183 ( .A(n5626), .B(n5650), .Z(n5628) );
  XNOR U7184 ( .A(q[5]), .B(DB[1790]), .Z(n5650) );
  XOR U7185 ( .A(q[4]), .B(DB[1789]), .Z(n5626) );
  XNOR U7186 ( .A(n5651), .B(n5652), .Z(n5639) );
  XNOR U7187 ( .A(n5635), .B(n5638), .Z(n5652) );
  XOR U7188 ( .A(q[0]), .B(DB[1785]), .Z(n5638) );
  XOR U7189 ( .A(q[3]), .B(DB[1788]), .Z(n5635) );
  IV U7190 ( .A(n5634), .Z(n5651) );
  XOR U7191 ( .A(n5632), .B(n5653), .Z(n5634) );
  XNOR U7192 ( .A(q[2]), .B(DB[1787]), .Z(n5653) );
  XOR U7193 ( .A(q[1]), .B(DB[1786]), .Z(n5632) );
  XOR U7194 ( .A(n5654), .B(n5655), .Z(n5647) );
  AND U7195 ( .A(n6), .B(n5656), .Z(n5654) );
  XOR U7196 ( .A(n5655), .B(n5657), .Z(n5656) );
  XOR U7197 ( .A(n5658), .B(n5659), .Z(n6) );
  AND U7198 ( .A(n5660), .B(n5661), .Z(n5658) );
  XNOR U7199 ( .A(n5659), .B(n5617), .Z(n5661) );
  XNOR U7200 ( .A(n5662), .B(n5663), .Z(n5617) );
  ANDN U7201 ( .B(n5664), .A(n5665), .Z(n5662) );
  XOR U7202 ( .A(n5663), .B(n5666), .Z(n5664) );
  XOR U7203 ( .A(n5659), .B(n5619), .Z(n5660) );
  XOR U7204 ( .A(n5667), .B(n5668), .Z(n5619) );
  AND U7205 ( .A(n10), .B(n5669), .Z(n5667) );
  XOR U7206 ( .A(n5670), .B(n5668), .Z(n5669) );
  XNOR U7207 ( .A(n5671), .B(n5672), .Z(n5659) );
  NAND U7208 ( .A(n5673), .B(n5674), .Z(n5672) );
  XOR U7209 ( .A(n5675), .B(n5642), .Z(n5674) );
  XNOR U7210 ( .A(n5676), .B(n5666), .Z(n5642) );
  XOR U7211 ( .A(n5677), .B(n5678), .Z(n5666) );
  ANDN U7212 ( .B(n5679), .A(n5680), .Z(n5677) );
  XOR U7213 ( .A(n5678), .B(n5681), .Z(n5679) );
  IV U7214 ( .A(n5665), .Z(n5676) );
  XOR U7215 ( .A(n5682), .B(n5683), .Z(n5665) );
  XOR U7216 ( .A(n5684), .B(n5685), .Z(n5683) );
  ANDN U7217 ( .B(n5686), .A(n5687), .Z(n5684) );
  XOR U7218 ( .A(n5688), .B(n5685), .Z(n5686) );
  IV U7219 ( .A(n5663), .Z(n5682) );
  XOR U7220 ( .A(n5689), .B(n5690), .Z(n5663) );
  ANDN U7221 ( .B(n5691), .A(n5692), .Z(n5689) );
  XOR U7222 ( .A(n5690), .B(n5693), .Z(n5691) );
  IV U7223 ( .A(n5671), .Z(n5675) );
  XOR U7224 ( .A(n5671), .B(n5646), .Z(n5673) );
  XOR U7225 ( .A(n5694), .B(n5695), .Z(n5646) );
  AND U7226 ( .A(n10), .B(n5696), .Z(n5694) );
  XOR U7227 ( .A(n5697), .B(n5695), .Z(n5696) );
  NANDN U7228 ( .A(n5655), .B(n5657), .Z(n5671) );
  XOR U7229 ( .A(n5698), .B(n5699), .Z(n5657) );
  AND U7230 ( .A(n10), .B(n5700), .Z(n5698) );
  XOR U7231 ( .A(n5699), .B(n5701), .Z(n5700) );
  XOR U7232 ( .A(n5702), .B(n5703), .Z(n10) );
  AND U7233 ( .A(n5704), .B(n5705), .Z(n5702) );
  XNOR U7234 ( .A(n5703), .B(n5668), .Z(n5705) );
  XNOR U7235 ( .A(n5706), .B(n5707), .Z(n5668) );
  ANDN U7236 ( .B(n5708), .A(n5709), .Z(n5706) );
  XOR U7237 ( .A(n5707), .B(n5710), .Z(n5708) );
  XOR U7238 ( .A(n5703), .B(n5670), .Z(n5704) );
  XOR U7239 ( .A(n5711), .B(n5712), .Z(n5670) );
  AND U7240 ( .A(n14), .B(n5713), .Z(n5711) );
  XOR U7241 ( .A(n5714), .B(n5712), .Z(n5713) );
  XNOR U7242 ( .A(n5715), .B(n5716), .Z(n5703) );
  NAND U7243 ( .A(n5717), .B(n5718), .Z(n5716) );
  XOR U7244 ( .A(n5719), .B(n5695), .Z(n5718) );
  XOR U7245 ( .A(n5709), .B(n5710), .Z(n5695) );
  XOR U7246 ( .A(n5720), .B(n5721), .Z(n5710) );
  ANDN U7247 ( .B(n5722), .A(n5723), .Z(n5720) );
  XOR U7248 ( .A(n5721), .B(n5724), .Z(n5722) );
  XOR U7249 ( .A(n5725), .B(n5726), .Z(n5709) );
  XOR U7250 ( .A(n5727), .B(n5728), .Z(n5726) );
  ANDN U7251 ( .B(n5729), .A(n5730), .Z(n5727) );
  XOR U7252 ( .A(n5731), .B(n5728), .Z(n5729) );
  IV U7253 ( .A(n5707), .Z(n5725) );
  XOR U7254 ( .A(n5732), .B(n5733), .Z(n5707) );
  ANDN U7255 ( .B(n5734), .A(n5735), .Z(n5732) );
  XOR U7256 ( .A(n5733), .B(n5736), .Z(n5734) );
  IV U7257 ( .A(n5715), .Z(n5719) );
  XOR U7258 ( .A(n5715), .B(n5697), .Z(n5717) );
  XOR U7259 ( .A(n5737), .B(n5738), .Z(n5697) );
  AND U7260 ( .A(n14), .B(n5739), .Z(n5737) );
  XOR U7261 ( .A(n5740), .B(n5738), .Z(n5739) );
  NANDN U7262 ( .A(n5699), .B(n5701), .Z(n5715) );
  XOR U7263 ( .A(n5741), .B(n5742), .Z(n5701) );
  AND U7264 ( .A(n14), .B(n5743), .Z(n5741) );
  XOR U7265 ( .A(n5742), .B(n5744), .Z(n5743) );
  XOR U7266 ( .A(n5745), .B(n5746), .Z(n14) );
  AND U7267 ( .A(n5747), .B(n5748), .Z(n5745) );
  XNOR U7268 ( .A(n5746), .B(n5712), .Z(n5748) );
  XNOR U7269 ( .A(n5749), .B(n5750), .Z(n5712) );
  ANDN U7270 ( .B(n5751), .A(n5752), .Z(n5749) );
  XOR U7271 ( .A(n5750), .B(n5753), .Z(n5751) );
  XOR U7272 ( .A(n5746), .B(n5714), .Z(n5747) );
  XOR U7273 ( .A(n5754), .B(n5755), .Z(n5714) );
  AND U7274 ( .A(n18), .B(n5756), .Z(n5754) );
  XOR U7275 ( .A(n5757), .B(n5755), .Z(n5756) );
  XNOR U7276 ( .A(n5758), .B(n5759), .Z(n5746) );
  NAND U7277 ( .A(n5760), .B(n5761), .Z(n5759) );
  XOR U7278 ( .A(n5762), .B(n5738), .Z(n5761) );
  XOR U7279 ( .A(n5752), .B(n5753), .Z(n5738) );
  XOR U7280 ( .A(n5763), .B(n5764), .Z(n5753) );
  ANDN U7281 ( .B(n5765), .A(n5766), .Z(n5763) );
  XOR U7282 ( .A(n5764), .B(n5767), .Z(n5765) );
  XOR U7283 ( .A(n5768), .B(n5769), .Z(n5752) );
  XOR U7284 ( .A(n5770), .B(n5771), .Z(n5769) );
  ANDN U7285 ( .B(n5772), .A(n5773), .Z(n5770) );
  XOR U7286 ( .A(n5774), .B(n5771), .Z(n5772) );
  IV U7287 ( .A(n5750), .Z(n5768) );
  XOR U7288 ( .A(n5775), .B(n5776), .Z(n5750) );
  ANDN U7289 ( .B(n5777), .A(n5778), .Z(n5775) );
  XOR U7290 ( .A(n5776), .B(n5779), .Z(n5777) );
  IV U7291 ( .A(n5758), .Z(n5762) );
  XOR U7292 ( .A(n5758), .B(n5740), .Z(n5760) );
  XOR U7293 ( .A(n5780), .B(n5781), .Z(n5740) );
  AND U7294 ( .A(n18), .B(n5782), .Z(n5780) );
  XOR U7295 ( .A(n5783), .B(n5781), .Z(n5782) );
  NANDN U7296 ( .A(n5742), .B(n5744), .Z(n5758) );
  XOR U7297 ( .A(n5784), .B(n5785), .Z(n5744) );
  AND U7298 ( .A(n18), .B(n5786), .Z(n5784) );
  XOR U7299 ( .A(n5785), .B(n5787), .Z(n5786) );
  XOR U7300 ( .A(n5788), .B(n5789), .Z(n18) );
  AND U7301 ( .A(n5790), .B(n5791), .Z(n5788) );
  XNOR U7302 ( .A(n5789), .B(n5755), .Z(n5791) );
  XNOR U7303 ( .A(n5792), .B(n5793), .Z(n5755) );
  ANDN U7304 ( .B(n5794), .A(n5795), .Z(n5792) );
  XOR U7305 ( .A(n5793), .B(n5796), .Z(n5794) );
  XOR U7306 ( .A(n5789), .B(n5757), .Z(n5790) );
  XOR U7307 ( .A(n5797), .B(n5798), .Z(n5757) );
  AND U7308 ( .A(n22), .B(n5799), .Z(n5797) );
  XOR U7309 ( .A(n5800), .B(n5798), .Z(n5799) );
  XNOR U7310 ( .A(n5801), .B(n5802), .Z(n5789) );
  NAND U7311 ( .A(n5803), .B(n5804), .Z(n5802) );
  XOR U7312 ( .A(n5805), .B(n5781), .Z(n5804) );
  XOR U7313 ( .A(n5795), .B(n5796), .Z(n5781) );
  XOR U7314 ( .A(n5806), .B(n5807), .Z(n5796) );
  ANDN U7315 ( .B(n5808), .A(n5809), .Z(n5806) );
  XOR U7316 ( .A(n5807), .B(n5810), .Z(n5808) );
  XOR U7317 ( .A(n5811), .B(n5812), .Z(n5795) );
  XOR U7318 ( .A(n5813), .B(n5814), .Z(n5812) );
  ANDN U7319 ( .B(n5815), .A(n5816), .Z(n5813) );
  XOR U7320 ( .A(n5817), .B(n5814), .Z(n5815) );
  IV U7321 ( .A(n5793), .Z(n5811) );
  XOR U7322 ( .A(n5818), .B(n5819), .Z(n5793) );
  ANDN U7323 ( .B(n5820), .A(n5821), .Z(n5818) );
  XOR U7324 ( .A(n5819), .B(n5822), .Z(n5820) );
  IV U7325 ( .A(n5801), .Z(n5805) );
  XOR U7326 ( .A(n5801), .B(n5783), .Z(n5803) );
  XOR U7327 ( .A(n5823), .B(n5824), .Z(n5783) );
  AND U7328 ( .A(n22), .B(n5825), .Z(n5823) );
  XOR U7329 ( .A(n5826), .B(n5824), .Z(n5825) );
  NANDN U7330 ( .A(n5785), .B(n5787), .Z(n5801) );
  XOR U7331 ( .A(n5827), .B(n5828), .Z(n5787) );
  AND U7332 ( .A(n22), .B(n5829), .Z(n5827) );
  XOR U7333 ( .A(n5828), .B(n5830), .Z(n5829) );
  XOR U7334 ( .A(n5831), .B(n5832), .Z(n22) );
  AND U7335 ( .A(n5833), .B(n5834), .Z(n5831) );
  XNOR U7336 ( .A(n5832), .B(n5798), .Z(n5834) );
  XNOR U7337 ( .A(n5835), .B(n5836), .Z(n5798) );
  ANDN U7338 ( .B(n5837), .A(n5838), .Z(n5835) );
  XOR U7339 ( .A(n5836), .B(n5839), .Z(n5837) );
  XOR U7340 ( .A(n5832), .B(n5800), .Z(n5833) );
  XOR U7341 ( .A(n5840), .B(n5841), .Z(n5800) );
  AND U7342 ( .A(n26), .B(n5842), .Z(n5840) );
  XOR U7343 ( .A(n5843), .B(n5841), .Z(n5842) );
  XNOR U7344 ( .A(n5844), .B(n5845), .Z(n5832) );
  NAND U7345 ( .A(n5846), .B(n5847), .Z(n5845) );
  XOR U7346 ( .A(n5848), .B(n5824), .Z(n5847) );
  XOR U7347 ( .A(n5838), .B(n5839), .Z(n5824) );
  XOR U7348 ( .A(n5849), .B(n5850), .Z(n5839) );
  ANDN U7349 ( .B(n5851), .A(n5852), .Z(n5849) );
  XOR U7350 ( .A(n5850), .B(n5853), .Z(n5851) );
  XOR U7351 ( .A(n5854), .B(n5855), .Z(n5838) );
  XOR U7352 ( .A(n5856), .B(n5857), .Z(n5855) );
  ANDN U7353 ( .B(n5858), .A(n5859), .Z(n5856) );
  XOR U7354 ( .A(n5860), .B(n5857), .Z(n5858) );
  IV U7355 ( .A(n5836), .Z(n5854) );
  XOR U7356 ( .A(n5861), .B(n5862), .Z(n5836) );
  ANDN U7357 ( .B(n5863), .A(n5864), .Z(n5861) );
  XOR U7358 ( .A(n5862), .B(n5865), .Z(n5863) );
  IV U7359 ( .A(n5844), .Z(n5848) );
  XOR U7360 ( .A(n5844), .B(n5826), .Z(n5846) );
  XOR U7361 ( .A(n5866), .B(n5867), .Z(n5826) );
  AND U7362 ( .A(n26), .B(n5868), .Z(n5866) );
  XOR U7363 ( .A(n5869), .B(n5867), .Z(n5868) );
  NANDN U7364 ( .A(n5828), .B(n5830), .Z(n5844) );
  XOR U7365 ( .A(n5870), .B(n5871), .Z(n5830) );
  AND U7366 ( .A(n26), .B(n5872), .Z(n5870) );
  XOR U7367 ( .A(n5871), .B(n5873), .Z(n5872) );
  XOR U7368 ( .A(n5874), .B(n5875), .Z(n26) );
  AND U7369 ( .A(n5876), .B(n5877), .Z(n5874) );
  XNOR U7370 ( .A(n5875), .B(n5841), .Z(n5877) );
  XNOR U7371 ( .A(n5878), .B(n5879), .Z(n5841) );
  ANDN U7372 ( .B(n5880), .A(n5881), .Z(n5878) );
  XOR U7373 ( .A(n5879), .B(n5882), .Z(n5880) );
  XOR U7374 ( .A(n5875), .B(n5843), .Z(n5876) );
  XOR U7375 ( .A(n5883), .B(n5884), .Z(n5843) );
  AND U7376 ( .A(n30), .B(n5885), .Z(n5883) );
  XOR U7377 ( .A(n5886), .B(n5884), .Z(n5885) );
  XNOR U7378 ( .A(n5887), .B(n5888), .Z(n5875) );
  NAND U7379 ( .A(n5889), .B(n5890), .Z(n5888) );
  XOR U7380 ( .A(n5891), .B(n5867), .Z(n5890) );
  XOR U7381 ( .A(n5881), .B(n5882), .Z(n5867) );
  XOR U7382 ( .A(n5892), .B(n5893), .Z(n5882) );
  ANDN U7383 ( .B(n5894), .A(n5895), .Z(n5892) );
  XOR U7384 ( .A(n5893), .B(n5896), .Z(n5894) );
  XOR U7385 ( .A(n5897), .B(n5898), .Z(n5881) );
  XOR U7386 ( .A(n5899), .B(n5900), .Z(n5898) );
  ANDN U7387 ( .B(n5901), .A(n5902), .Z(n5899) );
  XOR U7388 ( .A(n5903), .B(n5900), .Z(n5901) );
  IV U7389 ( .A(n5879), .Z(n5897) );
  XOR U7390 ( .A(n5904), .B(n5905), .Z(n5879) );
  ANDN U7391 ( .B(n5906), .A(n5907), .Z(n5904) );
  XOR U7392 ( .A(n5905), .B(n5908), .Z(n5906) );
  IV U7393 ( .A(n5887), .Z(n5891) );
  XOR U7394 ( .A(n5887), .B(n5869), .Z(n5889) );
  XOR U7395 ( .A(n5909), .B(n5910), .Z(n5869) );
  AND U7396 ( .A(n30), .B(n5911), .Z(n5909) );
  XOR U7397 ( .A(n5912), .B(n5910), .Z(n5911) );
  NANDN U7398 ( .A(n5871), .B(n5873), .Z(n5887) );
  XOR U7399 ( .A(n5913), .B(n5914), .Z(n5873) );
  AND U7400 ( .A(n30), .B(n5915), .Z(n5913) );
  XOR U7401 ( .A(n5914), .B(n5916), .Z(n5915) );
  XOR U7402 ( .A(n5917), .B(n5918), .Z(n30) );
  AND U7403 ( .A(n5919), .B(n5920), .Z(n5917) );
  XNOR U7404 ( .A(n5918), .B(n5884), .Z(n5920) );
  XNOR U7405 ( .A(n5921), .B(n5922), .Z(n5884) );
  ANDN U7406 ( .B(n5923), .A(n5924), .Z(n5921) );
  XOR U7407 ( .A(n5922), .B(n5925), .Z(n5923) );
  XOR U7408 ( .A(n5918), .B(n5886), .Z(n5919) );
  XOR U7409 ( .A(n5926), .B(n5927), .Z(n5886) );
  AND U7410 ( .A(n34), .B(n5928), .Z(n5926) );
  XOR U7411 ( .A(n5929), .B(n5927), .Z(n5928) );
  XNOR U7412 ( .A(n5930), .B(n5931), .Z(n5918) );
  NAND U7413 ( .A(n5932), .B(n5933), .Z(n5931) );
  XOR U7414 ( .A(n5934), .B(n5910), .Z(n5933) );
  XOR U7415 ( .A(n5924), .B(n5925), .Z(n5910) );
  XOR U7416 ( .A(n5935), .B(n5936), .Z(n5925) );
  ANDN U7417 ( .B(n5937), .A(n5938), .Z(n5935) );
  XOR U7418 ( .A(n5936), .B(n5939), .Z(n5937) );
  XOR U7419 ( .A(n5940), .B(n5941), .Z(n5924) );
  XOR U7420 ( .A(n5942), .B(n5943), .Z(n5941) );
  ANDN U7421 ( .B(n5944), .A(n5945), .Z(n5942) );
  XOR U7422 ( .A(n5946), .B(n5943), .Z(n5944) );
  IV U7423 ( .A(n5922), .Z(n5940) );
  XOR U7424 ( .A(n5947), .B(n5948), .Z(n5922) );
  ANDN U7425 ( .B(n5949), .A(n5950), .Z(n5947) );
  XOR U7426 ( .A(n5948), .B(n5951), .Z(n5949) );
  IV U7427 ( .A(n5930), .Z(n5934) );
  XOR U7428 ( .A(n5930), .B(n5912), .Z(n5932) );
  XOR U7429 ( .A(n5952), .B(n5953), .Z(n5912) );
  AND U7430 ( .A(n34), .B(n5954), .Z(n5952) );
  XOR U7431 ( .A(n5955), .B(n5953), .Z(n5954) );
  NANDN U7432 ( .A(n5914), .B(n5916), .Z(n5930) );
  XOR U7433 ( .A(n5956), .B(n5957), .Z(n5916) );
  AND U7434 ( .A(n34), .B(n5958), .Z(n5956) );
  XOR U7435 ( .A(n5957), .B(n5959), .Z(n5958) );
  XOR U7436 ( .A(n5960), .B(n5961), .Z(n34) );
  AND U7437 ( .A(n5962), .B(n5963), .Z(n5960) );
  XNOR U7438 ( .A(n5961), .B(n5927), .Z(n5963) );
  XNOR U7439 ( .A(n5964), .B(n5965), .Z(n5927) );
  ANDN U7440 ( .B(n5966), .A(n5967), .Z(n5964) );
  XOR U7441 ( .A(n5965), .B(n5968), .Z(n5966) );
  XOR U7442 ( .A(n5961), .B(n5929), .Z(n5962) );
  XOR U7443 ( .A(n5969), .B(n5970), .Z(n5929) );
  AND U7444 ( .A(n38), .B(n5971), .Z(n5969) );
  XOR U7445 ( .A(n5972), .B(n5970), .Z(n5971) );
  XNOR U7446 ( .A(n5973), .B(n5974), .Z(n5961) );
  NAND U7447 ( .A(n5975), .B(n5976), .Z(n5974) );
  XOR U7448 ( .A(n5977), .B(n5953), .Z(n5976) );
  XOR U7449 ( .A(n5967), .B(n5968), .Z(n5953) );
  XOR U7450 ( .A(n5978), .B(n5979), .Z(n5968) );
  ANDN U7451 ( .B(n5980), .A(n5981), .Z(n5978) );
  XOR U7452 ( .A(n5979), .B(n5982), .Z(n5980) );
  XOR U7453 ( .A(n5983), .B(n5984), .Z(n5967) );
  XOR U7454 ( .A(n5985), .B(n5986), .Z(n5984) );
  ANDN U7455 ( .B(n5987), .A(n5988), .Z(n5985) );
  XOR U7456 ( .A(n5989), .B(n5986), .Z(n5987) );
  IV U7457 ( .A(n5965), .Z(n5983) );
  XOR U7458 ( .A(n5990), .B(n5991), .Z(n5965) );
  ANDN U7459 ( .B(n5992), .A(n5993), .Z(n5990) );
  XOR U7460 ( .A(n5991), .B(n5994), .Z(n5992) );
  IV U7461 ( .A(n5973), .Z(n5977) );
  XOR U7462 ( .A(n5973), .B(n5955), .Z(n5975) );
  XOR U7463 ( .A(n5995), .B(n5996), .Z(n5955) );
  AND U7464 ( .A(n38), .B(n5997), .Z(n5995) );
  XOR U7465 ( .A(n5998), .B(n5996), .Z(n5997) );
  NANDN U7466 ( .A(n5957), .B(n5959), .Z(n5973) );
  XOR U7467 ( .A(n5999), .B(n6000), .Z(n5959) );
  AND U7468 ( .A(n38), .B(n6001), .Z(n5999) );
  XOR U7469 ( .A(n6000), .B(n6002), .Z(n6001) );
  XOR U7470 ( .A(n6003), .B(n6004), .Z(n38) );
  AND U7471 ( .A(n6005), .B(n6006), .Z(n6003) );
  XNOR U7472 ( .A(n6004), .B(n5970), .Z(n6006) );
  XNOR U7473 ( .A(n6007), .B(n6008), .Z(n5970) );
  ANDN U7474 ( .B(n6009), .A(n6010), .Z(n6007) );
  XOR U7475 ( .A(n6008), .B(n6011), .Z(n6009) );
  XOR U7476 ( .A(n6004), .B(n5972), .Z(n6005) );
  XOR U7477 ( .A(n6012), .B(n6013), .Z(n5972) );
  AND U7478 ( .A(n42), .B(n6014), .Z(n6012) );
  XOR U7479 ( .A(n6015), .B(n6013), .Z(n6014) );
  XNOR U7480 ( .A(n6016), .B(n6017), .Z(n6004) );
  NAND U7481 ( .A(n6018), .B(n6019), .Z(n6017) );
  XOR U7482 ( .A(n6020), .B(n5996), .Z(n6019) );
  XOR U7483 ( .A(n6010), .B(n6011), .Z(n5996) );
  XOR U7484 ( .A(n6021), .B(n6022), .Z(n6011) );
  ANDN U7485 ( .B(n6023), .A(n6024), .Z(n6021) );
  XOR U7486 ( .A(n6022), .B(n6025), .Z(n6023) );
  XOR U7487 ( .A(n6026), .B(n6027), .Z(n6010) );
  XOR U7488 ( .A(n6028), .B(n6029), .Z(n6027) );
  ANDN U7489 ( .B(n6030), .A(n6031), .Z(n6028) );
  XOR U7490 ( .A(n6032), .B(n6029), .Z(n6030) );
  IV U7491 ( .A(n6008), .Z(n6026) );
  XOR U7492 ( .A(n6033), .B(n6034), .Z(n6008) );
  ANDN U7493 ( .B(n6035), .A(n6036), .Z(n6033) );
  XOR U7494 ( .A(n6034), .B(n6037), .Z(n6035) );
  IV U7495 ( .A(n6016), .Z(n6020) );
  XOR U7496 ( .A(n6016), .B(n5998), .Z(n6018) );
  XOR U7497 ( .A(n6038), .B(n6039), .Z(n5998) );
  AND U7498 ( .A(n42), .B(n6040), .Z(n6038) );
  XOR U7499 ( .A(n6041), .B(n6039), .Z(n6040) );
  NANDN U7500 ( .A(n6000), .B(n6002), .Z(n6016) );
  XOR U7501 ( .A(n6042), .B(n6043), .Z(n6002) );
  AND U7502 ( .A(n42), .B(n6044), .Z(n6042) );
  XOR U7503 ( .A(n6043), .B(n6045), .Z(n6044) );
  XOR U7504 ( .A(n6046), .B(n6047), .Z(n42) );
  AND U7505 ( .A(n6048), .B(n6049), .Z(n6046) );
  XNOR U7506 ( .A(n6047), .B(n6013), .Z(n6049) );
  XNOR U7507 ( .A(n6050), .B(n6051), .Z(n6013) );
  ANDN U7508 ( .B(n6052), .A(n6053), .Z(n6050) );
  XOR U7509 ( .A(n6051), .B(n6054), .Z(n6052) );
  XOR U7510 ( .A(n6047), .B(n6015), .Z(n6048) );
  XOR U7511 ( .A(n6055), .B(n6056), .Z(n6015) );
  AND U7512 ( .A(n46), .B(n6057), .Z(n6055) );
  XOR U7513 ( .A(n6058), .B(n6056), .Z(n6057) );
  XNOR U7514 ( .A(n6059), .B(n6060), .Z(n6047) );
  NAND U7515 ( .A(n6061), .B(n6062), .Z(n6060) );
  XOR U7516 ( .A(n6063), .B(n6039), .Z(n6062) );
  XOR U7517 ( .A(n6053), .B(n6054), .Z(n6039) );
  XOR U7518 ( .A(n6064), .B(n6065), .Z(n6054) );
  ANDN U7519 ( .B(n6066), .A(n6067), .Z(n6064) );
  XOR U7520 ( .A(n6065), .B(n6068), .Z(n6066) );
  XOR U7521 ( .A(n6069), .B(n6070), .Z(n6053) );
  XOR U7522 ( .A(n6071), .B(n6072), .Z(n6070) );
  ANDN U7523 ( .B(n6073), .A(n6074), .Z(n6071) );
  XOR U7524 ( .A(n6075), .B(n6072), .Z(n6073) );
  IV U7525 ( .A(n6051), .Z(n6069) );
  XOR U7526 ( .A(n6076), .B(n6077), .Z(n6051) );
  ANDN U7527 ( .B(n6078), .A(n6079), .Z(n6076) );
  XOR U7528 ( .A(n6077), .B(n6080), .Z(n6078) );
  IV U7529 ( .A(n6059), .Z(n6063) );
  XOR U7530 ( .A(n6059), .B(n6041), .Z(n6061) );
  XOR U7531 ( .A(n6081), .B(n6082), .Z(n6041) );
  AND U7532 ( .A(n46), .B(n6083), .Z(n6081) );
  XOR U7533 ( .A(n6084), .B(n6082), .Z(n6083) );
  NANDN U7534 ( .A(n6043), .B(n6045), .Z(n6059) );
  XOR U7535 ( .A(n6085), .B(n6086), .Z(n6045) );
  AND U7536 ( .A(n46), .B(n6087), .Z(n6085) );
  XOR U7537 ( .A(n6086), .B(n6088), .Z(n6087) );
  XOR U7538 ( .A(n6089), .B(n6090), .Z(n46) );
  AND U7539 ( .A(n6091), .B(n6092), .Z(n6089) );
  XNOR U7540 ( .A(n6090), .B(n6056), .Z(n6092) );
  XNOR U7541 ( .A(n6093), .B(n6094), .Z(n6056) );
  ANDN U7542 ( .B(n6095), .A(n6096), .Z(n6093) );
  XOR U7543 ( .A(n6094), .B(n6097), .Z(n6095) );
  XOR U7544 ( .A(n6090), .B(n6058), .Z(n6091) );
  XOR U7545 ( .A(n6098), .B(n6099), .Z(n6058) );
  AND U7546 ( .A(n50), .B(n6100), .Z(n6098) );
  XOR U7547 ( .A(n6101), .B(n6099), .Z(n6100) );
  XNOR U7548 ( .A(n6102), .B(n6103), .Z(n6090) );
  NAND U7549 ( .A(n6104), .B(n6105), .Z(n6103) );
  XOR U7550 ( .A(n6106), .B(n6082), .Z(n6105) );
  XOR U7551 ( .A(n6096), .B(n6097), .Z(n6082) );
  XOR U7552 ( .A(n6107), .B(n6108), .Z(n6097) );
  ANDN U7553 ( .B(n6109), .A(n6110), .Z(n6107) );
  XOR U7554 ( .A(n6108), .B(n6111), .Z(n6109) );
  XOR U7555 ( .A(n6112), .B(n6113), .Z(n6096) );
  XOR U7556 ( .A(n6114), .B(n6115), .Z(n6113) );
  ANDN U7557 ( .B(n6116), .A(n6117), .Z(n6114) );
  XOR U7558 ( .A(n6118), .B(n6115), .Z(n6116) );
  IV U7559 ( .A(n6094), .Z(n6112) );
  XOR U7560 ( .A(n6119), .B(n6120), .Z(n6094) );
  ANDN U7561 ( .B(n6121), .A(n6122), .Z(n6119) );
  XOR U7562 ( .A(n6120), .B(n6123), .Z(n6121) );
  IV U7563 ( .A(n6102), .Z(n6106) );
  XOR U7564 ( .A(n6102), .B(n6084), .Z(n6104) );
  XOR U7565 ( .A(n6124), .B(n6125), .Z(n6084) );
  AND U7566 ( .A(n50), .B(n6126), .Z(n6124) );
  XOR U7567 ( .A(n6127), .B(n6125), .Z(n6126) );
  NANDN U7568 ( .A(n6086), .B(n6088), .Z(n6102) );
  XOR U7569 ( .A(n6128), .B(n6129), .Z(n6088) );
  AND U7570 ( .A(n50), .B(n6130), .Z(n6128) );
  XOR U7571 ( .A(n6129), .B(n6131), .Z(n6130) );
  XOR U7572 ( .A(n6132), .B(n6133), .Z(n50) );
  AND U7573 ( .A(n6134), .B(n6135), .Z(n6132) );
  XNOR U7574 ( .A(n6133), .B(n6099), .Z(n6135) );
  XNOR U7575 ( .A(n6136), .B(n6137), .Z(n6099) );
  ANDN U7576 ( .B(n6138), .A(n6139), .Z(n6136) );
  XOR U7577 ( .A(n6137), .B(n6140), .Z(n6138) );
  XOR U7578 ( .A(n6133), .B(n6101), .Z(n6134) );
  XOR U7579 ( .A(n6141), .B(n6142), .Z(n6101) );
  AND U7580 ( .A(n54), .B(n6143), .Z(n6141) );
  XOR U7581 ( .A(n6144), .B(n6142), .Z(n6143) );
  XNOR U7582 ( .A(n6145), .B(n6146), .Z(n6133) );
  NAND U7583 ( .A(n6147), .B(n6148), .Z(n6146) );
  XOR U7584 ( .A(n6149), .B(n6125), .Z(n6148) );
  XOR U7585 ( .A(n6139), .B(n6140), .Z(n6125) );
  XOR U7586 ( .A(n6150), .B(n6151), .Z(n6140) );
  ANDN U7587 ( .B(n6152), .A(n6153), .Z(n6150) );
  XOR U7588 ( .A(n6151), .B(n6154), .Z(n6152) );
  XOR U7589 ( .A(n6155), .B(n6156), .Z(n6139) );
  XOR U7590 ( .A(n6157), .B(n6158), .Z(n6156) );
  ANDN U7591 ( .B(n6159), .A(n6160), .Z(n6157) );
  XOR U7592 ( .A(n6161), .B(n6158), .Z(n6159) );
  IV U7593 ( .A(n6137), .Z(n6155) );
  XOR U7594 ( .A(n6162), .B(n6163), .Z(n6137) );
  ANDN U7595 ( .B(n6164), .A(n6165), .Z(n6162) );
  XOR U7596 ( .A(n6163), .B(n6166), .Z(n6164) );
  IV U7597 ( .A(n6145), .Z(n6149) );
  XOR U7598 ( .A(n6145), .B(n6127), .Z(n6147) );
  XOR U7599 ( .A(n6167), .B(n6168), .Z(n6127) );
  AND U7600 ( .A(n54), .B(n6169), .Z(n6167) );
  XOR U7601 ( .A(n6170), .B(n6168), .Z(n6169) );
  NANDN U7602 ( .A(n6129), .B(n6131), .Z(n6145) );
  XOR U7603 ( .A(n6171), .B(n6172), .Z(n6131) );
  AND U7604 ( .A(n54), .B(n6173), .Z(n6171) );
  XOR U7605 ( .A(n6172), .B(n6174), .Z(n6173) );
  XOR U7606 ( .A(n6175), .B(n6176), .Z(n54) );
  AND U7607 ( .A(n6177), .B(n6178), .Z(n6175) );
  XNOR U7608 ( .A(n6176), .B(n6142), .Z(n6178) );
  XNOR U7609 ( .A(n6179), .B(n6180), .Z(n6142) );
  ANDN U7610 ( .B(n6181), .A(n6182), .Z(n6179) );
  XOR U7611 ( .A(n6180), .B(n6183), .Z(n6181) );
  XOR U7612 ( .A(n6176), .B(n6144), .Z(n6177) );
  XOR U7613 ( .A(n6184), .B(n6185), .Z(n6144) );
  AND U7614 ( .A(n58), .B(n6186), .Z(n6184) );
  XOR U7615 ( .A(n6187), .B(n6185), .Z(n6186) );
  XNOR U7616 ( .A(n6188), .B(n6189), .Z(n6176) );
  NAND U7617 ( .A(n6190), .B(n6191), .Z(n6189) );
  XOR U7618 ( .A(n6192), .B(n6168), .Z(n6191) );
  XOR U7619 ( .A(n6182), .B(n6183), .Z(n6168) );
  XOR U7620 ( .A(n6193), .B(n6194), .Z(n6183) );
  ANDN U7621 ( .B(n6195), .A(n6196), .Z(n6193) );
  XOR U7622 ( .A(n6194), .B(n6197), .Z(n6195) );
  XOR U7623 ( .A(n6198), .B(n6199), .Z(n6182) );
  XOR U7624 ( .A(n6200), .B(n6201), .Z(n6199) );
  ANDN U7625 ( .B(n6202), .A(n6203), .Z(n6200) );
  XOR U7626 ( .A(n6204), .B(n6201), .Z(n6202) );
  IV U7627 ( .A(n6180), .Z(n6198) );
  XOR U7628 ( .A(n6205), .B(n6206), .Z(n6180) );
  ANDN U7629 ( .B(n6207), .A(n6208), .Z(n6205) );
  XOR U7630 ( .A(n6206), .B(n6209), .Z(n6207) );
  IV U7631 ( .A(n6188), .Z(n6192) );
  XOR U7632 ( .A(n6188), .B(n6170), .Z(n6190) );
  XOR U7633 ( .A(n6210), .B(n6211), .Z(n6170) );
  AND U7634 ( .A(n58), .B(n6212), .Z(n6210) );
  XOR U7635 ( .A(n6213), .B(n6211), .Z(n6212) );
  NANDN U7636 ( .A(n6172), .B(n6174), .Z(n6188) );
  XOR U7637 ( .A(n6214), .B(n6215), .Z(n6174) );
  AND U7638 ( .A(n58), .B(n6216), .Z(n6214) );
  XOR U7639 ( .A(n6215), .B(n6217), .Z(n6216) );
  XOR U7640 ( .A(n6218), .B(n6219), .Z(n58) );
  AND U7641 ( .A(n6220), .B(n6221), .Z(n6218) );
  XNOR U7642 ( .A(n6219), .B(n6185), .Z(n6221) );
  XNOR U7643 ( .A(n6222), .B(n6223), .Z(n6185) );
  ANDN U7644 ( .B(n6224), .A(n6225), .Z(n6222) );
  XOR U7645 ( .A(n6223), .B(n6226), .Z(n6224) );
  XOR U7646 ( .A(n6219), .B(n6187), .Z(n6220) );
  XOR U7647 ( .A(n6227), .B(n6228), .Z(n6187) );
  AND U7648 ( .A(n62), .B(n6229), .Z(n6227) );
  XOR U7649 ( .A(n6230), .B(n6228), .Z(n6229) );
  XNOR U7650 ( .A(n6231), .B(n6232), .Z(n6219) );
  NAND U7651 ( .A(n6233), .B(n6234), .Z(n6232) );
  XOR U7652 ( .A(n6235), .B(n6211), .Z(n6234) );
  XOR U7653 ( .A(n6225), .B(n6226), .Z(n6211) );
  XOR U7654 ( .A(n6236), .B(n6237), .Z(n6226) );
  ANDN U7655 ( .B(n6238), .A(n6239), .Z(n6236) );
  XOR U7656 ( .A(n6237), .B(n6240), .Z(n6238) );
  XOR U7657 ( .A(n6241), .B(n6242), .Z(n6225) );
  XOR U7658 ( .A(n6243), .B(n6244), .Z(n6242) );
  ANDN U7659 ( .B(n6245), .A(n6246), .Z(n6243) );
  XOR U7660 ( .A(n6247), .B(n6244), .Z(n6245) );
  IV U7661 ( .A(n6223), .Z(n6241) );
  XOR U7662 ( .A(n6248), .B(n6249), .Z(n6223) );
  ANDN U7663 ( .B(n6250), .A(n6251), .Z(n6248) );
  XOR U7664 ( .A(n6249), .B(n6252), .Z(n6250) );
  IV U7665 ( .A(n6231), .Z(n6235) );
  XOR U7666 ( .A(n6231), .B(n6213), .Z(n6233) );
  XOR U7667 ( .A(n6253), .B(n6254), .Z(n6213) );
  AND U7668 ( .A(n62), .B(n6255), .Z(n6253) );
  XOR U7669 ( .A(n6256), .B(n6254), .Z(n6255) );
  NANDN U7670 ( .A(n6215), .B(n6217), .Z(n6231) );
  XOR U7671 ( .A(n6257), .B(n6258), .Z(n6217) );
  AND U7672 ( .A(n62), .B(n6259), .Z(n6257) );
  XOR U7673 ( .A(n6258), .B(n6260), .Z(n6259) );
  XOR U7674 ( .A(n6261), .B(n6262), .Z(n62) );
  AND U7675 ( .A(n6263), .B(n6264), .Z(n6261) );
  XNOR U7676 ( .A(n6262), .B(n6228), .Z(n6264) );
  XNOR U7677 ( .A(n6265), .B(n6266), .Z(n6228) );
  ANDN U7678 ( .B(n6267), .A(n6268), .Z(n6265) );
  XOR U7679 ( .A(n6266), .B(n6269), .Z(n6267) );
  XOR U7680 ( .A(n6262), .B(n6230), .Z(n6263) );
  XOR U7681 ( .A(n6270), .B(n6271), .Z(n6230) );
  AND U7682 ( .A(n66), .B(n6272), .Z(n6270) );
  XOR U7683 ( .A(n6273), .B(n6271), .Z(n6272) );
  XNOR U7684 ( .A(n6274), .B(n6275), .Z(n6262) );
  NAND U7685 ( .A(n6276), .B(n6277), .Z(n6275) );
  XOR U7686 ( .A(n6278), .B(n6254), .Z(n6277) );
  XOR U7687 ( .A(n6268), .B(n6269), .Z(n6254) );
  XOR U7688 ( .A(n6279), .B(n6280), .Z(n6269) );
  ANDN U7689 ( .B(n6281), .A(n6282), .Z(n6279) );
  XOR U7690 ( .A(n6280), .B(n6283), .Z(n6281) );
  XOR U7691 ( .A(n6284), .B(n6285), .Z(n6268) );
  XOR U7692 ( .A(n6286), .B(n6287), .Z(n6285) );
  ANDN U7693 ( .B(n6288), .A(n6289), .Z(n6286) );
  XOR U7694 ( .A(n6290), .B(n6287), .Z(n6288) );
  IV U7695 ( .A(n6266), .Z(n6284) );
  XOR U7696 ( .A(n6291), .B(n6292), .Z(n6266) );
  ANDN U7697 ( .B(n6293), .A(n6294), .Z(n6291) );
  XOR U7698 ( .A(n6292), .B(n6295), .Z(n6293) );
  IV U7699 ( .A(n6274), .Z(n6278) );
  XOR U7700 ( .A(n6274), .B(n6256), .Z(n6276) );
  XOR U7701 ( .A(n6296), .B(n6297), .Z(n6256) );
  AND U7702 ( .A(n66), .B(n6298), .Z(n6296) );
  XOR U7703 ( .A(n6299), .B(n6297), .Z(n6298) );
  NANDN U7704 ( .A(n6258), .B(n6260), .Z(n6274) );
  XOR U7705 ( .A(n6300), .B(n6301), .Z(n6260) );
  AND U7706 ( .A(n66), .B(n6302), .Z(n6300) );
  XOR U7707 ( .A(n6301), .B(n6303), .Z(n6302) );
  XOR U7708 ( .A(n6304), .B(n6305), .Z(n66) );
  AND U7709 ( .A(n6306), .B(n6307), .Z(n6304) );
  XNOR U7710 ( .A(n6305), .B(n6271), .Z(n6307) );
  XNOR U7711 ( .A(n6308), .B(n6309), .Z(n6271) );
  ANDN U7712 ( .B(n6310), .A(n6311), .Z(n6308) );
  XOR U7713 ( .A(n6309), .B(n6312), .Z(n6310) );
  XOR U7714 ( .A(n6305), .B(n6273), .Z(n6306) );
  XOR U7715 ( .A(n6313), .B(n6314), .Z(n6273) );
  AND U7716 ( .A(n70), .B(n6315), .Z(n6313) );
  XOR U7717 ( .A(n6316), .B(n6314), .Z(n6315) );
  XNOR U7718 ( .A(n6317), .B(n6318), .Z(n6305) );
  NAND U7719 ( .A(n6319), .B(n6320), .Z(n6318) );
  XOR U7720 ( .A(n6321), .B(n6297), .Z(n6320) );
  XOR U7721 ( .A(n6311), .B(n6312), .Z(n6297) );
  XOR U7722 ( .A(n6322), .B(n6323), .Z(n6312) );
  ANDN U7723 ( .B(n6324), .A(n6325), .Z(n6322) );
  XOR U7724 ( .A(n6323), .B(n6326), .Z(n6324) );
  XOR U7725 ( .A(n6327), .B(n6328), .Z(n6311) );
  XOR U7726 ( .A(n6329), .B(n6330), .Z(n6328) );
  ANDN U7727 ( .B(n6331), .A(n6332), .Z(n6329) );
  XOR U7728 ( .A(n6333), .B(n6330), .Z(n6331) );
  IV U7729 ( .A(n6309), .Z(n6327) );
  XOR U7730 ( .A(n6334), .B(n6335), .Z(n6309) );
  ANDN U7731 ( .B(n6336), .A(n6337), .Z(n6334) );
  XOR U7732 ( .A(n6335), .B(n6338), .Z(n6336) );
  IV U7733 ( .A(n6317), .Z(n6321) );
  XOR U7734 ( .A(n6317), .B(n6299), .Z(n6319) );
  XOR U7735 ( .A(n6339), .B(n6340), .Z(n6299) );
  AND U7736 ( .A(n70), .B(n6341), .Z(n6339) );
  XOR U7737 ( .A(n6342), .B(n6340), .Z(n6341) );
  NANDN U7738 ( .A(n6301), .B(n6303), .Z(n6317) );
  XOR U7739 ( .A(n6343), .B(n6344), .Z(n6303) );
  AND U7740 ( .A(n70), .B(n6345), .Z(n6343) );
  XOR U7741 ( .A(n6344), .B(n6346), .Z(n6345) );
  XOR U7742 ( .A(n6347), .B(n6348), .Z(n70) );
  AND U7743 ( .A(n6349), .B(n6350), .Z(n6347) );
  XNOR U7744 ( .A(n6348), .B(n6314), .Z(n6350) );
  XNOR U7745 ( .A(n6351), .B(n6352), .Z(n6314) );
  ANDN U7746 ( .B(n6353), .A(n6354), .Z(n6351) );
  XOR U7747 ( .A(n6352), .B(n6355), .Z(n6353) );
  XOR U7748 ( .A(n6348), .B(n6316), .Z(n6349) );
  XOR U7749 ( .A(n6356), .B(n6357), .Z(n6316) );
  AND U7750 ( .A(n74), .B(n6358), .Z(n6356) );
  XOR U7751 ( .A(n6359), .B(n6357), .Z(n6358) );
  XNOR U7752 ( .A(n6360), .B(n6361), .Z(n6348) );
  NAND U7753 ( .A(n6362), .B(n6363), .Z(n6361) );
  XOR U7754 ( .A(n6364), .B(n6340), .Z(n6363) );
  XOR U7755 ( .A(n6354), .B(n6355), .Z(n6340) );
  XOR U7756 ( .A(n6365), .B(n6366), .Z(n6355) );
  ANDN U7757 ( .B(n6367), .A(n6368), .Z(n6365) );
  XOR U7758 ( .A(n6366), .B(n6369), .Z(n6367) );
  XOR U7759 ( .A(n6370), .B(n6371), .Z(n6354) );
  XOR U7760 ( .A(n6372), .B(n6373), .Z(n6371) );
  ANDN U7761 ( .B(n6374), .A(n6375), .Z(n6372) );
  XOR U7762 ( .A(n6376), .B(n6373), .Z(n6374) );
  IV U7763 ( .A(n6352), .Z(n6370) );
  XOR U7764 ( .A(n6377), .B(n6378), .Z(n6352) );
  ANDN U7765 ( .B(n6379), .A(n6380), .Z(n6377) );
  XOR U7766 ( .A(n6378), .B(n6381), .Z(n6379) );
  IV U7767 ( .A(n6360), .Z(n6364) );
  XOR U7768 ( .A(n6360), .B(n6342), .Z(n6362) );
  XOR U7769 ( .A(n6382), .B(n6383), .Z(n6342) );
  AND U7770 ( .A(n74), .B(n6384), .Z(n6382) );
  XOR U7771 ( .A(n6385), .B(n6383), .Z(n6384) );
  NANDN U7772 ( .A(n6344), .B(n6346), .Z(n6360) );
  XOR U7773 ( .A(n6386), .B(n6387), .Z(n6346) );
  AND U7774 ( .A(n74), .B(n6388), .Z(n6386) );
  XOR U7775 ( .A(n6387), .B(n6389), .Z(n6388) );
  XOR U7776 ( .A(n6390), .B(n6391), .Z(n74) );
  AND U7777 ( .A(n6392), .B(n6393), .Z(n6390) );
  XNOR U7778 ( .A(n6391), .B(n6357), .Z(n6393) );
  XNOR U7779 ( .A(n6394), .B(n6395), .Z(n6357) );
  ANDN U7780 ( .B(n6396), .A(n6397), .Z(n6394) );
  XOR U7781 ( .A(n6395), .B(n6398), .Z(n6396) );
  XOR U7782 ( .A(n6391), .B(n6359), .Z(n6392) );
  XOR U7783 ( .A(n6399), .B(n6400), .Z(n6359) );
  AND U7784 ( .A(n78), .B(n6401), .Z(n6399) );
  XOR U7785 ( .A(n6402), .B(n6400), .Z(n6401) );
  XNOR U7786 ( .A(n6403), .B(n6404), .Z(n6391) );
  NAND U7787 ( .A(n6405), .B(n6406), .Z(n6404) );
  XOR U7788 ( .A(n6407), .B(n6383), .Z(n6406) );
  XOR U7789 ( .A(n6397), .B(n6398), .Z(n6383) );
  XOR U7790 ( .A(n6408), .B(n6409), .Z(n6398) );
  ANDN U7791 ( .B(n6410), .A(n6411), .Z(n6408) );
  XOR U7792 ( .A(n6409), .B(n6412), .Z(n6410) );
  XOR U7793 ( .A(n6413), .B(n6414), .Z(n6397) );
  XOR U7794 ( .A(n6415), .B(n6416), .Z(n6414) );
  ANDN U7795 ( .B(n6417), .A(n6418), .Z(n6415) );
  XOR U7796 ( .A(n6419), .B(n6416), .Z(n6417) );
  IV U7797 ( .A(n6395), .Z(n6413) );
  XOR U7798 ( .A(n6420), .B(n6421), .Z(n6395) );
  ANDN U7799 ( .B(n6422), .A(n6423), .Z(n6420) );
  XOR U7800 ( .A(n6421), .B(n6424), .Z(n6422) );
  IV U7801 ( .A(n6403), .Z(n6407) );
  XOR U7802 ( .A(n6403), .B(n6385), .Z(n6405) );
  XOR U7803 ( .A(n6425), .B(n6426), .Z(n6385) );
  AND U7804 ( .A(n78), .B(n6427), .Z(n6425) );
  XOR U7805 ( .A(n6428), .B(n6426), .Z(n6427) );
  NANDN U7806 ( .A(n6387), .B(n6389), .Z(n6403) );
  XOR U7807 ( .A(n6429), .B(n6430), .Z(n6389) );
  AND U7808 ( .A(n78), .B(n6431), .Z(n6429) );
  XOR U7809 ( .A(n6430), .B(n6432), .Z(n6431) );
  XOR U7810 ( .A(n6433), .B(n6434), .Z(n78) );
  AND U7811 ( .A(n6435), .B(n6436), .Z(n6433) );
  XNOR U7812 ( .A(n6434), .B(n6400), .Z(n6436) );
  XNOR U7813 ( .A(n6437), .B(n6438), .Z(n6400) );
  ANDN U7814 ( .B(n6439), .A(n6440), .Z(n6437) );
  XOR U7815 ( .A(n6438), .B(n6441), .Z(n6439) );
  XOR U7816 ( .A(n6434), .B(n6402), .Z(n6435) );
  XOR U7817 ( .A(n6442), .B(n6443), .Z(n6402) );
  AND U7818 ( .A(n82), .B(n6444), .Z(n6442) );
  XOR U7819 ( .A(n6445), .B(n6443), .Z(n6444) );
  XNOR U7820 ( .A(n6446), .B(n6447), .Z(n6434) );
  NAND U7821 ( .A(n6448), .B(n6449), .Z(n6447) );
  XOR U7822 ( .A(n6450), .B(n6426), .Z(n6449) );
  XOR U7823 ( .A(n6440), .B(n6441), .Z(n6426) );
  XOR U7824 ( .A(n6451), .B(n6452), .Z(n6441) );
  ANDN U7825 ( .B(n6453), .A(n6454), .Z(n6451) );
  XOR U7826 ( .A(n6452), .B(n6455), .Z(n6453) );
  XOR U7827 ( .A(n6456), .B(n6457), .Z(n6440) );
  XOR U7828 ( .A(n6458), .B(n6459), .Z(n6457) );
  ANDN U7829 ( .B(n6460), .A(n6461), .Z(n6458) );
  XOR U7830 ( .A(n6462), .B(n6459), .Z(n6460) );
  IV U7831 ( .A(n6438), .Z(n6456) );
  XOR U7832 ( .A(n6463), .B(n6464), .Z(n6438) );
  ANDN U7833 ( .B(n6465), .A(n6466), .Z(n6463) );
  XOR U7834 ( .A(n6464), .B(n6467), .Z(n6465) );
  IV U7835 ( .A(n6446), .Z(n6450) );
  XOR U7836 ( .A(n6446), .B(n6428), .Z(n6448) );
  XOR U7837 ( .A(n6468), .B(n6469), .Z(n6428) );
  AND U7838 ( .A(n82), .B(n6470), .Z(n6468) );
  XOR U7839 ( .A(n6471), .B(n6469), .Z(n6470) );
  NANDN U7840 ( .A(n6430), .B(n6432), .Z(n6446) );
  XOR U7841 ( .A(n6472), .B(n6473), .Z(n6432) );
  AND U7842 ( .A(n82), .B(n6474), .Z(n6472) );
  XOR U7843 ( .A(n6473), .B(n6475), .Z(n6474) );
  XOR U7844 ( .A(n6476), .B(n6477), .Z(n82) );
  AND U7845 ( .A(n6478), .B(n6479), .Z(n6476) );
  XNOR U7846 ( .A(n6477), .B(n6443), .Z(n6479) );
  XNOR U7847 ( .A(n6480), .B(n6481), .Z(n6443) );
  ANDN U7848 ( .B(n6482), .A(n6483), .Z(n6480) );
  XOR U7849 ( .A(n6481), .B(n6484), .Z(n6482) );
  XOR U7850 ( .A(n6477), .B(n6445), .Z(n6478) );
  XOR U7851 ( .A(n6485), .B(n6486), .Z(n6445) );
  AND U7852 ( .A(n86), .B(n6487), .Z(n6485) );
  XOR U7853 ( .A(n6488), .B(n6486), .Z(n6487) );
  XNOR U7854 ( .A(n6489), .B(n6490), .Z(n6477) );
  NAND U7855 ( .A(n6491), .B(n6492), .Z(n6490) );
  XOR U7856 ( .A(n6493), .B(n6469), .Z(n6492) );
  XOR U7857 ( .A(n6483), .B(n6484), .Z(n6469) );
  XOR U7858 ( .A(n6494), .B(n6495), .Z(n6484) );
  ANDN U7859 ( .B(n6496), .A(n6497), .Z(n6494) );
  XOR U7860 ( .A(n6495), .B(n6498), .Z(n6496) );
  XOR U7861 ( .A(n6499), .B(n6500), .Z(n6483) );
  XOR U7862 ( .A(n6501), .B(n6502), .Z(n6500) );
  ANDN U7863 ( .B(n6503), .A(n6504), .Z(n6501) );
  XOR U7864 ( .A(n6505), .B(n6502), .Z(n6503) );
  IV U7865 ( .A(n6481), .Z(n6499) );
  XOR U7866 ( .A(n6506), .B(n6507), .Z(n6481) );
  ANDN U7867 ( .B(n6508), .A(n6509), .Z(n6506) );
  XOR U7868 ( .A(n6507), .B(n6510), .Z(n6508) );
  IV U7869 ( .A(n6489), .Z(n6493) );
  XOR U7870 ( .A(n6489), .B(n6471), .Z(n6491) );
  XOR U7871 ( .A(n6511), .B(n6512), .Z(n6471) );
  AND U7872 ( .A(n86), .B(n6513), .Z(n6511) );
  XOR U7873 ( .A(n6514), .B(n6512), .Z(n6513) );
  NANDN U7874 ( .A(n6473), .B(n6475), .Z(n6489) );
  XOR U7875 ( .A(n6515), .B(n6516), .Z(n6475) );
  AND U7876 ( .A(n86), .B(n6517), .Z(n6515) );
  XOR U7877 ( .A(n6516), .B(n6518), .Z(n6517) );
  XOR U7878 ( .A(n6519), .B(n6520), .Z(n86) );
  AND U7879 ( .A(n6521), .B(n6522), .Z(n6519) );
  XNOR U7880 ( .A(n6520), .B(n6486), .Z(n6522) );
  XNOR U7881 ( .A(n6523), .B(n6524), .Z(n6486) );
  ANDN U7882 ( .B(n6525), .A(n6526), .Z(n6523) );
  XOR U7883 ( .A(n6524), .B(n6527), .Z(n6525) );
  XOR U7884 ( .A(n6520), .B(n6488), .Z(n6521) );
  XOR U7885 ( .A(n6528), .B(n6529), .Z(n6488) );
  AND U7886 ( .A(n90), .B(n6530), .Z(n6528) );
  XOR U7887 ( .A(n6531), .B(n6529), .Z(n6530) );
  XNOR U7888 ( .A(n6532), .B(n6533), .Z(n6520) );
  NAND U7889 ( .A(n6534), .B(n6535), .Z(n6533) );
  XOR U7890 ( .A(n6536), .B(n6512), .Z(n6535) );
  XOR U7891 ( .A(n6526), .B(n6527), .Z(n6512) );
  XOR U7892 ( .A(n6537), .B(n6538), .Z(n6527) );
  ANDN U7893 ( .B(n6539), .A(n6540), .Z(n6537) );
  XOR U7894 ( .A(n6538), .B(n6541), .Z(n6539) );
  XOR U7895 ( .A(n6542), .B(n6543), .Z(n6526) );
  XOR U7896 ( .A(n6544), .B(n6545), .Z(n6543) );
  ANDN U7897 ( .B(n6546), .A(n6547), .Z(n6544) );
  XOR U7898 ( .A(n6548), .B(n6545), .Z(n6546) );
  IV U7899 ( .A(n6524), .Z(n6542) );
  XOR U7900 ( .A(n6549), .B(n6550), .Z(n6524) );
  ANDN U7901 ( .B(n6551), .A(n6552), .Z(n6549) );
  XOR U7902 ( .A(n6550), .B(n6553), .Z(n6551) );
  IV U7903 ( .A(n6532), .Z(n6536) );
  XOR U7904 ( .A(n6532), .B(n6514), .Z(n6534) );
  XOR U7905 ( .A(n6554), .B(n6555), .Z(n6514) );
  AND U7906 ( .A(n90), .B(n6556), .Z(n6554) );
  XOR U7907 ( .A(n6557), .B(n6555), .Z(n6556) );
  NANDN U7908 ( .A(n6516), .B(n6518), .Z(n6532) );
  XOR U7909 ( .A(n6558), .B(n6559), .Z(n6518) );
  AND U7910 ( .A(n90), .B(n6560), .Z(n6558) );
  XOR U7911 ( .A(n6559), .B(n6561), .Z(n6560) );
  XOR U7912 ( .A(n6562), .B(n6563), .Z(n90) );
  AND U7913 ( .A(n6564), .B(n6565), .Z(n6562) );
  XNOR U7914 ( .A(n6563), .B(n6529), .Z(n6565) );
  XNOR U7915 ( .A(n6566), .B(n6567), .Z(n6529) );
  ANDN U7916 ( .B(n6568), .A(n6569), .Z(n6566) );
  XOR U7917 ( .A(n6567), .B(n6570), .Z(n6568) );
  XOR U7918 ( .A(n6563), .B(n6531), .Z(n6564) );
  XOR U7919 ( .A(n6571), .B(n6572), .Z(n6531) );
  AND U7920 ( .A(n94), .B(n6573), .Z(n6571) );
  XOR U7921 ( .A(n6574), .B(n6572), .Z(n6573) );
  XNOR U7922 ( .A(n6575), .B(n6576), .Z(n6563) );
  NAND U7923 ( .A(n6577), .B(n6578), .Z(n6576) );
  XOR U7924 ( .A(n6579), .B(n6555), .Z(n6578) );
  XOR U7925 ( .A(n6569), .B(n6570), .Z(n6555) );
  XOR U7926 ( .A(n6580), .B(n6581), .Z(n6570) );
  ANDN U7927 ( .B(n6582), .A(n6583), .Z(n6580) );
  XOR U7928 ( .A(n6581), .B(n6584), .Z(n6582) );
  XOR U7929 ( .A(n6585), .B(n6586), .Z(n6569) );
  XOR U7930 ( .A(n6587), .B(n6588), .Z(n6586) );
  ANDN U7931 ( .B(n6589), .A(n6590), .Z(n6587) );
  XOR U7932 ( .A(n6591), .B(n6588), .Z(n6589) );
  IV U7933 ( .A(n6567), .Z(n6585) );
  XOR U7934 ( .A(n6592), .B(n6593), .Z(n6567) );
  ANDN U7935 ( .B(n6594), .A(n6595), .Z(n6592) );
  XOR U7936 ( .A(n6593), .B(n6596), .Z(n6594) );
  IV U7937 ( .A(n6575), .Z(n6579) );
  XOR U7938 ( .A(n6575), .B(n6557), .Z(n6577) );
  XOR U7939 ( .A(n6597), .B(n6598), .Z(n6557) );
  AND U7940 ( .A(n94), .B(n6599), .Z(n6597) );
  XOR U7941 ( .A(n6600), .B(n6598), .Z(n6599) );
  NANDN U7942 ( .A(n6559), .B(n6561), .Z(n6575) );
  XOR U7943 ( .A(n6601), .B(n6602), .Z(n6561) );
  AND U7944 ( .A(n94), .B(n6603), .Z(n6601) );
  XOR U7945 ( .A(n6602), .B(n6604), .Z(n6603) );
  XOR U7946 ( .A(n6605), .B(n6606), .Z(n94) );
  AND U7947 ( .A(n6607), .B(n6608), .Z(n6605) );
  XNOR U7948 ( .A(n6606), .B(n6572), .Z(n6608) );
  XNOR U7949 ( .A(n6609), .B(n6610), .Z(n6572) );
  ANDN U7950 ( .B(n6611), .A(n6612), .Z(n6609) );
  XOR U7951 ( .A(n6610), .B(n6613), .Z(n6611) );
  XOR U7952 ( .A(n6606), .B(n6574), .Z(n6607) );
  XOR U7953 ( .A(n6614), .B(n6615), .Z(n6574) );
  AND U7954 ( .A(n98), .B(n6616), .Z(n6614) );
  XOR U7955 ( .A(n6617), .B(n6615), .Z(n6616) );
  XNOR U7956 ( .A(n6618), .B(n6619), .Z(n6606) );
  NAND U7957 ( .A(n6620), .B(n6621), .Z(n6619) );
  XOR U7958 ( .A(n6622), .B(n6598), .Z(n6621) );
  XOR U7959 ( .A(n6612), .B(n6613), .Z(n6598) );
  XOR U7960 ( .A(n6623), .B(n6624), .Z(n6613) );
  ANDN U7961 ( .B(n6625), .A(n6626), .Z(n6623) );
  XOR U7962 ( .A(n6624), .B(n6627), .Z(n6625) );
  XOR U7963 ( .A(n6628), .B(n6629), .Z(n6612) );
  XOR U7964 ( .A(n6630), .B(n6631), .Z(n6629) );
  ANDN U7965 ( .B(n6632), .A(n6633), .Z(n6630) );
  XOR U7966 ( .A(n6634), .B(n6631), .Z(n6632) );
  IV U7967 ( .A(n6610), .Z(n6628) );
  XOR U7968 ( .A(n6635), .B(n6636), .Z(n6610) );
  ANDN U7969 ( .B(n6637), .A(n6638), .Z(n6635) );
  XOR U7970 ( .A(n6636), .B(n6639), .Z(n6637) );
  IV U7971 ( .A(n6618), .Z(n6622) );
  XOR U7972 ( .A(n6618), .B(n6600), .Z(n6620) );
  XOR U7973 ( .A(n6640), .B(n6641), .Z(n6600) );
  AND U7974 ( .A(n98), .B(n6642), .Z(n6640) );
  XOR U7975 ( .A(n6643), .B(n6641), .Z(n6642) );
  NANDN U7976 ( .A(n6602), .B(n6604), .Z(n6618) );
  XOR U7977 ( .A(n6644), .B(n6645), .Z(n6604) );
  AND U7978 ( .A(n98), .B(n6646), .Z(n6644) );
  XOR U7979 ( .A(n6645), .B(n6647), .Z(n6646) );
  XOR U7980 ( .A(n6648), .B(n6649), .Z(n98) );
  AND U7981 ( .A(n6650), .B(n6651), .Z(n6648) );
  XNOR U7982 ( .A(n6649), .B(n6615), .Z(n6651) );
  XNOR U7983 ( .A(n6652), .B(n6653), .Z(n6615) );
  ANDN U7984 ( .B(n6654), .A(n6655), .Z(n6652) );
  XOR U7985 ( .A(n6653), .B(n6656), .Z(n6654) );
  XOR U7986 ( .A(n6649), .B(n6617), .Z(n6650) );
  XOR U7987 ( .A(n6657), .B(n6658), .Z(n6617) );
  AND U7988 ( .A(n102), .B(n6659), .Z(n6657) );
  XOR U7989 ( .A(n6660), .B(n6658), .Z(n6659) );
  XNOR U7990 ( .A(n6661), .B(n6662), .Z(n6649) );
  NAND U7991 ( .A(n6663), .B(n6664), .Z(n6662) );
  XOR U7992 ( .A(n6665), .B(n6641), .Z(n6664) );
  XOR U7993 ( .A(n6655), .B(n6656), .Z(n6641) );
  XOR U7994 ( .A(n6666), .B(n6667), .Z(n6656) );
  ANDN U7995 ( .B(n6668), .A(n6669), .Z(n6666) );
  XOR U7996 ( .A(n6667), .B(n6670), .Z(n6668) );
  XOR U7997 ( .A(n6671), .B(n6672), .Z(n6655) );
  XOR U7998 ( .A(n6673), .B(n6674), .Z(n6672) );
  ANDN U7999 ( .B(n6675), .A(n6676), .Z(n6673) );
  XOR U8000 ( .A(n6677), .B(n6674), .Z(n6675) );
  IV U8001 ( .A(n6653), .Z(n6671) );
  XOR U8002 ( .A(n6678), .B(n6679), .Z(n6653) );
  ANDN U8003 ( .B(n6680), .A(n6681), .Z(n6678) );
  XOR U8004 ( .A(n6679), .B(n6682), .Z(n6680) );
  IV U8005 ( .A(n6661), .Z(n6665) );
  XOR U8006 ( .A(n6661), .B(n6643), .Z(n6663) );
  XOR U8007 ( .A(n6683), .B(n6684), .Z(n6643) );
  AND U8008 ( .A(n102), .B(n6685), .Z(n6683) );
  XOR U8009 ( .A(n6686), .B(n6684), .Z(n6685) );
  NANDN U8010 ( .A(n6645), .B(n6647), .Z(n6661) );
  XOR U8011 ( .A(n6687), .B(n6688), .Z(n6647) );
  AND U8012 ( .A(n102), .B(n6689), .Z(n6687) );
  XOR U8013 ( .A(n6688), .B(n6690), .Z(n6689) );
  XOR U8014 ( .A(n6691), .B(n6692), .Z(n102) );
  AND U8015 ( .A(n6693), .B(n6694), .Z(n6691) );
  XNOR U8016 ( .A(n6692), .B(n6658), .Z(n6694) );
  XNOR U8017 ( .A(n6695), .B(n6696), .Z(n6658) );
  ANDN U8018 ( .B(n6697), .A(n6698), .Z(n6695) );
  XOR U8019 ( .A(n6696), .B(n6699), .Z(n6697) );
  XOR U8020 ( .A(n6692), .B(n6660), .Z(n6693) );
  XOR U8021 ( .A(n6700), .B(n6701), .Z(n6660) );
  AND U8022 ( .A(n106), .B(n6702), .Z(n6700) );
  XOR U8023 ( .A(n6703), .B(n6701), .Z(n6702) );
  XNOR U8024 ( .A(n6704), .B(n6705), .Z(n6692) );
  NAND U8025 ( .A(n6706), .B(n6707), .Z(n6705) );
  XOR U8026 ( .A(n6708), .B(n6684), .Z(n6707) );
  XOR U8027 ( .A(n6698), .B(n6699), .Z(n6684) );
  XOR U8028 ( .A(n6709), .B(n6710), .Z(n6699) );
  ANDN U8029 ( .B(n6711), .A(n6712), .Z(n6709) );
  XOR U8030 ( .A(n6710), .B(n6713), .Z(n6711) );
  XOR U8031 ( .A(n6714), .B(n6715), .Z(n6698) );
  XOR U8032 ( .A(n6716), .B(n6717), .Z(n6715) );
  ANDN U8033 ( .B(n6718), .A(n6719), .Z(n6716) );
  XOR U8034 ( .A(n6720), .B(n6717), .Z(n6718) );
  IV U8035 ( .A(n6696), .Z(n6714) );
  XOR U8036 ( .A(n6721), .B(n6722), .Z(n6696) );
  ANDN U8037 ( .B(n6723), .A(n6724), .Z(n6721) );
  XOR U8038 ( .A(n6722), .B(n6725), .Z(n6723) );
  IV U8039 ( .A(n6704), .Z(n6708) );
  XOR U8040 ( .A(n6704), .B(n6686), .Z(n6706) );
  XOR U8041 ( .A(n6726), .B(n6727), .Z(n6686) );
  AND U8042 ( .A(n106), .B(n6728), .Z(n6726) );
  XOR U8043 ( .A(n6729), .B(n6727), .Z(n6728) );
  NANDN U8044 ( .A(n6688), .B(n6690), .Z(n6704) );
  XOR U8045 ( .A(n6730), .B(n6731), .Z(n6690) );
  AND U8046 ( .A(n106), .B(n6732), .Z(n6730) );
  XOR U8047 ( .A(n6731), .B(n6733), .Z(n6732) );
  XOR U8048 ( .A(n6734), .B(n6735), .Z(n106) );
  AND U8049 ( .A(n6736), .B(n6737), .Z(n6734) );
  XNOR U8050 ( .A(n6735), .B(n6701), .Z(n6737) );
  XNOR U8051 ( .A(n6738), .B(n6739), .Z(n6701) );
  ANDN U8052 ( .B(n6740), .A(n6741), .Z(n6738) );
  XOR U8053 ( .A(n6739), .B(n6742), .Z(n6740) );
  XOR U8054 ( .A(n6735), .B(n6703), .Z(n6736) );
  XOR U8055 ( .A(n6743), .B(n6744), .Z(n6703) );
  AND U8056 ( .A(n110), .B(n6745), .Z(n6743) );
  XOR U8057 ( .A(n6746), .B(n6744), .Z(n6745) );
  XNOR U8058 ( .A(n6747), .B(n6748), .Z(n6735) );
  NAND U8059 ( .A(n6749), .B(n6750), .Z(n6748) );
  XOR U8060 ( .A(n6751), .B(n6727), .Z(n6750) );
  XOR U8061 ( .A(n6741), .B(n6742), .Z(n6727) );
  XOR U8062 ( .A(n6752), .B(n6753), .Z(n6742) );
  ANDN U8063 ( .B(n6754), .A(n6755), .Z(n6752) );
  XOR U8064 ( .A(n6753), .B(n6756), .Z(n6754) );
  XOR U8065 ( .A(n6757), .B(n6758), .Z(n6741) );
  XOR U8066 ( .A(n6759), .B(n6760), .Z(n6758) );
  ANDN U8067 ( .B(n6761), .A(n6762), .Z(n6759) );
  XOR U8068 ( .A(n6763), .B(n6760), .Z(n6761) );
  IV U8069 ( .A(n6739), .Z(n6757) );
  XOR U8070 ( .A(n6764), .B(n6765), .Z(n6739) );
  ANDN U8071 ( .B(n6766), .A(n6767), .Z(n6764) );
  XOR U8072 ( .A(n6765), .B(n6768), .Z(n6766) );
  IV U8073 ( .A(n6747), .Z(n6751) );
  XOR U8074 ( .A(n6747), .B(n6729), .Z(n6749) );
  XOR U8075 ( .A(n6769), .B(n6770), .Z(n6729) );
  AND U8076 ( .A(n110), .B(n6771), .Z(n6769) );
  XOR U8077 ( .A(n6772), .B(n6770), .Z(n6771) );
  NANDN U8078 ( .A(n6731), .B(n6733), .Z(n6747) );
  XOR U8079 ( .A(n6773), .B(n6774), .Z(n6733) );
  AND U8080 ( .A(n110), .B(n6775), .Z(n6773) );
  XOR U8081 ( .A(n6774), .B(n6776), .Z(n6775) );
  XOR U8082 ( .A(n6777), .B(n6778), .Z(n110) );
  AND U8083 ( .A(n6779), .B(n6780), .Z(n6777) );
  XNOR U8084 ( .A(n6778), .B(n6744), .Z(n6780) );
  XNOR U8085 ( .A(n6781), .B(n6782), .Z(n6744) );
  ANDN U8086 ( .B(n6783), .A(n6784), .Z(n6781) );
  XOR U8087 ( .A(n6782), .B(n6785), .Z(n6783) );
  XOR U8088 ( .A(n6778), .B(n6746), .Z(n6779) );
  XOR U8089 ( .A(n6786), .B(n6787), .Z(n6746) );
  AND U8090 ( .A(n114), .B(n6788), .Z(n6786) );
  XOR U8091 ( .A(n6789), .B(n6787), .Z(n6788) );
  XNOR U8092 ( .A(n6790), .B(n6791), .Z(n6778) );
  NAND U8093 ( .A(n6792), .B(n6793), .Z(n6791) );
  XOR U8094 ( .A(n6794), .B(n6770), .Z(n6793) );
  XOR U8095 ( .A(n6784), .B(n6785), .Z(n6770) );
  XOR U8096 ( .A(n6795), .B(n6796), .Z(n6785) );
  ANDN U8097 ( .B(n6797), .A(n6798), .Z(n6795) );
  XOR U8098 ( .A(n6796), .B(n6799), .Z(n6797) );
  XOR U8099 ( .A(n6800), .B(n6801), .Z(n6784) );
  XOR U8100 ( .A(n6802), .B(n6803), .Z(n6801) );
  ANDN U8101 ( .B(n6804), .A(n6805), .Z(n6802) );
  XOR U8102 ( .A(n6806), .B(n6803), .Z(n6804) );
  IV U8103 ( .A(n6782), .Z(n6800) );
  XOR U8104 ( .A(n6807), .B(n6808), .Z(n6782) );
  ANDN U8105 ( .B(n6809), .A(n6810), .Z(n6807) );
  XOR U8106 ( .A(n6808), .B(n6811), .Z(n6809) );
  IV U8107 ( .A(n6790), .Z(n6794) );
  XOR U8108 ( .A(n6790), .B(n6772), .Z(n6792) );
  XOR U8109 ( .A(n6812), .B(n6813), .Z(n6772) );
  AND U8110 ( .A(n114), .B(n6814), .Z(n6812) );
  XOR U8111 ( .A(n6815), .B(n6813), .Z(n6814) );
  NANDN U8112 ( .A(n6774), .B(n6776), .Z(n6790) );
  XOR U8113 ( .A(n6816), .B(n6817), .Z(n6776) );
  AND U8114 ( .A(n114), .B(n6818), .Z(n6816) );
  XOR U8115 ( .A(n6817), .B(n6819), .Z(n6818) );
  XOR U8116 ( .A(n6820), .B(n6821), .Z(n114) );
  AND U8117 ( .A(n6822), .B(n6823), .Z(n6820) );
  XNOR U8118 ( .A(n6821), .B(n6787), .Z(n6823) );
  XNOR U8119 ( .A(n6824), .B(n6825), .Z(n6787) );
  ANDN U8120 ( .B(n6826), .A(n6827), .Z(n6824) );
  XOR U8121 ( .A(n6825), .B(n6828), .Z(n6826) );
  XOR U8122 ( .A(n6821), .B(n6789), .Z(n6822) );
  XOR U8123 ( .A(n6829), .B(n6830), .Z(n6789) );
  AND U8124 ( .A(n118), .B(n6831), .Z(n6829) );
  XOR U8125 ( .A(n6832), .B(n6830), .Z(n6831) );
  XNOR U8126 ( .A(n6833), .B(n6834), .Z(n6821) );
  NAND U8127 ( .A(n6835), .B(n6836), .Z(n6834) );
  XOR U8128 ( .A(n6837), .B(n6813), .Z(n6836) );
  XOR U8129 ( .A(n6827), .B(n6828), .Z(n6813) );
  XOR U8130 ( .A(n6838), .B(n6839), .Z(n6828) );
  ANDN U8131 ( .B(n6840), .A(n6841), .Z(n6838) );
  XOR U8132 ( .A(n6839), .B(n6842), .Z(n6840) );
  XOR U8133 ( .A(n6843), .B(n6844), .Z(n6827) );
  XOR U8134 ( .A(n6845), .B(n6846), .Z(n6844) );
  ANDN U8135 ( .B(n6847), .A(n6848), .Z(n6845) );
  XOR U8136 ( .A(n6849), .B(n6846), .Z(n6847) );
  IV U8137 ( .A(n6825), .Z(n6843) );
  XOR U8138 ( .A(n6850), .B(n6851), .Z(n6825) );
  ANDN U8139 ( .B(n6852), .A(n6853), .Z(n6850) );
  XOR U8140 ( .A(n6851), .B(n6854), .Z(n6852) );
  IV U8141 ( .A(n6833), .Z(n6837) );
  XOR U8142 ( .A(n6833), .B(n6815), .Z(n6835) );
  XOR U8143 ( .A(n6855), .B(n6856), .Z(n6815) );
  AND U8144 ( .A(n118), .B(n6857), .Z(n6855) );
  XOR U8145 ( .A(n6858), .B(n6856), .Z(n6857) );
  NANDN U8146 ( .A(n6817), .B(n6819), .Z(n6833) );
  XOR U8147 ( .A(n6859), .B(n6860), .Z(n6819) );
  AND U8148 ( .A(n118), .B(n6861), .Z(n6859) );
  XOR U8149 ( .A(n6860), .B(n6862), .Z(n6861) );
  XOR U8150 ( .A(n6863), .B(n6864), .Z(n118) );
  AND U8151 ( .A(n6865), .B(n6866), .Z(n6863) );
  XNOR U8152 ( .A(n6864), .B(n6830), .Z(n6866) );
  XNOR U8153 ( .A(n6867), .B(n6868), .Z(n6830) );
  ANDN U8154 ( .B(n6869), .A(n6870), .Z(n6867) );
  XOR U8155 ( .A(n6868), .B(n6871), .Z(n6869) );
  XOR U8156 ( .A(n6864), .B(n6832), .Z(n6865) );
  XOR U8157 ( .A(n6872), .B(n6873), .Z(n6832) );
  AND U8158 ( .A(n122), .B(n6874), .Z(n6872) );
  XOR U8159 ( .A(n6875), .B(n6873), .Z(n6874) );
  XNOR U8160 ( .A(n6876), .B(n6877), .Z(n6864) );
  NAND U8161 ( .A(n6878), .B(n6879), .Z(n6877) );
  XOR U8162 ( .A(n6880), .B(n6856), .Z(n6879) );
  XOR U8163 ( .A(n6870), .B(n6871), .Z(n6856) );
  XOR U8164 ( .A(n6881), .B(n6882), .Z(n6871) );
  ANDN U8165 ( .B(n6883), .A(n6884), .Z(n6881) );
  XOR U8166 ( .A(n6882), .B(n6885), .Z(n6883) );
  XOR U8167 ( .A(n6886), .B(n6887), .Z(n6870) );
  XOR U8168 ( .A(n6888), .B(n6889), .Z(n6887) );
  ANDN U8169 ( .B(n6890), .A(n6891), .Z(n6888) );
  XOR U8170 ( .A(n6892), .B(n6889), .Z(n6890) );
  IV U8171 ( .A(n6868), .Z(n6886) );
  XOR U8172 ( .A(n6893), .B(n6894), .Z(n6868) );
  ANDN U8173 ( .B(n6895), .A(n6896), .Z(n6893) );
  XOR U8174 ( .A(n6894), .B(n6897), .Z(n6895) );
  IV U8175 ( .A(n6876), .Z(n6880) );
  XOR U8176 ( .A(n6876), .B(n6858), .Z(n6878) );
  XOR U8177 ( .A(n6898), .B(n6899), .Z(n6858) );
  AND U8178 ( .A(n122), .B(n6900), .Z(n6898) );
  XOR U8179 ( .A(n6901), .B(n6899), .Z(n6900) );
  NANDN U8180 ( .A(n6860), .B(n6862), .Z(n6876) );
  XOR U8181 ( .A(n6902), .B(n6903), .Z(n6862) );
  AND U8182 ( .A(n122), .B(n6904), .Z(n6902) );
  XOR U8183 ( .A(n6903), .B(n6905), .Z(n6904) );
  XOR U8184 ( .A(n6906), .B(n6907), .Z(n122) );
  AND U8185 ( .A(n6908), .B(n6909), .Z(n6906) );
  XNOR U8186 ( .A(n6907), .B(n6873), .Z(n6909) );
  XNOR U8187 ( .A(n6910), .B(n6911), .Z(n6873) );
  ANDN U8188 ( .B(n6912), .A(n6913), .Z(n6910) );
  XOR U8189 ( .A(n6911), .B(n6914), .Z(n6912) );
  XOR U8190 ( .A(n6907), .B(n6875), .Z(n6908) );
  XOR U8191 ( .A(n6915), .B(n6916), .Z(n6875) );
  AND U8192 ( .A(n126), .B(n6917), .Z(n6915) );
  XOR U8193 ( .A(n6918), .B(n6916), .Z(n6917) );
  XNOR U8194 ( .A(n6919), .B(n6920), .Z(n6907) );
  NAND U8195 ( .A(n6921), .B(n6922), .Z(n6920) );
  XOR U8196 ( .A(n6923), .B(n6899), .Z(n6922) );
  XOR U8197 ( .A(n6913), .B(n6914), .Z(n6899) );
  XOR U8198 ( .A(n6924), .B(n6925), .Z(n6914) );
  ANDN U8199 ( .B(n6926), .A(n6927), .Z(n6924) );
  XOR U8200 ( .A(n6925), .B(n6928), .Z(n6926) );
  XOR U8201 ( .A(n6929), .B(n6930), .Z(n6913) );
  XOR U8202 ( .A(n6931), .B(n6932), .Z(n6930) );
  ANDN U8203 ( .B(n6933), .A(n6934), .Z(n6931) );
  XOR U8204 ( .A(n6935), .B(n6932), .Z(n6933) );
  IV U8205 ( .A(n6911), .Z(n6929) );
  XOR U8206 ( .A(n6936), .B(n6937), .Z(n6911) );
  ANDN U8207 ( .B(n6938), .A(n6939), .Z(n6936) );
  XOR U8208 ( .A(n6937), .B(n6940), .Z(n6938) );
  IV U8209 ( .A(n6919), .Z(n6923) );
  XOR U8210 ( .A(n6919), .B(n6901), .Z(n6921) );
  XOR U8211 ( .A(n6941), .B(n6942), .Z(n6901) );
  AND U8212 ( .A(n126), .B(n6943), .Z(n6941) );
  XOR U8213 ( .A(n6944), .B(n6942), .Z(n6943) );
  NANDN U8214 ( .A(n6903), .B(n6905), .Z(n6919) );
  XOR U8215 ( .A(n6945), .B(n6946), .Z(n6905) );
  AND U8216 ( .A(n126), .B(n6947), .Z(n6945) );
  XOR U8217 ( .A(n6946), .B(n6948), .Z(n6947) );
  XOR U8218 ( .A(n6949), .B(n6950), .Z(n126) );
  AND U8219 ( .A(n6951), .B(n6952), .Z(n6949) );
  XNOR U8220 ( .A(n6950), .B(n6916), .Z(n6952) );
  XNOR U8221 ( .A(n6953), .B(n6954), .Z(n6916) );
  ANDN U8222 ( .B(n6955), .A(n6956), .Z(n6953) );
  XOR U8223 ( .A(n6954), .B(n6957), .Z(n6955) );
  XOR U8224 ( .A(n6950), .B(n6918), .Z(n6951) );
  XOR U8225 ( .A(n6958), .B(n6959), .Z(n6918) );
  AND U8226 ( .A(n130), .B(n6960), .Z(n6958) );
  XOR U8227 ( .A(n6961), .B(n6959), .Z(n6960) );
  XNOR U8228 ( .A(n6962), .B(n6963), .Z(n6950) );
  NAND U8229 ( .A(n6964), .B(n6965), .Z(n6963) );
  XOR U8230 ( .A(n6966), .B(n6942), .Z(n6965) );
  XOR U8231 ( .A(n6956), .B(n6957), .Z(n6942) );
  XOR U8232 ( .A(n6967), .B(n6968), .Z(n6957) );
  ANDN U8233 ( .B(n6969), .A(n6970), .Z(n6967) );
  XOR U8234 ( .A(n6968), .B(n6971), .Z(n6969) );
  XOR U8235 ( .A(n6972), .B(n6973), .Z(n6956) );
  XOR U8236 ( .A(n6974), .B(n6975), .Z(n6973) );
  ANDN U8237 ( .B(n6976), .A(n6977), .Z(n6974) );
  XOR U8238 ( .A(n6978), .B(n6975), .Z(n6976) );
  IV U8239 ( .A(n6954), .Z(n6972) );
  XOR U8240 ( .A(n6979), .B(n6980), .Z(n6954) );
  ANDN U8241 ( .B(n6981), .A(n6982), .Z(n6979) );
  XOR U8242 ( .A(n6980), .B(n6983), .Z(n6981) );
  IV U8243 ( .A(n6962), .Z(n6966) );
  XOR U8244 ( .A(n6962), .B(n6944), .Z(n6964) );
  XOR U8245 ( .A(n6984), .B(n6985), .Z(n6944) );
  AND U8246 ( .A(n130), .B(n6986), .Z(n6984) );
  XOR U8247 ( .A(n6987), .B(n6985), .Z(n6986) );
  NANDN U8248 ( .A(n6946), .B(n6948), .Z(n6962) );
  XOR U8249 ( .A(n6988), .B(n6989), .Z(n6948) );
  AND U8250 ( .A(n130), .B(n6990), .Z(n6988) );
  XOR U8251 ( .A(n6989), .B(n6991), .Z(n6990) );
  XOR U8252 ( .A(n6992), .B(n6993), .Z(n130) );
  AND U8253 ( .A(n6994), .B(n6995), .Z(n6992) );
  XNOR U8254 ( .A(n6993), .B(n6959), .Z(n6995) );
  XNOR U8255 ( .A(n6996), .B(n6997), .Z(n6959) );
  ANDN U8256 ( .B(n6998), .A(n6999), .Z(n6996) );
  XOR U8257 ( .A(n6997), .B(n7000), .Z(n6998) );
  XOR U8258 ( .A(n6993), .B(n6961), .Z(n6994) );
  XOR U8259 ( .A(n7001), .B(n7002), .Z(n6961) );
  AND U8260 ( .A(n134), .B(n7003), .Z(n7001) );
  XOR U8261 ( .A(n7004), .B(n7002), .Z(n7003) );
  XNOR U8262 ( .A(n7005), .B(n7006), .Z(n6993) );
  NAND U8263 ( .A(n7007), .B(n7008), .Z(n7006) );
  XOR U8264 ( .A(n7009), .B(n6985), .Z(n7008) );
  XOR U8265 ( .A(n6999), .B(n7000), .Z(n6985) );
  XOR U8266 ( .A(n7010), .B(n7011), .Z(n7000) );
  ANDN U8267 ( .B(n7012), .A(n7013), .Z(n7010) );
  XOR U8268 ( .A(n7011), .B(n7014), .Z(n7012) );
  XOR U8269 ( .A(n7015), .B(n7016), .Z(n6999) );
  XOR U8270 ( .A(n7017), .B(n7018), .Z(n7016) );
  ANDN U8271 ( .B(n7019), .A(n7020), .Z(n7017) );
  XOR U8272 ( .A(n7021), .B(n7018), .Z(n7019) );
  IV U8273 ( .A(n6997), .Z(n7015) );
  XOR U8274 ( .A(n7022), .B(n7023), .Z(n6997) );
  ANDN U8275 ( .B(n7024), .A(n7025), .Z(n7022) );
  XOR U8276 ( .A(n7023), .B(n7026), .Z(n7024) );
  IV U8277 ( .A(n7005), .Z(n7009) );
  XOR U8278 ( .A(n7005), .B(n6987), .Z(n7007) );
  XOR U8279 ( .A(n7027), .B(n7028), .Z(n6987) );
  AND U8280 ( .A(n134), .B(n7029), .Z(n7027) );
  XOR U8281 ( .A(n7030), .B(n7028), .Z(n7029) );
  NANDN U8282 ( .A(n6989), .B(n6991), .Z(n7005) );
  XOR U8283 ( .A(n7031), .B(n7032), .Z(n6991) );
  AND U8284 ( .A(n134), .B(n7033), .Z(n7031) );
  XOR U8285 ( .A(n7032), .B(n7034), .Z(n7033) );
  XOR U8286 ( .A(n7035), .B(n7036), .Z(n134) );
  AND U8287 ( .A(n7037), .B(n7038), .Z(n7035) );
  XNOR U8288 ( .A(n7036), .B(n7002), .Z(n7038) );
  XNOR U8289 ( .A(n7039), .B(n7040), .Z(n7002) );
  ANDN U8290 ( .B(n7041), .A(n7042), .Z(n7039) );
  XOR U8291 ( .A(n7040), .B(n7043), .Z(n7041) );
  XOR U8292 ( .A(n7036), .B(n7004), .Z(n7037) );
  XOR U8293 ( .A(n7044), .B(n7045), .Z(n7004) );
  AND U8294 ( .A(n138), .B(n7046), .Z(n7044) );
  XOR U8295 ( .A(n7047), .B(n7045), .Z(n7046) );
  XNOR U8296 ( .A(n7048), .B(n7049), .Z(n7036) );
  NAND U8297 ( .A(n7050), .B(n7051), .Z(n7049) );
  XOR U8298 ( .A(n7052), .B(n7028), .Z(n7051) );
  XOR U8299 ( .A(n7042), .B(n7043), .Z(n7028) );
  XOR U8300 ( .A(n7053), .B(n7054), .Z(n7043) );
  ANDN U8301 ( .B(n7055), .A(n7056), .Z(n7053) );
  XOR U8302 ( .A(n7054), .B(n7057), .Z(n7055) );
  XOR U8303 ( .A(n7058), .B(n7059), .Z(n7042) );
  XOR U8304 ( .A(n7060), .B(n7061), .Z(n7059) );
  ANDN U8305 ( .B(n7062), .A(n7063), .Z(n7060) );
  XOR U8306 ( .A(n7064), .B(n7061), .Z(n7062) );
  IV U8307 ( .A(n7040), .Z(n7058) );
  XOR U8308 ( .A(n7065), .B(n7066), .Z(n7040) );
  ANDN U8309 ( .B(n7067), .A(n7068), .Z(n7065) );
  XOR U8310 ( .A(n7066), .B(n7069), .Z(n7067) );
  IV U8311 ( .A(n7048), .Z(n7052) );
  XOR U8312 ( .A(n7048), .B(n7030), .Z(n7050) );
  XOR U8313 ( .A(n7070), .B(n7071), .Z(n7030) );
  AND U8314 ( .A(n138), .B(n7072), .Z(n7070) );
  XOR U8315 ( .A(n7073), .B(n7071), .Z(n7072) );
  NANDN U8316 ( .A(n7032), .B(n7034), .Z(n7048) );
  XOR U8317 ( .A(n7074), .B(n7075), .Z(n7034) );
  AND U8318 ( .A(n138), .B(n7076), .Z(n7074) );
  XOR U8319 ( .A(n7075), .B(n7077), .Z(n7076) );
  XOR U8320 ( .A(n7078), .B(n7079), .Z(n138) );
  AND U8321 ( .A(n7080), .B(n7081), .Z(n7078) );
  XNOR U8322 ( .A(n7079), .B(n7045), .Z(n7081) );
  XNOR U8323 ( .A(n7082), .B(n7083), .Z(n7045) );
  ANDN U8324 ( .B(n7084), .A(n7085), .Z(n7082) );
  XOR U8325 ( .A(n7083), .B(n7086), .Z(n7084) );
  XOR U8326 ( .A(n7079), .B(n7047), .Z(n7080) );
  XOR U8327 ( .A(n7087), .B(n7088), .Z(n7047) );
  AND U8328 ( .A(n142), .B(n7089), .Z(n7087) );
  XOR U8329 ( .A(n7090), .B(n7088), .Z(n7089) );
  XNOR U8330 ( .A(n7091), .B(n7092), .Z(n7079) );
  NAND U8331 ( .A(n7093), .B(n7094), .Z(n7092) );
  XOR U8332 ( .A(n7095), .B(n7071), .Z(n7094) );
  XOR U8333 ( .A(n7085), .B(n7086), .Z(n7071) );
  XOR U8334 ( .A(n7096), .B(n7097), .Z(n7086) );
  ANDN U8335 ( .B(n7098), .A(n7099), .Z(n7096) );
  XOR U8336 ( .A(n7097), .B(n7100), .Z(n7098) );
  XOR U8337 ( .A(n7101), .B(n7102), .Z(n7085) );
  XOR U8338 ( .A(n7103), .B(n7104), .Z(n7102) );
  ANDN U8339 ( .B(n7105), .A(n7106), .Z(n7103) );
  XOR U8340 ( .A(n7107), .B(n7104), .Z(n7105) );
  IV U8341 ( .A(n7083), .Z(n7101) );
  XOR U8342 ( .A(n7108), .B(n7109), .Z(n7083) );
  ANDN U8343 ( .B(n7110), .A(n7111), .Z(n7108) );
  XOR U8344 ( .A(n7109), .B(n7112), .Z(n7110) );
  IV U8345 ( .A(n7091), .Z(n7095) );
  XOR U8346 ( .A(n7091), .B(n7073), .Z(n7093) );
  XOR U8347 ( .A(n7113), .B(n7114), .Z(n7073) );
  AND U8348 ( .A(n142), .B(n7115), .Z(n7113) );
  XOR U8349 ( .A(n7116), .B(n7114), .Z(n7115) );
  NANDN U8350 ( .A(n7075), .B(n7077), .Z(n7091) );
  XOR U8351 ( .A(n7117), .B(n7118), .Z(n7077) );
  AND U8352 ( .A(n142), .B(n7119), .Z(n7117) );
  XOR U8353 ( .A(n7118), .B(n7120), .Z(n7119) );
  XOR U8354 ( .A(n7121), .B(n7122), .Z(n142) );
  AND U8355 ( .A(n7123), .B(n7124), .Z(n7121) );
  XNOR U8356 ( .A(n7122), .B(n7088), .Z(n7124) );
  XNOR U8357 ( .A(n7125), .B(n7126), .Z(n7088) );
  ANDN U8358 ( .B(n7127), .A(n7128), .Z(n7125) );
  XOR U8359 ( .A(n7126), .B(n7129), .Z(n7127) );
  XOR U8360 ( .A(n7122), .B(n7090), .Z(n7123) );
  XOR U8361 ( .A(n7130), .B(n7131), .Z(n7090) );
  AND U8362 ( .A(n146), .B(n7132), .Z(n7130) );
  XOR U8363 ( .A(n7133), .B(n7131), .Z(n7132) );
  XNOR U8364 ( .A(n7134), .B(n7135), .Z(n7122) );
  NAND U8365 ( .A(n7136), .B(n7137), .Z(n7135) );
  XOR U8366 ( .A(n7138), .B(n7114), .Z(n7137) );
  XOR U8367 ( .A(n7128), .B(n7129), .Z(n7114) );
  XOR U8368 ( .A(n7139), .B(n7140), .Z(n7129) );
  ANDN U8369 ( .B(n7141), .A(n7142), .Z(n7139) );
  XOR U8370 ( .A(n7140), .B(n7143), .Z(n7141) );
  XOR U8371 ( .A(n7144), .B(n7145), .Z(n7128) );
  XOR U8372 ( .A(n7146), .B(n7147), .Z(n7145) );
  ANDN U8373 ( .B(n7148), .A(n7149), .Z(n7146) );
  XOR U8374 ( .A(n7150), .B(n7147), .Z(n7148) );
  IV U8375 ( .A(n7126), .Z(n7144) );
  XOR U8376 ( .A(n7151), .B(n7152), .Z(n7126) );
  ANDN U8377 ( .B(n7153), .A(n7154), .Z(n7151) );
  XOR U8378 ( .A(n7152), .B(n7155), .Z(n7153) );
  IV U8379 ( .A(n7134), .Z(n7138) );
  XOR U8380 ( .A(n7134), .B(n7116), .Z(n7136) );
  XOR U8381 ( .A(n7156), .B(n7157), .Z(n7116) );
  AND U8382 ( .A(n146), .B(n7158), .Z(n7156) );
  XOR U8383 ( .A(n7159), .B(n7157), .Z(n7158) );
  NANDN U8384 ( .A(n7118), .B(n7120), .Z(n7134) );
  XOR U8385 ( .A(n7160), .B(n7161), .Z(n7120) );
  AND U8386 ( .A(n146), .B(n7162), .Z(n7160) );
  XOR U8387 ( .A(n7161), .B(n7163), .Z(n7162) );
  XOR U8388 ( .A(n7164), .B(n7165), .Z(n146) );
  AND U8389 ( .A(n7166), .B(n7167), .Z(n7164) );
  XNOR U8390 ( .A(n7165), .B(n7131), .Z(n7167) );
  XNOR U8391 ( .A(n7168), .B(n7169), .Z(n7131) );
  ANDN U8392 ( .B(n7170), .A(n7171), .Z(n7168) );
  XOR U8393 ( .A(n7169), .B(n7172), .Z(n7170) );
  XOR U8394 ( .A(n7165), .B(n7133), .Z(n7166) );
  XOR U8395 ( .A(n7173), .B(n7174), .Z(n7133) );
  AND U8396 ( .A(n150), .B(n7175), .Z(n7173) );
  XOR U8397 ( .A(n7176), .B(n7174), .Z(n7175) );
  XNOR U8398 ( .A(n7177), .B(n7178), .Z(n7165) );
  NAND U8399 ( .A(n7179), .B(n7180), .Z(n7178) );
  XOR U8400 ( .A(n7181), .B(n7157), .Z(n7180) );
  XOR U8401 ( .A(n7171), .B(n7172), .Z(n7157) );
  XOR U8402 ( .A(n7182), .B(n7183), .Z(n7172) );
  ANDN U8403 ( .B(n7184), .A(n7185), .Z(n7182) );
  XOR U8404 ( .A(n7183), .B(n7186), .Z(n7184) );
  XOR U8405 ( .A(n7187), .B(n7188), .Z(n7171) );
  XOR U8406 ( .A(n7189), .B(n7190), .Z(n7188) );
  ANDN U8407 ( .B(n7191), .A(n7192), .Z(n7189) );
  XOR U8408 ( .A(n7193), .B(n7190), .Z(n7191) );
  IV U8409 ( .A(n7169), .Z(n7187) );
  XOR U8410 ( .A(n7194), .B(n7195), .Z(n7169) );
  ANDN U8411 ( .B(n7196), .A(n7197), .Z(n7194) );
  XOR U8412 ( .A(n7195), .B(n7198), .Z(n7196) );
  IV U8413 ( .A(n7177), .Z(n7181) );
  XOR U8414 ( .A(n7177), .B(n7159), .Z(n7179) );
  XOR U8415 ( .A(n7199), .B(n7200), .Z(n7159) );
  AND U8416 ( .A(n150), .B(n7201), .Z(n7199) );
  XOR U8417 ( .A(n7202), .B(n7200), .Z(n7201) );
  NANDN U8418 ( .A(n7161), .B(n7163), .Z(n7177) );
  XOR U8419 ( .A(n7203), .B(n7204), .Z(n7163) );
  AND U8420 ( .A(n150), .B(n7205), .Z(n7203) );
  XOR U8421 ( .A(n7204), .B(n7206), .Z(n7205) );
  XOR U8422 ( .A(n7207), .B(n7208), .Z(n150) );
  AND U8423 ( .A(n7209), .B(n7210), .Z(n7207) );
  XNOR U8424 ( .A(n7208), .B(n7174), .Z(n7210) );
  XNOR U8425 ( .A(n7211), .B(n7212), .Z(n7174) );
  ANDN U8426 ( .B(n7213), .A(n7214), .Z(n7211) );
  XOR U8427 ( .A(n7212), .B(n7215), .Z(n7213) );
  XOR U8428 ( .A(n7208), .B(n7176), .Z(n7209) );
  XOR U8429 ( .A(n7216), .B(n7217), .Z(n7176) );
  AND U8430 ( .A(n154), .B(n7218), .Z(n7216) );
  XOR U8431 ( .A(n7219), .B(n7217), .Z(n7218) );
  XNOR U8432 ( .A(n7220), .B(n7221), .Z(n7208) );
  NAND U8433 ( .A(n7222), .B(n7223), .Z(n7221) );
  XOR U8434 ( .A(n7224), .B(n7200), .Z(n7223) );
  XOR U8435 ( .A(n7214), .B(n7215), .Z(n7200) );
  XOR U8436 ( .A(n7225), .B(n7226), .Z(n7215) );
  ANDN U8437 ( .B(n7227), .A(n7228), .Z(n7225) );
  XOR U8438 ( .A(n7226), .B(n7229), .Z(n7227) );
  XOR U8439 ( .A(n7230), .B(n7231), .Z(n7214) );
  XOR U8440 ( .A(n7232), .B(n7233), .Z(n7231) );
  ANDN U8441 ( .B(n7234), .A(n7235), .Z(n7232) );
  XOR U8442 ( .A(n7236), .B(n7233), .Z(n7234) );
  IV U8443 ( .A(n7212), .Z(n7230) );
  XOR U8444 ( .A(n7237), .B(n7238), .Z(n7212) );
  ANDN U8445 ( .B(n7239), .A(n7240), .Z(n7237) );
  XOR U8446 ( .A(n7238), .B(n7241), .Z(n7239) );
  IV U8447 ( .A(n7220), .Z(n7224) );
  XOR U8448 ( .A(n7220), .B(n7202), .Z(n7222) );
  XOR U8449 ( .A(n7242), .B(n7243), .Z(n7202) );
  AND U8450 ( .A(n154), .B(n7244), .Z(n7242) );
  XOR U8451 ( .A(n7245), .B(n7243), .Z(n7244) );
  NANDN U8452 ( .A(n7204), .B(n7206), .Z(n7220) );
  XOR U8453 ( .A(n7246), .B(n7247), .Z(n7206) );
  AND U8454 ( .A(n154), .B(n7248), .Z(n7246) );
  XOR U8455 ( .A(n7247), .B(n7249), .Z(n7248) );
  XOR U8456 ( .A(n7250), .B(n7251), .Z(n154) );
  AND U8457 ( .A(n7252), .B(n7253), .Z(n7250) );
  XNOR U8458 ( .A(n7251), .B(n7217), .Z(n7253) );
  XNOR U8459 ( .A(n7254), .B(n7255), .Z(n7217) );
  ANDN U8460 ( .B(n7256), .A(n7257), .Z(n7254) );
  XOR U8461 ( .A(n7255), .B(n7258), .Z(n7256) );
  XOR U8462 ( .A(n7251), .B(n7219), .Z(n7252) );
  XOR U8463 ( .A(n7259), .B(n7260), .Z(n7219) );
  AND U8464 ( .A(n158), .B(n7261), .Z(n7259) );
  XOR U8465 ( .A(n7262), .B(n7260), .Z(n7261) );
  XNOR U8466 ( .A(n7263), .B(n7264), .Z(n7251) );
  NAND U8467 ( .A(n7265), .B(n7266), .Z(n7264) );
  XOR U8468 ( .A(n7267), .B(n7243), .Z(n7266) );
  XOR U8469 ( .A(n7257), .B(n7258), .Z(n7243) );
  XOR U8470 ( .A(n7268), .B(n7269), .Z(n7258) );
  ANDN U8471 ( .B(n7270), .A(n7271), .Z(n7268) );
  XOR U8472 ( .A(n7269), .B(n7272), .Z(n7270) );
  XOR U8473 ( .A(n7273), .B(n7274), .Z(n7257) );
  XOR U8474 ( .A(n7275), .B(n7276), .Z(n7274) );
  ANDN U8475 ( .B(n7277), .A(n7278), .Z(n7275) );
  XOR U8476 ( .A(n7279), .B(n7276), .Z(n7277) );
  IV U8477 ( .A(n7255), .Z(n7273) );
  XOR U8478 ( .A(n7280), .B(n7281), .Z(n7255) );
  ANDN U8479 ( .B(n7282), .A(n7283), .Z(n7280) );
  XOR U8480 ( .A(n7281), .B(n7284), .Z(n7282) );
  IV U8481 ( .A(n7263), .Z(n7267) );
  XOR U8482 ( .A(n7263), .B(n7245), .Z(n7265) );
  XOR U8483 ( .A(n7285), .B(n7286), .Z(n7245) );
  AND U8484 ( .A(n158), .B(n7287), .Z(n7285) );
  XOR U8485 ( .A(n7288), .B(n7286), .Z(n7287) );
  NANDN U8486 ( .A(n7247), .B(n7249), .Z(n7263) );
  XOR U8487 ( .A(n7289), .B(n7290), .Z(n7249) );
  AND U8488 ( .A(n158), .B(n7291), .Z(n7289) );
  XOR U8489 ( .A(n7290), .B(n7292), .Z(n7291) );
  XOR U8490 ( .A(n7293), .B(n7294), .Z(n158) );
  AND U8491 ( .A(n7295), .B(n7296), .Z(n7293) );
  XNOR U8492 ( .A(n7294), .B(n7260), .Z(n7296) );
  XNOR U8493 ( .A(n7297), .B(n7298), .Z(n7260) );
  ANDN U8494 ( .B(n7299), .A(n7300), .Z(n7297) );
  XOR U8495 ( .A(n7298), .B(n7301), .Z(n7299) );
  XOR U8496 ( .A(n7294), .B(n7262), .Z(n7295) );
  XOR U8497 ( .A(n7302), .B(n7303), .Z(n7262) );
  AND U8498 ( .A(n162), .B(n7304), .Z(n7302) );
  XOR U8499 ( .A(n7305), .B(n7303), .Z(n7304) );
  XNOR U8500 ( .A(n7306), .B(n7307), .Z(n7294) );
  NAND U8501 ( .A(n7308), .B(n7309), .Z(n7307) );
  XOR U8502 ( .A(n7310), .B(n7286), .Z(n7309) );
  XOR U8503 ( .A(n7300), .B(n7301), .Z(n7286) );
  XOR U8504 ( .A(n7311), .B(n7312), .Z(n7301) );
  ANDN U8505 ( .B(n7313), .A(n7314), .Z(n7311) );
  XOR U8506 ( .A(n7312), .B(n7315), .Z(n7313) );
  XOR U8507 ( .A(n7316), .B(n7317), .Z(n7300) );
  XOR U8508 ( .A(n7318), .B(n7319), .Z(n7317) );
  ANDN U8509 ( .B(n7320), .A(n7321), .Z(n7318) );
  XOR U8510 ( .A(n7322), .B(n7319), .Z(n7320) );
  IV U8511 ( .A(n7298), .Z(n7316) );
  XOR U8512 ( .A(n7323), .B(n7324), .Z(n7298) );
  ANDN U8513 ( .B(n7325), .A(n7326), .Z(n7323) );
  XOR U8514 ( .A(n7324), .B(n7327), .Z(n7325) );
  IV U8515 ( .A(n7306), .Z(n7310) );
  XOR U8516 ( .A(n7306), .B(n7288), .Z(n7308) );
  XOR U8517 ( .A(n7328), .B(n7329), .Z(n7288) );
  AND U8518 ( .A(n162), .B(n7330), .Z(n7328) );
  XOR U8519 ( .A(n7331), .B(n7329), .Z(n7330) );
  NANDN U8520 ( .A(n7290), .B(n7292), .Z(n7306) );
  XOR U8521 ( .A(n7332), .B(n7333), .Z(n7292) );
  AND U8522 ( .A(n162), .B(n7334), .Z(n7332) );
  XOR U8523 ( .A(n7333), .B(n7335), .Z(n7334) );
  XOR U8524 ( .A(n7336), .B(n7337), .Z(n162) );
  AND U8525 ( .A(n7338), .B(n7339), .Z(n7336) );
  XNOR U8526 ( .A(n7337), .B(n7303), .Z(n7339) );
  XNOR U8527 ( .A(n7340), .B(n7341), .Z(n7303) );
  ANDN U8528 ( .B(n7342), .A(n7343), .Z(n7340) );
  XOR U8529 ( .A(n7341), .B(n7344), .Z(n7342) );
  XOR U8530 ( .A(n7337), .B(n7305), .Z(n7338) );
  XOR U8531 ( .A(n7345), .B(n7346), .Z(n7305) );
  AND U8532 ( .A(n166), .B(n7347), .Z(n7345) );
  XOR U8533 ( .A(n7348), .B(n7346), .Z(n7347) );
  XNOR U8534 ( .A(n7349), .B(n7350), .Z(n7337) );
  NAND U8535 ( .A(n7351), .B(n7352), .Z(n7350) );
  XOR U8536 ( .A(n7353), .B(n7329), .Z(n7352) );
  XOR U8537 ( .A(n7343), .B(n7344), .Z(n7329) );
  XOR U8538 ( .A(n7354), .B(n7355), .Z(n7344) );
  ANDN U8539 ( .B(n7356), .A(n7357), .Z(n7354) );
  XOR U8540 ( .A(n7355), .B(n7358), .Z(n7356) );
  XOR U8541 ( .A(n7359), .B(n7360), .Z(n7343) );
  XOR U8542 ( .A(n7361), .B(n7362), .Z(n7360) );
  ANDN U8543 ( .B(n7363), .A(n7364), .Z(n7361) );
  XOR U8544 ( .A(n7365), .B(n7362), .Z(n7363) );
  IV U8545 ( .A(n7341), .Z(n7359) );
  XOR U8546 ( .A(n7366), .B(n7367), .Z(n7341) );
  ANDN U8547 ( .B(n7368), .A(n7369), .Z(n7366) );
  XOR U8548 ( .A(n7367), .B(n7370), .Z(n7368) );
  IV U8549 ( .A(n7349), .Z(n7353) );
  XOR U8550 ( .A(n7349), .B(n7331), .Z(n7351) );
  XOR U8551 ( .A(n7371), .B(n7372), .Z(n7331) );
  AND U8552 ( .A(n166), .B(n7373), .Z(n7371) );
  XOR U8553 ( .A(n7374), .B(n7372), .Z(n7373) );
  NANDN U8554 ( .A(n7333), .B(n7335), .Z(n7349) );
  XOR U8555 ( .A(n7375), .B(n7376), .Z(n7335) );
  AND U8556 ( .A(n166), .B(n7377), .Z(n7375) );
  XOR U8557 ( .A(n7376), .B(n7378), .Z(n7377) );
  XOR U8558 ( .A(n7379), .B(n7380), .Z(n166) );
  AND U8559 ( .A(n7381), .B(n7382), .Z(n7379) );
  XNOR U8560 ( .A(n7380), .B(n7346), .Z(n7382) );
  XNOR U8561 ( .A(n7383), .B(n7384), .Z(n7346) );
  ANDN U8562 ( .B(n7385), .A(n7386), .Z(n7383) );
  XOR U8563 ( .A(n7384), .B(n7387), .Z(n7385) );
  XOR U8564 ( .A(n7380), .B(n7348), .Z(n7381) );
  XOR U8565 ( .A(n7388), .B(n7389), .Z(n7348) );
  AND U8566 ( .A(n170), .B(n7390), .Z(n7388) );
  XOR U8567 ( .A(n7391), .B(n7389), .Z(n7390) );
  XNOR U8568 ( .A(n7392), .B(n7393), .Z(n7380) );
  NAND U8569 ( .A(n7394), .B(n7395), .Z(n7393) );
  XOR U8570 ( .A(n7396), .B(n7372), .Z(n7395) );
  XOR U8571 ( .A(n7386), .B(n7387), .Z(n7372) );
  XOR U8572 ( .A(n7397), .B(n7398), .Z(n7387) );
  ANDN U8573 ( .B(n7399), .A(n7400), .Z(n7397) );
  XOR U8574 ( .A(n7398), .B(n7401), .Z(n7399) );
  XOR U8575 ( .A(n7402), .B(n7403), .Z(n7386) );
  XOR U8576 ( .A(n7404), .B(n7405), .Z(n7403) );
  ANDN U8577 ( .B(n7406), .A(n7407), .Z(n7404) );
  XOR U8578 ( .A(n7408), .B(n7405), .Z(n7406) );
  IV U8579 ( .A(n7384), .Z(n7402) );
  XOR U8580 ( .A(n7409), .B(n7410), .Z(n7384) );
  ANDN U8581 ( .B(n7411), .A(n7412), .Z(n7409) );
  XOR U8582 ( .A(n7410), .B(n7413), .Z(n7411) );
  IV U8583 ( .A(n7392), .Z(n7396) );
  XOR U8584 ( .A(n7392), .B(n7374), .Z(n7394) );
  XOR U8585 ( .A(n7414), .B(n7415), .Z(n7374) );
  AND U8586 ( .A(n170), .B(n7416), .Z(n7414) );
  XOR U8587 ( .A(n7417), .B(n7415), .Z(n7416) );
  NANDN U8588 ( .A(n7376), .B(n7378), .Z(n7392) );
  XOR U8589 ( .A(n7418), .B(n7419), .Z(n7378) );
  AND U8590 ( .A(n170), .B(n7420), .Z(n7418) );
  XOR U8591 ( .A(n7419), .B(n7421), .Z(n7420) );
  XOR U8592 ( .A(n7422), .B(n7423), .Z(n170) );
  AND U8593 ( .A(n7424), .B(n7425), .Z(n7422) );
  XNOR U8594 ( .A(n7423), .B(n7389), .Z(n7425) );
  XNOR U8595 ( .A(n7426), .B(n7427), .Z(n7389) );
  ANDN U8596 ( .B(n7428), .A(n7429), .Z(n7426) );
  XOR U8597 ( .A(n7427), .B(n7430), .Z(n7428) );
  XOR U8598 ( .A(n7423), .B(n7391), .Z(n7424) );
  XOR U8599 ( .A(n7431), .B(n7432), .Z(n7391) );
  AND U8600 ( .A(n174), .B(n7433), .Z(n7431) );
  XOR U8601 ( .A(n7434), .B(n7432), .Z(n7433) );
  XNOR U8602 ( .A(n7435), .B(n7436), .Z(n7423) );
  NAND U8603 ( .A(n7437), .B(n7438), .Z(n7436) );
  XOR U8604 ( .A(n7439), .B(n7415), .Z(n7438) );
  XOR U8605 ( .A(n7429), .B(n7430), .Z(n7415) );
  XOR U8606 ( .A(n7440), .B(n7441), .Z(n7430) );
  ANDN U8607 ( .B(n7442), .A(n7443), .Z(n7440) );
  XOR U8608 ( .A(n7441), .B(n7444), .Z(n7442) );
  XOR U8609 ( .A(n7445), .B(n7446), .Z(n7429) );
  XOR U8610 ( .A(n7447), .B(n7448), .Z(n7446) );
  ANDN U8611 ( .B(n7449), .A(n7450), .Z(n7447) );
  XOR U8612 ( .A(n7451), .B(n7448), .Z(n7449) );
  IV U8613 ( .A(n7427), .Z(n7445) );
  XOR U8614 ( .A(n7452), .B(n7453), .Z(n7427) );
  ANDN U8615 ( .B(n7454), .A(n7455), .Z(n7452) );
  XOR U8616 ( .A(n7453), .B(n7456), .Z(n7454) );
  IV U8617 ( .A(n7435), .Z(n7439) );
  XOR U8618 ( .A(n7435), .B(n7417), .Z(n7437) );
  XOR U8619 ( .A(n7457), .B(n7458), .Z(n7417) );
  AND U8620 ( .A(n174), .B(n7459), .Z(n7457) );
  XOR U8621 ( .A(n7460), .B(n7458), .Z(n7459) );
  NANDN U8622 ( .A(n7419), .B(n7421), .Z(n7435) );
  XOR U8623 ( .A(n7461), .B(n7462), .Z(n7421) );
  AND U8624 ( .A(n174), .B(n7463), .Z(n7461) );
  XOR U8625 ( .A(n7462), .B(n7464), .Z(n7463) );
  XOR U8626 ( .A(n7465), .B(n7466), .Z(n174) );
  AND U8627 ( .A(n7467), .B(n7468), .Z(n7465) );
  XNOR U8628 ( .A(n7466), .B(n7432), .Z(n7468) );
  XNOR U8629 ( .A(n7469), .B(n7470), .Z(n7432) );
  ANDN U8630 ( .B(n7471), .A(n7472), .Z(n7469) );
  XOR U8631 ( .A(n7470), .B(n7473), .Z(n7471) );
  XOR U8632 ( .A(n7466), .B(n7434), .Z(n7467) );
  XOR U8633 ( .A(n7474), .B(n7475), .Z(n7434) );
  AND U8634 ( .A(n178), .B(n7476), .Z(n7474) );
  XOR U8635 ( .A(n7477), .B(n7475), .Z(n7476) );
  XNOR U8636 ( .A(n7478), .B(n7479), .Z(n7466) );
  NAND U8637 ( .A(n7480), .B(n7481), .Z(n7479) );
  XOR U8638 ( .A(n7482), .B(n7458), .Z(n7481) );
  XOR U8639 ( .A(n7472), .B(n7473), .Z(n7458) );
  XOR U8640 ( .A(n7483), .B(n7484), .Z(n7473) );
  ANDN U8641 ( .B(n7485), .A(n7486), .Z(n7483) );
  XOR U8642 ( .A(n7484), .B(n7487), .Z(n7485) );
  XOR U8643 ( .A(n7488), .B(n7489), .Z(n7472) );
  XOR U8644 ( .A(n7490), .B(n7491), .Z(n7489) );
  ANDN U8645 ( .B(n7492), .A(n7493), .Z(n7490) );
  XOR U8646 ( .A(n7494), .B(n7491), .Z(n7492) );
  IV U8647 ( .A(n7470), .Z(n7488) );
  XOR U8648 ( .A(n7495), .B(n7496), .Z(n7470) );
  ANDN U8649 ( .B(n7497), .A(n7498), .Z(n7495) );
  XOR U8650 ( .A(n7496), .B(n7499), .Z(n7497) );
  IV U8651 ( .A(n7478), .Z(n7482) );
  XOR U8652 ( .A(n7478), .B(n7460), .Z(n7480) );
  XOR U8653 ( .A(n7500), .B(n7501), .Z(n7460) );
  AND U8654 ( .A(n178), .B(n7502), .Z(n7500) );
  XOR U8655 ( .A(n7503), .B(n7501), .Z(n7502) );
  NANDN U8656 ( .A(n7462), .B(n7464), .Z(n7478) );
  XOR U8657 ( .A(n7504), .B(n7505), .Z(n7464) );
  AND U8658 ( .A(n178), .B(n7506), .Z(n7504) );
  XOR U8659 ( .A(n7505), .B(n7507), .Z(n7506) );
  XOR U8660 ( .A(n7508), .B(n7509), .Z(n178) );
  AND U8661 ( .A(n7510), .B(n7511), .Z(n7508) );
  XNOR U8662 ( .A(n7509), .B(n7475), .Z(n7511) );
  XNOR U8663 ( .A(n7512), .B(n7513), .Z(n7475) );
  ANDN U8664 ( .B(n7514), .A(n7515), .Z(n7512) );
  XOR U8665 ( .A(n7513), .B(n7516), .Z(n7514) );
  XOR U8666 ( .A(n7509), .B(n7477), .Z(n7510) );
  XOR U8667 ( .A(n7517), .B(n7518), .Z(n7477) );
  AND U8668 ( .A(n182), .B(n7519), .Z(n7517) );
  XOR U8669 ( .A(n7520), .B(n7518), .Z(n7519) );
  XNOR U8670 ( .A(n7521), .B(n7522), .Z(n7509) );
  NAND U8671 ( .A(n7523), .B(n7524), .Z(n7522) );
  XOR U8672 ( .A(n7525), .B(n7501), .Z(n7524) );
  XOR U8673 ( .A(n7515), .B(n7516), .Z(n7501) );
  XOR U8674 ( .A(n7526), .B(n7527), .Z(n7516) );
  ANDN U8675 ( .B(n7528), .A(n7529), .Z(n7526) );
  XOR U8676 ( .A(n7527), .B(n7530), .Z(n7528) );
  XOR U8677 ( .A(n7531), .B(n7532), .Z(n7515) );
  XOR U8678 ( .A(n7533), .B(n7534), .Z(n7532) );
  ANDN U8679 ( .B(n7535), .A(n7536), .Z(n7533) );
  XOR U8680 ( .A(n7537), .B(n7534), .Z(n7535) );
  IV U8681 ( .A(n7513), .Z(n7531) );
  XOR U8682 ( .A(n7538), .B(n7539), .Z(n7513) );
  ANDN U8683 ( .B(n7540), .A(n7541), .Z(n7538) );
  XOR U8684 ( .A(n7539), .B(n7542), .Z(n7540) );
  IV U8685 ( .A(n7521), .Z(n7525) );
  XOR U8686 ( .A(n7521), .B(n7503), .Z(n7523) );
  XOR U8687 ( .A(n7543), .B(n7544), .Z(n7503) );
  AND U8688 ( .A(n182), .B(n7545), .Z(n7543) );
  XOR U8689 ( .A(n7546), .B(n7544), .Z(n7545) );
  NANDN U8690 ( .A(n7505), .B(n7507), .Z(n7521) );
  XOR U8691 ( .A(n7547), .B(n7548), .Z(n7507) );
  AND U8692 ( .A(n182), .B(n7549), .Z(n7547) );
  XOR U8693 ( .A(n7548), .B(n7550), .Z(n7549) );
  XOR U8694 ( .A(n7551), .B(n7552), .Z(n182) );
  AND U8695 ( .A(n7553), .B(n7554), .Z(n7551) );
  XNOR U8696 ( .A(n7552), .B(n7518), .Z(n7554) );
  XNOR U8697 ( .A(n7555), .B(n7556), .Z(n7518) );
  ANDN U8698 ( .B(n7557), .A(n7558), .Z(n7555) );
  XOR U8699 ( .A(n7556), .B(n7559), .Z(n7557) );
  XOR U8700 ( .A(n7552), .B(n7520), .Z(n7553) );
  XOR U8701 ( .A(n7560), .B(n7561), .Z(n7520) );
  AND U8702 ( .A(n186), .B(n7562), .Z(n7560) );
  XOR U8703 ( .A(n7563), .B(n7561), .Z(n7562) );
  XNOR U8704 ( .A(n7564), .B(n7565), .Z(n7552) );
  NAND U8705 ( .A(n7566), .B(n7567), .Z(n7565) );
  XOR U8706 ( .A(n7568), .B(n7544), .Z(n7567) );
  XOR U8707 ( .A(n7558), .B(n7559), .Z(n7544) );
  XOR U8708 ( .A(n7569), .B(n7570), .Z(n7559) );
  ANDN U8709 ( .B(n7571), .A(n7572), .Z(n7569) );
  XOR U8710 ( .A(n7570), .B(n7573), .Z(n7571) );
  XOR U8711 ( .A(n7574), .B(n7575), .Z(n7558) );
  XOR U8712 ( .A(n7576), .B(n7577), .Z(n7575) );
  ANDN U8713 ( .B(n7578), .A(n7579), .Z(n7576) );
  XOR U8714 ( .A(n7580), .B(n7577), .Z(n7578) );
  IV U8715 ( .A(n7556), .Z(n7574) );
  XOR U8716 ( .A(n7581), .B(n7582), .Z(n7556) );
  ANDN U8717 ( .B(n7583), .A(n7584), .Z(n7581) );
  XOR U8718 ( .A(n7582), .B(n7585), .Z(n7583) );
  IV U8719 ( .A(n7564), .Z(n7568) );
  XOR U8720 ( .A(n7564), .B(n7546), .Z(n7566) );
  XOR U8721 ( .A(n7586), .B(n7587), .Z(n7546) );
  AND U8722 ( .A(n186), .B(n7588), .Z(n7586) );
  XOR U8723 ( .A(n7589), .B(n7587), .Z(n7588) );
  NANDN U8724 ( .A(n7548), .B(n7550), .Z(n7564) );
  XOR U8725 ( .A(n7590), .B(n7591), .Z(n7550) );
  AND U8726 ( .A(n186), .B(n7592), .Z(n7590) );
  XOR U8727 ( .A(n7591), .B(n7593), .Z(n7592) );
  XOR U8728 ( .A(n7594), .B(n7595), .Z(n186) );
  AND U8729 ( .A(n7596), .B(n7597), .Z(n7594) );
  XNOR U8730 ( .A(n7595), .B(n7561), .Z(n7597) );
  XNOR U8731 ( .A(n7598), .B(n7599), .Z(n7561) );
  ANDN U8732 ( .B(n7600), .A(n7601), .Z(n7598) );
  XOR U8733 ( .A(n7599), .B(n7602), .Z(n7600) );
  XOR U8734 ( .A(n7595), .B(n7563), .Z(n7596) );
  XOR U8735 ( .A(n7603), .B(n7604), .Z(n7563) );
  AND U8736 ( .A(n190), .B(n7605), .Z(n7603) );
  XOR U8737 ( .A(n7606), .B(n7604), .Z(n7605) );
  XNOR U8738 ( .A(n7607), .B(n7608), .Z(n7595) );
  NAND U8739 ( .A(n7609), .B(n7610), .Z(n7608) );
  XOR U8740 ( .A(n7611), .B(n7587), .Z(n7610) );
  XOR U8741 ( .A(n7601), .B(n7602), .Z(n7587) );
  XOR U8742 ( .A(n7612), .B(n7613), .Z(n7602) );
  ANDN U8743 ( .B(n7614), .A(n7615), .Z(n7612) );
  XOR U8744 ( .A(n7613), .B(n7616), .Z(n7614) );
  XOR U8745 ( .A(n7617), .B(n7618), .Z(n7601) );
  XOR U8746 ( .A(n7619), .B(n7620), .Z(n7618) );
  ANDN U8747 ( .B(n7621), .A(n7622), .Z(n7619) );
  XOR U8748 ( .A(n7623), .B(n7620), .Z(n7621) );
  IV U8749 ( .A(n7599), .Z(n7617) );
  XOR U8750 ( .A(n7624), .B(n7625), .Z(n7599) );
  ANDN U8751 ( .B(n7626), .A(n7627), .Z(n7624) );
  XOR U8752 ( .A(n7625), .B(n7628), .Z(n7626) );
  IV U8753 ( .A(n7607), .Z(n7611) );
  XOR U8754 ( .A(n7607), .B(n7589), .Z(n7609) );
  XOR U8755 ( .A(n7629), .B(n7630), .Z(n7589) );
  AND U8756 ( .A(n190), .B(n7631), .Z(n7629) );
  XOR U8757 ( .A(n7632), .B(n7630), .Z(n7631) );
  NANDN U8758 ( .A(n7591), .B(n7593), .Z(n7607) );
  XOR U8759 ( .A(n7633), .B(n7634), .Z(n7593) );
  AND U8760 ( .A(n190), .B(n7635), .Z(n7633) );
  XOR U8761 ( .A(n7634), .B(n7636), .Z(n7635) );
  XOR U8762 ( .A(n7637), .B(n7638), .Z(n190) );
  AND U8763 ( .A(n7639), .B(n7640), .Z(n7637) );
  XNOR U8764 ( .A(n7638), .B(n7604), .Z(n7640) );
  XNOR U8765 ( .A(n7641), .B(n7642), .Z(n7604) );
  ANDN U8766 ( .B(n7643), .A(n7644), .Z(n7641) );
  XOR U8767 ( .A(n7642), .B(n7645), .Z(n7643) );
  XOR U8768 ( .A(n7638), .B(n7606), .Z(n7639) );
  XOR U8769 ( .A(n7646), .B(n7647), .Z(n7606) );
  AND U8770 ( .A(n194), .B(n7648), .Z(n7646) );
  XOR U8771 ( .A(n7649), .B(n7647), .Z(n7648) );
  XNOR U8772 ( .A(n7650), .B(n7651), .Z(n7638) );
  NAND U8773 ( .A(n7652), .B(n7653), .Z(n7651) );
  XOR U8774 ( .A(n7654), .B(n7630), .Z(n7653) );
  XOR U8775 ( .A(n7644), .B(n7645), .Z(n7630) );
  XOR U8776 ( .A(n7655), .B(n7656), .Z(n7645) );
  ANDN U8777 ( .B(n7657), .A(n7658), .Z(n7655) );
  XOR U8778 ( .A(n7656), .B(n7659), .Z(n7657) );
  XOR U8779 ( .A(n7660), .B(n7661), .Z(n7644) );
  XOR U8780 ( .A(n7662), .B(n7663), .Z(n7661) );
  ANDN U8781 ( .B(n7664), .A(n7665), .Z(n7662) );
  XOR U8782 ( .A(n7666), .B(n7663), .Z(n7664) );
  IV U8783 ( .A(n7642), .Z(n7660) );
  XOR U8784 ( .A(n7667), .B(n7668), .Z(n7642) );
  ANDN U8785 ( .B(n7669), .A(n7670), .Z(n7667) );
  XOR U8786 ( .A(n7668), .B(n7671), .Z(n7669) );
  IV U8787 ( .A(n7650), .Z(n7654) );
  XOR U8788 ( .A(n7650), .B(n7632), .Z(n7652) );
  XOR U8789 ( .A(n7672), .B(n7673), .Z(n7632) );
  AND U8790 ( .A(n194), .B(n7674), .Z(n7672) );
  XOR U8791 ( .A(n7675), .B(n7673), .Z(n7674) );
  NANDN U8792 ( .A(n7634), .B(n7636), .Z(n7650) );
  XOR U8793 ( .A(n7676), .B(n7677), .Z(n7636) );
  AND U8794 ( .A(n194), .B(n7678), .Z(n7676) );
  XOR U8795 ( .A(n7677), .B(n7679), .Z(n7678) );
  XOR U8796 ( .A(n7680), .B(n7681), .Z(n194) );
  AND U8797 ( .A(n7682), .B(n7683), .Z(n7680) );
  XNOR U8798 ( .A(n7681), .B(n7647), .Z(n7683) );
  XNOR U8799 ( .A(n7684), .B(n7685), .Z(n7647) );
  ANDN U8800 ( .B(n7686), .A(n7687), .Z(n7684) );
  XOR U8801 ( .A(n7685), .B(n7688), .Z(n7686) );
  XOR U8802 ( .A(n7681), .B(n7649), .Z(n7682) );
  XOR U8803 ( .A(n7689), .B(n7690), .Z(n7649) );
  AND U8804 ( .A(n198), .B(n7691), .Z(n7689) );
  XOR U8805 ( .A(n7692), .B(n7690), .Z(n7691) );
  XNOR U8806 ( .A(n7693), .B(n7694), .Z(n7681) );
  NAND U8807 ( .A(n7695), .B(n7696), .Z(n7694) );
  XOR U8808 ( .A(n7697), .B(n7673), .Z(n7696) );
  XOR U8809 ( .A(n7687), .B(n7688), .Z(n7673) );
  XOR U8810 ( .A(n7698), .B(n7699), .Z(n7688) );
  ANDN U8811 ( .B(n7700), .A(n7701), .Z(n7698) );
  XOR U8812 ( .A(n7699), .B(n7702), .Z(n7700) );
  XOR U8813 ( .A(n7703), .B(n7704), .Z(n7687) );
  XOR U8814 ( .A(n7705), .B(n7706), .Z(n7704) );
  ANDN U8815 ( .B(n7707), .A(n7708), .Z(n7705) );
  XOR U8816 ( .A(n7709), .B(n7706), .Z(n7707) );
  IV U8817 ( .A(n7685), .Z(n7703) );
  XOR U8818 ( .A(n7710), .B(n7711), .Z(n7685) );
  ANDN U8819 ( .B(n7712), .A(n7713), .Z(n7710) );
  XOR U8820 ( .A(n7711), .B(n7714), .Z(n7712) );
  IV U8821 ( .A(n7693), .Z(n7697) );
  XOR U8822 ( .A(n7693), .B(n7675), .Z(n7695) );
  XOR U8823 ( .A(n7715), .B(n7716), .Z(n7675) );
  AND U8824 ( .A(n198), .B(n7717), .Z(n7715) );
  XOR U8825 ( .A(n7718), .B(n7716), .Z(n7717) );
  NANDN U8826 ( .A(n7677), .B(n7679), .Z(n7693) );
  XOR U8827 ( .A(n7719), .B(n7720), .Z(n7679) );
  AND U8828 ( .A(n198), .B(n7721), .Z(n7719) );
  XOR U8829 ( .A(n7720), .B(n7722), .Z(n7721) );
  XOR U8830 ( .A(n7723), .B(n7724), .Z(n198) );
  AND U8831 ( .A(n7725), .B(n7726), .Z(n7723) );
  XNOR U8832 ( .A(n7724), .B(n7690), .Z(n7726) );
  XNOR U8833 ( .A(n7727), .B(n7728), .Z(n7690) );
  ANDN U8834 ( .B(n7729), .A(n7730), .Z(n7727) );
  XOR U8835 ( .A(n7728), .B(n7731), .Z(n7729) );
  XOR U8836 ( .A(n7724), .B(n7692), .Z(n7725) );
  XOR U8837 ( .A(n7732), .B(n7733), .Z(n7692) );
  AND U8838 ( .A(n202), .B(n7734), .Z(n7732) );
  XOR U8839 ( .A(n7735), .B(n7733), .Z(n7734) );
  XNOR U8840 ( .A(n7736), .B(n7737), .Z(n7724) );
  NAND U8841 ( .A(n7738), .B(n7739), .Z(n7737) );
  XOR U8842 ( .A(n7740), .B(n7716), .Z(n7739) );
  XOR U8843 ( .A(n7730), .B(n7731), .Z(n7716) );
  XOR U8844 ( .A(n7741), .B(n7742), .Z(n7731) );
  ANDN U8845 ( .B(n7743), .A(n7744), .Z(n7741) );
  XOR U8846 ( .A(n7742), .B(n7745), .Z(n7743) );
  XOR U8847 ( .A(n7746), .B(n7747), .Z(n7730) );
  XOR U8848 ( .A(n7748), .B(n7749), .Z(n7747) );
  ANDN U8849 ( .B(n7750), .A(n7751), .Z(n7748) );
  XOR U8850 ( .A(n7752), .B(n7749), .Z(n7750) );
  IV U8851 ( .A(n7728), .Z(n7746) );
  XOR U8852 ( .A(n7753), .B(n7754), .Z(n7728) );
  ANDN U8853 ( .B(n7755), .A(n7756), .Z(n7753) );
  XOR U8854 ( .A(n7754), .B(n7757), .Z(n7755) );
  IV U8855 ( .A(n7736), .Z(n7740) );
  XOR U8856 ( .A(n7736), .B(n7718), .Z(n7738) );
  XOR U8857 ( .A(n7758), .B(n7759), .Z(n7718) );
  AND U8858 ( .A(n202), .B(n7760), .Z(n7758) );
  XOR U8859 ( .A(n7761), .B(n7759), .Z(n7760) );
  NANDN U8860 ( .A(n7720), .B(n7722), .Z(n7736) );
  XOR U8861 ( .A(n7762), .B(n7763), .Z(n7722) );
  AND U8862 ( .A(n202), .B(n7764), .Z(n7762) );
  XOR U8863 ( .A(n7763), .B(n7765), .Z(n7764) );
  XOR U8864 ( .A(n7766), .B(n7767), .Z(n202) );
  AND U8865 ( .A(n7768), .B(n7769), .Z(n7766) );
  XNOR U8866 ( .A(n7767), .B(n7733), .Z(n7769) );
  XNOR U8867 ( .A(n7770), .B(n7771), .Z(n7733) );
  ANDN U8868 ( .B(n7772), .A(n7773), .Z(n7770) );
  XOR U8869 ( .A(n7771), .B(n7774), .Z(n7772) );
  XOR U8870 ( .A(n7767), .B(n7735), .Z(n7768) );
  XOR U8871 ( .A(n7775), .B(n7776), .Z(n7735) );
  AND U8872 ( .A(n206), .B(n7777), .Z(n7775) );
  XOR U8873 ( .A(n7778), .B(n7776), .Z(n7777) );
  XNOR U8874 ( .A(n7779), .B(n7780), .Z(n7767) );
  NAND U8875 ( .A(n7781), .B(n7782), .Z(n7780) );
  XOR U8876 ( .A(n7783), .B(n7759), .Z(n7782) );
  XOR U8877 ( .A(n7773), .B(n7774), .Z(n7759) );
  XOR U8878 ( .A(n7784), .B(n7785), .Z(n7774) );
  ANDN U8879 ( .B(n7786), .A(n7787), .Z(n7784) );
  XOR U8880 ( .A(n7785), .B(n7788), .Z(n7786) );
  XOR U8881 ( .A(n7789), .B(n7790), .Z(n7773) );
  XOR U8882 ( .A(n7791), .B(n7792), .Z(n7790) );
  ANDN U8883 ( .B(n7793), .A(n7794), .Z(n7791) );
  XOR U8884 ( .A(n7795), .B(n7792), .Z(n7793) );
  IV U8885 ( .A(n7771), .Z(n7789) );
  XOR U8886 ( .A(n7796), .B(n7797), .Z(n7771) );
  ANDN U8887 ( .B(n7798), .A(n7799), .Z(n7796) );
  XOR U8888 ( .A(n7797), .B(n7800), .Z(n7798) );
  IV U8889 ( .A(n7779), .Z(n7783) );
  XOR U8890 ( .A(n7779), .B(n7761), .Z(n7781) );
  XOR U8891 ( .A(n7801), .B(n7802), .Z(n7761) );
  AND U8892 ( .A(n206), .B(n7803), .Z(n7801) );
  XOR U8893 ( .A(n7804), .B(n7802), .Z(n7803) );
  NANDN U8894 ( .A(n7763), .B(n7765), .Z(n7779) );
  XOR U8895 ( .A(n7805), .B(n7806), .Z(n7765) );
  AND U8896 ( .A(n206), .B(n7807), .Z(n7805) );
  XOR U8897 ( .A(n7806), .B(n7808), .Z(n7807) );
  XOR U8898 ( .A(n7809), .B(n7810), .Z(n206) );
  AND U8899 ( .A(n7811), .B(n7812), .Z(n7809) );
  XNOR U8900 ( .A(n7810), .B(n7776), .Z(n7812) );
  XNOR U8901 ( .A(n7813), .B(n7814), .Z(n7776) );
  ANDN U8902 ( .B(n7815), .A(n7816), .Z(n7813) );
  XOR U8903 ( .A(n7814), .B(n7817), .Z(n7815) );
  XOR U8904 ( .A(n7810), .B(n7778), .Z(n7811) );
  XOR U8905 ( .A(n7818), .B(n7819), .Z(n7778) );
  AND U8906 ( .A(n210), .B(n7820), .Z(n7818) );
  XOR U8907 ( .A(n7821), .B(n7819), .Z(n7820) );
  XNOR U8908 ( .A(n7822), .B(n7823), .Z(n7810) );
  NAND U8909 ( .A(n7824), .B(n7825), .Z(n7823) );
  XOR U8910 ( .A(n7826), .B(n7802), .Z(n7825) );
  XOR U8911 ( .A(n7816), .B(n7817), .Z(n7802) );
  XOR U8912 ( .A(n7827), .B(n7828), .Z(n7817) );
  ANDN U8913 ( .B(n7829), .A(n7830), .Z(n7827) );
  XOR U8914 ( .A(n7828), .B(n7831), .Z(n7829) );
  XOR U8915 ( .A(n7832), .B(n7833), .Z(n7816) );
  XOR U8916 ( .A(n7834), .B(n7835), .Z(n7833) );
  ANDN U8917 ( .B(n7836), .A(n7837), .Z(n7834) );
  XOR U8918 ( .A(n7838), .B(n7835), .Z(n7836) );
  IV U8919 ( .A(n7814), .Z(n7832) );
  XOR U8920 ( .A(n7839), .B(n7840), .Z(n7814) );
  ANDN U8921 ( .B(n7841), .A(n7842), .Z(n7839) );
  XOR U8922 ( .A(n7840), .B(n7843), .Z(n7841) );
  IV U8923 ( .A(n7822), .Z(n7826) );
  XOR U8924 ( .A(n7822), .B(n7804), .Z(n7824) );
  XOR U8925 ( .A(n7844), .B(n7845), .Z(n7804) );
  AND U8926 ( .A(n210), .B(n7846), .Z(n7844) );
  XOR U8927 ( .A(n7847), .B(n7845), .Z(n7846) );
  NANDN U8928 ( .A(n7806), .B(n7808), .Z(n7822) );
  XOR U8929 ( .A(n7848), .B(n7849), .Z(n7808) );
  AND U8930 ( .A(n210), .B(n7850), .Z(n7848) );
  XOR U8931 ( .A(n7849), .B(n7851), .Z(n7850) );
  XOR U8932 ( .A(n7852), .B(n7853), .Z(n210) );
  AND U8933 ( .A(n7854), .B(n7855), .Z(n7852) );
  XNOR U8934 ( .A(n7853), .B(n7819), .Z(n7855) );
  XNOR U8935 ( .A(n7856), .B(n7857), .Z(n7819) );
  ANDN U8936 ( .B(n7858), .A(n7859), .Z(n7856) );
  XOR U8937 ( .A(n7857), .B(n7860), .Z(n7858) );
  XOR U8938 ( .A(n7853), .B(n7821), .Z(n7854) );
  XOR U8939 ( .A(n7861), .B(n7862), .Z(n7821) );
  AND U8940 ( .A(n214), .B(n7863), .Z(n7861) );
  XOR U8941 ( .A(n7864), .B(n7862), .Z(n7863) );
  XNOR U8942 ( .A(n7865), .B(n7866), .Z(n7853) );
  NAND U8943 ( .A(n7867), .B(n7868), .Z(n7866) );
  XOR U8944 ( .A(n7869), .B(n7845), .Z(n7868) );
  XOR U8945 ( .A(n7859), .B(n7860), .Z(n7845) );
  XOR U8946 ( .A(n7870), .B(n7871), .Z(n7860) );
  ANDN U8947 ( .B(n7872), .A(n7873), .Z(n7870) );
  XOR U8948 ( .A(n7871), .B(n7874), .Z(n7872) );
  XOR U8949 ( .A(n7875), .B(n7876), .Z(n7859) );
  XOR U8950 ( .A(n7877), .B(n7878), .Z(n7876) );
  ANDN U8951 ( .B(n7879), .A(n7880), .Z(n7877) );
  XOR U8952 ( .A(n7881), .B(n7878), .Z(n7879) );
  IV U8953 ( .A(n7857), .Z(n7875) );
  XOR U8954 ( .A(n7882), .B(n7883), .Z(n7857) );
  ANDN U8955 ( .B(n7884), .A(n7885), .Z(n7882) );
  XOR U8956 ( .A(n7883), .B(n7886), .Z(n7884) );
  IV U8957 ( .A(n7865), .Z(n7869) );
  XOR U8958 ( .A(n7865), .B(n7847), .Z(n7867) );
  XOR U8959 ( .A(n7887), .B(n7888), .Z(n7847) );
  AND U8960 ( .A(n214), .B(n7889), .Z(n7887) );
  XOR U8961 ( .A(n7890), .B(n7888), .Z(n7889) );
  NANDN U8962 ( .A(n7849), .B(n7851), .Z(n7865) );
  XOR U8963 ( .A(n7891), .B(n7892), .Z(n7851) );
  AND U8964 ( .A(n214), .B(n7893), .Z(n7891) );
  XOR U8965 ( .A(n7892), .B(n7894), .Z(n7893) );
  XOR U8966 ( .A(n7895), .B(n7896), .Z(n214) );
  AND U8967 ( .A(n7897), .B(n7898), .Z(n7895) );
  XNOR U8968 ( .A(n7896), .B(n7862), .Z(n7898) );
  XNOR U8969 ( .A(n7899), .B(n7900), .Z(n7862) );
  ANDN U8970 ( .B(n7901), .A(n7902), .Z(n7899) );
  XOR U8971 ( .A(n7900), .B(n7903), .Z(n7901) );
  XOR U8972 ( .A(n7896), .B(n7864), .Z(n7897) );
  XOR U8973 ( .A(n7904), .B(n7905), .Z(n7864) );
  AND U8974 ( .A(n218), .B(n7906), .Z(n7904) );
  XOR U8975 ( .A(n7907), .B(n7905), .Z(n7906) );
  XNOR U8976 ( .A(n7908), .B(n7909), .Z(n7896) );
  NAND U8977 ( .A(n7910), .B(n7911), .Z(n7909) );
  XOR U8978 ( .A(n7912), .B(n7888), .Z(n7911) );
  XOR U8979 ( .A(n7902), .B(n7903), .Z(n7888) );
  XOR U8980 ( .A(n7913), .B(n7914), .Z(n7903) );
  ANDN U8981 ( .B(n7915), .A(n7916), .Z(n7913) );
  XOR U8982 ( .A(n7914), .B(n7917), .Z(n7915) );
  XOR U8983 ( .A(n7918), .B(n7919), .Z(n7902) );
  XOR U8984 ( .A(n7920), .B(n7921), .Z(n7919) );
  ANDN U8985 ( .B(n7922), .A(n7923), .Z(n7920) );
  XOR U8986 ( .A(n7924), .B(n7921), .Z(n7922) );
  IV U8987 ( .A(n7900), .Z(n7918) );
  XOR U8988 ( .A(n7925), .B(n7926), .Z(n7900) );
  ANDN U8989 ( .B(n7927), .A(n7928), .Z(n7925) );
  XOR U8990 ( .A(n7926), .B(n7929), .Z(n7927) );
  IV U8991 ( .A(n7908), .Z(n7912) );
  XOR U8992 ( .A(n7908), .B(n7890), .Z(n7910) );
  XOR U8993 ( .A(n7930), .B(n7931), .Z(n7890) );
  AND U8994 ( .A(n218), .B(n7932), .Z(n7930) );
  XOR U8995 ( .A(n7933), .B(n7931), .Z(n7932) );
  NANDN U8996 ( .A(n7892), .B(n7894), .Z(n7908) );
  XOR U8997 ( .A(n7934), .B(n7935), .Z(n7894) );
  AND U8998 ( .A(n218), .B(n7936), .Z(n7934) );
  XOR U8999 ( .A(n7935), .B(n7937), .Z(n7936) );
  XOR U9000 ( .A(n7938), .B(n7939), .Z(n218) );
  AND U9001 ( .A(n7940), .B(n7941), .Z(n7938) );
  XNOR U9002 ( .A(n7939), .B(n7905), .Z(n7941) );
  XNOR U9003 ( .A(n7942), .B(n7943), .Z(n7905) );
  ANDN U9004 ( .B(n7944), .A(n7945), .Z(n7942) );
  XOR U9005 ( .A(n7943), .B(n7946), .Z(n7944) );
  XOR U9006 ( .A(n7939), .B(n7907), .Z(n7940) );
  XOR U9007 ( .A(n7947), .B(n7948), .Z(n7907) );
  AND U9008 ( .A(n222), .B(n7949), .Z(n7947) );
  XOR U9009 ( .A(n7950), .B(n7948), .Z(n7949) );
  XNOR U9010 ( .A(n7951), .B(n7952), .Z(n7939) );
  NAND U9011 ( .A(n7953), .B(n7954), .Z(n7952) );
  XOR U9012 ( .A(n7955), .B(n7931), .Z(n7954) );
  XOR U9013 ( .A(n7945), .B(n7946), .Z(n7931) );
  XOR U9014 ( .A(n7956), .B(n7957), .Z(n7946) );
  ANDN U9015 ( .B(n7958), .A(n7959), .Z(n7956) );
  XOR U9016 ( .A(n7957), .B(n7960), .Z(n7958) );
  XOR U9017 ( .A(n7961), .B(n7962), .Z(n7945) );
  XOR U9018 ( .A(n7963), .B(n7964), .Z(n7962) );
  ANDN U9019 ( .B(n7965), .A(n7966), .Z(n7963) );
  XOR U9020 ( .A(n7967), .B(n7964), .Z(n7965) );
  IV U9021 ( .A(n7943), .Z(n7961) );
  XOR U9022 ( .A(n7968), .B(n7969), .Z(n7943) );
  ANDN U9023 ( .B(n7970), .A(n7971), .Z(n7968) );
  XOR U9024 ( .A(n7969), .B(n7972), .Z(n7970) );
  IV U9025 ( .A(n7951), .Z(n7955) );
  XOR U9026 ( .A(n7951), .B(n7933), .Z(n7953) );
  XOR U9027 ( .A(n7973), .B(n7974), .Z(n7933) );
  AND U9028 ( .A(n222), .B(n7975), .Z(n7973) );
  XOR U9029 ( .A(n7976), .B(n7974), .Z(n7975) );
  NANDN U9030 ( .A(n7935), .B(n7937), .Z(n7951) );
  XOR U9031 ( .A(n7977), .B(n7978), .Z(n7937) );
  AND U9032 ( .A(n222), .B(n7979), .Z(n7977) );
  XOR U9033 ( .A(n7978), .B(n7980), .Z(n7979) );
  XOR U9034 ( .A(n7981), .B(n7982), .Z(n222) );
  AND U9035 ( .A(n7983), .B(n7984), .Z(n7981) );
  XNOR U9036 ( .A(n7982), .B(n7948), .Z(n7984) );
  XNOR U9037 ( .A(n7985), .B(n7986), .Z(n7948) );
  ANDN U9038 ( .B(n7987), .A(n7988), .Z(n7985) );
  XOR U9039 ( .A(n7986), .B(n7989), .Z(n7987) );
  XOR U9040 ( .A(n7982), .B(n7950), .Z(n7983) );
  XOR U9041 ( .A(n7990), .B(n7991), .Z(n7950) );
  AND U9042 ( .A(n226), .B(n7992), .Z(n7990) );
  XOR U9043 ( .A(n7993), .B(n7991), .Z(n7992) );
  XNOR U9044 ( .A(n7994), .B(n7995), .Z(n7982) );
  NAND U9045 ( .A(n7996), .B(n7997), .Z(n7995) );
  XOR U9046 ( .A(n7998), .B(n7974), .Z(n7997) );
  XOR U9047 ( .A(n7988), .B(n7989), .Z(n7974) );
  XOR U9048 ( .A(n7999), .B(n8000), .Z(n7989) );
  ANDN U9049 ( .B(n8001), .A(n8002), .Z(n7999) );
  XOR U9050 ( .A(n8000), .B(n8003), .Z(n8001) );
  XOR U9051 ( .A(n8004), .B(n8005), .Z(n7988) );
  XOR U9052 ( .A(n8006), .B(n8007), .Z(n8005) );
  ANDN U9053 ( .B(n8008), .A(n8009), .Z(n8006) );
  XOR U9054 ( .A(n8010), .B(n8007), .Z(n8008) );
  IV U9055 ( .A(n7986), .Z(n8004) );
  XOR U9056 ( .A(n8011), .B(n8012), .Z(n7986) );
  ANDN U9057 ( .B(n8013), .A(n8014), .Z(n8011) );
  XOR U9058 ( .A(n8012), .B(n8015), .Z(n8013) );
  IV U9059 ( .A(n7994), .Z(n7998) );
  XOR U9060 ( .A(n7994), .B(n7976), .Z(n7996) );
  XOR U9061 ( .A(n8016), .B(n8017), .Z(n7976) );
  AND U9062 ( .A(n226), .B(n8018), .Z(n8016) );
  XOR U9063 ( .A(n8019), .B(n8017), .Z(n8018) );
  NANDN U9064 ( .A(n7978), .B(n7980), .Z(n7994) );
  XOR U9065 ( .A(n8020), .B(n8021), .Z(n7980) );
  AND U9066 ( .A(n226), .B(n8022), .Z(n8020) );
  XOR U9067 ( .A(n8021), .B(n8023), .Z(n8022) );
  XOR U9068 ( .A(n8024), .B(n8025), .Z(n226) );
  AND U9069 ( .A(n8026), .B(n8027), .Z(n8024) );
  XNOR U9070 ( .A(n8025), .B(n7991), .Z(n8027) );
  XNOR U9071 ( .A(n8028), .B(n8029), .Z(n7991) );
  ANDN U9072 ( .B(n8030), .A(n8031), .Z(n8028) );
  XOR U9073 ( .A(n8029), .B(n8032), .Z(n8030) );
  XOR U9074 ( .A(n8025), .B(n7993), .Z(n8026) );
  XOR U9075 ( .A(n8033), .B(n8034), .Z(n7993) );
  AND U9076 ( .A(n230), .B(n8035), .Z(n8033) );
  XOR U9077 ( .A(n8036), .B(n8034), .Z(n8035) );
  XNOR U9078 ( .A(n8037), .B(n8038), .Z(n8025) );
  NAND U9079 ( .A(n8039), .B(n8040), .Z(n8038) );
  XOR U9080 ( .A(n8041), .B(n8017), .Z(n8040) );
  XOR U9081 ( .A(n8031), .B(n8032), .Z(n8017) );
  XOR U9082 ( .A(n8042), .B(n8043), .Z(n8032) );
  ANDN U9083 ( .B(n8044), .A(n8045), .Z(n8042) );
  XOR U9084 ( .A(n8043), .B(n8046), .Z(n8044) );
  XOR U9085 ( .A(n8047), .B(n8048), .Z(n8031) );
  XOR U9086 ( .A(n8049), .B(n8050), .Z(n8048) );
  ANDN U9087 ( .B(n8051), .A(n8052), .Z(n8049) );
  XOR U9088 ( .A(n8053), .B(n8050), .Z(n8051) );
  IV U9089 ( .A(n8029), .Z(n8047) );
  XOR U9090 ( .A(n8054), .B(n8055), .Z(n8029) );
  ANDN U9091 ( .B(n8056), .A(n8057), .Z(n8054) );
  XOR U9092 ( .A(n8055), .B(n8058), .Z(n8056) );
  IV U9093 ( .A(n8037), .Z(n8041) );
  XOR U9094 ( .A(n8037), .B(n8019), .Z(n8039) );
  XOR U9095 ( .A(n8059), .B(n8060), .Z(n8019) );
  AND U9096 ( .A(n230), .B(n8061), .Z(n8059) );
  XOR U9097 ( .A(n8062), .B(n8060), .Z(n8061) );
  NANDN U9098 ( .A(n8021), .B(n8023), .Z(n8037) );
  XOR U9099 ( .A(n8063), .B(n8064), .Z(n8023) );
  AND U9100 ( .A(n230), .B(n8065), .Z(n8063) );
  XOR U9101 ( .A(n8064), .B(n8066), .Z(n8065) );
  XOR U9102 ( .A(n8067), .B(n8068), .Z(n230) );
  AND U9103 ( .A(n8069), .B(n8070), .Z(n8067) );
  XNOR U9104 ( .A(n8068), .B(n8034), .Z(n8070) );
  XNOR U9105 ( .A(n8071), .B(n8072), .Z(n8034) );
  ANDN U9106 ( .B(n8073), .A(n8074), .Z(n8071) );
  XOR U9107 ( .A(n8072), .B(n8075), .Z(n8073) );
  XOR U9108 ( .A(n8068), .B(n8036), .Z(n8069) );
  XOR U9109 ( .A(n8076), .B(n8077), .Z(n8036) );
  AND U9110 ( .A(n234), .B(n8078), .Z(n8076) );
  XOR U9111 ( .A(n8079), .B(n8077), .Z(n8078) );
  XNOR U9112 ( .A(n8080), .B(n8081), .Z(n8068) );
  NAND U9113 ( .A(n8082), .B(n8083), .Z(n8081) );
  XOR U9114 ( .A(n8084), .B(n8060), .Z(n8083) );
  XOR U9115 ( .A(n8074), .B(n8075), .Z(n8060) );
  XOR U9116 ( .A(n8085), .B(n8086), .Z(n8075) );
  ANDN U9117 ( .B(n8087), .A(n8088), .Z(n8085) );
  XOR U9118 ( .A(n8086), .B(n8089), .Z(n8087) );
  XOR U9119 ( .A(n8090), .B(n8091), .Z(n8074) );
  XOR U9120 ( .A(n8092), .B(n8093), .Z(n8091) );
  ANDN U9121 ( .B(n8094), .A(n8095), .Z(n8092) );
  XOR U9122 ( .A(n8096), .B(n8093), .Z(n8094) );
  IV U9123 ( .A(n8072), .Z(n8090) );
  XOR U9124 ( .A(n8097), .B(n8098), .Z(n8072) );
  ANDN U9125 ( .B(n8099), .A(n8100), .Z(n8097) );
  XOR U9126 ( .A(n8098), .B(n8101), .Z(n8099) );
  IV U9127 ( .A(n8080), .Z(n8084) );
  XOR U9128 ( .A(n8080), .B(n8062), .Z(n8082) );
  XOR U9129 ( .A(n8102), .B(n8103), .Z(n8062) );
  AND U9130 ( .A(n234), .B(n8104), .Z(n8102) );
  XOR U9131 ( .A(n8105), .B(n8103), .Z(n8104) );
  NANDN U9132 ( .A(n8064), .B(n8066), .Z(n8080) );
  XOR U9133 ( .A(n8106), .B(n8107), .Z(n8066) );
  AND U9134 ( .A(n234), .B(n8108), .Z(n8106) );
  XOR U9135 ( .A(n8107), .B(n8109), .Z(n8108) );
  XOR U9136 ( .A(n8110), .B(n8111), .Z(n234) );
  AND U9137 ( .A(n8112), .B(n8113), .Z(n8110) );
  XNOR U9138 ( .A(n8111), .B(n8077), .Z(n8113) );
  XNOR U9139 ( .A(n8114), .B(n8115), .Z(n8077) );
  ANDN U9140 ( .B(n8116), .A(n8117), .Z(n8114) );
  XOR U9141 ( .A(n8115), .B(n8118), .Z(n8116) );
  XOR U9142 ( .A(n8111), .B(n8079), .Z(n8112) );
  XOR U9143 ( .A(n8119), .B(n8120), .Z(n8079) );
  AND U9144 ( .A(n238), .B(n8121), .Z(n8119) );
  XOR U9145 ( .A(n8122), .B(n8120), .Z(n8121) );
  XNOR U9146 ( .A(n8123), .B(n8124), .Z(n8111) );
  NAND U9147 ( .A(n8125), .B(n8126), .Z(n8124) );
  XOR U9148 ( .A(n8127), .B(n8103), .Z(n8126) );
  XOR U9149 ( .A(n8117), .B(n8118), .Z(n8103) );
  XOR U9150 ( .A(n8128), .B(n8129), .Z(n8118) );
  ANDN U9151 ( .B(n8130), .A(n8131), .Z(n8128) );
  XOR U9152 ( .A(n8129), .B(n8132), .Z(n8130) );
  XOR U9153 ( .A(n8133), .B(n8134), .Z(n8117) );
  XOR U9154 ( .A(n8135), .B(n8136), .Z(n8134) );
  ANDN U9155 ( .B(n8137), .A(n8138), .Z(n8135) );
  XOR U9156 ( .A(n8139), .B(n8136), .Z(n8137) );
  IV U9157 ( .A(n8115), .Z(n8133) );
  XOR U9158 ( .A(n8140), .B(n8141), .Z(n8115) );
  ANDN U9159 ( .B(n8142), .A(n8143), .Z(n8140) );
  XOR U9160 ( .A(n8141), .B(n8144), .Z(n8142) );
  IV U9161 ( .A(n8123), .Z(n8127) );
  XOR U9162 ( .A(n8123), .B(n8105), .Z(n8125) );
  XOR U9163 ( .A(n8145), .B(n8146), .Z(n8105) );
  AND U9164 ( .A(n238), .B(n8147), .Z(n8145) );
  XOR U9165 ( .A(n8148), .B(n8146), .Z(n8147) );
  NANDN U9166 ( .A(n8107), .B(n8109), .Z(n8123) );
  XOR U9167 ( .A(n8149), .B(n8150), .Z(n8109) );
  AND U9168 ( .A(n238), .B(n8151), .Z(n8149) );
  XOR U9169 ( .A(n8150), .B(n8152), .Z(n8151) );
  XOR U9170 ( .A(n8153), .B(n8154), .Z(n238) );
  AND U9171 ( .A(n8155), .B(n8156), .Z(n8153) );
  XNOR U9172 ( .A(n8154), .B(n8120), .Z(n8156) );
  XNOR U9173 ( .A(n8157), .B(n8158), .Z(n8120) );
  ANDN U9174 ( .B(n8159), .A(n8160), .Z(n8157) );
  XOR U9175 ( .A(n8158), .B(n8161), .Z(n8159) );
  XOR U9176 ( .A(n8154), .B(n8122), .Z(n8155) );
  XOR U9177 ( .A(n8162), .B(n8163), .Z(n8122) );
  AND U9178 ( .A(n242), .B(n8164), .Z(n8162) );
  XOR U9179 ( .A(n8165), .B(n8163), .Z(n8164) );
  XNOR U9180 ( .A(n8166), .B(n8167), .Z(n8154) );
  NAND U9181 ( .A(n8168), .B(n8169), .Z(n8167) );
  XOR U9182 ( .A(n8170), .B(n8146), .Z(n8169) );
  XOR U9183 ( .A(n8160), .B(n8161), .Z(n8146) );
  XOR U9184 ( .A(n8171), .B(n8172), .Z(n8161) );
  ANDN U9185 ( .B(n8173), .A(n8174), .Z(n8171) );
  XOR U9186 ( .A(n8172), .B(n8175), .Z(n8173) );
  XOR U9187 ( .A(n8176), .B(n8177), .Z(n8160) );
  XOR U9188 ( .A(n8178), .B(n8179), .Z(n8177) );
  ANDN U9189 ( .B(n8180), .A(n8181), .Z(n8178) );
  XOR U9190 ( .A(n8182), .B(n8179), .Z(n8180) );
  IV U9191 ( .A(n8158), .Z(n8176) );
  XOR U9192 ( .A(n8183), .B(n8184), .Z(n8158) );
  ANDN U9193 ( .B(n8185), .A(n8186), .Z(n8183) );
  XOR U9194 ( .A(n8184), .B(n8187), .Z(n8185) );
  IV U9195 ( .A(n8166), .Z(n8170) );
  XOR U9196 ( .A(n8166), .B(n8148), .Z(n8168) );
  XOR U9197 ( .A(n8188), .B(n8189), .Z(n8148) );
  AND U9198 ( .A(n242), .B(n8190), .Z(n8188) );
  XOR U9199 ( .A(n8191), .B(n8189), .Z(n8190) );
  NANDN U9200 ( .A(n8150), .B(n8152), .Z(n8166) );
  XOR U9201 ( .A(n8192), .B(n8193), .Z(n8152) );
  AND U9202 ( .A(n242), .B(n8194), .Z(n8192) );
  XOR U9203 ( .A(n8193), .B(n8195), .Z(n8194) );
  XOR U9204 ( .A(n8196), .B(n8197), .Z(n242) );
  AND U9205 ( .A(n8198), .B(n8199), .Z(n8196) );
  XNOR U9206 ( .A(n8197), .B(n8163), .Z(n8199) );
  XNOR U9207 ( .A(n8200), .B(n8201), .Z(n8163) );
  ANDN U9208 ( .B(n8202), .A(n8203), .Z(n8200) );
  XOR U9209 ( .A(n8201), .B(n8204), .Z(n8202) );
  XOR U9210 ( .A(n8197), .B(n8165), .Z(n8198) );
  XOR U9211 ( .A(n8205), .B(n8206), .Z(n8165) );
  AND U9212 ( .A(n246), .B(n8207), .Z(n8205) );
  XOR U9213 ( .A(n8208), .B(n8206), .Z(n8207) );
  XNOR U9214 ( .A(n8209), .B(n8210), .Z(n8197) );
  NAND U9215 ( .A(n8211), .B(n8212), .Z(n8210) );
  XOR U9216 ( .A(n8213), .B(n8189), .Z(n8212) );
  XOR U9217 ( .A(n8203), .B(n8204), .Z(n8189) );
  XOR U9218 ( .A(n8214), .B(n8215), .Z(n8204) );
  ANDN U9219 ( .B(n8216), .A(n8217), .Z(n8214) );
  XOR U9220 ( .A(n8215), .B(n8218), .Z(n8216) );
  XOR U9221 ( .A(n8219), .B(n8220), .Z(n8203) );
  XOR U9222 ( .A(n8221), .B(n8222), .Z(n8220) );
  ANDN U9223 ( .B(n8223), .A(n8224), .Z(n8221) );
  XOR U9224 ( .A(n8225), .B(n8222), .Z(n8223) );
  IV U9225 ( .A(n8201), .Z(n8219) );
  XOR U9226 ( .A(n8226), .B(n8227), .Z(n8201) );
  ANDN U9227 ( .B(n8228), .A(n8229), .Z(n8226) );
  XOR U9228 ( .A(n8227), .B(n8230), .Z(n8228) );
  IV U9229 ( .A(n8209), .Z(n8213) );
  XOR U9230 ( .A(n8209), .B(n8191), .Z(n8211) );
  XOR U9231 ( .A(n8231), .B(n8232), .Z(n8191) );
  AND U9232 ( .A(n246), .B(n8233), .Z(n8231) );
  XOR U9233 ( .A(n8234), .B(n8232), .Z(n8233) );
  NANDN U9234 ( .A(n8193), .B(n8195), .Z(n8209) );
  XOR U9235 ( .A(n8235), .B(n8236), .Z(n8195) );
  AND U9236 ( .A(n246), .B(n8237), .Z(n8235) );
  XOR U9237 ( .A(n8236), .B(n8238), .Z(n8237) );
  XOR U9238 ( .A(n8239), .B(n8240), .Z(n246) );
  AND U9239 ( .A(n8241), .B(n8242), .Z(n8239) );
  XNOR U9240 ( .A(n8240), .B(n8206), .Z(n8242) );
  XNOR U9241 ( .A(n8243), .B(n8244), .Z(n8206) );
  ANDN U9242 ( .B(n8245), .A(n8246), .Z(n8243) );
  XOR U9243 ( .A(n8244), .B(n8247), .Z(n8245) );
  XOR U9244 ( .A(n8240), .B(n8208), .Z(n8241) );
  XOR U9245 ( .A(n8248), .B(n8249), .Z(n8208) );
  AND U9246 ( .A(n250), .B(n8250), .Z(n8248) );
  XOR U9247 ( .A(n8251), .B(n8249), .Z(n8250) );
  XNOR U9248 ( .A(n8252), .B(n8253), .Z(n8240) );
  NAND U9249 ( .A(n8254), .B(n8255), .Z(n8253) );
  XOR U9250 ( .A(n8256), .B(n8232), .Z(n8255) );
  XOR U9251 ( .A(n8246), .B(n8247), .Z(n8232) );
  XOR U9252 ( .A(n8257), .B(n8258), .Z(n8247) );
  ANDN U9253 ( .B(n8259), .A(n8260), .Z(n8257) );
  XOR U9254 ( .A(n8258), .B(n8261), .Z(n8259) );
  XOR U9255 ( .A(n8262), .B(n8263), .Z(n8246) );
  XOR U9256 ( .A(n8264), .B(n8265), .Z(n8263) );
  ANDN U9257 ( .B(n8266), .A(n8267), .Z(n8264) );
  XOR U9258 ( .A(n8268), .B(n8265), .Z(n8266) );
  IV U9259 ( .A(n8244), .Z(n8262) );
  XOR U9260 ( .A(n8269), .B(n8270), .Z(n8244) );
  ANDN U9261 ( .B(n8271), .A(n8272), .Z(n8269) );
  XOR U9262 ( .A(n8270), .B(n8273), .Z(n8271) );
  IV U9263 ( .A(n8252), .Z(n8256) );
  XOR U9264 ( .A(n8252), .B(n8234), .Z(n8254) );
  XOR U9265 ( .A(n8274), .B(n8275), .Z(n8234) );
  AND U9266 ( .A(n250), .B(n8276), .Z(n8274) );
  XOR U9267 ( .A(n8277), .B(n8275), .Z(n8276) );
  NANDN U9268 ( .A(n8236), .B(n8238), .Z(n8252) );
  XOR U9269 ( .A(n8278), .B(n8279), .Z(n8238) );
  AND U9270 ( .A(n250), .B(n8280), .Z(n8278) );
  XOR U9271 ( .A(n8279), .B(n8281), .Z(n8280) );
  XOR U9272 ( .A(n8282), .B(n8283), .Z(n250) );
  AND U9273 ( .A(n8284), .B(n8285), .Z(n8282) );
  XNOR U9274 ( .A(n8283), .B(n8249), .Z(n8285) );
  XNOR U9275 ( .A(n8286), .B(n8287), .Z(n8249) );
  ANDN U9276 ( .B(n8288), .A(n8289), .Z(n8286) );
  XOR U9277 ( .A(n8287), .B(n8290), .Z(n8288) );
  XOR U9278 ( .A(n8283), .B(n8251), .Z(n8284) );
  XOR U9279 ( .A(n8291), .B(n8292), .Z(n8251) );
  AND U9280 ( .A(n254), .B(n8293), .Z(n8291) );
  XOR U9281 ( .A(n8294), .B(n8292), .Z(n8293) );
  XNOR U9282 ( .A(n8295), .B(n8296), .Z(n8283) );
  NAND U9283 ( .A(n8297), .B(n8298), .Z(n8296) );
  XOR U9284 ( .A(n8299), .B(n8275), .Z(n8298) );
  XOR U9285 ( .A(n8289), .B(n8290), .Z(n8275) );
  XOR U9286 ( .A(n8300), .B(n8301), .Z(n8290) );
  ANDN U9287 ( .B(n8302), .A(n8303), .Z(n8300) );
  XOR U9288 ( .A(n8301), .B(n8304), .Z(n8302) );
  XOR U9289 ( .A(n8305), .B(n8306), .Z(n8289) );
  XOR U9290 ( .A(n8307), .B(n8308), .Z(n8306) );
  ANDN U9291 ( .B(n8309), .A(n8310), .Z(n8307) );
  XOR U9292 ( .A(n8311), .B(n8308), .Z(n8309) );
  IV U9293 ( .A(n8287), .Z(n8305) );
  XOR U9294 ( .A(n8312), .B(n8313), .Z(n8287) );
  ANDN U9295 ( .B(n8314), .A(n8315), .Z(n8312) );
  XOR U9296 ( .A(n8313), .B(n8316), .Z(n8314) );
  IV U9297 ( .A(n8295), .Z(n8299) );
  XOR U9298 ( .A(n8295), .B(n8277), .Z(n8297) );
  XOR U9299 ( .A(n8317), .B(n8318), .Z(n8277) );
  AND U9300 ( .A(n254), .B(n8319), .Z(n8317) );
  XOR U9301 ( .A(n8320), .B(n8318), .Z(n8319) );
  NANDN U9302 ( .A(n8279), .B(n8281), .Z(n8295) );
  XOR U9303 ( .A(n8321), .B(n8322), .Z(n8281) );
  AND U9304 ( .A(n254), .B(n8323), .Z(n8321) );
  XOR U9305 ( .A(n8322), .B(n8324), .Z(n8323) );
  XOR U9306 ( .A(n8325), .B(n8326), .Z(n254) );
  AND U9307 ( .A(n8327), .B(n8328), .Z(n8325) );
  XNOR U9308 ( .A(n8326), .B(n8292), .Z(n8328) );
  XNOR U9309 ( .A(n8329), .B(n8330), .Z(n8292) );
  ANDN U9310 ( .B(n8331), .A(n8332), .Z(n8329) );
  XOR U9311 ( .A(n8330), .B(n8333), .Z(n8331) );
  XOR U9312 ( .A(n8326), .B(n8294), .Z(n8327) );
  XOR U9313 ( .A(n8334), .B(n8335), .Z(n8294) );
  AND U9314 ( .A(n258), .B(n8336), .Z(n8334) );
  XOR U9315 ( .A(n8337), .B(n8335), .Z(n8336) );
  XNOR U9316 ( .A(n8338), .B(n8339), .Z(n8326) );
  NAND U9317 ( .A(n8340), .B(n8341), .Z(n8339) );
  XOR U9318 ( .A(n8342), .B(n8318), .Z(n8341) );
  XOR U9319 ( .A(n8332), .B(n8333), .Z(n8318) );
  XOR U9320 ( .A(n8343), .B(n8344), .Z(n8333) );
  ANDN U9321 ( .B(n8345), .A(n8346), .Z(n8343) );
  XOR U9322 ( .A(n8344), .B(n8347), .Z(n8345) );
  XOR U9323 ( .A(n8348), .B(n8349), .Z(n8332) );
  XOR U9324 ( .A(n8350), .B(n8351), .Z(n8349) );
  ANDN U9325 ( .B(n8352), .A(n8353), .Z(n8350) );
  XOR U9326 ( .A(n8354), .B(n8351), .Z(n8352) );
  IV U9327 ( .A(n8330), .Z(n8348) );
  XOR U9328 ( .A(n8355), .B(n8356), .Z(n8330) );
  ANDN U9329 ( .B(n8357), .A(n8358), .Z(n8355) );
  XOR U9330 ( .A(n8356), .B(n8359), .Z(n8357) );
  IV U9331 ( .A(n8338), .Z(n8342) );
  XOR U9332 ( .A(n8338), .B(n8320), .Z(n8340) );
  XOR U9333 ( .A(n8360), .B(n8361), .Z(n8320) );
  AND U9334 ( .A(n258), .B(n8362), .Z(n8360) );
  XOR U9335 ( .A(n8363), .B(n8361), .Z(n8362) );
  NANDN U9336 ( .A(n8322), .B(n8324), .Z(n8338) );
  XOR U9337 ( .A(n8364), .B(n8365), .Z(n8324) );
  AND U9338 ( .A(n258), .B(n8366), .Z(n8364) );
  XOR U9339 ( .A(n8365), .B(n8367), .Z(n8366) );
  XOR U9340 ( .A(n8368), .B(n8369), .Z(n258) );
  AND U9341 ( .A(n8370), .B(n8371), .Z(n8368) );
  XNOR U9342 ( .A(n8369), .B(n8335), .Z(n8371) );
  XNOR U9343 ( .A(n8372), .B(n8373), .Z(n8335) );
  ANDN U9344 ( .B(n8374), .A(n8375), .Z(n8372) );
  XOR U9345 ( .A(n8373), .B(n8376), .Z(n8374) );
  XOR U9346 ( .A(n8369), .B(n8337), .Z(n8370) );
  XOR U9347 ( .A(n8377), .B(n8378), .Z(n8337) );
  AND U9348 ( .A(n262), .B(n8379), .Z(n8377) );
  XOR U9349 ( .A(n8380), .B(n8378), .Z(n8379) );
  XNOR U9350 ( .A(n8381), .B(n8382), .Z(n8369) );
  NAND U9351 ( .A(n8383), .B(n8384), .Z(n8382) );
  XOR U9352 ( .A(n8385), .B(n8361), .Z(n8384) );
  XOR U9353 ( .A(n8375), .B(n8376), .Z(n8361) );
  XOR U9354 ( .A(n8386), .B(n8387), .Z(n8376) );
  ANDN U9355 ( .B(n8388), .A(n8389), .Z(n8386) );
  XOR U9356 ( .A(n8387), .B(n8390), .Z(n8388) );
  XOR U9357 ( .A(n8391), .B(n8392), .Z(n8375) );
  XOR U9358 ( .A(n8393), .B(n8394), .Z(n8392) );
  ANDN U9359 ( .B(n8395), .A(n8396), .Z(n8393) );
  XOR U9360 ( .A(n8397), .B(n8394), .Z(n8395) );
  IV U9361 ( .A(n8373), .Z(n8391) );
  XOR U9362 ( .A(n8398), .B(n8399), .Z(n8373) );
  ANDN U9363 ( .B(n8400), .A(n8401), .Z(n8398) );
  XOR U9364 ( .A(n8399), .B(n8402), .Z(n8400) );
  IV U9365 ( .A(n8381), .Z(n8385) );
  XOR U9366 ( .A(n8381), .B(n8363), .Z(n8383) );
  XOR U9367 ( .A(n8403), .B(n8404), .Z(n8363) );
  AND U9368 ( .A(n262), .B(n8405), .Z(n8403) );
  XOR U9369 ( .A(n8406), .B(n8404), .Z(n8405) );
  NANDN U9370 ( .A(n8365), .B(n8367), .Z(n8381) );
  XOR U9371 ( .A(n8407), .B(n8408), .Z(n8367) );
  AND U9372 ( .A(n262), .B(n8409), .Z(n8407) );
  XOR U9373 ( .A(n8408), .B(n8410), .Z(n8409) );
  XOR U9374 ( .A(n8411), .B(n8412), .Z(n262) );
  AND U9375 ( .A(n8413), .B(n8414), .Z(n8411) );
  XNOR U9376 ( .A(n8412), .B(n8378), .Z(n8414) );
  XNOR U9377 ( .A(n8415), .B(n8416), .Z(n8378) );
  ANDN U9378 ( .B(n8417), .A(n8418), .Z(n8415) );
  XOR U9379 ( .A(n8416), .B(n8419), .Z(n8417) );
  XOR U9380 ( .A(n8412), .B(n8380), .Z(n8413) );
  XOR U9381 ( .A(n8420), .B(n8421), .Z(n8380) );
  AND U9382 ( .A(n266), .B(n8422), .Z(n8420) );
  XOR U9383 ( .A(n8423), .B(n8421), .Z(n8422) );
  XNOR U9384 ( .A(n8424), .B(n8425), .Z(n8412) );
  NAND U9385 ( .A(n8426), .B(n8427), .Z(n8425) );
  XOR U9386 ( .A(n8428), .B(n8404), .Z(n8427) );
  XOR U9387 ( .A(n8418), .B(n8419), .Z(n8404) );
  XOR U9388 ( .A(n8429), .B(n8430), .Z(n8419) );
  ANDN U9389 ( .B(n8431), .A(n8432), .Z(n8429) );
  XOR U9390 ( .A(n8430), .B(n8433), .Z(n8431) );
  XOR U9391 ( .A(n8434), .B(n8435), .Z(n8418) );
  XOR U9392 ( .A(n8436), .B(n8437), .Z(n8435) );
  ANDN U9393 ( .B(n8438), .A(n8439), .Z(n8436) );
  XOR U9394 ( .A(n8440), .B(n8437), .Z(n8438) );
  IV U9395 ( .A(n8416), .Z(n8434) );
  XOR U9396 ( .A(n8441), .B(n8442), .Z(n8416) );
  ANDN U9397 ( .B(n8443), .A(n8444), .Z(n8441) );
  XOR U9398 ( .A(n8442), .B(n8445), .Z(n8443) );
  IV U9399 ( .A(n8424), .Z(n8428) );
  XOR U9400 ( .A(n8424), .B(n8406), .Z(n8426) );
  XOR U9401 ( .A(n8446), .B(n8447), .Z(n8406) );
  AND U9402 ( .A(n266), .B(n8448), .Z(n8446) );
  XOR U9403 ( .A(n8449), .B(n8447), .Z(n8448) );
  NANDN U9404 ( .A(n8408), .B(n8410), .Z(n8424) );
  XOR U9405 ( .A(n8450), .B(n8451), .Z(n8410) );
  AND U9406 ( .A(n266), .B(n8452), .Z(n8450) );
  XOR U9407 ( .A(n8451), .B(n8453), .Z(n8452) );
  XOR U9408 ( .A(n8454), .B(n8455), .Z(n266) );
  AND U9409 ( .A(n8456), .B(n8457), .Z(n8454) );
  XNOR U9410 ( .A(n8455), .B(n8421), .Z(n8457) );
  XNOR U9411 ( .A(n8458), .B(n8459), .Z(n8421) );
  ANDN U9412 ( .B(n8460), .A(n8461), .Z(n8458) );
  XOR U9413 ( .A(n8459), .B(n8462), .Z(n8460) );
  XOR U9414 ( .A(n8455), .B(n8423), .Z(n8456) );
  XOR U9415 ( .A(n8463), .B(n8464), .Z(n8423) );
  AND U9416 ( .A(n270), .B(n8465), .Z(n8463) );
  XOR U9417 ( .A(n8466), .B(n8464), .Z(n8465) );
  XNOR U9418 ( .A(n8467), .B(n8468), .Z(n8455) );
  NAND U9419 ( .A(n8469), .B(n8470), .Z(n8468) );
  XOR U9420 ( .A(n8471), .B(n8447), .Z(n8470) );
  XOR U9421 ( .A(n8461), .B(n8462), .Z(n8447) );
  XOR U9422 ( .A(n8472), .B(n8473), .Z(n8462) );
  ANDN U9423 ( .B(n8474), .A(n8475), .Z(n8472) );
  XOR U9424 ( .A(n8473), .B(n8476), .Z(n8474) );
  XOR U9425 ( .A(n8477), .B(n8478), .Z(n8461) );
  XOR U9426 ( .A(n8479), .B(n8480), .Z(n8478) );
  ANDN U9427 ( .B(n8481), .A(n8482), .Z(n8479) );
  XOR U9428 ( .A(n8483), .B(n8480), .Z(n8481) );
  IV U9429 ( .A(n8459), .Z(n8477) );
  XOR U9430 ( .A(n8484), .B(n8485), .Z(n8459) );
  ANDN U9431 ( .B(n8486), .A(n8487), .Z(n8484) );
  XOR U9432 ( .A(n8485), .B(n8488), .Z(n8486) );
  IV U9433 ( .A(n8467), .Z(n8471) );
  XOR U9434 ( .A(n8467), .B(n8449), .Z(n8469) );
  XOR U9435 ( .A(n8489), .B(n8490), .Z(n8449) );
  AND U9436 ( .A(n270), .B(n8491), .Z(n8489) );
  XOR U9437 ( .A(n8492), .B(n8490), .Z(n8491) );
  NANDN U9438 ( .A(n8451), .B(n8453), .Z(n8467) );
  XOR U9439 ( .A(n8493), .B(n8494), .Z(n8453) );
  AND U9440 ( .A(n270), .B(n8495), .Z(n8493) );
  XOR U9441 ( .A(n8494), .B(n8496), .Z(n8495) );
  XOR U9442 ( .A(n8497), .B(n8498), .Z(n270) );
  AND U9443 ( .A(n8499), .B(n8500), .Z(n8497) );
  XNOR U9444 ( .A(n8498), .B(n8464), .Z(n8500) );
  XNOR U9445 ( .A(n8501), .B(n8502), .Z(n8464) );
  ANDN U9446 ( .B(n8503), .A(n8504), .Z(n8501) );
  XOR U9447 ( .A(n8502), .B(n8505), .Z(n8503) );
  XOR U9448 ( .A(n8498), .B(n8466), .Z(n8499) );
  XOR U9449 ( .A(n8506), .B(n8507), .Z(n8466) );
  AND U9450 ( .A(n274), .B(n8508), .Z(n8506) );
  XOR U9451 ( .A(n8509), .B(n8507), .Z(n8508) );
  XNOR U9452 ( .A(n8510), .B(n8511), .Z(n8498) );
  NAND U9453 ( .A(n8512), .B(n8513), .Z(n8511) );
  XOR U9454 ( .A(n8514), .B(n8490), .Z(n8513) );
  XOR U9455 ( .A(n8504), .B(n8505), .Z(n8490) );
  XOR U9456 ( .A(n8515), .B(n8516), .Z(n8505) );
  ANDN U9457 ( .B(n8517), .A(n8518), .Z(n8515) );
  XOR U9458 ( .A(n8516), .B(n8519), .Z(n8517) );
  XOR U9459 ( .A(n8520), .B(n8521), .Z(n8504) );
  XOR U9460 ( .A(n8522), .B(n8523), .Z(n8521) );
  ANDN U9461 ( .B(n8524), .A(n8525), .Z(n8522) );
  XOR U9462 ( .A(n8526), .B(n8523), .Z(n8524) );
  IV U9463 ( .A(n8502), .Z(n8520) );
  XOR U9464 ( .A(n8527), .B(n8528), .Z(n8502) );
  ANDN U9465 ( .B(n8529), .A(n8530), .Z(n8527) );
  XOR U9466 ( .A(n8528), .B(n8531), .Z(n8529) );
  IV U9467 ( .A(n8510), .Z(n8514) );
  XOR U9468 ( .A(n8510), .B(n8492), .Z(n8512) );
  XOR U9469 ( .A(n8532), .B(n8533), .Z(n8492) );
  AND U9470 ( .A(n274), .B(n8534), .Z(n8532) );
  XOR U9471 ( .A(n8535), .B(n8533), .Z(n8534) );
  NANDN U9472 ( .A(n8494), .B(n8496), .Z(n8510) );
  XOR U9473 ( .A(n8536), .B(n8537), .Z(n8496) );
  AND U9474 ( .A(n274), .B(n8538), .Z(n8536) );
  XOR U9475 ( .A(n8537), .B(n8539), .Z(n8538) );
  XOR U9476 ( .A(n8540), .B(n8541), .Z(n274) );
  AND U9477 ( .A(n8542), .B(n8543), .Z(n8540) );
  XNOR U9478 ( .A(n8541), .B(n8507), .Z(n8543) );
  XNOR U9479 ( .A(n8544), .B(n8545), .Z(n8507) );
  ANDN U9480 ( .B(n8546), .A(n8547), .Z(n8544) );
  XOR U9481 ( .A(n8545), .B(n8548), .Z(n8546) );
  XOR U9482 ( .A(n8541), .B(n8509), .Z(n8542) );
  XOR U9483 ( .A(n8549), .B(n8550), .Z(n8509) );
  AND U9484 ( .A(n278), .B(n8551), .Z(n8549) );
  XOR U9485 ( .A(n8552), .B(n8550), .Z(n8551) );
  XNOR U9486 ( .A(n8553), .B(n8554), .Z(n8541) );
  NAND U9487 ( .A(n8555), .B(n8556), .Z(n8554) );
  XOR U9488 ( .A(n8557), .B(n8533), .Z(n8556) );
  XOR U9489 ( .A(n8547), .B(n8548), .Z(n8533) );
  XOR U9490 ( .A(n8558), .B(n8559), .Z(n8548) );
  ANDN U9491 ( .B(n8560), .A(n8561), .Z(n8558) );
  XOR U9492 ( .A(n8559), .B(n8562), .Z(n8560) );
  XOR U9493 ( .A(n8563), .B(n8564), .Z(n8547) );
  XOR U9494 ( .A(n8565), .B(n8566), .Z(n8564) );
  ANDN U9495 ( .B(n8567), .A(n8568), .Z(n8565) );
  XOR U9496 ( .A(n8569), .B(n8566), .Z(n8567) );
  IV U9497 ( .A(n8545), .Z(n8563) );
  XOR U9498 ( .A(n8570), .B(n8571), .Z(n8545) );
  ANDN U9499 ( .B(n8572), .A(n8573), .Z(n8570) );
  XOR U9500 ( .A(n8571), .B(n8574), .Z(n8572) );
  IV U9501 ( .A(n8553), .Z(n8557) );
  XOR U9502 ( .A(n8553), .B(n8535), .Z(n8555) );
  XOR U9503 ( .A(n8575), .B(n8576), .Z(n8535) );
  AND U9504 ( .A(n278), .B(n8577), .Z(n8575) );
  XOR U9505 ( .A(n8578), .B(n8576), .Z(n8577) );
  NANDN U9506 ( .A(n8537), .B(n8539), .Z(n8553) );
  XOR U9507 ( .A(n8579), .B(n8580), .Z(n8539) );
  AND U9508 ( .A(n278), .B(n8581), .Z(n8579) );
  XOR U9509 ( .A(n8580), .B(n8582), .Z(n8581) );
  XOR U9510 ( .A(n8583), .B(n8584), .Z(n278) );
  AND U9511 ( .A(n8585), .B(n8586), .Z(n8583) );
  XNOR U9512 ( .A(n8584), .B(n8550), .Z(n8586) );
  XNOR U9513 ( .A(n8587), .B(n8588), .Z(n8550) );
  ANDN U9514 ( .B(n8589), .A(n8590), .Z(n8587) );
  XOR U9515 ( .A(n8588), .B(n8591), .Z(n8589) );
  XOR U9516 ( .A(n8584), .B(n8552), .Z(n8585) );
  XOR U9517 ( .A(n8592), .B(n8593), .Z(n8552) );
  AND U9518 ( .A(n282), .B(n8594), .Z(n8592) );
  XOR U9519 ( .A(n8595), .B(n8593), .Z(n8594) );
  XNOR U9520 ( .A(n8596), .B(n8597), .Z(n8584) );
  NAND U9521 ( .A(n8598), .B(n8599), .Z(n8597) );
  XOR U9522 ( .A(n8600), .B(n8576), .Z(n8599) );
  XOR U9523 ( .A(n8590), .B(n8591), .Z(n8576) );
  XOR U9524 ( .A(n8601), .B(n8602), .Z(n8591) );
  ANDN U9525 ( .B(n8603), .A(n8604), .Z(n8601) );
  XOR U9526 ( .A(n8602), .B(n8605), .Z(n8603) );
  XOR U9527 ( .A(n8606), .B(n8607), .Z(n8590) );
  XOR U9528 ( .A(n8608), .B(n8609), .Z(n8607) );
  ANDN U9529 ( .B(n8610), .A(n8611), .Z(n8608) );
  XOR U9530 ( .A(n8612), .B(n8609), .Z(n8610) );
  IV U9531 ( .A(n8588), .Z(n8606) );
  XOR U9532 ( .A(n8613), .B(n8614), .Z(n8588) );
  ANDN U9533 ( .B(n8615), .A(n8616), .Z(n8613) );
  XOR U9534 ( .A(n8614), .B(n8617), .Z(n8615) );
  IV U9535 ( .A(n8596), .Z(n8600) );
  XOR U9536 ( .A(n8596), .B(n8578), .Z(n8598) );
  XOR U9537 ( .A(n8618), .B(n8619), .Z(n8578) );
  AND U9538 ( .A(n282), .B(n8620), .Z(n8618) );
  XOR U9539 ( .A(n8621), .B(n8619), .Z(n8620) );
  NANDN U9540 ( .A(n8580), .B(n8582), .Z(n8596) );
  XOR U9541 ( .A(n8622), .B(n8623), .Z(n8582) );
  AND U9542 ( .A(n282), .B(n8624), .Z(n8622) );
  XOR U9543 ( .A(n8623), .B(n8625), .Z(n8624) );
  XOR U9544 ( .A(n8626), .B(n8627), .Z(n282) );
  AND U9545 ( .A(n8628), .B(n8629), .Z(n8626) );
  XNOR U9546 ( .A(n8627), .B(n8593), .Z(n8629) );
  XNOR U9547 ( .A(n8630), .B(n8631), .Z(n8593) );
  ANDN U9548 ( .B(n8632), .A(n8633), .Z(n8630) );
  XOR U9549 ( .A(n8631), .B(n8634), .Z(n8632) );
  XOR U9550 ( .A(n8627), .B(n8595), .Z(n8628) );
  XOR U9551 ( .A(n8635), .B(n8636), .Z(n8595) );
  AND U9552 ( .A(n286), .B(n8637), .Z(n8635) );
  XOR U9553 ( .A(n8638), .B(n8636), .Z(n8637) );
  XNOR U9554 ( .A(n8639), .B(n8640), .Z(n8627) );
  NAND U9555 ( .A(n8641), .B(n8642), .Z(n8640) );
  XOR U9556 ( .A(n8643), .B(n8619), .Z(n8642) );
  XOR U9557 ( .A(n8633), .B(n8634), .Z(n8619) );
  XOR U9558 ( .A(n8644), .B(n8645), .Z(n8634) );
  ANDN U9559 ( .B(n8646), .A(n8647), .Z(n8644) );
  XOR U9560 ( .A(n8645), .B(n8648), .Z(n8646) );
  XOR U9561 ( .A(n8649), .B(n8650), .Z(n8633) );
  XOR U9562 ( .A(n8651), .B(n8652), .Z(n8650) );
  ANDN U9563 ( .B(n8653), .A(n8654), .Z(n8651) );
  XOR U9564 ( .A(n8655), .B(n8652), .Z(n8653) );
  IV U9565 ( .A(n8631), .Z(n8649) );
  XOR U9566 ( .A(n8656), .B(n8657), .Z(n8631) );
  ANDN U9567 ( .B(n8658), .A(n8659), .Z(n8656) );
  XOR U9568 ( .A(n8657), .B(n8660), .Z(n8658) );
  IV U9569 ( .A(n8639), .Z(n8643) );
  XOR U9570 ( .A(n8639), .B(n8621), .Z(n8641) );
  XOR U9571 ( .A(n8661), .B(n8662), .Z(n8621) );
  AND U9572 ( .A(n286), .B(n8663), .Z(n8661) );
  XOR U9573 ( .A(n8664), .B(n8662), .Z(n8663) );
  NANDN U9574 ( .A(n8623), .B(n8625), .Z(n8639) );
  XOR U9575 ( .A(n8665), .B(n8666), .Z(n8625) );
  AND U9576 ( .A(n286), .B(n8667), .Z(n8665) );
  XOR U9577 ( .A(n8666), .B(n8668), .Z(n8667) );
  XOR U9578 ( .A(n8669), .B(n8670), .Z(n286) );
  AND U9579 ( .A(n8671), .B(n8672), .Z(n8669) );
  XNOR U9580 ( .A(n8670), .B(n8636), .Z(n8672) );
  XNOR U9581 ( .A(n8673), .B(n8674), .Z(n8636) );
  ANDN U9582 ( .B(n8675), .A(n8676), .Z(n8673) );
  XOR U9583 ( .A(n8674), .B(n8677), .Z(n8675) );
  XOR U9584 ( .A(n8670), .B(n8638), .Z(n8671) );
  XOR U9585 ( .A(n8678), .B(n8679), .Z(n8638) );
  AND U9586 ( .A(n290), .B(n8680), .Z(n8678) );
  XOR U9587 ( .A(n8681), .B(n8679), .Z(n8680) );
  XNOR U9588 ( .A(n8682), .B(n8683), .Z(n8670) );
  NAND U9589 ( .A(n8684), .B(n8685), .Z(n8683) );
  XOR U9590 ( .A(n8686), .B(n8662), .Z(n8685) );
  XOR U9591 ( .A(n8676), .B(n8677), .Z(n8662) );
  XOR U9592 ( .A(n8687), .B(n8688), .Z(n8677) );
  ANDN U9593 ( .B(n8689), .A(n8690), .Z(n8687) );
  XOR U9594 ( .A(n8688), .B(n8691), .Z(n8689) );
  XOR U9595 ( .A(n8692), .B(n8693), .Z(n8676) );
  XOR U9596 ( .A(n8694), .B(n8695), .Z(n8693) );
  ANDN U9597 ( .B(n8696), .A(n8697), .Z(n8694) );
  XOR U9598 ( .A(n8698), .B(n8695), .Z(n8696) );
  IV U9599 ( .A(n8674), .Z(n8692) );
  XOR U9600 ( .A(n8699), .B(n8700), .Z(n8674) );
  ANDN U9601 ( .B(n8701), .A(n8702), .Z(n8699) );
  XOR U9602 ( .A(n8700), .B(n8703), .Z(n8701) );
  IV U9603 ( .A(n8682), .Z(n8686) );
  XOR U9604 ( .A(n8682), .B(n8664), .Z(n8684) );
  XOR U9605 ( .A(n8704), .B(n8705), .Z(n8664) );
  AND U9606 ( .A(n290), .B(n8706), .Z(n8704) );
  XOR U9607 ( .A(n8707), .B(n8705), .Z(n8706) );
  NANDN U9608 ( .A(n8666), .B(n8668), .Z(n8682) );
  XOR U9609 ( .A(n8708), .B(n8709), .Z(n8668) );
  AND U9610 ( .A(n290), .B(n8710), .Z(n8708) );
  XOR U9611 ( .A(n8709), .B(n8711), .Z(n8710) );
  XOR U9612 ( .A(n8712), .B(n8713), .Z(n290) );
  AND U9613 ( .A(n8714), .B(n8715), .Z(n8712) );
  XNOR U9614 ( .A(n8713), .B(n8679), .Z(n8715) );
  XNOR U9615 ( .A(n8716), .B(n8717), .Z(n8679) );
  ANDN U9616 ( .B(n8718), .A(n8719), .Z(n8716) );
  XOR U9617 ( .A(n8717), .B(n8720), .Z(n8718) );
  XOR U9618 ( .A(n8713), .B(n8681), .Z(n8714) );
  XOR U9619 ( .A(n8721), .B(n8722), .Z(n8681) );
  AND U9620 ( .A(n294), .B(n8723), .Z(n8721) );
  XOR U9621 ( .A(n8724), .B(n8722), .Z(n8723) );
  XNOR U9622 ( .A(n8725), .B(n8726), .Z(n8713) );
  NAND U9623 ( .A(n8727), .B(n8728), .Z(n8726) );
  XOR U9624 ( .A(n8729), .B(n8705), .Z(n8728) );
  XOR U9625 ( .A(n8719), .B(n8720), .Z(n8705) );
  XOR U9626 ( .A(n8730), .B(n8731), .Z(n8720) );
  ANDN U9627 ( .B(n8732), .A(n8733), .Z(n8730) );
  XOR U9628 ( .A(n8731), .B(n8734), .Z(n8732) );
  XOR U9629 ( .A(n8735), .B(n8736), .Z(n8719) );
  XOR U9630 ( .A(n8737), .B(n8738), .Z(n8736) );
  ANDN U9631 ( .B(n8739), .A(n8740), .Z(n8737) );
  XOR U9632 ( .A(n8741), .B(n8738), .Z(n8739) );
  IV U9633 ( .A(n8717), .Z(n8735) );
  XOR U9634 ( .A(n8742), .B(n8743), .Z(n8717) );
  ANDN U9635 ( .B(n8744), .A(n8745), .Z(n8742) );
  XOR U9636 ( .A(n8743), .B(n8746), .Z(n8744) );
  IV U9637 ( .A(n8725), .Z(n8729) );
  XOR U9638 ( .A(n8725), .B(n8707), .Z(n8727) );
  XOR U9639 ( .A(n8747), .B(n8748), .Z(n8707) );
  AND U9640 ( .A(n294), .B(n8749), .Z(n8747) );
  XOR U9641 ( .A(n8750), .B(n8748), .Z(n8749) );
  NANDN U9642 ( .A(n8709), .B(n8711), .Z(n8725) );
  XOR U9643 ( .A(n8751), .B(n8752), .Z(n8711) );
  AND U9644 ( .A(n294), .B(n8753), .Z(n8751) );
  XOR U9645 ( .A(n8752), .B(n8754), .Z(n8753) );
  XOR U9646 ( .A(n8755), .B(n8756), .Z(n294) );
  AND U9647 ( .A(n8757), .B(n8758), .Z(n8755) );
  XNOR U9648 ( .A(n8756), .B(n8722), .Z(n8758) );
  XNOR U9649 ( .A(n8759), .B(n8760), .Z(n8722) );
  ANDN U9650 ( .B(n8761), .A(n8762), .Z(n8759) );
  XOR U9651 ( .A(n8760), .B(n8763), .Z(n8761) );
  XOR U9652 ( .A(n8756), .B(n8724), .Z(n8757) );
  XOR U9653 ( .A(n8764), .B(n8765), .Z(n8724) );
  AND U9654 ( .A(n298), .B(n8766), .Z(n8764) );
  XOR U9655 ( .A(n8767), .B(n8765), .Z(n8766) );
  XNOR U9656 ( .A(n8768), .B(n8769), .Z(n8756) );
  NAND U9657 ( .A(n8770), .B(n8771), .Z(n8769) );
  XOR U9658 ( .A(n8772), .B(n8748), .Z(n8771) );
  XOR U9659 ( .A(n8762), .B(n8763), .Z(n8748) );
  XOR U9660 ( .A(n8773), .B(n8774), .Z(n8763) );
  ANDN U9661 ( .B(n8775), .A(n8776), .Z(n8773) );
  XOR U9662 ( .A(n8774), .B(n8777), .Z(n8775) );
  XOR U9663 ( .A(n8778), .B(n8779), .Z(n8762) );
  XOR U9664 ( .A(n8780), .B(n8781), .Z(n8779) );
  ANDN U9665 ( .B(n8782), .A(n8783), .Z(n8780) );
  XOR U9666 ( .A(n8784), .B(n8781), .Z(n8782) );
  IV U9667 ( .A(n8760), .Z(n8778) );
  XOR U9668 ( .A(n8785), .B(n8786), .Z(n8760) );
  ANDN U9669 ( .B(n8787), .A(n8788), .Z(n8785) );
  XOR U9670 ( .A(n8786), .B(n8789), .Z(n8787) );
  IV U9671 ( .A(n8768), .Z(n8772) );
  XOR U9672 ( .A(n8768), .B(n8750), .Z(n8770) );
  XOR U9673 ( .A(n8790), .B(n8791), .Z(n8750) );
  AND U9674 ( .A(n298), .B(n8792), .Z(n8790) );
  XOR U9675 ( .A(n8793), .B(n8791), .Z(n8792) );
  NANDN U9676 ( .A(n8752), .B(n8754), .Z(n8768) );
  XOR U9677 ( .A(n8794), .B(n8795), .Z(n8754) );
  AND U9678 ( .A(n298), .B(n8796), .Z(n8794) );
  XOR U9679 ( .A(n8795), .B(n8797), .Z(n8796) );
  XOR U9680 ( .A(n8798), .B(n8799), .Z(n298) );
  AND U9681 ( .A(n8800), .B(n8801), .Z(n8798) );
  XNOR U9682 ( .A(n8799), .B(n8765), .Z(n8801) );
  XNOR U9683 ( .A(n8802), .B(n8803), .Z(n8765) );
  ANDN U9684 ( .B(n8804), .A(n8805), .Z(n8802) );
  XOR U9685 ( .A(n8803), .B(n8806), .Z(n8804) );
  XOR U9686 ( .A(n8799), .B(n8767), .Z(n8800) );
  XOR U9687 ( .A(n8807), .B(n8808), .Z(n8767) );
  AND U9688 ( .A(n302), .B(n8809), .Z(n8807) );
  XOR U9689 ( .A(n8810), .B(n8808), .Z(n8809) );
  XNOR U9690 ( .A(n8811), .B(n8812), .Z(n8799) );
  NAND U9691 ( .A(n8813), .B(n8814), .Z(n8812) );
  XOR U9692 ( .A(n8815), .B(n8791), .Z(n8814) );
  XOR U9693 ( .A(n8805), .B(n8806), .Z(n8791) );
  XOR U9694 ( .A(n8816), .B(n8817), .Z(n8806) );
  ANDN U9695 ( .B(n8818), .A(n8819), .Z(n8816) );
  XOR U9696 ( .A(n8817), .B(n8820), .Z(n8818) );
  XOR U9697 ( .A(n8821), .B(n8822), .Z(n8805) );
  XOR U9698 ( .A(n8823), .B(n8824), .Z(n8822) );
  ANDN U9699 ( .B(n8825), .A(n8826), .Z(n8823) );
  XOR U9700 ( .A(n8827), .B(n8824), .Z(n8825) );
  IV U9701 ( .A(n8803), .Z(n8821) );
  XOR U9702 ( .A(n8828), .B(n8829), .Z(n8803) );
  ANDN U9703 ( .B(n8830), .A(n8831), .Z(n8828) );
  XOR U9704 ( .A(n8829), .B(n8832), .Z(n8830) );
  IV U9705 ( .A(n8811), .Z(n8815) );
  XOR U9706 ( .A(n8811), .B(n8793), .Z(n8813) );
  XOR U9707 ( .A(n8833), .B(n8834), .Z(n8793) );
  AND U9708 ( .A(n302), .B(n8835), .Z(n8833) );
  XOR U9709 ( .A(n8836), .B(n8834), .Z(n8835) );
  NANDN U9710 ( .A(n8795), .B(n8797), .Z(n8811) );
  XOR U9711 ( .A(n8837), .B(n8838), .Z(n8797) );
  AND U9712 ( .A(n302), .B(n8839), .Z(n8837) );
  XOR U9713 ( .A(n8838), .B(n8840), .Z(n8839) );
  XOR U9714 ( .A(n8841), .B(n8842), .Z(n302) );
  AND U9715 ( .A(n8843), .B(n8844), .Z(n8841) );
  XNOR U9716 ( .A(n8842), .B(n8808), .Z(n8844) );
  XNOR U9717 ( .A(n8845), .B(n8846), .Z(n8808) );
  ANDN U9718 ( .B(n8847), .A(n8848), .Z(n8845) );
  XOR U9719 ( .A(n8846), .B(n8849), .Z(n8847) );
  XOR U9720 ( .A(n8842), .B(n8810), .Z(n8843) );
  XOR U9721 ( .A(n8850), .B(n8851), .Z(n8810) );
  AND U9722 ( .A(n306), .B(n8852), .Z(n8850) );
  XOR U9723 ( .A(n8853), .B(n8851), .Z(n8852) );
  XNOR U9724 ( .A(n8854), .B(n8855), .Z(n8842) );
  NAND U9725 ( .A(n8856), .B(n8857), .Z(n8855) );
  XOR U9726 ( .A(n8858), .B(n8834), .Z(n8857) );
  XOR U9727 ( .A(n8848), .B(n8849), .Z(n8834) );
  XOR U9728 ( .A(n8859), .B(n8860), .Z(n8849) );
  ANDN U9729 ( .B(n8861), .A(n8862), .Z(n8859) );
  XOR U9730 ( .A(n8860), .B(n8863), .Z(n8861) );
  XOR U9731 ( .A(n8864), .B(n8865), .Z(n8848) );
  XOR U9732 ( .A(n8866), .B(n8867), .Z(n8865) );
  ANDN U9733 ( .B(n8868), .A(n8869), .Z(n8866) );
  XOR U9734 ( .A(n8870), .B(n8867), .Z(n8868) );
  IV U9735 ( .A(n8846), .Z(n8864) );
  XOR U9736 ( .A(n8871), .B(n8872), .Z(n8846) );
  ANDN U9737 ( .B(n8873), .A(n8874), .Z(n8871) );
  XOR U9738 ( .A(n8872), .B(n8875), .Z(n8873) );
  IV U9739 ( .A(n8854), .Z(n8858) );
  XOR U9740 ( .A(n8854), .B(n8836), .Z(n8856) );
  XOR U9741 ( .A(n8876), .B(n8877), .Z(n8836) );
  AND U9742 ( .A(n306), .B(n8878), .Z(n8876) );
  XOR U9743 ( .A(n8879), .B(n8877), .Z(n8878) );
  NANDN U9744 ( .A(n8838), .B(n8840), .Z(n8854) );
  XOR U9745 ( .A(n8880), .B(n8881), .Z(n8840) );
  AND U9746 ( .A(n306), .B(n8882), .Z(n8880) );
  XOR U9747 ( .A(n8881), .B(n8883), .Z(n8882) );
  XOR U9748 ( .A(n8884), .B(n8885), .Z(n306) );
  AND U9749 ( .A(n8886), .B(n8887), .Z(n8884) );
  XNOR U9750 ( .A(n8885), .B(n8851), .Z(n8887) );
  XNOR U9751 ( .A(n8888), .B(n8889), .Z(n8851) );
  ANDN U9752 ( .B(n8890), .A(n8891), .Z(n8888) );
  XOR U9753 ( .A(n8889), .B(n8892), .Z(n8890) );
  XOR U9754 ( .A(n8885), .B(n8853), .Z(n8886) );
  XOR U9755 ( .A(n8893), .B(n8894), .Z(n8853) );
  AND U9756 ( .A(n310), .B(n8895), .Z(n8893) );
  XOR U9757 ( .A(n8896), .B(n8894), .Z(n8895) );
  XNOR U9758 ( .A(n8897), .B(n8898), .Z(n8885) );
  NAND U9759 ( .A(n8899), .B(n8900), .Z(n8898) );
  XOR U9760 ( .A(n8901), .B(n8877), .Z(n8900) );
  XOR U9761 ( .A(n8891), .B(n8892), .Z(n8877) );
  XOR U9762 ( .A(n8902), .B(n8903), .Z(n8892) );
  ANDN U9763 ( .B(n8904), .A(n8905), .Z(n8902) );
  XOR U9764 ( .A(n8903), .B(n8906), .Z(n8904) );
  XOR U9765 ( .A(n8907), .B(n8908), .Z(n8891) );
  XOR U9766 ( .A(n8909), .B(n8910), .Z(n8908) );
  ANDN U9767 ( .B(n8911), .A(n8912), .Z(n8909) );
  XOR U9768 ( .A(n8913), .B(n8910), .Z(n8911) );
  IV U9769 ( .A(n8889), .Z(n8907) );
  XOR U9770 ( .A(n8914), .B(n8915), .Z(n8889) );
  ANDN U9771 ( .B(n8916), .A(n8917), .Z(n8914) );
  XOR U9772 ( .A(n8915), .B(n8918), .Z(n8916) );
  IV U9773 ( .A(n8897), .Z(n8901) );
  XOR U9774 ( .A(n8897), .B(n8879), .Z(n8899) );
  XOR U9775 ( .A(n8919), .B(n8920), .Z(n8879) );
  AND U9776 ( .A(n310), .B(n8921), .Z(n8919) );
  XOR U9777 ( .A(n8922), .B(n8920), .Z(n8921) );
  NANDN U9778 ( .A(n8881), .B(n8883), .Z(n8897) );
  XOR U9779 ( .A(n8923), .B(n8924), .Z(n8883) );
  AND U9780 ( .A(n310), .B(n8925), .Z(n8923) );
  XOR U9781 ( .A(n8924), .B(n8926), .Z(n8925) );
  XOR U9782 ( .A(n8927), .B(n8928), .Z(n310) );
  AND U9783 ( .A(n8929), .B(n8930), .Z(n8927) );
  XNOR U9784 ( .A(n8928), .B(n8894), .Z(n8930) );
  XNOR U9785 ( .A(n8931), .B(n8932), .Z(n8894) );
  ANDN U9786 ( .B(n8933), .A(n8934), .Z(n8931) );
  XOR U9787 ( .A(n8932), .B(n8935), .Z(n8933) );
  XOR U9788 ( .A(n8928), .B(n8896), .Z(n8929) );
  XOR U9789 ( .A(n8936), .B(n8937), .Z(n8896) );
  AND U9790 ( .A(n314), .B(n8938), .Z(n8936) );
  XOR U9791 ( .A(n8939), .B(n8937), .Z(n8938) );
  XNOR U9792 ( .A(n8940), .B(n8941), .Z(n8928) );
  NAND U9793 ( .A(n8942), .B(n8943), .Z(n8941) );
  XOR U9794 ( .A(n8944), .B(n8920), .Z(n8943) );
  XOR U9795 ( .A(n8934), .B(n8935), .Z(n8920) );
  XOR U9796 ( .A(n8945), .B(n8946), .Z(n8935) );
  ANDN U9797 ( .B(n8947), .A(n8948), .Z(n8945) );
  XOR U9798 ( .A(n8946), .B(n8949), .Z(n8947) );
  XOR U9799 ( .A(n8950), .B(n8951), .Z(n8934) );
  XOR U9800 ( .A(n8952), .B(n8953), .Z(n8951) );
  ANDN U9801 ( .B(n8954), .A(n8955), .Z(n8952) );
  XOR U9802 ( .A(n8956), .B(n8953), .Z(n8954) );
  IV U9803 ( .A(n8932), .Z(n8950) );
  XOR U9804 ( .A(n8957), .B(n8958), .Z(n8932) );
  ANDN U9805 ( .B(n8959), .A(n8960), .Z(n8957) );
  XOR U9806 ( .A(n8958), .B(n8961), .Z(n8959) );
  IV U9807 ( .A(n8940), .Z(n8944) );
  XOR U9808 ( .A(n8940), .B(n8922), .Z(n8942) );
  XOR U9809 ( .A(n8962), .B(n8963), .Z(n8922) );
  AND U9810 ( .A(n314), .B(n8964), .Z(n8962) );
  XOR U9811 ( .A(n8965), .B(n8963), .Z(n8964) );
  NANDN U9812 ( .A(n8924), .B(n8926), .Z(n8940) );
  XOR U9813 ( .A(n8966), .B(n8967), .Z(n8926) );
  AND U9814 ( .A(n314), .B(n8968), .Z(n8966) );
  XOR U9815 ( .A(n8967), .B(n8969), .Z(n8968) );
  XOR U9816 ( .A(n8970), .B(n8971), .Z(n314) );
  AND U9817 ( .A(n8972), .B(n8973), .Z(n8970) );
  XNOR U9818 ( .A(n8971), .B(n8937), .Z(n8973) );
  XNOR U9819 ( .A(n8974), .B(n8975), .Z(n8937) );
  ANDN U9820 ( .B(n8976), .A(n8977), .Z(n8974) );
  XOR U9821 ( .A(n8975), .B(n8978), .Z(n8976) );
  XOR U9822 ( .A(n8971), .B(n8939), .Z(n8972) );
  XOR U9823 ( .A(n8979), .B(n8980), .Z(n8939) );
  AND U9824 ( .A(n318), .B(n8981), .Z(n8979) );
  XOR U9825 ( .A(n8982), .B(n8980), .Z(n8981) );
  XNOR U9826 ( .A(n8983), .B(n8984), .Z(n8971) );
  NAND U9827 ( .A(n8985), .B(n8986), .Z(n8984) );
  XOR U9828 ( .A(n8987), .B(n8963), .Z(n8986) );
  XOR U9829 ( .A(n8977), .B(n8978), .Z(n8963) );
  XOR U9830 ( .A(n8988), .B(n8989), .Z(n8978) );
  ANDN U9831 ( .B(n8990), .A(n8991), .Z(n8988) );
  XOR U9832 ( .A(n8989), .B(n8992), .Z(n8990) );
  XOR U9833 ( .A(n8993), .B(n8994), .Z(n8977) );
  XOR U9834 ( .A(n8995), .B(n8996), .Z(n8994) );
  ANDN U9835 ( .B(n8997), .A(n8998), .Z(n8995) );
  XOR U9836 ( .A(n8999), .B(n8996), .Z(n8997) );
  IV U9837 ( .A(n8975), .Z(n8993) );
  XOR U9838 ( .A(n9000), .B(n9001), .Z(n8975) );
  ANDN U9839 ( .B(n9002), .A(n9003), .Z(n9000) );
  XOR U9840 ( .A(n9001), .B(n9004), .Z(n9002) );
  IV U9841 ( .A(n8983), .Z(n8987) );
  XOR U9842 ( .A(n8983), .B(n8965), .Z(n8985) );
  XOR U9843 ( .A(n9005), .B(n9006), .Z(n8965) );
  AND U9844 ( .A(n318), .B(n9007), .Z(n9005) );
  XOR U9845 ( .A(n9008), .B(n9006), .Z(n9007) );
  NANDN U9846 ( .A(n8967), .B(n8969), .Z(n8983) );
  XOR U9847 ( .A(n9009), .B(n9010), .Z(n8969) );
  AND U9848 ( .A(n318), .B(n9011), .Z(n9009) );
  XOR U9849 ( .A(n9010), .B(n9012), .Z(n9011) );
  XOR U9850 ( .A(n9013), .B(n9014), .Z(n318) );
  AND U9851 ( .A(n9015), .B(n9016), .Z(n9013) );
  XNOR U9852 ( .A(n9014), .B(n8980), .Z(n9016) );
  XNOR U9853 ( .A(n9017), .B(n9018), .Z(n8980) );
  ANDN U9854 ( .B(n9019), .A(n9020), .Z(n9017) );
  XOR U9855 ( .A(n9018), .B(n9021), .Z(n9019) );
  XOR U9856 ( .A(n9014), .B(n8982), .Z(n9015) );
  XOR U9857 ( .A(n9022), .B(n9023), .Z(n8982) );
  AND U9858 ( .A(n322), .B(n9024), .Z(n9022) );
  XOR U9859 ( .A(n9025), .B(n9023), .Z(n9024) );
  XNOR U9860 ( .A(n9026), .B(n9027), .Z(n9014) );
  NAND U9861 ( .A(n9028), .B(n9029), .Z(n9027) );
  XOR U9862 ( .A(n9030), .B(n9006), .Z(n9029) );
  XOR U9863 ( .A(n9020), .B(n9021), .Z(n9006) );
  XOR U9864 ( .A(n9031), .B(n9032), .Z(n9021) );
  ANDN U9865 ( .B(n9033), .A(n9034), .Z(n9031) );
  XOR U9866 ( .A(n9032), .B(n9035), .Z(n9033) );
  XOR U9867 ( .A(n9036), .B(n9037), .Z(n9020) );
  XOR U9868 ( .A(n9038), .B(n9039), .Z(n9037) );
  ANDN U9869 ( .B(n9040), .A(n9041), .Z(n9038) );
  XOR U9870 ( .A(n9042), .B(n9039), .Z(n9040) );
  IV U9871 ( .A(n9018), .Z(n9036) );
  XOR U9872 ( .A(n9043), .B(n9044), .Z(n9018) );
  ANDN U9873 ( .B(n9045), .A(n9046), .Z(n9043) );
  XOR U9874 ( .A(n9044), .B(n9047), .Z(n9045) );
  IV U9875 ( .A(n9026), .Z(n9030) );
  XOR U9876 ( .A(n9026), .B(n9008), .Z(n9028) );
  XOR U9877 ( .A(n9048), .B(n9049), .Z(n9008) );
  AND U9878 ( .A(n322), .B(n9050), .Z(n9048) );
  XOR U9879 ( .A(n9051), .B(n9049), .Z(n9050) );
  NANDN U9880 ( .A(n9010), .B(n9012), .Z(n9026) );
  XOR U9881 ( .A(n9052), .B(n9053), .Z(n9012) );
  AND U9882 ( .A(n322), .B(n9054), .Z(n9052) );
  XOR U9883 ( .A(n9053), .B(n9055), .Z(n9054) );
  XOR U9884 ( .A(n9056), .B(n9057), .Z(n322) );
  AND U9885 ( .A(n9058), .B(n9059), .Z(n9056) );
  XNOR U9886 ( .A(n9057), .B(n9023), .Z(n9059) );
  XNOR U9887 ( .A(n9060), .B(n9061), .Z(n9023) );
  ANDN U9888 ( .B(n9062), .A(n9063), .Z(n9060) );
  XOR U9889 ( .A(n9061), .B(n9064), .Z(n9062) );
  XOR U9890 ( .A(n9057), .B(n9025), .Z(n9058) );
  XOR U9891 ( .A(n9065), .B(n9066), .Z(n9025) );
  AND U9892 ( .A(n326), .B(n9067), .Z(n9065) );
  XOR U9893 ( .A(n9068), .B(n9066), .Z(n9067) );
  XNOR U9894 ( .A(n9069), .B(n9070), .Z(n9057) );
  NAND U9895 ( .A(n9071), .B(n9072), .Z(n9070) );
  XOR U9896 ( .A(n9073), .B(n9049), .Z(n9072) );
  XOR U9897 ( .A(n9063), .B(n9064), .Z(n9049) );
  XOR U9898 ( .A(n9074), .B(n9075), .Z(n9064) );
  ANDN U9899 ( .B(n9076), .A(n9077), .Z(n9074) );
  XOR U9900 ( .A(n9075), .B(n9078), .Z(n9076) );
  XOR U9901 ( .A(n9079), .B(n9080), .Z(n9063) );
  XOR U9902 ( .A(n9081), .B(n9082), .Z(n9080) );
  ANDN U9903 ( .B(n9083), .A(n9084), .Z(n9081) );
  XOR U9904 ( .A(n9085), .B(n9082), .Z(n9083) );
  IV U9905 ( .A(n9061), .Z(n9079) );
  XOR U9906 ( .A(n9086), .B(n9087), .Z(n9061) );
  ANDN U9907 ( .B(n9088), .A(n9089), .Z(n9086) );
  XOR U9908 ( .A(n9087), .B(n9090), .Z(n9088) );
  IV U9909 ( .A(n9069), .Z(n9073) );
  XOR U9910 ( .A(n9069), .B(n9051), .Z(n9071) );
  XOR U9911 ( .A(n9091), .B(n9092), .Z(n9051) );
  AND U9912 ( .A(n326), .B(n9093), .Z(n9091) );
  XOR U9913 ( .A(n9094), .B(n9092), .Z(n9093) );
  NANDN U9914 ( .A(n9053), .B(n9055), .Z(n9069) );
  XOR U9915 ( .A(n9095), .B(n9096), .Z(n9055) );
  AND U9916 ( .A(n326), .B(n9097), .Z(n9095) );
  XOR U9917 ( .A(n9096), .B(n9098), .Z(n9097) );
  XOR U9918 ( .A(n9099), .B(n9100), .Z(n326) );
  AND U9919 ( .A(n9101), .B(n9102), .Z(n9099) );
  XNOR U9920 ( .A(n9100), .B(n9066), .Z(n9102) );
  XNOR U9921 ( .A(n9103), .B(n9104), .Z(n9066) );
  ANDN U9922 ( .B(n9105), .A(n9106), .Z(n9103) );
  XOR U9923 ( .A(n9104), .B(n9107), .Z(n9105) );
  XOR U9924 ( .A(n9100), .B(n9068), .Z(n9101) );
  XOR U9925 ( .A(n9108), .B(n9109), .Z(n9068) );
  AND U9926 ( .A(n330), .B(n9110), .Z(n9108) );
  XOR U9927 ( .A(n9111), .B(n9109), .Z(n9110) );
  XNOR U9928 ( .A(n9112), .B(n9113), .Z(n9100) );
  NAND U9929 ( .A(n9114), .B(n9115), .Z(n9113) );
  XOR U9930 ( .A(n9116), .B(n9092), .Z(n9115) );
  XOR U9931 ( .A(n9106), .B(n9107), .Z(n9092) );
  XOR U9932 ( .A(n9117), .B(n9118), .Z(n9107) );
  ANDN U9933 ( .B(n9119), .A(n9120), .Z(n9117) );
  XOR U9934 ( .A(n9118), .B(n9121), .Z(n9119) );
  XOR U9935 ( .A(n9122), .B(n9123), .Z(n9106) );
  XOR U9936 ( .A(n9124), .B(n9125), .Z(n9123) );
  ANDN U9937 ( .B(n9126), .A(n9127), .Z(n9124) );
  XOR U9938 ( .A(n9128), .B(n9125), .Z(n9126) );
  IV U9939 ( .A(n9104), .Z(n9122) );
  XOR U9940 ( .A(n9129), .B(n9130), .Z(n9104) );
  ANDN U9941 ( .B(n9131), .A(n9132), .Z(n9129) );
  XOR U9942 ( .A(n9130), .B(n9133), .Z(n9131) );
  IV U9943 ( .A(n9112), .Z(n9116) );
  XOR U9944 ( .A(n9112), .B(n9094), .Z(n9114) );
  XOR U9945 ( .A(n9134), .B(n9135), .Z(n9094) );
  AND U9946 ( .A(n330), .B(n9136), .Z(n9134) );
  XOR U9947 ( .A(n9137), .B(n9135), .Z(n9136) );
  NANDN U9948 ( .A(n9096), .B(n9098), .Z(n9112) );
  XOR U9949 ( .A(n9138), .B(n9139), .Z(n9098) );
  AND U9950 ( .A(n330), .B(n9140), .Z(n9138) );
  XOR U9951 ( .A(n9139), .B(n9141), .Z(n9140) );
  XOR U9952 ( .A(n9142), .B(n9143), .Z(n330) );
  AND U9953 ( .A(n9144), .B(n9145), .Z(n9142) );
  XNOR U9954 ( .A(n9143), .B(n9109), .Z(n9145) );
  XNOR U9955 ( .A(n9146), .B(n9147), .Z(n9109) );
  ANDN U9956 ( .B(n9148), .A(n9149), .Z(n9146) );
  XOR U9957 ( .A(n9147), .B(n9150), .Z(n9148) );
  XOR U9958 ( .A(n9143), .B(n9111), .Z(n9144) );
  XOR U9959 ( .A(n9151), .B(n9152), .Z(n9111) );
  AND U9960 ( .A(n334), .B(n9153), .Z(n9151) );
  XOR U9961 ( .A(n9154), .B(n9152), .Z(n9153) );
  XNOR U9962 ( .A(n9155), .B(n9156), .Z(n9143) );
  NAND U9963 ( .A(n9157), .B(n9158), .Z(n9156) );
  XOR U9964 ( .A(n9159), .B(n9135), .Z(n9158) );
  XOR U9965 ( .A(n9149), .B(n9150), .Z(n9135) );
  XOR U9966 ( .A(n9160), .B(n9161), .Z(n9150) );
  ANDN U9967 ( .B(n9162), .A(n9163), .Z(n9160) );
  XOR U9968 ( .A(n9161), .B(n9164), .Z(n9162) );
  XOR U9969 ( .A(n9165), .B(n9166), .Z(n9149) );
  XOR U9970 ( .A(n9167), .B(n9168), .Z(n9166) );
  ANDN U9971 ( .B(n9169), .A(n9170), .Z(n9167) );
  XOR U9972 ( .A(n9171), .B(n9168), .Z(n9169) );
  IV U9973 ( .A(n9147), .Z(n9165) );
  XOR U9974 ( .A(n9172), .B(n9173), .Z(n9147) );
  ANDN U9975 ( .B(n9174), .A(n9175), .Z(n9172) );
  XOR U9976 ( .A(n9173), .B(n9176), .Z(n9174) );
  IV U9977 ( .A(n9155), .Z(n9159) );
  XOR U9978 ( .A(n9155), .B(n9137), .Z(n9157) );
  XOR U9979 ( .A(n9177), .B(n9178), .Z(n9137) );
  AND U9980 ( .A(n334), .B(n9179), .Z(n9177) );
  XOR U9981 ( .A(n9180), .B(n9178), .Z(n9179) );
  NANDN U9982 ( .A(n9139), .B(n9141), .Z(n9155) );
  XOR U9983 ( .A(n9181), .B(n9182), .Z(n9141) );
  AND U9984 ( .A(n334), .B(n9183), .Z(n9181) );
  XOR U9985 ( .A(n9182), .B(n9184), .Z(n9183) );
  XOR U9986 ( .A(n9185), .B(n9186), .Z(n334) );
  AND U9987 ( .A(n9187), .B(n9188), .Z(n9185) );
  XNOR U9988 ( .A(n9186), .B(n9152), .Z(n9188) );
  XNOR U9989 ( .A(n9189), .B(n9190), .Z(n9152) );
  ANDN U9990 ( .B(n9191), .A(n9192), .Z(n9189) );
  XOR U9991 ( .A(n9190), .B(n9193), .Z(n9191) );
  XOR U9992 ( .A(n9186), .B(n9154), .Z(n9187) );
  XOR U9993 ( .A(n9194), .B(n9195), .Z(n9154) );
  AND U9994 ( .A(n338), .B(n9196), .Z(n9194) );
  XOR U9995 ( .A(n9197), .B(n9195), .Z(n9196) );
  XNOR U9996 ( .A(n9198), .B(n9199), .Z(n9186) );
  NAND U9997 ( .A(n9200), .B(n9201), .Z(n9199) );
  XOR U9998 ( .A(n9202), .B(n9178), .Z(n9201) );
  XOR U9999 ( .A(n9192), .B(n9193), .Z(n9178) );
  XOR U10000 ( .A(n9203), .B(n9204), .Z(n9193) );
  ANDN U10001 ( .B(n9205), .A(n9206), .Z(n9203) );
  XOR U10002 ( .A(n9204), .B(n9207), .Z(n9205) );
  XOR U10003 ( .A(n9208), .B(n9209), .Z(n9192) );
  XOR U10004 ( .A(n9210), .B(n9211), .Z(n9209) );
  ANDN U10005 ( .B(n9212), .A(n9213), .Z(n9210) );
  XOR U10006 ( .A(n9214), .B(n9211), .Z(n9212) );
  IV U10007 ( .A(n9190), .Z(n9208) );
  XOR U10008 ( .A(n9215), .B(n9216), .Z(n9190) );
  ANDN U10009 ( .B(n9217), .A(n9218), .Z(n9215) );
  XOR U10010 ( .A(n9216), .B(n9219), .Z(n9217) );
  IV U10011 ( .A(n9198), .Z(n9202) );
  XOR U10012 ( .A(n9198), .B(n9180), .Z(n9200) );
  XOR U10013 ( .A(n9220), .B(n9221), .Z(n9180) );
  AND U10014 ( .A(n338), .B(n9222), .Z(n9220) );
  XOR U10015 ( .A(n9223), .B(n9221), .Z(n9222) );
  NANDN U10016 ( .A(n9182), .B(n9184), .Z(n9198) );
  XOR U10017 ( .A(n9224), .B(n9225), .Z(n9184) );
  AND U10018 ( .A(n338), .B(n9226), .Z(n9224) );
  XOR U10019 ( .A(n9225), .B(n9227), .Z(n9226) );
  XOR U10020 ( .A(n9228), .B(n9229), .Z(n338) );
  AND U10021 ( .A(n9230), .B(n9231), .Z(n9228) );
  XNOR U10022 ( .A(n9229), .B(n9195), .Z(n9231) );
  XNOR U10023 ( .A(n9232), .B(n9233), .Z(n9195) );
  ANDN U10024 ( .B(n9234), .A(n9235), .Z(n9232) );
  XOR U10025 ( .A(n9233), .B(n9236), .Z(n9234) );
  XOR U10026 ( .A(n9229), .B(n9197), .Z(n9230) );
  XOR U10027 ( .A(n9237), .B(n9238), .Z(n9197) );
  AND U10028 ( .A(n342), .B(n9239), .Z(n9237) );
  XOR U10029 ( .A(n9240), .B(n9238), .Z(n9239) );
  XNOR U10030 ( .A(n9241), .B(n9242), .Z(n9229) );
  NAND U10031 ( .A(n9243), .B(n9244), .Z(n9242) );
  XOR U10032 ( .A(n9245), .B(n9221), .Z(n9244) );
  XOR U10033 ( .A(n9235), .B(n9236), .Z(n9221) );
  XOR U10034 ( .A(n9246), .B(n9247), .Z(n9236) );
  ANDN U10035 ( .B(n9248), .A(n9249), .Z(n9246) );
  XOR U10036 ( .A(n9247), .B(n9250), .Z(n9248) );
  XOR U10037 ( .A(n9251), .B(n9252), .Z(n9235) );
  XOR U10038 ( .A(n9253), .B(n9254), .Z(n9252) );
  ANDN U10039 ( .B(n9255), .A(n9256), .Z(n9253) );
  XOR U10040 ( .A(n9257), .B(n9254), .Z(n9255) );
  IV U10041 ( .A(n9233), .Z(n9251) );
  XOR U10042 ( .A(n9258), .B(n9259), .Z(n9233) );
  ANDN U10043 ( .B(n9260), .A(n9261), .Z(n9258) );
  XOR U10044 ( .A(n9259), .B(n9262), .Z(n9260) );
  IV U10045 ( .A(n9241), .Z(n9245) );
  XOR U10046 ( .A(n9241), .B(n9223), .Z(n9243) );
  XOR U10047 ( .A(n9263), .B(n9264), .Z(n9223) );
  AND U10048 ( .A(n342), .B(n9265), .Z(n9263) );
  XOR U10049 ( .A(n9266), .B(n9264), .Z(n9265) );
  NANDN U10050 ( .A(n9225), .B(n9227), .Z(n9241) );
  XOR U10051 ( .A(n9267), .B(n9268), .Z(n9227) );
  AND U10052 ( .A(n342), .B(n9269), .Z(n9267) );
  XOR U10053 ( .A(n9268), .B(n9270), .Z(n9269) );
  XOR U10054 ( .A(n9271), .B(n9272), .Z(n342) );
  AND U10055 ( .A(n9273), .B(n9274), .Z(n9271) );
  XNOR U10056 ( .A(n9272), .B(n9238), .Z(n9274) );
  XNOR U10057 ( .A(n9275), .B(n9276), .Z(n9238) );
  ANDN U10058 ( .B(n9277), .A(n9278), .Z(n9275) );
  XOR U10059 ( .A(n9276), .B(n9279), .Z(n9277) );
  XOR U10060 ( .A(n9272), .B(n9240), .Z(n9273) );
  XOR U10061 ( .A(n9280), .B(n9281), .Z(n9240) );
  AND U10062 ( .A(n346), .B(n9282), .Z(n9280) );
  XOR U10063 ( .A(n9283), .B(n9281), .Z(n9282) );
  XNOR U10064 ( .A(n9284), .B(n9285), .Z(n9272) );
  NAND U10065 ( .A(n9286), .B(n9287), .Z(n9285) );
  XOR U10066 ( .A(n9288), .B(n9264), .Z(n9287) );
  XOR U10067 ( .A(n9278), .B(n9279), .Z(n9264) );
  XOR U10068 ( .A(n9289), .B(n9290), .Z(n9279) );
  ANDN U10069 ( .B(n9291), .A(n9292), .Z(n9289) );
  XOR U10070 ( .A(n9290), .B(n9293), .Z(n9291) );
  XOR U10071 ( .A(n9294), .B(n9295), .Z(n9278) );
  XOR U10072 ( .A(n9296), .B(n9297), .Z(n9295) );
  ANDN U10073 ( .B(n9298), .A(n9299), .Z(n9296) );
  XOR U10074 ( .A(n9300), .B(n9297), .Z(n9298) );
  IV U10075 ( .A(n9276), .Z(n9294) );
  XOR U10076 ( .A(n9301), .B(n9302), .Z(n9276) );
  ANDN U10077 ( .B(n9303), .A(n9304), .Z(n9301) );
  XOR U10078 ( .A(n9302), .B(n9305), .Z(n9303) );
  IV U10079 ( .A(n9284), .Z(n9288) );
  XOR U10080 ( .A(n9284), .B(n9266), .Z(n9286) );
  XOR U10081 ( .A(n9306), .B(n9307), .Z(n9266) );
  AND U10082 ( .A(n346), .B(n9308), .Z(n9306) );
  XOR U10083 ( .A(n9309), .B(n9307), .Z(n9308) );
  NANDN U10084 ( .A(n9268), .B(n9270), .Z(n9284) );
  XOR U10085 ( .A(n9310), .B(n9311), .Z(n9270) );
  AND U10086 ( .A(n346), .B(n9312), .Z(n9310) );
  XOR U10087 ( .A(n9311), .B(n9313), .Z(n9312) );
  XOR U10088 ( .A(n9314), .B(n9315), .Z(n346) );
  AND U10089 ( .A(n9316), .B(n9317), .Z(n9314) );
  XNOR U10090 ( .A(n9315), .B(n9281), .Z(n9317) );
  XNOR U10091 ( .A(n9318), .B(n9319), .Z(n9281) );
  ANDN U10092 ( .B(n9320), .A(n9321), .Z(n9318) );
  XOR U10093 ( .A(n9319), .B(n9322), .Z(n9320) );
  XOR U10094 ( .A(n9315), .B(n9283), .Z(n9316) );
  XOR U10095 ( .A(n9323), .B(n9324), .Z(n9283) );
  AND U10096 ( .A(n350), .B(n9325), .Z(n9323) );
  XOR U10097 ( .A(n9326), .B(n9324), .Z(n9325) );
  XNOR U10098 ( .A(n9327), .B(n9328), .Z(n9315) );
  NAND U10099 ( .A(n9329), .B(n9330), .Z(n9328) );
  XOR U10100 ( .A(n9331), .B(n9307), .Z(n9330) );
  XOR U10101 ( .A(n9321), .B(n9322), .Z(n9307) );
  XOR U10102 ( .A(n9332), .B(n9333), .Z(n9322) );
  ANDN U10103 ( .B(n9334), .A(n9335), .Z(n9332) );
  XOR U10104 ( .A(n9333), .B(n9336), .Z(n9334) );
  XOR U10105 ( .A(n9337), .B(n9338), .Z(n9321) );
  XOR U10106 ( .A(n9339), .B(n9340), .Z(n9338) );
  ANDN U10107 ( .B(n9341), .A(n9342), .Z(n9339) );
  XOR U10108 ( .A(n9343), .B(n9340), .Z(n9341) );
  IV U10109 ( .A(n9319), .Z(n9337) );
  XOR U10110 ( .A(n9344), .B(n9345), .Z(n9319) );
  ANDN U10111 ( .B(n9346), .A(n9347), .Z(n9344) );
  XOR U10112 ( .A(n9345), .B(n9348), .Z(n9346) );
  IV U10113 ( .A(n9327), .Z(n9331) );
  XOR U10114 ( .A(n9327), .B(n9309), .Z(n9329) );
  XOR U10115 ( .A(n9349), .B(n9350), .Z(n9309) );
  AND U10116 ( .A(n350), .B(n9351), .Z(n9349) );
  XOR U10117 ( .A(n9352), .B(n9350), .Z(n9351) );
  NANDN U10118 ( .A(n9311), .B(n9313), .Z(n9327) );
  XOR U10119 ( .A(n9353), .B(n9354), .Z(n9313) );
  AND U10120 ( .A(n350), .B(n9355), .Z(n9353) );
  XOR U10121 ( .A(n9354), .B(n9356), .Z(n9355) );
  XOR U10122 ( .A(n9357), .B(n9358), .Z(n350) );
  AND U10123 ( .A(n9359), .B(n9360), .Z(n9357) );
  XNOR U10124 ( .A(n9358), .B(n9324), .Z(n9360) );
  XNOR U10125 ( .A(n9361), .B(n9362), .Z(n9324) );
  ANDN U10126 ( .B(n9363), .A(n9364), .Z(n9361) );
  XOR U10127 ( .A(n9362), .B(n9365), .Z(n9363) );
  XOR U10128 ( .A(n9358), .B(n9326), .Z(n9359) );
  XOR U10129 ( .A(n9366), .B(n9367), .Z(n9326) );
  AND U10130 ( .A(n354), .B(n9368), .Z(n9366) );
  XOR U10131 ( .A(n9369), .B(n9367), .Z(n9368) );
  XNOR U10132 ( .A(n9370), .B(n9371), .Z(n9358) );
  NAND U10133 ( .A(n9372), .B(n9373), .Z(n9371) );
  XOR U10134 ( .A(n9374), .B(n9350), .Z(n9373) );
  XOR U10135 ( .A(n9364), .B(n9365), .Z(n9350) );
  XOR U10136 ( .A(n9375), .B(n9376), .Z(n9365) );
  ANDN U10137 ( .B(n9377), .A(n9378), .Z(n9375) );
  XOR U10138 ( .A(n9376), .B(n9379), .Z(n9377) );
  XOR U10139 ( .A(n9380), .B(n9381), .Z(n9364) );
  XOR U10140 ( .A(n9382), .B(n9383), .Z(n9381) );
  ANDN U10141 ( .B(n9384), .A(n9385), .Z(n9382) );
  XOR U10142 ( .A(n9386), .B(n9383), .Z(n9384) );
  IV U10143 ( .A(n9362), .Z(n9380) );
  XOR U10144 ( .A(n9387), .B(n9388), .Z(n9362) );
  ANDN U10145 ( .B(n9389), .A(n9390), .Z(n9387) );
  XOR U10146 ( .A(n9388), .B(n9391), .Z(n9389) );
  IV U10147 ( .A(n9370), .Z(n9374) );
  XOR U10148 ( .A(n9370), .B(n9352), .Z(n9372) );
  XOR U10149 ( .A(n9392), .B(n9393), .Z(n9352) );
  AND U10150 ( .A(n354), .B(n9394), .Z(n9392) );
  XOR U10151 ( .A(n9395), .B(n9393), .Z(n9394) );
  NANDN U10152 ( .A(n9354), .B(n9356), .Z(n9370) );
  XOR U10153 ( .A(n9396), .B(n9397), .Z(n9356) );
  AND U10154 ( .A(n354), .B(n9398), .Z(n9396) );
  XOR U10155 ( .A(n9397), .B(n9399), .Z(n9398) );
  XOR U10156 ( .A(n9400), .B(n9401), .Z(n354) );
  AND U10157 ( .A(n9402), .B(n9403), .Z(n9400) );
  XNOR U10158 ( .A(n9401), .B(n9367), .Z(n9403) );
  XNOR U10159 ( .A(n9404), .B(n9405), .Z(n9367) );
  ANDN U10160 ( .B(n9406), .A(n9407), .Z(n9404) );
  XOR U10161 ( .A(n9405), .B(n9408), .Z(n9406) );
  XOR U10162 ( .A(n9401), .B(n9369), .Z(n9402) );
  XOR U10163 ( .A(n9409), .B(n9410), .Z(n9369) );
  AND U10164 ( .A(n358), .B(n9411), .Z(n9409) );
  XOR U10165 ( .A(n9412), .B(n9410), .Z(n9411) );
  XNOR U10166 ( .A(n9413), .B(n9414), .Z(n9401) );
  NAND U10167 ( .A(n9415), .B(n9416), .Z(n9414) );
  XOR U10168 ( .A(n9417), .B(n9393), .Z(n9416) );
  XOR U10169 ( .A(n9407), .B(n9408), .Z(n9393) );
  XOR U10170 ( .A(n9418), .B(n9419), .Z(n9408) );
  ANDN U10171 ( .B(n9420), .A(n9421), .Z(n9418) );
  XOR U10172 ( .A(n9419), .B(n9422), .Z(n9420) );
  XOR U10173 ( .A(n9423), .B(n9424), .Z(n9407) );
  XOR U10174 ( .A(n9425), .B(n9426), .Z(n9424) );
  ANDN U10175 ( .B(n9427), .A(n9428), .Z(n9425) );
  XOR U10176 ( .A(n9429), .B(n9426), .Z(n9427) );
  IV U10177 ( .A(n9405), .Z(n9423) );
  XOR U10178 ( .A(n9430), .B(n9431), .Z(n9405) );
  ANDN U10179 ( .B(n9432), .A(n9433), .Z(n9430) );
  XOR U10180 ( .A(n9431), .B(n9434), .Z(n9432) );
  IV U10181 ( .A(n9413), .Z(n9417) );
  XOR U10182 ( .A(n9413), .B(n9395), .Z(n9415) );
  XOR U10183 ( .A(n9435), .B(n9436), .Z(n9395) );
  AND U10184 ( .A(n358), .B(n9437), .Z(n9435) );
  XOR U10185 ( .A(n9438), .B(n9436), .Z(n9437) );
  NANDN U10186 ( .A(n9397), .B(n9399), .Z(n9413) );
  XOR U10187 ( .A(n9439), .B(n9440), .Z(n9399) );
  AND U10188 ( .A(n358), .B(n9441), .Z(n9439) );
  XOR U10189 ( .A(n9440), .B(n9442), .Z(n9441) );
  XOR U10190 ( .A(n9443), .B(n9444), .Z(n358) );
  AND U10191 ( .A(n9445), .B(n9446), .Z(n9443) );
  XNOR U10192 ( .A(n9444), .B(n9410), .Z(n9446) );
  XNOR U10193 ( .A(n9447), .B(n9448), .Z(n9410) );
  ANDN U10194 ( .B(n9449), .A(n9450), .Z(n9447) );
  XOR U10195 ( .A(n9448), .B(n9451), .Z(n9449) );
  XOR U10196 ( .A(n9444), .B(n9412), .Z(n9445) );
  XOR U10197 ( .A(n9452), .B(n9453), .Z(n9412) );
  AND U10198 ( .A(n362), .B(n9454), .Z(n9452) );
  XOR U10199 ( .A(n9455), .B(n9453), .Z(n9454) );
  XNOR U10200 ( .A(n9456), .B(n9457), .Z(n9444) );
  NAND U10201 ( .A(n9458), .B(n9459), .Z(n9457) );
  XOR U10202 ( .A(n9460), .B(n9436), .Z(n9459) );
  XOR U10203 ( .A(n9450), .B(n9451), .Z(n9436) );
  XOR U10204 ( .A(n9461), .B(n9462), .Z(n9451) );
  ANDN U10205 ( .B(n9463), .A(n9464), .Z(n9461) );
  XOR U10206 ( .A(n9462), .B(n9465), .Z(n9463) );
  XOR U10207 ( .A(n9466), .B(n9467), .Z(n9450) );
  XOR U10208 ( .A(n9468), .B(n9469), .Z(n9467) );
  ANDN U10209 ( .B(n9470), .A(n9471), .Z(n9468) );
  XOR U10210 ( .A(n9472), .B(n9469), .Z(n9470) );
  IV U10211 ( .A(n9448), .Z(n9466) );
  XOR U10212 ( .A(n9473), .B(n9474), .Z(n9448) );
  ANDN U10213 ( .B(n9475), .A(n9476), .Z(n9473) );
  XOR U10214 ( .A(n9474), .B(n9477), .Z(n9475) );
  IV U10215 ( .A(n9456), .Z(n9460) );
  XOR U10216 ( .A(n9456), .B(n9438), .Z(n9458) );
  XOR U10217 ( .A(n9478), .B(n9479), .Z(n9438) );
  AND U10218 ( .A(n362), .B(n9480), .Z(n9478) );
  XOR U10219 ( .A(n9481), .B(n9479), .Z(n9480) );
  NANDN U10220 ( .A(n9440), .B(n9442), .Z(n9456) );
  XOR U10221 ( .A(n9482), .B(n9483), .Z(n9442) );
  AND U10222 ( .A(n362), .B(n9484), .Z(n9482) );
  XOR U10223 ( .A(n9483), .B(n9485), .Z(n9484) );
  XOR U10224 ( .A(n9486), .B(n9487), .Z(n362) );
  AND U10225 ( .A(n9488), .B(n9489), .Z(n9486) );
  XNOR U10226 ( .A(n9487), .B(n9453), .Z(n9489) );
  XNOR U10227 ( .A(n9490), .B(n9491), .Z(n9453) );
  ANDN U10228 ( .B(n9492), .A(n9493), .Z(n9490) );
  XOR U10229 ( .A(n9491), .B(n9494), .Z(n9492) );
  XOR U10230 ( .A(n9487), .B(n9455), .Z(n9488) );
  XOR U10231 ( .A(n9495), .B(n9496), .Z(n9455) );
  AND U10232 ( .A(n366), .B(n9497), .Z(n9495) );
  XOR U10233 ( .A(n9498), .B(n9496), .Z(n9497) );
  XNOR U10234 ( .A(n9499), .B(n9500), .Z(n9487) );
  NAND U10235 ( .A(n9501), .B(n9502), .Z(n9500) );
  XOR U10236 ( .A(n9503), .B(n9479), .Z(n9502) );
  XOR U10237 ( .A(n9493), .B(n9494), .Z(n9479) );
  XOR U10238 ( .A(n9504), .B(n9505), .Z(n9494) );
  ANDN U10239 ( .B(n9506), .A(n9507), .Z(n9504) );
  XOR U10240 ( .A(n9505), .B(n9508), .Z(n9506) );
  XOR U10241 ( .A(n9509), .B(n9510), .Z(n9493) );
  XOR U10242 ( .A(n9511), .B(n9512), .Z(n9510) );
  ANDN U10243 ( .B(n9513), .A(n9514), .Z(n9511) );
  XOR U10244 ( .A(n9515), .B(n9512), .Z(n9513) );
  IV U10245 ( .A(n9491), .Z(n9509) );
  XOR U10246 ( .A(n9516), .B(n9517), .Z(n9491) );
  ANDN U10247 ( .B(n9518), .A(n9519), .Z(n9516) );
  XOR U10248 ( .A(n9517), .B(n9520), .Z(n9518) );
  IV U10249 ( .A(n9499), .Z(n9503) );
  XOR U10250 ( .A(n9499), .B(n9481), .Z(n9501) );
  XOR U10251 ( .A(n9521), .B(n9522), .Z(n9481) );
  AND U10252 ( .A(n366), .B(n9523), .Z(n9521) );
  XOR U10253 ( .A(n9524), .B(n9522), .Z(n9523) );
  NANDN U10254 ( .A(n9483), .B(n9485), .Z(n9499) );
  XOR U10255 ( .A(n9525), .B(n9526), .Z(n9485) );
  AND U10256 ( .A(n366), .B(n9527), .Z(n9525) );
  XOR U10257 ( .A(n9526), .B(n9528), .Z(n9527) );
  XOR U10258 ( .A(n9529), .B(n9530), .Z(n366) );
  AND U10259 ( .A(n9531), .B(n9532), .Z(n9529) );
  XNOR U10260 ( .A(n9530), .B(n9496), .Z(n9532) );
  XNOR U10261 ( .A(n9533), .B(n9534), .Z(n9496) );
  ANDN U10262 ( .B(n9535), .A(n9536), .Z(n9533) );
  XOR U10263 ( .A(n9534), .B(n9537), .Z(n9535) );
  XOR U10264 ( .A(n9530), .B(n9498), .Z(n9531) );
  XOR U10265 ( .A(n9538), .B(n9539), .Z(n9498) );
  AND U10266 ( .A(n370), .B(n9540), .Z(n9538) );
  XOR U10267 ( .A(n9541), .B(n9539), .Z(n9540) );
  XNOR U10268 ( .A(n9542), .B(n9543), .Z(n9530) );
  NAND U10269 ( .A(n9544), .B(n9545), .Z(n9543) );
  XOR U10270 ( .A(n9546), .B(n9522), .Z(n9545) );
  XOR U10271 ( .A(n9536), .B(n9537), .Z(n9522) );
  XOR U10272 ( .A(n9547), .B(n9548), .Z(n9537) );
  ANDN U10273 ( .B(n9549), .A(n9550), .Z(n9547) );
  XOR U10274 ( .A(n9548), .B(n9551), .Z(n9549) );
  XOR U10275 ( .A(n9552), .B(n9553), .Z(n9536) );
  XOR U10276 ( .A(n9554), .B(n9555), .Z(n9553) );
  ANDN U10277 ( .B(n9556), .A(n9557), .Z(n9554) );
  XOR U10278 ( .A(n9558), .B(n9555), .Z(n9556) );
  IV U10279 ( .A(n9534), .Z(n9552) );
  XOR U10280 ( .A(n9559), .B(n9560), .Z(n9534) );
  ANDN U10281 ( .B(n9561), .A(n9562), .Z(n9559) );
  XOR U10282 ( .A(n9560), .B(n9563), .Z(n9561) );
  IV U10283 ( .A(n9542), .Z(n9546) );
  XOR U10284 ( .A(n9542), .B(n9524), .Z(n9544) );
  XOR U10285 ( .A(n9564), .B(n9565), .Z(n9524) );
  AND U10286 ( .A(n370), .B(n9566), .Z(n9564) );
  XOR U10287 ( .A(n9567), .B(n9565), .Z(n9566) );
  NANDN U10288 ( .A(n9526), .B(n9528), .Z(n9542) );
  XOR U10289 ( .A(n9568), .B(n9569), .Z(n9528) );
  AND U10290 ( .A(n370), .B(n9570), .Z(n9568) );
  XOR U10291 ( .A(n9569), .B(n9571), .Z(n9570) );
  XOR U10292 ( .A(n9572), .B(n9573), .Z(n370) );
  AND U10293 ( .A(n9574), .B(n9575), .Z(n9572) );
  XNOR U10294 ( .A(n9573), .B(n9539), .Z(n9575) );
  XNOR U10295 ( .A(n9576), .B(n9577), .Z(n9539) );
  ANDN U10296 ( .B(n9578), .A(n9579), .Z(n9576) );
  XOR U10297 ( .A(n9577), .B(n9580), .Z(n9578) );
  XOR U10298 ( .A(n9573), .B(n9541), .Z(n9574) );
  XOR U10299 ( .A(n9581), .B(n9582), .Z(n9541) );
  AND U10300 ( .A(n374), .B(n9583), .Z(n9581) );
  XOR U10301 ( .A(n9584), .B(n9582), .Z(n9583) );
  XNOR U10302 ( .A(n9585), .B(n9586), .Z(n9573) );
  NAND U10303 ( .A(n9587), .B(n9588), .Z(n9586) );
  XOR U10304 ( .A(n9589), .B(n9565), .Z(n9588) );
  XOR U10305 ( .A(n9579), .B(n9580), .Z(n9565) );
  XOR U10306 ( .A(n9590), .B(n9591), .Z(n9580) );
  ANDN U10307 ( .B(n9592), .A(n9593), .Z(n9590) );
  XOR U10308 ( .A(n9591), .B(n9594), .Z(n9592) );
  XOR U10309 ( .A(n9595), .B(n9596), .Z(n9579) );
  XOR U10310 ( .A(n9597), .B(n9598), .Z(n9596) );
  ANDN U10311 ( .B(n9599), .A(n9600), .Z(n9597) );
  XOR U10312 ( .A(n9601), .B(n9598), .Z(n9599) );
  IV U10313 ( .A(n9577), .Z(n9595) );
  XOR U10314 ( .A(n9602), .B(n9603), .Z(n9577) );
  ANDN U10315 ( .B(n9604), .A(n9605), .Z(n9602) );
  XOR U10316 ( .A(n9603), .B(n9606), .Z(n9604) );
  IV U10317 ( .A(n9585), .Z(n9589) );
  XOR U10318 ( .A(n9585), .B(n9567), .Z(n9587) );
  XOR U10319 ( .A(n9607), .B(n9608), .Z(n9567) );
  AND U10320 ( .A(n374), .B(n9609), .Z(n9607) );
  XOR U10321 ( .A(n9610), .B(n9608), .Z(n9609) );
  NANDN U10322 ( .A(n9569), .B(n9571), .Z(n9585) );
  XOR U10323 ( .A(n9611), .B(n9612), .Z(n9571) );
  AND U10324 ( .A(n374), .B(n9613), .Z(n9611) );
  XOR U10325 ( .A(n9612), .B(n9614), .Z(n9613) );
  XOR U10326 ( .A(n9615), .B(n9616), .Z(n374) );
  AND U10327 ( .A(n9617), .B(n9618), .Z(n9615) );
  XNOR U10328 ( .A(n9616), .B(n9582), .Z(n9618) );
  XNOR U10329 ( .A(n9619), .B(n9620), .Z(n9582) );
  ANDN U10330 ( .B(n9621), .A(n9622), .Z(n9619) );
  XOR U10331 ( .A(n9620), .B(n9623), .Z(n9621) );
  XOR U10332 ( .A(n9616), .B(n9584), .Z(n9617) );
  XOR U10333 ( .A(n9624), .B(n9625), .Z(n9584) );
  AND U10334 ( .A(n378), .B(n9626), .Z(n9624) );
  XOR U10335 ( .A(n9627), .B(n9625), .Z(n9626) );
  XNOR U10336 ( .A(n9628), .B(n9629), .Z(n9616) );
  NAND U10337 ( .A(n9630), .B(n9631), .Z(n9629) );
  XOR U10338 ( .A(n9632), .B(n9608), .Z(n9631) );
  XOR U10339 ( .A(n9622), .B(n9623), .Z(n9608) );
  XOR U10340 ( .A(n9633), .B(n9634), .Z(n9623) );
  ANDN U10341 ( .B(n9635), .A(n9636), .Z(n9633) );
  XOR U10342 ( .A(n9634), .B(n9637), .Z(n9635) );
  XOR U10343 ( .A(n9638), .B(n9639), .Z(n9622) );
  XOR U10344 ( .A(n9640), .B(n9641), .Z(n9639) );
  ANDN U10345 ( .B(n9642), .A(n9643), .Z(n9640) );
  XOR U10346 ( .A(n9644), .B(n9641), .Z(n9642) );
  IV U10347 ( .A(n9620), .Z(n9638) );
  XOR U10348 ( .A(n9645), .B(n9646), .Z(n9620) );
  ANDN U10349 ( .B(n9647), .A(n9648), .Z(n9645) );
  XOR U10350 ( .A(n9646), .B(n9649), .Z(n9647) );
  IV U10351 ( .A(n9628), .Z(n9632) );
  XOR U10352 ( .A(n9628), .B(n9610), .Z(n9630) );
  XOR U10353 ( .A(n9650), .B(n9651), .Z(n9610) );
  AND U10354 ( .A(n378), .B(n9652), .Z(n9650) );
  XOR U10355 ( .A(n9653), .B(n9651), .Z(n9652) );
  NANDN U10356 ( .A(n9612), .B(n9614), .Z(n9628) );
  XOR U10357 ( .A(n9654), .B(n9655), .Z(n9614) );
  AND U10358 ( .A(n378), .B(n9656), .Z(n9654) );
  XOR U10359 ( .A(n9655), .B(n9657), .Z(n9656) );
  XOR U10360 ( .A(n9658), .B(n9659), .Z(n378) );
  AND U10361 ( .A(n9660), .B(n9661), .Z(n9658) );
  XNOR U10362 ( .A(n9659), .B(n9625), .Z(n9661) );
  XNOR U10363 ( .A(n9662), .B(n9663), .Z(n9625) );
  ANDN U10364 ( .B(n9664), .A(n9665), .Z(n9662) );
  XOR U10365 ( .A(n9663), .B(n9666), .Z(n9664) );
  XOR U10366 ( .A(n9659), .B(n9627), .Z(n9660) );
  XOR U10367 ( .A(n9667), .B(n9668), .Z(n9627) );
  AND U10368 ( .A(n382), .B(n9669), .Z(n9667) );
  XOR U10369 ( .A(n9670), .B(n9668), .Z(n9669) );
  XNOR U10370 ( .A(n9671), .B(n9672), .Z(n9659) );
  NAND U10371 ( .A(n9673), .B(n9674), .Z(n9672) );
  XOR U10372 ( .A(n9675), .B(n9651), .Z(n9674) );
  XOR U10373 ( .A(n9665), .B(n9666), .Z(n9651) );
  XOR U10374 ( .A(n9676), .B(n9677), .Z(n9666) );
  ANDN U10375 ( .B(n9678), .A(n9679), .Z(n9676) );
  XOR U10376 ( .A(n9677), .B(n9680), .Z(n9678) );
  XOR U10377 ( .A(n9681), .B(n9682), .Z(n9665) );
  XOR U10378 ( .A(n9683), .B(n9684), .Z(n9682) );
  ANDN U10379 ( .B(n9685), .A(n9686), .Z(n9683) );
  XOR U10380 ( .A(n9687), .B(n9684), .Z(n9685) );
  IV U10381 ( .A(n9663), .Z(n9681) );
  XOR U10382 ( .A(n9688), .B(n9689), .Z(n9663) );
  ANDN U10383 ( .B(n9690), .A(n9691), .Z(n9688) );
  XOR U10384 ( .A(n9689), .B(n9692), .Z(n9690) );
  IV U10385 ( .A(n9671), .Z(n9675) );
  XOR U10386 ( .A(n9671), .B(n9653), .Z(n9673) );
  XOR U10387 ( .A(n9693), .B(n9694), .Z(n9653) );
  AND U10388 ( .A(n382), .B(n9695), .Z(n9693) );
  XOR U10389 ( .A(n9696), .B(n9694), .Z(n9695) );
  NANDN U10390 ( .A(n9655), .B(n9657), .Z(n9671) );
  XOR U10391 ( .A(n9697), .B(n9698), .Z(n9657) );
  AND U10392 ( .A(n382), .B(n9699), .Z(n9697) );
  XOR U10393 ( .A(n9698), .B(n9700), .Z(n9699) );
  XOR U10394 ( .A(n9701), .B(n9702), .Z(n382) );
  AND U10395 ( .A(n9703), .B(n9704), .Z(n9701) );
  XNOR U10396 ( .A(n9702), .B(n9668), .Z(n9704) );
  XNOR U10397 ( .A(n9705), .B(n9706), .Z(n9668) );
  ANDN U10398 ( .B(n9707), .A(n9708), .Z(n9705) );
  XOR U10399 ( .A(n9706), .B(n9709), .Z(n9707) );
  XOR U10400 ( .A(n9702), .B(n9670), .Z(n9703) );
  XOR U10401 ( .A(n9710), .B(n9711), .Z(n9670) );
  AND U10402 ( .A(n386), .B(n9712), .Z(n9710) );
  XOR U10403 ( .A(n9713), .B(n9711), .Z(n9712) );
  XNOR U10404 ( .A(n9714), .B(n9715), .Z(n9702) );
  NAND U10405 ( .A(n9716), .B(n9717), .Z(n9715) );
  XOR U10406 ( .A(n9718), .B(n9694), .Z(n9717) );
  XOR U10407 ( .A(n9708), .B(n9709), .Z(n9694) );
  XOR U10408 ( .A(n9719), .B(n9720), .Z(n9709) );
  ANDN U10409 ( .B(n9721), .A(n9722), .Z(n9719) );
  XOR U10410 ( .A(n9720), .B(n9723), .Z(n9721) );
  XOR U10411 ( .A(n9724), .B(n9725), .Z(n9708) );
  XOR U10412 ( .A(n9726), .B(n9727), .Z(n9725) );
  ANDN U10413 ( .B(n9728), .A(n9729), .Z(n9726) );
  XOR U10414 ( .A(n9730), .B(n9727), .Z(n9728) );
  IV U10415 ( .A(n9706), .Z(n9724) );
  XOR U10416 ( .A(n9731), .B(n9732), .Z(n9706) );
  ANDN U10417 ( .B(n9733), .A(n9734), .Z(n9731) );
  XOR U10418 ( .A(n9732), .B(n9735), .Z(n9733) );
  IV U10419 ( .A(n9714), .Z(n9718) );
  XOR U10420 ( .A(n9714), .B(n9696), .Z(n9716) );
  XOR U10421 ( .A(n9736), .B(n9737), .Z(n9696) );
  AND U10422 ( .A(n386), .B(n9738), .Z(n9736) );
  XOR U10423 ( .A(n9739), .B(n9737), .Z(n9738) );
  NANDN U10424 ( .A(n9698), .B(n9700), .Z(n9714) );
  XOR U10425 ( .A(n9740), .B(n9741), .Z(n9700) );
  AND U10426 ( .A(n386), .B(n9742), .Z(n9740) );
  XOR U10427 ( .A(n9741), .B(n9743), .Z(n9742) );
  XOR U10428 ( .A(n9744), .B(n9745), .Z(n386) );
  AND U10429 ( .A(n9746), .B(n9747), .Z(n9744) );
  XNOR U10430 ( .A(n9745), .B(n9711), .Z(n9747) );
  XNOR U10431 ( .A(n9748), .B(n9749), .Z(n9711) );
  ANDN U10432 ( .B(n9750), .A(n9751), .Z(n9748) );
  XOR U10433 ( .A(n9749), .B(n9752), .Z(n9750) );
  XOR U10434 ( .A(n9745), .B(n9713), .Z(n9746) );
  XOR U10435 ( .A(n9753), .B(n9754), .Z(n9713) );
  AND U10436 ( .A(n390), .B(n9755), .Z(n9753) );
  XOR U10437 ( .A(n9756), .B(n9754), .Z(n9755) );
  XNOR U10438 ( .A(n9757), .B(n9758), .Z(n9745) );
  NAND U10439 ( .A(n9759), .B(n9760), .Z(n9758) );
  XOR U10440 ( .A(n9761), .B(n9737), .Z(n9760) );
  XOR U10441 ( .A(n9751), .B(n9752), .Z(n9737) );
  XOR U10442 ( .A(n9762), .B(n9763), .Z(n9752) );
  ANDN U10443 ( .B(n9764), .A(n9765), .Z(n9762) );
  XOR U10444 ( .A(n9763), .B(n9766), .Z(n9764) );
  XOR U10445 ( .A(n9767), .B(n9768), .Z(n9751) );
  XOR U10446 ( .A(n9769), .B(n9770), .Z(n9768) );
  ANDN U10447 ( .B(n9771), .A(n9772), .Z(n9769) );
  XOR U10448 ( .A(n9773), .B(n9770), .Z(n9771) );
  IV U10449 ( .A(n9749), .Z(n9767) );
  XOR U10450 ( .A(n9774), .B(n9775), .Z(n9749) );
  ANDN U10451 ( .B(n9776), .A(n9777), .Z(n9774) );
  XOR U10452 ( .A(n9775), .B(n9778), .Z(n9776) );
  IV U10453 ( .A(n9757), .Z(n9761) );
  XOR U10454 ( .A(n9757), .B(n9739), .Z(n9759) );
  XOR U10455 ( .A(n9779), .B(n9780), .Z(n9739) );
  AND U10456 ( .A(n390), .B(n9781), .Z(n9779) );
  XOR U10457 ( .A(n9782), .B(n9780), .Z(n9781) );
  NANDN U10458 ( .A(n9741), .B(n9743), .Z(n9757) );
  XOR U10459 ( .A(n9783), .B(n9784), .Z(n9743) );
  AND U10460 ( .A(n390), .B(n9785), .Z(n9783) );
  XOR U10461 ( .A(n9784), .B(n9786), .Z(n9785) );
  XOR U10462 ( .A(n9787), .B(n9788), .Z(n390) );
  AND U10463 ( .A(n9789), .B(n9790), .Z(n9787) );
  XNOR U10464 ( .A(n9788), .B(n9754), .Z(n9790) );
  XNOR U10465 ( .A(n9791), .B(n9792), .Z(n9754) );
  ANDN U10466 ( .B(n9793), .A(n9794), .Z(n9791) );
  XOR U10467 ( .A(n9792), .B(n9795), .Z(n9793) );
  XOR U10468 ( .A(n9788), .B(n9756), .Z(n9789) );
  XOR U10469 ( .A(n9796), .B(n9797), .Z(n9756) );
  AND U10470 ( .A(n394), .B(n9798), .Z(n9796) );
  XOR U10471 ( .A(n9799), .B(n9797), .Z(n9798) );
  XNOR U10472 ( .A(n9800), .B(n9801), .Z(n9788) );
  NAND U10473 ( .A(n9802), .B(n9803), .Z(n9801) );
  XOR U10474 ( .A(n9804), .B(n9780), .Z(n9803) );
  XOR U10475 ( .A(n9794), .B(n9795), .Z(n9780) );
  XOR U10476 ( .A(n9805), .B(n9806), .Z(n9795) );
  ANDN U10477 ( .B(n9807), .A(n9808), .Z(n9805) );
  XOR U10478 ( .A(n9806), .B(n9809), .Z(n9807) );
  XOR U10479 ( .A(n9810), .B(n9811), .Z(n9794) );
  XOR U10480 ( .A(n9812), .B(n9813), .Z(n9811) );
  ANDN U10481 ( .B(n9814), .A(n9815), .Z(n9812) );
  XOR U10482 ( .A(n9816), .B(n9813), .Z(n9814) );
  IV U10483 ( .A(n9792), .Z(n9810) );
  XOR U10484 ( .A(n9817), .B(n9818), .Z(n9792) );
  ANDN U10485 ( .B(n9819), .A(n9820), .Z(n9817) );
  XOR U10486 ( .A(n9818), .B(n9821), .Z(n9819) );
  IV U10487 ( .A(n9800), .Z(n9804) );
  XOR U10488 ( .A(n9800), .B(n9782), .Z(n9802) );
  XOR U10489 ( .A(n9822), .B(n9823), .Z(n9782) );
  AND U10490 ( .A(n394), .B(n9824), .Z(n9822) );
  XOR U10491 ( .A(n9825), .B(n9823), .Z(n9824) );
  NANDN U10492 ( .A(n9784), .B(n9786), .Z(n9800) );
  XOR U10493 ( .A(n9826), .B(n9827), .Z(n9786) );
  AND U10494 ( .A(n394), .B(n9828), .Z(n9826) );
  XOR U10495 ( .A(n9827), .B(n9829), .Z(n9828) );
  XOR U10496 ( .A(n9830), .B(n9831), .Z(n394) );
  AND U10497 ( .A(n9832), .B(n9833), .Z(n9830) );
  XNOR U10498 ( .A(n9831), .B(n9797), .Z(n9833) );
  XNOR U10499 ( .A(n9834), .B(n9835), .Z(n9797) );
  ANDN U10500 ( .B(n9836), .A(n9837), .Z(n9834) );
  XOR U10501 ( .A(n9835), .B(n9838), .Z(n9836) );
  XOR U10502 ( .A(n9831), .B(n9799), .Z(n9832) );
  XOR U10503 ( .A(n9839), .B(n9840), .Z(n9799) );
  AND U10504 ( .A(n398), .B(n9841), .Z(n9839) );
  XOR U10505 ( .A(n9842), .B(n9840), .Z(n9841) );
  XNOR U10506 ( .A(n9843), .B(n9844), .Z(n9831) );
  NAND U10507 ( .A(n9845), .B(n9846), .Z(n9844) );
  XOR U10508 ( .A(n9847), .B(n9823), .Z(n9846) );
  XOR U10509 ( .A(n9837), .B(n9838), .Z(n9823) );
  XOR U10510 ( .A(n9848), .B(n9849), .Z(n9838) );
  ANDN U10511 ( .B(n9850), .A(n9851), .Z(n9848) );
  XOR U10512 ( .A(n9849), .B(n9852), .Z(n9850) );
  XOR U10513 ( .A(n9853), .B(n9854), .Z(n9837) );
  XOR U10514 ( .A(n9855), .B(n9856), .Z(n9854) );
  ANDN U10515 ( .B(n9857), .A(n9858), .Z(n9855) );
  XOR U10516 ( .A(n9859), .B(n9856), .Z(n9857) );
  IV U10517 ( .A(n9835), .Z(n9853) );
  XOR U10518 ( .A(n9860), .B(n9861), .Z(n9835) );
  ANDN U10519 ( .B(n9862), .A(n9863), .Z(n9860) );
  XOR U10520 ( .A(n9861), .B(n9864), .Z(n9862) );
  IV U10521 ( .A(n9843), .Z(n9847) );
  XOR U10522 ( .A(n9843), .B(n9825), .Z(n9845) );
  XOR U10523 ( .A(n9865), .B(n9866), .Z(n9825) );
  AND U10524 ( .A(n398), .B(n9867), .Z(n9865) );
  XOR U10525 ( .A(n9868), .B(n9866), .Z(n9867) );
  NANDN U10526 ( .A(n9827), .B(n9829), .Z(n9843) );
  XOR U10527 ( .A(n9869), .B(n9870), .Z(n9829) );
  AND U10528 ( .A(n398), .B(n9871), .Z(n9869) );
  XOR U10529 ( .A(n9870), .B(n9872), .Z(n9871) );
  XOR U10530 ( .A(n9873), .B(n9874), .Z(n398) );
  AND U10531 ( .A(n9875), .B(n9876), .Z(n9873) );
  XNOR U10532 ( .A(n9874), .B(n9840), .Z(n9876) );
  XNOR U10533 ( .A(n9877), .B(n9878), .Z(n9840) );
  ANDN U10534 ( .B(n9879), .A(n9880), .Z(n9877) );
  XOR U10535 ( .A(n9878), .B(n9881), .Z(n9879) );
  XOR U10536 ( .A(n9874), .B(n9842), .Z(n9875) );
  XOR U10537 ( .A(n9882), .B(n9883), .Z(n9842) );
  AND U10538 ( .A(n402), .B(n9884), .Z(n9882) );
  XOR U10539 ( .A(n9885), .B(n9883), .Z(n9884) );
  XNOR U10540 ( .A(n9886), .B(n9887), .Z(n9874) );
  NAND U10541 ( .A(n9888), .B(n9889), .Z(n9887) );
  XOR U10542 ( .A(n9890), .B(n9866), .Z(n9889) );
  XOR U10543 ( .A(n9880), .B(n9881), .Z(n9866) );
  XOR U10544 ( .A(n9891), .B(n9892), .Z(n9881) );
  ANDN U10545 ( .B(n9893), .A(n9894), .Z(n9891) );
  XOR U10546 ( .A(n9892), .B(n9895), .Z(n9893) );
  XOR U10547 ( .A(n9896), .B(n9897), .Z(n9880) );
  XOR U10548 ( .A(n9898), .B(n9899), .Z(n9897) );
  ANDN U10549 ( .B(n9900), .A(n9901), .Z(n9898) );
  XOR U10550 ( .A(n9902), .B(n9899), .Z(n9900) );
  IV U10551 ( .A(n9878), .Z(n9896) );
  XOR U10552 ( .A(n9903), .B(n9904), .Z(n9878) );
  ANDN U10553 ( .B(n9905), .A(n9906), .Z(n9903) );
  XOR U10554 ( .A(n9904), .B(n9907), .Z(n9905) );
  IV U10555 ( .A(n9886), .Z(n9890) );
  XOR U10556 ( .A(n9886), .B(n9868), .Z(n9888) );
  XOR U10557 ( .A(n9908), .B(n9909), .Z(n9868) );
  AND U10558 ( .A(n402), .B(n9910), .Z(n9908) );
  XOR U10559 ( .A(n9911), .B(n9909), .Z(n9910) );
  NANDN U10560 ( .A(n9870), .B(n9872), .Z(n9886) );
  XOR U10561 ( .A(n9912), .B(n9913), .Z(n9872) );
  AND U10562 ( .A(n402), .B(n9914), .Z(n9912) );
  XOR U10563 ( .A(n9913), .B(n9915), .Z(n9914) );
  XOR U10564 ( .A(n9916), .B(n9917), .Z(n402) );
  AND U10565 ( .A(n9918), .B(n9919), .Z(n9916) );
  XNOR U10566 ( .A(n9917), .B(n9883), .Z(n9919) );
  XNOR U10567 ( .A(n9920), .B(n9921), .Z(n9883) );
  ANDN U10568 ( .B(n9922), .A(n9923), .Z(n9920) );
  XOR U10569 ( .A(n9921), .B(n9924), .Z(n9922) );
  XOR U10570 ( .A(n9917), .B(n9885), .Z(n9918) );
  XOR U10571 ( .A(n9925), .B(n9926), .Z(n9885) );
  AND U10572 ( .A(n406), .B(n9927), .Z(n9925) );
  XOR U10573 ( .A(n9928), .B(n9926), .Z(n9927) );
  XNOR U10574 ( .A(n9929), .B(n9930), .Z(n9917) );
  NAND U10575 ( .A(n9931), .B(n9932), .Z(n9930) );
  XOR U10576 ( .A(n9933), .B(n9909), .Z(n9932) );
  XOR U10577 ( .A(n9923), .B(n9924), .Z(n9909) );
  XOR U10578 ( .A(n9934), .B(n9935), .Z(n9924) );
  ANDN U10579 ( .B(n9936), .A(n9937), .Z(n9934) );
  XOR U10580 ( .A(n9935), .B(n9938), .Z(n9936) );
  XOR U10581 ( .A(n9939), .B(n9940), .Z(n9923) );
  XOR U10582 ( .A(n9941), .B(n9942), .Z(n9940) );
  ANDN U10583 ( .B(n9943), .A(n9944), .Z(n9941) );
  XOR U10584 ( .A(n9945), .B(n9942), .Z(n9943) );
  IV U10585 ( .A(n9921), .Z(n9939) );
  XOR U10586 ( .A(n9946), .B(n9947), .Z(n9921) );
  ANDN U10587 ( .B(n9948), .A(n9949), .Z(n9946) );
  XOR U10588 ( .A(n9947), .B(n9950), .Z(n9948) );
  IV U10589 ( .A(n9929), .Z(n9933) );
  XOR U10590 ( .A(n9929), .B(n9911), .Z(n9931) );
  XOR U10591 ( .A(n9951), .B(n9952), .Z(n9911) );
  AND U10592 ( .A(n406), .B(n9953), .Z(n9951) );
  XOR U10593 ( .A(n9954), .B(n9952), .Z(n9953) );
  NANDN U10594 ( .A(n9913), .B(n9915), .Z(n9929) );
  XOR U10595 ( .A(n9955), .B(n9956), .Z(n9915) );
  AND U10596 ( .A(n406), .B(n9957), .Z(n9955) );
  XOR U10597 ( .A(n9956), .B(n9958), .Z(n9957) );
  XOR U10598 ( .A(n9959), .B(n9960), .Z(n406) );
  AND U10599 ( .A(n9961), .B(n9962), .Z(n9959) );
  XNOR U10600 ( .A(n9960), .B(n9926), .Z(n9962) );
  XNOR U10601 ( .A(n9963), .B(n9964), .Z(n9926) );
  ANDN U10602 ( .B(n9965), .A(n9966), .Z(n9963) );
  XOR U10603 ( .A(n9964), .B(n9967), .Z(n9965) );
  XOR U10604 ( .A(n9960), .B(n9928), .Z(n9961) );
  XOR U10605 ( .A(n9968), .B(n9969), .Z(n9928) );
  AND U10606 ( .A(n410), .B(n9970), .Z(n9968) );
  XOR U10607 ( .A(n9971), .B(n9969), .Z(n9970) );
  XNOR U10608 ( .A(n9972), .B(n9973), .Z(n9960) );
  NAND U10609 ( .A(n9974), .B(n9975), .Z(n9973) );
  XOR U10610 ( .A(n9976), .B(n9952), .Z(n9975) );
  XOR U10611 ( .A(n9966), .B(n9967), .Z(n9952) );
  XOR U10612 ( .A(n9977), .B(n9978), .Z(n9967) );
  ANDN U10613 ( .B(n9979), .A(n9980), .Z(n9977) );
  XOR U10614 ( .A(n9978), .B(n9981), .Z(n9979) );
  XOR U10615 ( .A(n9982), .B(n9983), .Z(n9966) );
  XOR U10616 ( .A(n9984), .B(n9985), .Z(n9983) );
  ANDN U10617 ( .B(n9986), .A(n9987), .Z(n9984) );
  XOR U10618 ( .A(n9988), .B(n9985), .Z(n9986) );
  IV U10619 ( .A(n9964), .Z(n9982) );
  XOR U10620 ( .A(n9989), .B(n9990), .Z(n9964) );
  ANDN U10621 ( .B(n9991), .A(n9992), .Z(n9989) );
  XOR U10622 ( .A(n9990), .B(n9993), .Z(n9991) );
  IV U10623 ( .A(n9972), .Z(n9976) );
  XOR U10624 ( .A(n9972), .B(n9954), .Z(n9974) );
  XOR U10625 ( .A(n9994), .B(n9995), .Z(n9954) );
  AND U10626 ( .A(n410), .B(n9996), .Z(n9994) );
  XOR U10627 ( .A(n9997), .B(n9995), .Z(n9996) );
  NANDN U10628 ( .A(n9956), .B(n9958), .Z(n9972) );
  XOR U10629 ( .A(n9998), .B(n9999), .Z(n9958) );
  AND U10630 ( .A(n410), .B(n10000), .Z(n9998) );
  XOR U10631 ( .A(n9999), .B(n10001), .Z(n10000) );
  XOR U10632 ( .A(n10002), .B(n10003), .Z(n410) );
  AND U10633 ( .A(n10004), .B(n10005), .Z(n10002) );
  XNOR U10634 ( .A(n10003), .B(n9969), .Z(n10005) );
  XNOR U10635 ( .A(n10006), .B(n10007), .Z(n9969) );
  ANDN U10636 ( .B(n10008), .A(n10009), .Z(n10006) );
  XOR U10637 ( .A(n10007), .B(n10010), .Z(n10008) );
  XOR U10638 ( .A(n10003), .B(n9971), .Z(n10004) );
  XOR U10639 ( .A(n10011), .B(n10012), .Z(n9971) );
  AND U10640 ( .A(n414), .B(n10013), .Z(n10011) );
  XOR U10641 ( .A(n10014), .B(n10012), .Z(n10013) );
  XNOR U10642 ( .A(n10015), .B(n10016), .Z(n10003) );
  NAND U10643 ( .A(n10017), .B(n10018), .Z(n10016) );
  XOR U10644 ( .A(n10019), .B(n9995), .Z(n10018) );
  XOR U10645 ( .A(n10009), .B(n10010), .Z(n9995) );
  XOR U10646 ( .A(n10020), .B(n10021), .Z(n10010) );
  ANDN U10647 ( .B(n10022), .A(n10023), .Z(n10020) );
  XOR U10648 ( .A(n10021), .B(n10024), .Z(n10022) );
  XOR U10649 ( .A(n10025), .B(n10026), .Z(n10009) );
  XOR U10650 ( .A(n10027), .B(n10028), .Z(n10026) );
  ANDN U10651 ( .B(n10029), .A(n10030), .Z(n10027) );
  XOR U10652 ( .A(n10031), .B(n10028), .Z(n10029) );
  IV U10653 ( .A(n10007), .Z(n10025) );
  XOR U10654 ( .A(n10032), .B(n10033), .Z(n10007) );
  ANDN U10655 ( .B(n10034), .A(n10035), .Z(n10032) );
  XOR U10656 ( .A(n10033), .B(n10036), .Z(n10034) );
  IV U10657 ( .A(n10015), .Z(n10019) );
  XOR U10658 ( .A(n10015), .B(n9997), .Z(n10017) );
  XOR U10659 ( .A(n10037), .B(n10038), .Z(n9997) );
  AND U10660 ( .A(n414), .B(n10039), .Z(n10037) );
  XOR U10661 ( .A(n10040), .B(n10038), .Z(n10039) );
  NANDN U10662 ( .A(n9999), .B(n10001), .Z(n10015) );
  XOR U10663 ( .A(n10041), .B(n10042), .Z(n10001) );
  AND U10664 ( .A(n414), .B(n10043), .Z(n10041) );
  XOR U10665 ( .A(n10042), .B(n10044), .Z(n10043) );
  XOR U10666 ( .A(n10045), .B(n10046), .Z(n414) );
  AND U10667 ( .A(n10047), .B(n10048), .Z(n10045) );
  XNOR U10668 ( .A(n10046), .B(n10012), .Z(n10048) );
  XNOR U10669 ( .A(n10049), .B(n10050), .Z(n10012) );
  ANDN U10670 ( .B(n10051), .A(n10052), .Z(n10049) );
  XOR U10671 ( .A(n10050), .B(n10053), .Z(n10051) );
  XOR U10672 ( .A(n10046), .B(n10014), .Z(n10047) );
  XOR U10673 ( .A(n10054), .B(n10055), .Z(n10014) );
  AND U10674 ( .A(n418), .B(n10056), .Z(n10054) );
  XOR U10675 ( .A(n10057), .B(n10055), .Z(n10056) );
  XNOR U10676 ( .A(n10058), .B(n10059), .Z(n10046) );
  NAND U10677 ( .A(n10060), .B(n10061), .Z(n10059) );
  XOR U10678 ( .A(n10062), .B(n10038), .Z(n10061) );
  XOR U10679 ( .A(n10052), .B(n10053), .Z(n10038) );
  XOR U10680 ( .A(n10063), .B(n10064), .Z(n10053) );
  ANDN U10681 ( .B(n10065), .A(n10066), .Z(n10063) );
  XOR U10682 ( .A(n10064), .B(n10067), .Z(n10065) );
  XOR U10683 ( .A(n10068), .B(n10069), .Z(n10052) );
  XOR U10684 ( .A(n10070), .B(n10071), .Z(n10069) );
  ANDN U10685 ( .B(n10072), .A(n10073), .Z(n10070) );
  XOR U10686 ( .A(n10074), .B(n10071), .Z(n10072) );
  IV U10687 ( .A(n10050), .Z(n10068) );
  XOR U10688 ( .A(n10075), .B(n10076), .Z(n10050) );
  ANDN U10689 ( .B(n10077), .A(n10078), .Z(n10075) );
  XOR U10690 ( .A(n10076), .B(n10079), .Z(n10077) );
  IV U10691 ( .A(n10058), .Z(n10062) );
  XOR U10692 ( .A(n10058), .B(n10040), .Z(n10060) );
  XOR U10693 ( .A(n10080), .B(n10081), .Z(n10040) );
  AND U10694 ( .A(n418), .B(n10082), .Z(n10080) );
  XOR U10695 ( .A(n10083), .B(n10081), .Z(n10082) );
  NANDN U10696 ( .A(n10042), .B(n10044), .Z(n10058) );
  XOR U10697 ( .A(n10084), .B(n10085), .Z(n10044) );
  AND U10698 ( .A(n418), .B(n10086), .Z(n10084) );
  XOR U10699 ( .A(n10085), .B(n10087), .Z(n10086) );
  XOR U10700 ( .A(n10088), .B(n10089), .Z(n418) );
  AND U10701 ( .A(n10090), .B(n10091), .Z(n10088) );
  XNOR U10702 ( .A(n10089), .B(n10055), .Z(n10091) );
  XNOR U10703 ( .A(n10092), .B(n10093), .Z(n10055) );
  ANDN U10704 ( .B(n10094), .A(n10095), .Z(n10092) );
  XOR U10705 ( .A(n10093), .B(n10096), .Z(n10094) );
  XOR U10706 ( .A(n10089), .B(n10057), .Z(n10090) );
  XOR U10707 ( .A(n10097), .B(n10098), .Z(n10057) );
  AND U10708 ( .A(n422), .B(n10099), .Z(n10097) );
  XOR U10709 ( .A(n10100), .B(n10098), .Z(n10099) );
  XNOR U10710 ( .A(n10101), .B(n10102), .Z(n10089) );
  NAND U10711 ( .A(n10103), .B(n10104), .Z(n10102) );
  XOR U10712 ( .A(n10105), .B(n10081), .Z(n10104) );
  XOR U10713 ( .A(n10095), .B(n10096), .Z(n10081) );
  XOR U10714 ( .A(n10106), .B(n10107), .Z(n10096) );
  ANDN U10715 ( .B(n10108), .A(n10109), .Z(n10106) );
  XOR U10716 ( .A(n10107), .B(n10110), .Z(n10108) );
  XOR U10717 ( .A(n10111), .B(n10112), .Z(n10095) );
  XOR U10718 ( .A(n10113), .B(n10114), .Z(n10112) );
  ANDN U10719 ( .B(n10115), .A(n10116), .Z(n10113) );
  XOR U10720 ( .A(n10117), .B(n10114), .Z(n10115) );
  IV U10721 ( .A(n10093), .Z(n10111) );
  XOR U10722 ( .A(n10118), .B(n10119), .Z(n10093) );
  ANDN U10723 ( .B(n10120), .A(n10121), .Z(n10118) );
  XOR U10724 ( .A(n10119), .B(n10122), .Z(n10120) );
  IV U10725 ( .A(n10101), .Z(n10105) );
  XOR U10726 ( .A(n10101), .B(n10083), .Z(n10103) );
  XOR U10727 ( .A(n10123), .B(n10124), .Z(n10083) );
  AND U10728 ( .A(n422), .B(n10125), .Z(n10123) );
  XOR U10729 ( .A(n10126), .B(n10124), .Z(n10125) );
  NANDN U10730 ( .A(n10085), .B(n10087), .Z(n10101) );
  XOR U10731 ( .A(n10127), .B(n10128), .Z(n10087) );
  AND U10732 ( .A(n422), .B(n10129), .Z(n10127) );
  XOR U10733 ( .A(n10128), .B(n10130), .Z(n10129) );
  XOR U10734 ( .A(n10131), .B(n10132), .Z(n422) );
  AND U10735 ( .A(n10133), .B(n10134), .Z(n10131) );
  XNOR U10736 ( .A(n10132), .B(n10098), .Z(n10134) );
  XNOR U10737 ( .A(n10135), .B(n10136), .Z(n10098) );
  ANDN U10738 ( .B(n10137), .A(n10138), .Z(n10135) );
  XOR U10739 ( .A(n10136), .B(n10139), .Z(n10137) );
  XOR U10740 ( .A(n10132), .B(n10100), .Z(n10133) );
  XOR U10741 ( .A(n10140), .B(n10141), .Z(n10100) );
  AND U10742 ( .A(n426), .B(n10142), .Z(n10140) );
  XOR U10743 ( .A(n10143), .B(n10141), .Z(n10142) );
  XNOR U10744 ( .A(n10144), .B(n10145), .Z(n10132) );
  NAND U10745 ( .A(n10146), .B(n10147), .Z(n10145) );
  XOR U10746 ( .A(n10148), .B(n10124), .Z(n10147) );
  XOR U10747 ( .A(n10138), .B(n10139), .Z(n10124) );
  XOR U10748 ( .A(n10149), .B(n10150), .Z(n10139) );
  ANDN U10749 ( .B(n10151), .A(n10152), .Z(n10149) );
  XOR U10750 ( .A(n10150), .B(n10153), .Z(n10151) );
  XOR U10751 ( .A(n10154), .B(n10155), .Z(n10138) );
  XOR U10752 ( .A(n10156), .B(n10157), .Z(n10155) );
  ANDN U10753 ( .B(n10158), .A(n10159), .Z(n10156) );
  XOR U10754 ( .A(n10160), .B(n10157), .Z(n10158) );
  IV U10755 ( .A(n10136), .Z(n10154) );
  XOR U10756 ( .A(n10161), .B(n10162), .Z(n10136) );
  ANDN U10757 ( .B(n10163), .A(n10164), .Z(n10161) );
  XOR U10758 ( .A(n10162), .B(n10165), .Z(n10163) );
  IV U10759 ( .A(n10144), .Z(n10148) );
  XOR U10760 ( .A(n10144), .B(n10126), .Z(n10146) );
  XOR U10761 ( .A(n10166), .B(n10167), .Z(n10126) );
  AND U10762 ( .A(n426), .B(n10168), .Z(n10166) );
  XOR U10763 ( .A(n10169), .B(n10167), .Z(n10168) );
  NANDN U10764 ( .A(n10128), .B(n10130), .Z(n10144) );
  XOR U10765 ( .A(n10170), .B(n10171), .Z(n10130) );
  AND U10766 ( .A(n426), .B(n10172), .Z(n10170) );
  XOR U10767 ( .A(n10171), .B(n10173), .Z(n10172) );
  XOR U10768 ( .A(n10174), .B(n10175), .Z(n426) );
  AND U10769 ( .A(n10176), .B(n10177), .Z(n10174) );
  XNOR U10770 ( .A(n10175), .B(n10141), .Z(n10177) );
  XNOR U10771 ( .A(n10178), .B(n10179), .Z(n10141) );
  ANDN U10772 ( .B(n10180), .A(n10181), .Z(n10178) );
  XOR U10773 ( .A(n10179), .B(n10182), .Z(n10180) );
  XOR U10774 ( .A(n10175), .B(n10143), .Z(n10176) );
  XOR U10775 ( .A(n10183), .B(n10184), .Z(n10143) );
  AND U10776 ( .A(n430), .B(n10185), .Z(n10183) );
  XOR U10777 ( .A(n10186), .B(n10184), .Z(n10185) );
  XNOR U10778 ( .A(n10187), .B(n10188), .Z(n10175) );
  NAND U10779 ( .A(n10189), .B(n10190), .Z(n10188) );
  XOR U10780 ( .A(n10191), .B(n10167), .Z(n10190) );
  XOR U10781 ( .A(n10181), .B(n10182), .Z(n10167) );
  XOR U10782 ( .A(n10192), .B(n10193), .Z(n10182) );
  ANDN U10783 ( .B(n10194), .A(n10195), .Z(n10192) );
  XOR U10784 ( .A(n10193), .B(n10196), .Z(n10194) );
  XOR U10785 ( .A(n10197), .B(n10198), .Z(n10181) );
  XOR U10786 ( .A(n10199), .B(n10200), .Z(n10198) );
  ANDN U10787 ( .B(n10201), .A(n10202), .Z(n10199) );
  XOR U10788 ( .A(n10203), .B(n10200), .Z(n10201) );
  IV U10789 ( .A(n10179), .Z(n10197) );
  XOR U10790 ( .A(n10204), .B(n10205), .Z(n10179) );
  ANDN U10791 ( .B(n10206), .A(n10207), .Z(n10204) );
  XOR U10792 ( .A(n10205), .B(n10208), .Z(n10206) );
  IV U10793 ( .A(n10187), .Z(n10191) );
  XOR U10794 ( .A(n10187), .B(n10169), .Z(n10189) );
  XOR U10795 ( .A(n10209), .B(n10210), .Z(n10169) );
  AND U10796 ( .A(n430), .B(n10211), .Z(n10209) );
  XOR U10797 ( .A(n10212), .B(n10210), .Z(n10211) );
  NANDN U10798 ( .A(n10171), .B(n10173), .Z(n10187) );
  XOR U10799 ( .A(n10213), .B(n10214), .Z(n10173) );
  AND U10800 ( .A(n430), .B(n10215), .Z(n10213) );
  XOR U10801 ( .A(n10214), .B(n10216), .Z(n10215) );
  XOR U10802 ( .A(n10217), .B(n10218), .Z(n430) );
  AND U10803 ( .A(n10219), .B(n10220), .Z(n10217) );
  XNOR U10804 ( .A(n10218), .B(n10184), .Z(n10220) );
  XNOR U10805 ( .A(n10221), .B(n10222), .Z(n10184) );
  ANDN U10806 ( .B(n10223), .A(n10224), .Z(n10221) );
  XOR U10807 ( .A(n10222), .B(n10225), .Z(n10223) );
  XOR U10808 ( .A(n10218), .B(n10186), .Z(n10219) );
  XOR U10809 ( .A(n10226), .B(n10227), .Z(n10186) );
  AND U10810 ( .A(n434), .B(n10228), .Z(n10226) );
  XOR U10811 ( .A(n10229), .B(n10227), .Z(n10228) );
  XNOR U10812 ( .A(n10230), .B(n10231), .Z(n10218) );
  NAND U10813 ( .A(n10232), .B(n10233), .Z(n10231) );
  XOR U10814 ( .A(n10234), .B(n10210), .Z(n10233) );
  XOR U10815 ( .A(n10224), .B(n10225), .Z(n10210) );
  XOR U10816 ( .A(n10235), .B(n10236), .Z(n10225) );
  ANDN U10817 ( .B(n10237), .A(n10238), .Z(n10235) );
  XOR U10818 ( .A(n10236), .B(n10239), .Z(n10237) );
  XOR U10819 ( .A(n10240), .B(n10241), .Z(n10224) );
  XOR U10820 ( .A(n10242), .B(n10243), .Z(n10241) );
  ANDN U10821 ( .B(n10244), .A(n10245), .Z(n10242) );
  XOR U10822 ( .A(n10246), .B(n10243), .Z(n10244) );
  IV U10823 ( .A(n10222), .Z(n10240) );
  XOR U10824 ( .A(n10247), .B(n10248), .Z(n10222) );
  ANDN U10825 ( .B(n10249), .A(n10250), .Z(n10247) );
  XOR U10826 ( .A(n10248), .B(n10251), .Z(n10249) );
  IV U10827 ( .A(n10230), .Z(n10234) );
  XOR U10828 ( .A(n10230), .B(n10212), .Z(n10232) );
  XOR U10829 ( .A(n10252), .B(n10253), .Z(n10212) );
  AND U10830 ( .A(n434), .B(n10254), .Z(n10252) );
  XOR U10831 ( .A(n10255), .B(n10253), .Z(n10254) );
  NANDN U10832 ( .A(n10214), .B(n10216), .Z(n10230) );
  XOR U10833 ( .A(n10256), .B(n10257), .Z(n10216) );
  AND U10834 ( .A(n434), .B(n10258), .Z(n10256) );
  XOR U10835 ( .A(n10257), .B(n10259), .Z(n10258) );
  XOR U10836 ( .A(n10260), .B(n10261), .Z(n434) );
  AND U10837 ( .A(n10262), .B(n10263), .Z(n10260) );
  XNOR U10838 ( .A(n10261), .B(n10227), .Z(n10263) );
  XNOR U10839 ( .A(n10264), .B(n10265), .Z(n10227) );
  ANDN U10840 ( .B(n10266), .A(n10267), .Z(n10264) );
  XOR U10841 ( .A(n10265), .B(n10268), .Z(n10266) );
  XOR U10842 ( .A(n10261), .B(n10229), .Z(n10262) );
  XOR U10843 ( .A(n10269), .B(n10270), .Z(n10229) );
  AND U10844 ( .A(n438), .B(n10271), .Z(n10269) );
  XOR U10845 ( .A(n10272), .B(n10270), .Z(n10271) );
  XNOR U10846 ( .A(n10273), .B(n10274), .Z(n10261) );
  NAND U10847 ( .A(n10275), .B(n10276), .Z(n10274) );
  XOR U10848 ( .A(n10277), .B(n10253), .Z(n10276) );
  XOR U10849 ( .A(n10267), .B(n10268), .Z(n10253) );
  XOR U10850 ( .A(n10278), .B(n10279), .Z(n10268) );
  ANDN U10851 ( .B(n10280), .A(n10281), .Z(n10278) );
  XOR U10852 ( .A(n10279), .B(n10282), .Z(n10280) );
  XOR U10853 ( .A(n10283), .B(n10284), .Z(n10267) );
  XOR U10854 ( .A(n10285), .B(n10286), .Z(n10284) );
  ANDN U10855 ( .B(n10287), .A(n10288), .Z(n10285) );
  XOR U10856 ( .A(n10289), .B(n10286), .Z(n10287) );
  IV U10857 ( .A(n10265), .Z(n10283) );
  XOR U10858 ( .A(n10290), .B(n10291), .Z(n10265) );
  ANDN U10859 ( .B(n10292), .A(n10293), .Z(n10290) );
  XOR U10860 ( .A(n10291), .B(n10294), .Z(n10292) );
  IV U10861 ( .A(n10273), .Z(n10277) );
  XOR U10862 ( .A(n10273), .B(n10255), .Z(n10275) );
  XOR U10863 ( .A(n10295), .B(n10296), .Z(n10255) );
  AND U10864 ( .A(n438), .B(n10297), .Z(n10295) );
  XOR U10865 ( .A(n10298), .B(n10296), .Z(n10297) );
  NANDN U10866 ( .A(n10257), .B(n10259), .Z(n10273) );
  XOR U10867 ( .A(n10299), .B(n10300), .Z(n10259) );
  AND U10868 ( .A(n438), .B(n10301), .Z(n10299) );
  XOR U10869 ( .A(n10300), .B(n10302), .Z(n10301) );
  XOR U10870 ( .A(n10303), .B(n10304), .Z(n438) );
  AND U10871 ( .A(n10305), .B(n10306), .Z(n10303) );
  XNOR U10872 ( .A(n10304), .B(n10270), .Z(n10306) );
  XNOR U10873 ( .A(n10307), .B(n10308), .Z(n10270) );
  ANDN U10874 ( .B(n10309), .A(n10310), .Z(n10307) );
  XOR U10875 ( .A(n10308), .B(n10311), .Z(n10309) );
  XOR U10876 ( .A(n10304), .B(n10272), .Z(n10305) );
  XOR U10877 ( .A(n10312), .B(n10313), .Z(n10272) );
  AND U10878 ( .A(n442), .B(n10314), .Z(n10312) );
  XOR U10879 ( .A(n10315), .B(n10313), .Z(n10314) );
  XNOR U10880 ( .A(n10316), .B(n10317), .Z(n10304) );
  NAND U10881 ( .A(n10318), .B(n10319), .Z(n10317) );
  XOR U10882 ( .A(n10320), .B(n10296), .Z(n10319) );
  XOR U10883 ( .A(n10310), .B(n10311), .Z(n10296) );
  XOR U10884 ( .A(n10321), .B(n10322), .Z(n10311) );
  ANDN U10885 ( .B(n10323), .A(n10324), .Z(n10321) );
  XOR U10886 ( .A(n10322), .B(n10325), .Z(n10323) );
  XOR U10887 ( .A(n10326), .B(n10327), .Z(n10310) );
  XOR U10888 ( .A(n10328), .B(n10329), .Z(n10327) );
  ANDN U10889 ( .B(n10330), .A(n10331), .Z(n10328) );
  XOR U10890 ( .A(n10332), .B(n10329), .Z(n10330) );
  IV U10891 ( .A(n10308), .Z(n10326) );
  XOR U10892 ( .A(n10333), .B(n10334), .Z(n10308) );
  ANDN U10893 ( .B(n10335), .A(n10336), .Z(n10333) );
  XOR U10894 ( .A(n10334), .B(n10337), .Z(n10335) );
  IV U10895 ( .A(n10316), .Z(n10320) );
  XOR U10896 ( .A(n10316), .B(n10298), .Z(n10318) );
  XOR U10897 ( .A(n10338), .B(n10339), .Z(n10298) );
  AND U10898 ( .A(n442), .B(n10340), .Z(n10338) );
  XOR U10899 ( .A(n10341), .B(n10339), .Z(n10340) );
  NANDN U10900 ( .A(n10300), .B(n10302), .Z(n10316) );
  XOR U10901 ( .A(n10342), .B(n10343), .Z(n10302) );
  AND U10902 ( .A(n442), .B(n10344), .Z(n10342) );
  XOR U10903 ( .A(n10343), .B(n10345), .Z(n10344) );
  XOR U10904 ( .A(n10346), .B(n10347), .Z(n442) );
  AND U10905 ( .A(n10348), .B(n10349), .Z(n10346) );
  XNOR U10906 ( .A(n10347), .B(n10313), .Z(n10349) );
  XNOR U10907 ( .A(n10350), .B(n10351), .Z(n10313) );
  ANDN U10908 ( .B(n10352), .A(n10353), .Z(n10350) );
  XOR U10909 ( .A(n10351), .B(n10354), .Z(n10352) );
  XOR U10910 ( .A(n10347), .B(n10315), .Z(n10348) );
  XOR U10911 ( .A(n10355), .B(n10356), .Z(n10315) );
  AND U10912 ( .A(n446), .B(n10357), .Z(n10355) );
  XOR U10913 ( .A(n10358), .B(n10356), .Z(n10357) );
  XNOR U10914 ( .A(n10359), .B(n10360), .Z(n10347) );
  NAND U10915 ( .A(n10361), .B(n10362), .Z(n10360) );
  XOR U10916 ( .A(n10363), .B(n10339), .Z(n10362) );
  XOR U10917 ( .A(n10353), .B(n10354), .Z(n10339) );
  XOR U10918 ( .A(n10364), .B(n10365), .Z(n10354) );
  ANDN U10919 ( .B(n10366), .A(n10367), .Z(n10364) );
  XOR U10920 ( .A(n10365), .B(n10368), .Z(n10366) );
  XOR U10921 ( .A(n10369), .B(n10370), .Z(n10353) );
  XOR U10922 ( .A(n10371), .B(n10372), .Z(n10370) );
  ANDN U10923 ( .B(n10373), .A(n10374), .Z(n10371) );
  XOR U10924 ( .A(n10375), .B(n10372), .Z(n10373) );
  IV U10925 ( .A(n10351), .Z(n10369) );
  XOR U10926 ( .A(n10376), .B(n10377), .Z(n10351) );
  ANDN U10927 ( .B(n10378), .A(n10379), .Z(n10376) );
  XOR U10928 ( .A(n10377), .B(n10380), .Z(n10378) );
  IV U10929 ( .A(n10359), .Z(n10363) );
  XOR U10930 ( .A(n10359), .B(n10341), .Z(n10361) );
  XOR U10931 ( .A(n10381), .B(n10382), .Z(n10341) );
  AND U10932 ( .A(n446), .B(n10383), .Z(n10381) );
  XOR U10933 ( .A(n10384), .B(n10382), .Z(n10383) );
  NANDN U10934 ( .A(n10343), .B(n10345), .Z(n10359) );
  XOR U10935 ( .A(n10385), .B(n10386), .Z(n10345) );
  AND U10936 ( .A(n446), .B(n10387), .Z(n10385) );
  XOR U10937 ( .A(n10386), .B(n10388), .Z(n10387) );
  XOR U10938 ( .A(n10389), .B(n10390), .Z(n446) );
  AND U10939 ( .A(n10391), .B(n10392), .Z(n10389) );
  XNOR U10940 ( .A(n10390), .B(n10356), .Z(n10392) );
  XNOR U10941 ( .A(n10393), .B(n10394), .Z(n10356) );
  ANDN U10942 ( .B(n10395), .A(n10396), .Z(n10393) );
  XOR U10943 ( .A(n10394), .B(n10397), .Z(n10395) );
  XOR U10944 ( .A(n10390), .B(n10358), .Z(n10391) );
  XOR U10945 ( .A(n10398), .B(n10399), .Z(n10358) );
  AND U10946 ( .A(n450), .B(n10400), .Z(n10398) );
  XOR U10947 ( .A(n10401), .B(n10399), .Z(n10400) );
  XNOR U10948 ( .A(n10402), .B(n10403), .Z(n10390) );
  NAND U10949 ( .A(n10404), .B(n10405), .Z(n10403) );
  XOR U10950 ( .A(n10406), .B(n10382), .Z(n10405) );
  XOR U10951 ( .A(n10396), .B(n10397), .Z(n10382) );
  XOR U10952 ( .A(n10407), .B(n10408), .Z(n10397) );
  ANDN U10953 ( .B(n10409), .A(n10410), .Z(n10407) );
  XOR U10954 ( .A(n10408), .B(n10411), .Z(n10409) );
  XOR U10955 ( .A(n10412), .B(n10413), .Z(n10396) );
  XOR U10956 ( .A(n10414), .B(n10415), .Z(n10413) );
  ANDN U10957 ( .B(n10416), .A(n10417), .Z(n10414) );
  XOR U10958 ( .A(n10418), .B(n10415), .Z(n10416) );
  IV U10959 ( .A(n10394), .Z(n10412) );
  XOR U10960 ( .A(n10419), .B(n10420), .Z(n10394) );
  ANDN U10961 ( .B(n10421), .A(n10422), .Z(n10419) );
  XOR U10962 ( .A(n10420), .B(n10423), .Z(n10421) );
  IV U10963 ( .A(n10402), .Z(n10406) );
  XOR U10964 ( .A(n10402), .B(n10384), .Z(n10404) );
  XOR U10965 ( .A(n10424), .B(n10425), .Z(n10384) );
  AND U10966 ( .A(n450), .B(n10426), .Z(n10424) );
  XOR U10967 ( .A(n10427), .B(n10425), .Z(n10426) );
  NANDN U10968 ( .A(n10386), .B(n10388), .Z(n10402) );
  XOR U10969 ( .A(n10428), .B(n10429), .Z(n10388) );
  AND U10970 ( .A(n450), .B(n10430), .Z(n10428) );
  XOR U10971 ( .A(n10429), .B(n10431), .Z(n10430) );
  XOR U10972 ( .A(n10432), .B(n10433), .Z(n450) );
  AND U10973 ( .A(n10434), .B(n10435), .Z(n10432) );
  XNOR U10974 ( .A(n10433), .B(n10399), .Z(n10435) );
  XNOR U10975 ( .A(n10436), .B(n10437), .Z(n10399) );
  ANDN U10976 ( .B(n10438), .A(n10439), .Z(n10436) );
  XOR U10977 ( .A(n10437), .B(n10440), .Z(n10438) );
  XOR U10978 ( .A(n10433), .B(n10401), .Z(n10434) );
  XOR U10979 ( .A(n10441), .B(n10442), .Z(n10401) );
  AND U10980 ( .A(n454), .B(n10443), .Z(n10441) );
  XOR U10981 ( .A(n10444), .B(n10442), .Z(n10443) );
  XNOR U10982 ( .A(n10445), .B(n10446), .Z(n10433) );
  NAND U10983 ( .A(n10447), .B(n10448), .Z(n10446) );
  XOR U10984 ( .A(n10449), .B(n10425), .Z(n10448) );
  XOR U10985 ( .A(n10439), .B(n10440), .Z(n10425) );
  XOR U10986 ( .A(n10450), .B(n10451), .Z(n10440) );
  ANDN U10987 ( .B(n10452), .A(n10453), .Z(n10450) );
  XOR U10988 ( .A(n10451), .B(n10454), .Z(n10452) );
  XOR U10989 ( .A(n10455), .B(n10456), .Z(n10439) );
  XOR U10990 ( .A(n10457), .B(n10458), .Z(n10456) );
  ANDN U10991 ( .B(n10459), .A(n10460), .Z(n10457) );
  XOR U10992 ( .A(n10461), .B(n10458), .Z(n10459) );
  IV U10993 ( .A(n10437), .Z(n10455) );
  XOR U10994 ( .A(n10462), .B(n10463), .Z(n10437) );
  ANDN U10995 ( .B(n10464), .A(n10465), .Z(n10462) );
  XOR U10996 ( .A(n10463), .B(n10466), .Z(n10464) );
  IV U10997 ( .A(n10445), .Z(n10449) );
  XOR U10998 ( .A(n10445), .B(n10427), .Z(n10447) );
  XOR U10999 ( .A(n10467), .B(n10468), .Z(n10427) );
  AND U11000 ( .A(n454), .B(n10469), .Z(n10467) );
  XOR U11001 ( .A(n10470), .B(n10468), .Z(n10469) );
  NANDN U11002 ( .A(n10429), .B(n10431), .Z(n10445) );
  XOR U11003 ( .A(n10471), .B(n10472), .Z(n10431) );
  AND U11004 ( .A(n454), .B(n10473), .Z(n10471) );
  XOR U11005 ( .A(n10472), .B(n10474), .Z(n10473) );
  XOR U11006 ( .A(n10475), .B(n10476), .Z(n454) );
  AND U11007 ( .A(n10477), .B(n10478), .Z(n10475) );
  XNOR U11008 ( .A(n10476), .B(n10442), .Z(n10478) );
  XNOR U11009 ( .A(n10479), .B(n10480), .Z(n10442) );
  ANDN U11010 ( .B(n10481), .A(n10482), .Z(n10479) );
  XOR U11011 ( .A(n10480), .B(n10483), .Z(n10481) );
  XOR U11012 ( .A(n10476), .B(n10444), .Z(n10477) );
  XOR U11013 ( .A(n10484), .B(n10485), .Z(n10444) );
  AND U11014 ( .A(n458), .B(n10486), .Z(n10484) );
  XOR U11015 ( .A(n10487), .B(n10485), .Z(n10486) );
  XNOR U11016 ( .A(n10488), .B(n10489), .Z(n10476) );
  NAND U11017 ( .A(n10490), .B(n10491), .Z(n10489) );
  XOR U11018 ( .A(n10492), .B(n10468), .Z(n10491) );
  XOR U11019 ( .A(n10482), .B(n10483), .Z(n10468) );
  XOR U11020 ( .A(n10493), .B(n10494), .Z(n10483) );
  ANDN U11021 ( .B(n10495), .A(n10496), .Z(n10493) );
  XOR U11022 ( .A(n10494), .B(n10497), .Z(n10495) );
  XOR U11023 ( .A(n10498), .B(n10499), .Z(n10482) );
  XOR U11024 ( .A(n10500), .B(n10501), .Z(n10499) );
  ANDN U11025 ( .B(n10502), .A(n10503), .Z(n10500) );
  XOR U11026 ( .A(n10504), .B(n10501), .Z(n10502) );
  IV U11027 ( .A(n10480), .Z(n10498) );
  XOR U11028 ( .A(n10505), .B(n10506), .Z(n10480) );
  ANDN U11029 ( .B(n10507), .A(n10508), .Z(n10505) );
  XOR U11030 ( .A(n10506), .B(n10509), .Z(n10507) );
  IV U11031 ( .A(n10488), .Z(n10492) );
  XOR U11032 ( .A(n10488), .B(n10470), .Z(n10490) );
  XOR U11033 ( .A(n10510), .B(n10511), .Z(n10470) );
  AND U11034 ( .A(n458), .B(n10512), .Z(n10510) );
  XOR U11035 ( .A(n10513), .B(n10511), .Z(n10512) );
  NANDN U11036 ( .A(n10472), .B(n10474), .Z(n10488) );
  XOR U11037 ( .A(n10514), .B(n10515), .Z(n10474) );
  AND U11038 ( .A(n458), .B(n10516), .Z(n10514) );
  XOR U11039 ( .A(n10515), .B(n10517), .Z(n10516) );
  XOR U11040 ( .A(n10518), .B(n10519), .Z(n458) );
  AND U11041 ( .A(n10520), .B(n10521), .Z(n10518) );
  XNOR U11042 ( .A(n10519), .B(n10485), .Z(n10521) );
  XNOR U11043 ( .A(n10522), .B(n10523), .Z(n10485) );
  ANDN U11044 ( .B(n10524), .A(n10525), .Z(n10522) );
  XOR U11045 ( .A(n10523), .B(n10526), .Z(n10524) );
  XOR U11046 ( .A(n10519), .B(n10487), .Z(n10520) );
  XOR U11047 ( .A(n10527), .B(n10528), .Z(n10487) );
  AND U11048 ( .A(n462), .B(n10529), .Z(n10527) );
  XOR U11049 ( .A(n10530), .B(n10528), .Z(n10529) );
  XNOR U11050 ( .A(n10531), .B(n10532), .Z(n10519) );
  NAND U11051 ( .A(n10533), .B(n10534), .Z(n10532) );
  XOR U11052 ( .A(n10535), .B(n10511), .Z(n10534) );
  XOR U11053 ( .A(n10525), .B(n10526), .Z(n10511) );
  XOR U11054 ( .A(n10536), .B(n10537), .Z(n10526) );
  ANDN U11055 ( .B(n10538), .A(n10539), .Z(n10536) );
  XOR U11056 ( .A(n10537), .B(n10540), .Z(n10538) );
  XOR U11057 ( .A(n10541), .B(n10542), .Z(n10525) );
  XOR U11058 ( .A(n10543), .B(n10544), .Z(n10542) );
  ANDN U11059 ( .B(n10545), .A(n10546), .Z(n10543) );
  XOR U11060 ( .A(n10547), .B(n10544), .Z(n10545) );
  IV U11061 ( .A(n10523), .Z(n10541) );
  XOR U11062 ( .A(n10548), .B(n10549), .Z(n10523) );
  ANDN U11063 ( .B(n10550), .A(n10551), .Z(n10548) );
  XOR U11064 ( .A(n10549), .B(n10552), .Z(n10550) );
  IV U11065 ( .A(n10531), .Z(n10535) );
  XOR U11066 ( .A(n10531), .B(n10513), .Z(n10533) );
  XOR U11067 ( .A(n10553), .B(n10554), .Z(n10513) );
  AND U11068 ( .A(n462), .B(n10555), .Z(n10553) );
  XOR U11069 ( .A(n10556), .B(n10554), .Z(n10555) );
  NANDN U11070 ( .A(n10515), .B(n10517), .Z(n10531) );
  XOR U11071 ( .A(n10557), .B(n10558), .Z(n10517) );
  AND U11072 ( .A(n462), .B(n10559), .Z(n10557) );
  XOR U11073 ( .A(n10558), .B(n10560), .Z(n10559) );
  XOR U11074 ( .A(n10561), .B(n10562), .Z(n462) );
  AND U11075 ( .A(n10563), .B(n10564), .Z(n10561) );
  XNOR U11076 ( .A(n10562), .B(n10528), .Z(n10564) );
  XNOR U11077 ( .A(n10565), .B(n10566), .Z(n10528) );
  ANDN U11078 ( .B(n10567), .A(n10568), .Z(n10565) );
  XOR U11079 ( .A(n10566), .B(n10569), .Z(n10567) );
  XOR U11080 ( .A(n10562), .B(n10530), .Z(n10563) );
  XOR U11081 ( .A(n10570), .B(n10571), .Z(n10530) );
  AND U11082 ( .A(n466), .B(n10572), .Z(n10570) );
  XOR U11083 ( .A(n10573), .B(n10571), .Z(n10572) );
  XNOR U11084 ( .A(n10574), .B(n10575), .Z(n10562) );
  NAND U11085 ( .A(n10576), .B(n10577), .Z(n10575) );
  XOR U11086 ( .A(n10578), .B(n10554), .Z(n10577) );
  XOR U11087 ( .A(n10568), .B(n10569), .Z(n10554) );
  XOR U11088 ( .A(n10579), .B(n10580), .Z(n10569) );
  ANDN U11089 ( .B(n10581), .A(n10582), .Z(n10579) );
  XOR U11090 ( .A(n10580), .B(n10583), .Z(n10581) );
  XOR U11091 ( .A(n10584), .B(n10585), .Z(n10568) );
  XOR U11092 ( .A(n10586), .B(n10587), .Z(n10585) );
  ANDN U11093 ( .B(n10588), .A(n10589), .Z(n10586) );
  XOR U11094 ( .A(n10590), .B(n10587), .Z(n10588) );
  IV U11095 ( .A(n10566), .Z(n10584) );
  XOR U11096 ( .A(n10591), .B(n10592), .Z(n10566) );
  ANDN U11097 ( .B(n10593), .A(n10594), .Z(n10591) );
  XOR U11098 ( .A(n10592), .B(n10595), .Z(n10593) );
  IV U11099 ( .A(n10574), .Z(n10578) );
  XOR U11100 ( .A(n10574), .B(n10556), .Z(n10576) );
  XOR U11101 ( .A(n10596), .B(n10597), .Z(n10556) );
  AND U11102 ( .A(n466), .B(n10598), .Z(n10596) );
  XOR U11103 ( .A(n10599), .B(n10597), .Z(n10598) );
  NANDN U11104 ( .A(n10558), .B(n10560), .Z(n10574) );
  XOR U11105 ( .A(n10600), .B(n10601), .Z(n10560) );
  AND U11106 ( .A(n466), .B(n10602), .Z(n10600) );
  XOR U11107 ( .A(n10601), .B(n10603), .Z(n10602) );
  XOR U11108 ( .A(n10604), .B(n10605), .Z(n466) );
  AND U11109 ( .A(n10606), .B(n10607), .Z(n10604) );
  XNOR U11110 ( .A(n10605), .B(n10571), .Z(n10607) );
  XNOR U11111 ( .A(n10608), .B(n10609), .Z(n10571) );
  ANDN U11112 ( .B(n10610), .A(n10611), .Z(n10608) );
  XOR U11113 ( .A(n10609), .B(n10612), .Z(n10610) );
  XOR U11114 ( .A(n10605), .B(n10573), .Z(n10606) );
  XOR U11115 ( .A(n10613), .B(n10614), .Z(n10573) );
  AND U11116 ( .A(n470), .B(n10615), .Z(n10613) );
  XOR U11117 ( .A(n10616), .B(n10614), .Z(n10615) );
  XNOR U11118 ( .A(n10617), .B(n10618), .Z(n10605) );
  NAND U11119 ( .A(n10619), .B(n10620), .Z(n10618) );
  XOR U11120 ( .A(n10621), .B(n10597), .Z(n10620) );
  XOR U11121 ( .A(n10611), .B(n10612), .Z(n10597) );
  XOR U11122 ( .A(n10622), .B(n10623), .Z(n10612) );
  ANDN U11123 ( .B(n10624), .A(n10625), .Z(n10622) );
  XOR U11124 ( .A(n10623), .B(n10626), .Z(n10624) );
  XOR U11125 ( .A(n10627), .B(n10628), .Z(n10611) );
  XOR U11126 ( .A(n10629), .B(n10630), .Z(n10628) );
  ANDN U11127 ( .B(n10631), .A(n10632), .Z(n10629) );
  XOR U11128 ( .A(n10633), .B(n10630), .Z(n10631) );
  IV U11129 ( .A(n10609), .Z(n10627) );
  XOR U11130 ( .A(n10634), .B(n10635), .Z(n10609) );
  ANDN U11131 ( .B(n10636), .A(n10637), .Z(n10634) );
  XOR U11132 ( .A(n10635), .B(n10638), .Z(n10636) );
  IV U11133 ( .A(n10617), .Z(n10621) );
  XOR U11134 ( .A(n10617), .B(n10599), .Z(n10619) );
  XOR U11135 ( .A(n10639), .B(n10640), .Z(n10599) );
  AND U11136 ( .A(n470), .B(n10641), .Z(n10639) );
  XOR U11137 ( .A(n10642), .B(n10640), .Z(n10641) );
  NANDN U11138 ( .A(n10601), .B(n10603), .Z(n10617) );
  XOR U11139 ( .A(n10643), .B(n10644), .Z(n10603) );
  AND U11140 ( .A(n470), .B(n10645), .Z(n10643) );
  XOR U11141 ( .A(n10644), .B(n10646), .Z(n10645) );
  XOR U11142 ( .A(n10647), .B(n10648), .Z(n470) );
  AND U11143 ( .A(n10649), .B(n10650), .Z(n10647) );
  XNOR U11144 ( .A(n10648), .B(n10614), .Z(n10650) );
  XNOR U11145 ( .A(n10651), .B(n10652), .Z(n10614) );
  ANDN U11146 ( .B(n10653), .A(n10654), .Z(n10651) );
  XOR U11147 ( .A(n10652), .B(n10655), .Z(n10653) );
  XOR U11148 ( .A(n10648), .B(n10616), .Z(n10649) );
  XOR U11149 ( .A(n10656), .B(n10657), .Z(n10616) );
  AND U11150 ( .A(n474), .B(n10658), .Z(n10656) );
  XOR U11151 ( .A(n10659), .B(n10657), .Z(n10658) );
  XNOR U11152 ( .A(n10660), .B(n10661), .Z(n10648) );
  NAND U11153 ( .A(n10662), .B(n10663), .Z(n10661) );
  XOR U11154 ( .A(n10664), .B(n10640), .Z(n10663) );
  XOR U11155 ( .A(n10654), .B(n10655), .Z(n10640) );
  XOR U11156 ( .A(n10665), .B(n10666), .Z(n10655) );
  ANDN U11157 ( .B(n10667), .A(n10668), .Z(n10665) );
  XOR U11158 ( .A(n10666), .B(n10669), .Z(n10667) );
  XOR U11159 ( .A(n10670), .B(n10671), .Z(n10654) );
  XOR U11160 ( .A(n10672), .B(n10673), .Z(n10671) );
  ANDN U11161 ( .B(n10674), .A(n10675), .Z(n10672) );
  XOR U11162 ( .A(n10676), .B(n10673), .Z(n10674) );
  IV U11163 ( .A(n10652), .Z(n10670) );
  XOR U11164 ( .A(n10677), .B(n10678), .Z(n10652) );
  ANDN U11165 ( .B(n10679), .A(n10680), .Z(n10677) );
  XOR U11166 ( .A(n10678), .B(n10681), .Z(n10679) );
  IV U11167 ( .A(n10660), .Z(n10664) );
  XOR U11168 ( .A(n10660), .B(n10642), .Z(n10662) );
  XOR U11169 ( .A(n10682), .B(n10683), .Z(n10642) );
  AND U11170 ( .A(n474), .B(n10684), .Z(n10682) );
  XOR U11171 ( .A(n10685), .B(n10683), .Z(n10684) );
  NANDN U11172 ( .A(n10644), .B(n10646), .Z(n10660) );
  XOR U11173 ( .A(n10686), .B(n10687), .Z(n10646) );
  AND U11174 ( .A(n474), .B(n10688), .Z(n10686) );
  XOR U11175 ( .A(n10687), .B(n10689), .Z(n10688) );
  XOR U11176 ( .A(n10690), .B(n10691), .Z(n474) );
  AND U11177 ( .A(n10692), .B(n10693), .Z(n10690) );
  XNOR U11178 ( .A(n10691), .B(n10657), .Z(n10693) );
  XNOR U11179 ( .A(n10694), .B(n10695), .Z(n10657) );
  ANDN U11180 ( .B(n10696), .A(n10697), .Z(n10694) );
  XOR U11181 ( .A(n10695), .B(n10698), .Z(n10696) );
  XOR U11182 ( .A(n10691), .B(n10659), .Z(n10692) );
  XOR U11183 ( .A(n10699), .B(n10700), .Z(n10659) );
  AND U11184 ( .A(n478), .B(n10701), .Z(n10699) );
  XOR U11185 ( .A(n10702), .B(n10700), .Z(n10701) );
  XNOR U11186 ( .A(n10703), .B(n10704), .Z(n10691) );
  NAND U11187 ( .A(n10705), .B(n10706), .Z(n10704) );
  XOR U11188 ( .A(n10707), .B(n10683), .Z(n10706) );
  XOR U11189 ( .A(n10697), .B(n10698), .Z(n10683) );
  XOR U11190 ( .A(n10708), .B(n10709), .Z(n10698) );
  ANDN U11191 ( .B(n10710), .A(n10711), .Z(n10708) );
  XOR U11192 ( .A(n10709), .B(n10712), .Z(n10710) );
  XOR U11193 ( .A(n10713), .B(n10714), .Z(n10697) );
  XOR U11194 ( .A(n10715), .B(n10716), .Z(n10714) );
  ANDN U11195 ( .B(n10717), .A(n10718), .Z(n10715) );
  XOR U11196 ( .A(n10719), .B(n10716), .Z(n10717) );
  IV U11197 ( .A(n10695), .Z(n10713) );
  XOR U11198 ( .A(n10720), .B(n10721), .Z(n10695) );
  ANDN U11199 ( .B(n10722), .A(n10723), .Z(n10720) );
  XOR U11200 ( .A(n10721), .B(n10724), .Z(n10722) );
  IV U11201 ( .A(n10703), .Z(n10707) );
  XOR U11202 ( .A(n10703), .B(n10685), .Z(n10705) );
  XOR U11203 ( .A(n10725), .B(n10726), .Z(n10685) );
  AND U11204 ( .A(n478), .B(n10727), .Z(n10725) );
  XOR U11205 ( .A(n10728), .B(n10726), .Z(n10727) );
  NANDN U11206 ( .A(n10687), .B(n10689), .Z(n10703) );
  XOR U11207 ( .A(n10729), .B(n10730), .Z(n10689) );
  AND U11208 ( .A(n478), .B(n10731), .Z(n10729) );
  XOR U11209 ( .A(n10730), .B(n10732), .Z(n10731) );
  XOR U11210 ( .A(n10733), .B(n10734), .Z(n478) );
  AND U11211 ( .A(n10735), .B(n10736), .Z(n10733) );
  XNOR U11212 ( .A(n10734), .B(n10700), .Z(n10736) );
  XNOR U11213 ( .A(n10737), .B(n10738), .Z(n10700) );
  ANDN U11214 ( .B(n10739), .A(n10740), .Z(n10737) );
  XOR U11215 ( .A(n10738), .B(n10741), .Z(n10739) );
  XOR U11216 ( .A(n10734), .B(n10702), .Z(n10735) );
  XOR U11217 ( .A(n10742), .B(n10743), .Z(n10702) );
  AND U11218 ( .A(n482), .B(n10744), .Z(n10742) );
  XOR U11219 ( .A(n10745), .B(n10743), .Z(n10744) );
  XNOR U11220 ( .A(n10746), .B(n10747), .Z(n10734) );
  NAND U11221 ( .A(n10748), .B(n10749), .Z(n10747) );
  XOR U11222 ( .A(n10750), .B(n10726), .Z(n10749) );
  XOR U11223 ( .A(n10740), .B(n10741), .Z(n10726) );
  XOR U11224 ( .A(n10751), .B(n10752), .Z(n10741) );
  ANDN U11225 ( .B(n10753), .A(n10754), .Z(n10751) );
  XOR U11226 ( .A(n10752), .B(n10755), .Z(n10753) );
  XOR U11227 ( .A(n10756), .B(n10757), .Z(n10740) );
  XOR U11228 ( .A(n10758), .B(n10759), .Z(n10757) );
  ANDN U11229 ( .B(n10760), .A(n10761), .Z(n10758) );
  XOR U11230 ( .A(n10762), .B(n10759), .Z(n10760) );
  IV U11231 ( .A(n10738), .Z(n10756) );
  XOR U11232 ( .A(n10763), .B(n10764), .Z(n10738) );
  ANDN U11233 ( .B(n10765), .A(n10766), .Z(n10763) );
  XOR U11234 ( .A(n10764), .B(n10767), .Z(n10765) );
  IV U11235 ( .A(n10746), .Z(n10750) );
  XOR U11236 ( .A(n10746), .B(n10728), .Z(n10748) );
  XOR U11237 ( .A(n10768), .B(n10769), .Z(n10728) );
  AND U11238 ( .A(n482), .B(n10770), .Z(n10768) );
  XOR U11239 ( .A(n10771), .B(n10769), .Z(n10770) );
  NANDN U11240 ( .A(n10730), .B(n10732), .Z(n10746) );
  XOR U11241 ( .A(n10772), .B(n10773), .Z(n10732) );
  AND U11242 ( .A(n482), .B(n10774), .Z(n10772) );
  XOR U11243 ( .A(n10773), .B(n10775), .Z(n10774) );
  XOR U11244 ( .A(n10776), .B(n10777), .Z(n482) );
  AND U11245 ( .A(n10778), .B(n10779), .Z(n10776) );
  XNOR U11246 ( .A(n10777), .B(n10743), .Z(n10779) );
  XNOR U11247 ( .A(n10780), .B(n10781), .Z(n10743) );
  ANDN U11248 ( .B(n10782), .A(n10783), .Z(n10780) );
  XOR U11249 ( .A(n10781), .B(n10784), .Z(n10782) );
  XOR U11250 ( .A(n10777), .B(n10745), .Z(n10778) );
  XOR U11251 ( .A(n10785), .B(n10786), .Z(n10745) );
  AND U11252 ( .A(n486), .B(n10787), .Z(n10785) );
  XOR U11253 ( .A(n10788), .B(n10786), .Z(n10787) );
  XNOR U11254 ( .A(n10789), .B(n10790), .Z(n10777) );
  NAND U11255 ( .A(n10791), .B(n10792), .Z(n10790) );
  XOR U11256 ( .A(n10793), .B(n10769), .Z(n10792) );
  XOR U11257 ( .A(n10783), .B(n10784), .Z(n10769) );
  XOR U11258 ( .A(n10794), .B(n10795), .Z(n10784) );
  ANDN U11259 ( .B(n10796), .A(n10797), .Z(n10794) );
  XOR U11260 ( .A(n10795), .B(n10798), .Z(n10796) );
  XOR U11261 ( .A(n10799), .B(n10800), .Z(n10783) );
  XOR U11262 ( .A(n10801), .B(n10802), .Z(n10800) );
  ANDN U11263 ( .B(n10803), .A(n10804), .Z(n10801) );
  XOR U11264 ( .A(n10805), .B(n10802), .Z(n10803) );
  IV U11265 ( .A(n10781), .Z(n10799) );
  XOR U11266 ( .A(n10806), .B(n10807), .Z(n10781) );
  ANDN U11267 ( .B(n10808), .A(n10809), .Z(n10806) );
  XOR U11268 ( .A(n10807), .B(n10810), .Z(n10808) );
  IV U11269 ( .A(n10789), .Z(n10793) );
  XOR U11270 ( .A(n10789), .B(n10771), .Z(n10791) );
  XOR U11271 ( .A(n10811), .B(n10812), .Z(n10771) );
  AND U11272 ( .A(n486), .B(n10813), .Z(n10811) );
  XOR U11273 ( .A(n10814), .B(n10812), .Z(n10813) );
  NANDN U11274 ( .A(n10773), .B(n10775), .Z(n10789) );
  XOR U11275 ( .A(n10815), .B(n10816), .Z(n10775) );
  AND U11276 ( .A(n486), .B(n10817), .Z(n10815) );
  XOR U11277 ( .A(n10816), .B(n10818), .Z(n10817) );
  XOR U11278 ( .A(n10819), .B(n10820), .Z(n486) );
  AND U11279 ( .A(n10821), .B(n10822), .Z(n10819) );
  XNOR U11280 ( .A(n10820), .B(n10786), .Z(n10822) );
  XNOR U11281 ( .A(n10823), .B(n10824), .Z(n10786) );
  ANDN U11282 ( .B(n10825), .A(n10826), .Z(n10823) );
  XOR U11283 ( .A(n10824), .B(n10827), .Z(n10825) );
  XOR U11284 ( .A(n10820), .B(n10788), .Z(n10821) );
  XOR U11285 ( .A(n10828), .B(n10829), .Z(n10788) );
  AND U11286 ( .A(n490), .B(n10830), .Z(n10828) );
  XOR U11287 ( .A(n10831), .B(n10829), .Z(n10830) );
  XNOR U11288 ( .A(n10832), .B(n10833), .Z(n10820) );
  NAND U11289 ( .A(n10834), .B(n10835), .Z(n10833) );
  XOR U11290 ( .A(n10836), .B(n10812), .Z(n10835) );
  XOR U11291 ( .A(n10826), .B(n10827), .Z(n10812) );
  XOR U11292 ( .A(n10837), .B(n10838), .Z(n10827) );
  ANDN U11293 ( .B(n10839), .A(n10840), .Z(n10837) );
  XOR U11294 ( .A(n10838), .B(n10841), .Z(n10839) );
  XOR U11295 ( .A(n10842), .B(n10843), .Z(n10826) );
  XOR U11296 ( .A(n10844), .B(n10845), .Z(n10843) );
  ANDN U11297 ( .B(n10846), .A(n10847), .Z(n10844) );
  XOR U11298 ( .A(n10848), .B(n10845), .Z(n10846) );
  IV U11299 ( .A(n10824), .Z(n10842) );
  XOR U11300 ( .A(n10849), .B(n10850), .Z(n10824) );
  ANDN U11301 ( .B(n10851), .A(n10852), .Z(n10849) );
  XOR U11302 ( .A(n10850), .B(n10853), .Z(n10851) );
  IV U11303 ( .A(n10832), .Z(n10836) );
  XOR U11304 ( .A(n10832), .B(n10814), .Z(n10834) );
  XOR U11305 ( .A(n10854), .B(n10855), .Z(n10814) );
  AND U11306 ( .A(n490), .B(n10856), .Z(n10854) );
  XOR U11307 ( .A(n10857), .B(n10855), .Z(n10856) );
  NANDN U11308 ( .A(n10816), .B(n10818), .Z(n10832) );
  XOR U11309 ( .A(n10858), .B(n10859), .Z(n10818) );
  AND U11310 ( .A(n490), .B(n10860), .Z(n10858) );
  XOR U11311 ( .A(n10859), .B(n10861), .Z(n10860) );
  XOR U11312 ( .A(n10862), .B(n10863), .Z(n490) );
  AND U11313 ( .A(n10864), .B(n10865), .Z(n10862) );
  XNOR U11314 ( .A(n10863), .B(n10829), .Z(n10865) );
  XNOR U11315 ( .A(n10866), .B(n10867), .Z(n10829) );
  ANDN U11316 ( .B(n10868), .A(n10869), .Z(n10866) );
  XOR U11317 ( .A(n10867), .B(n10870), .Z(n10868) );
  XOR U11318 ( .A(n10863), .B(n10831), .Z(n10864) );
  XOR U11319 ( .A(n10871), .B(n10872), .Z(n10831) );
  AND U11320 ( .A(n494), .B(n10873), .Z(n10871) );
  XOR U11321 ( .A(n10874), .B(n10872), .Z(n10873) );
  XNOR U11322 ( .A(n10875), .B(n10876), .Z(n10863) );
  NAND U11323 ( .A(n10877), .B(n10878), .Z(n10876) );
  XOR U11324 ( .A(n10879), .B(n10855), .Z(n10878) );
  XOR U11325 ( .A(n10869), .B(n10870), .Z(n10855) );
  XOR U11326 ( .A(n10880), .B(n10881), .Z(n10870) );
  ANDN U11327 ( .B(n10882), .A(n10883), .Z(n10880) );
  XOR U11328 ( .A(n10881), .B(n10884), .Z(n10882) );
  XOR U11329 ( .A(n10885), .B(n10886), .Z(n10869) );
  XOR U11330 ( .A(n10887), .B(n10888), .Z(n10886) );
  ANDN U11331 ( .B(n10889), .A(n10890), .Z(n10887) );
  XOR U11332 ( .A(n10891), .B(n10888), .Z(n10889) );
  IV U11333 ( .A(n10867), .Z(n10885) );
  XOR U11334 ( .A(n10892), .B(n10893), .Z(n10867) );
  ANDN U11335 ( .B(n10894), .A(n10895), .Z(n10892) );
  XOR U11336 ( .A(n10893), .B(n10896), .Z(n10894) );
  IV U11337 ( .A(n10875), .Z(n10879) );
  XOR U11338 ( .A(n10875), .B(n10857), .Z(n10877) );
  XOR U11339 ( .A(n10897), .B(n10898), .Z(n10857) );
  AND U11340 ( .A(n494), .B(n10899), .Z(n10897) );
  XOR U11341 ( .A(n10900), .B(n10898), .Z(n10899) );
  NANDN U11342 ( .A(n10859), .B(n10861), .Z(n10875) );
  XOR U11343 ( .A(n10901), .B(n10902), .Z(n10861) );
  AND U11344 ( .A(n494), .B(n10903), .Z(n10901) );
  XOR U11345 ( .A(n10902), .B(n10904), .Z(n10903) );
  XOR U11346 ( .A(n10905), .B(n10906), .Z(n494) );
  AND U11347 ( .A(n10907), .B(n10908), .Z(n10905) );
  XNOR U11348 ( .A(n10906), .B(n10872), .Z(n10908) );
  XNOR U11349 ( .A(n10909), .B(n10910), .Z(n10872) );
  ANDN U11350 ( .B(n10911), .A(n10912), .Z(n10909) );
  XOR U11351 ( .A(n10910), .B(n10913), .Z(n10911) );
  XOR U11352 ( .A(n10906), .B(n10874), .Z(n10907) );
  XOR U11353 ( .A(n10914), .B(n10915), .Z(n10874) );
  AND U11354 ( .A(n498), .B(n10916), .Z(n10914) );
  XOR U11355 ( .A(n10917), .B(n10915), .Z(n10916) );
  XNOR U11356 ( .A(n10918), .B(n10919), .Z(n10906) );
  NAND U11357 ( .A(n10920), .B(n10921), .Z(n10919) );
  XOR U11358 ( .A(n10922), .B(n10898), .Z(n10921) );
  XOR U11359 ( .A(n10912), .B(n10913), .Z(n10898) );
  XOR U11360 ( .A(n10923), .B(n10924), .Z(n10913) );
  ANDN U11361 ( .B(n10925), .A(n10926), .Z(n10923) );
  XOR U11362 ( .A(n10924), .B(n10927), .Z(n10925) );
  XOR U11363 ( .A(n10928), .B(n10929), .Z(n10912) );
  XOR U11364 ( .A(n10930), .B(n10931), .Z(n10929) );
  ANDN U11365 ( .B(n10932), .A(n10933), .Z(n10930) );
  XOR U11366 ( .A(n10934), .B(n10931), .Z(n10932) );
  IV U11367 ( .A(n10910), .Z(n10928) );
  XOR U11368 ( .A(n10935), .B(n10936), .Z(n10910) );
  ANDN U11369 ( .B(n10937), .A(n10938), .Z(n10935) );
  XOR U11370 ( .A(n10936), .B(n10939), .Z(n10937) );
  IV U11371 ( .A(n10918), .Z(n10922) );
  XOR U11372 ( .A(n10918), .B(n10900), .Z(n10920) );
  XOR U11373 ( .A(n10940), .B(n10941), .Z(n10900) );
  AND U11374 ( .A(n498), .B(n10942), .Z(n10940) );
  XOR U11375 ( .A(n10943), .B(n10941), .Z(n10942) );
  NANDN U11376 ( .A(n10902), .B(n10904), .Z(n10918) );
  XOR U11377 ( .A(n10944), .B(n10945), .Z(n10904) );
  AND U11378 ( .A(n498), .B(n10946), .Z(n10944) );
  XOR U11379 ( .A(n10945), .B(n10947), .Z(n10946) );
  XOR U11380 ( .A(n10948), .B(n10949), .Z(n498) );
  AND U11381 ( .A(n10950), .B(n10951), .Z(n10948) );
  XNOR U11382 ( .A(n10949), .B(n10915), .Z(n10951) );
  XNOR U11383 ( .A(n10952), .B(n10953), .Z(n10915) );
  ANDN U11384 ( .B(n10954), .A(n10955), .Z(n10952) );
  XOR U11385 ( .A(n10953), .B(n10956), .Z(n10954) );
  XOR U11386 ( .A(n10949), .B(n10917), .Z(n10950) );
  XOR U11387 ( .A(n10957), .B(n10958), .Z(n10917) );
  AND U11388 ( .A(n502), .B(n10959), .Z(n10957) );
  XOR U11389 ( .A(n10960), .B(n10958), .Z(n10959) );
  XNOR U11390 ( .A(n10961), .B(n10962), .Z(n10949) );
  NAND U11391 ( .A(n10963), .B(n10964), .Z(n10962) );
  XOR U11392 ( .A(n10965), .B(n10941), .Z(n10964) );
  XOR U11393 ( .A(n10955), .B(n10956), .Z(n10941) );
  XOR U11394 ( .A(n10966), .B(n10967), .Z(n10956) );
  ANDN U11395 ( .B(n10968), .A(n10969), .Z(n10966) );
  XOR U11396 ( .A(n10967), .B(n10970), .Z(n10968) );
  XOR U11397 ( .A(n10971), .B(n10972), .Z(n10955) );
  XOR U11398 ( .A(n10973), .B(n10974), .Z(n10972) );
  ANDN U11399 ( .B(n10975), .A(n10976), .Z(n10973) );
  XOR U11400 ( .A(n10977), .B(n10974), .Z(n10975) );
  IV U11401 ( .A(n10953), .Z(n10971) );
  XOR U11402 ( .A(n10978), .B(n10979), .Z(n10953) );
  ANDN U11403 ( .B(n10980), .A(n10981), .Z(n10978) );
  XOR U11404 ( .A(n10979), .B(n10982), .Z(n10980) );
  IV U11405 ( .A(n10961), .Z(n10965) );
  XOR U11406 ( .A(n10961), .B(n10943), .Z(n10963) );
  XOR U11407 ( .A(n10983), .B(n10984), .Z(n10943) );
  AND U11408 ( .A(n502), .B(n10985), .Z(n10983) );
  XOR U11409 ( .A(n10986), .B(n10984), .Z(n10985) );
  NANDN U11410 ( .A(n10945), .B(n10947), .Z(n10961) );
  XOR U11411 ( .A(n10987), .B(n10988), .Z(n10947) );
  AND U11412 ( .A(n502), .B(n10989), .Z(n10987) );
  XOR U11413 ( .A(n10988), .B(n10990), .Z(n10989) );
  XOR U11414 ( .A(n10991), .B(n10992), .Z(n502) );
  AND U11415 ( .A(n10993), .B(n10994), .Z(n10991) );
  XNOR U11416 ( .A(n10992), .B(n10958), .Z(n10994) );
  XNOR U11417 ( .A(n10995), .B(n10996), .Z(n10958) );
  ANDN U11418 ( .B(n10997), .A(n10998), .Z(n10995) );
  XOR U11419 ( .A(n10996), .B(n10999), .Z(n10997) );
  XOR U11420 ( .A(n10992), .B(n10960), .Z(n10993) );
  XOR U11421 ( .A(n11000), .B(n11001), .Z(n10960) );
  AND U11422 ( .A(n506), .B(n11002), .Z(n11000) );
  XOR U11423 ( .A(n11003), .B(n11001), .Z(n11002) );
  XNOR U11424 ( .A(n11004), .B(n11005), .Z(n10992) );
  NAND U11425 ( .A(n11006), .B(n11007), .Z(n11005) );
  XOR U11426 ( .A(n11008), .B(n10984), .Z(n11007) );
  XOR U11427 ( .A(n10998), .B(n10999), .Z(n10984) );
  XOR U11428 ( .A(n11009), .B(n11010), .Z(n10999) );
  ANDN U11429 ( .B(n11011), .A(n11012), .Z(n11009) );
  XOR U11430 ( .A(n11010), .B(n11013), .Z(n11011) );
  XOR U11431 ( .A(n11014), .B(n11015), .Z(n10998) );
  XOR U11432 ( .A(n11016), .B(n11017), .Z(n11015) );
  ANDN U11433 ( .B(n11018), .A(n11019), .Z(n11016) );
  XOR U11434 ( .A(n11020), .B(n11017), .Z(n11018) );
  IV U11435 ( .A(n10996), .Z(n11014) );
  XOR U11436 ( .A(n11021), .B(n11022), .Z(n10996) );
  ANDN U11437 ( .B(n11023), .A(n11024), .Z(n11021) );
  XOR U11438 ( .A(n11022), .B(n11025), .Z(n11023) );
  IV U11439 ( .A(n11004), .Z(n11008) );
  XOR U11440 ( .A(n11004), .B(n10986), .Z(n11006) );
  XOR U11441 ( .A(n11026), .B(n11027), .Z(n10986) );
  AND U11442 ( .A(n506), .B(n11028), .Z(n11026) );
  XOR U11443 ( .A(n11029), .B(n11027), .Z(n11028) );
  NANDN U11444 ( .A(n10988), .B(n10990), .Z(n11004) );
  XOR U11445 ( .A(n11030), .B(n11031), .Z(n10990) );
  AND U11446 ( .A(n506), .B(n11032), .Z(n11030) );
  XOR U11447 ( .A(n11031), .B(n11033), .Z(n11032) );
  XOR U11448 ( .A(n11034), .B(n11035), .Z(n506) );
  AND U11449 ( .A(n11036), .B(n11037), .Z(n11034) );
  XNOR U11450 ( .A(n11035), .B(n11001), .Z(n11037) );
  XNOR U11451 ( .A(n11038), .B(n11039), .Z(n11001) );
  ANDN U11452 ( .B(n11040), .A(n11041), .Z(n11038) );
  XOR U11453 ( .A(n11039), .B(n11042), .Z(n11040) );
  XOR U11454 ( .A(n11035), .B(n11003), .Z(n11036) );
  XOR U11455 ( .A(n11043), .B(n11044), .Z(n11003) );
  AND U11456 ( .A(n510), .B(n11045), .Z(n11043) );
  XOR U11457 ( .A(n11046), .B(n11044), .Z(n11045) );
  XNOR U11458 ( .A(n11047), .B(n11048), .Z(n11035) );
  NAND U11459 ( .A(n11049), .B(n11050), .Z(n11048) );
  XOR U11460 ( .A(n11051), .B(n11027), .Z(n11050) );
  XOR U11461 ( .A(n11041), .B(n11042), .Z(n11027) );
  XOR U11462 ( .A(n11052), .B(n11053), .Z(n11042) );
  ANDN U11463 ( .B(n11054), .A(n11055), .Z(n11052) );
  XOR U11464 ( .A(n11053), .B(n11056), .Z(n11054) );
  XOR U11465 ( .A(n11057), .B(n11058), .Z(n11041) );
  XOR U11466 ( .A(n11059), .B(n11060), .Z(n11058) );
  ANDN U11467 ( .B(n11061), .A(n11062), .Z(n11059) );
  XOR U11468 ( .A(n11063), .B(n11060), .Z(n11061) );
  IV U11469 ( .A(n11039), .Z(n11057) );
  XOR U11470 ( .A(n11064), .B(n11065), .Z(n11039) );
  ANDN U11471 ( .B(n11066), .A(n11067), .Z(n11064) );
  XOR U11472 ( .A(n11065), .B(n11068), .Z(n11066) );
  IV U11473 ( .A(n11047), .Z(n11051) );
  XOR U11474 ( .A(n11047), .B(n11029), .Z(n11049) );
  XOR U11475 ( .A(n11069), .B(n11070), .Z(n11029) );
  AND U11476 ( .A(n510), .B(n11071), .Z(n11069) );
  XOR U11477 ( .A(n11072), .B(n11070), .Z(n11071) );
  NANDN U11478 ( .A(n11031), .B(n11033), .Z(n11047) );
  XOR U11479 ( .A(n11073), .B(n11074), .Z(n11033) );
  AND U11480 ( .A(n510), .B(n11075), .Z(n11073) );
  XOR U11481 ( .A(n11074), .B(n11076), .Z(n11075) );
  XOR U11482 ( .A(n11077), .B(n11078), .Z(n510) );
  AND U11483 ( .A(n11079), .B(n11080), .Z(n11077) );
  XNOR U11484 ( .A(n11078), .B(n11044), .Z(n11080) );
  XNOR U11485 ( .A(n11081), .B(n11082), .Z(n11044) );
  ANDN U11486 ( .B(n11083), .A(n11084), .Z(n11081) );
  XOR U11487 ( .A(n11082), .B(n11085), .Z(n11083) );
  XOR U11488 ( .A(n11078), .B(n11046), .Z(n11079) );
  XOR U11489 ( .A(n11086), .B(n11087), .Z(n11046) );
  AND U11490 ( .A(n514), .B(n11088), .Z(n11086) );
  XOR U11491 ( .A(n11089), .B(n11087), .Z(n11088) );
  XNOR U11492 ( .A(n11090), .B(n11091), .Z(n11078) );
  NAND U11493 ( .A(n11092), .B(n11093), .Z(n11091) );
  XOR U11494 ( .A(n11094), .B(n11070), .Z(n11093) );
  XOR U11495 ( .A(n11084), .B(n11085), .Z(n11070) );
  XOR U11496 ( .A(n11095), .B(n11096), .Z(n11085) );
  ANDN U11497 ( .B(n11097), .A(n11098), .Z(n11095) );
  XOR U11498 ( .A(n11096), .B(n11099), .Z(n11097) );
  XOR U11499 ( .A(n11100), .B(n11101), .Z(n11084) );
  XOR U11500 ( .A(n11102), .B(n11103), .Z(n11101) );
  ANDN U11501 ( .B(n11104), .A(n11105), .Z(n11102) );
  XOR U11502 ( .A(n11106), .B(n11103), .Z(n11104) );
  IV U11503 ( .A(n11082), .Z(n11100) );
  XOR U11504 ( .A(n11107), .B(n11108), .Z(n11082) );
  ANDN U11505 ( .B(n11109), .A(n11110), .Z(n11107) );
  XOR U11506 ( .A(n11108), .B(n11111), .Z(n11109) );
  IV U11507 ( .A(n11090), .Z(n11094) );
  XOR U11508 ( .A(n11090), .B(n11072), .Z(n11092) );
  XOR U11509 ( .A(n11112), .B(n11113), .Z(n11072) );
  AND U11510 ( .A(n514), .B(n11114), .Z(n11112) );
  XOR U11511 ( .A(n11115), .B(n11113), .Z(n11114) );
  NANDN U11512 ( .A(n11074), .B(n11076), .Z(n11090) );
  XOR U11513 ( .A(n11116), .B(n11117), .Z(n11076) );
  AND U11514 ( .A(n514), .B(n11118), .Z(n11116) );
  XOR U11515 ( .A(n11117), .B(n11119), .Z(n11118) );
  XOR U11516 ( .A(n11120), .B(n11121), .Z(n514) );
  AND U11517 ( .A(n11122), .B(n11123), .Z(n11120) );
  XNOR U11518 ( .A(n11121), .B(n11087), .Z(n11123) );
  XNOR U11519 ( .A(n11124), .B(n11125), .Z(n11087) );
  ANDN U11520 ( .B(n11126), .A(n11127), .Z(n11124) );
  XOR U11521 ( .A(n11125), .B(n11128), .Z(n11126) );
  XOR U11522 ( .A(n11121), .B(n11089), .Z(n11122) );
  XOR U11523 ( .A(n11129), .B(n11130), .Z(n11089) );
  AND U11524 ( .A(n518), .B(n11131), .Z(n11129) );
  XOR U11525 ( .A(n11132), .B(n11130), .Z(n11131) );
  XNOR U11526 ( .A(n11133), .B(n11134), .Z(n11121) );
  NAND U11527 ( .A(n11135), .B(n11136), .Z(n11134) );
  XOR U11528 ( .A(n11137), .B(n11113), .Z(n11136) );
  XOR U11529 ( .A(n11127), .B(n11128), .Z(n11113) );
  XOR U11530 ( .A(n11138), .B(n11139), .Z(n11128) );
  ANDN U11531 ( .B(n11140), .A(n11141), .Z(n11138) );
  XOR U11532 ( .A(n11139), .B(n11142), .Z(n11140) );
  XOR U11533 ( .A(n11143), .B(n11144), .Z(n11127) );
  XOR U11534 ( .A(n11145), .B(n11146), .Z(n11144) );
  ANDN U11535 ( .B(n11147), .A(n11148), .Z(n11145) );
  XOR U11536 ( .A(n11149), .B(n11146), .Z(n11147) );
  IV U11537 ( .A(n11125), .Z(n11143) );
  XOR U11538 ( .A(n11150), .B(n11151), .Z(n11125) );
  ANDN U11539 ( .B(n11152), .A(n11153), .Z(n11150) );
  XOR U11540 ( .A(n11151), .B(n11154), .Z(n11152) );
  IV U11541 ( .A(n11133), .Z(n11137) );
  XOR U11542 ( .A(n11133), .B(n11115), .Z(n11135) );
  XOR U11543 ( .A(n11155), .B(n11156), .Z(n11115) );
  AND U11544 ( .A(n518), .B(n11157), .Z(n11155) );
  XOR U11545 ( .A(n11158), .B(n11156), .Z(n11157) );
  NANDN U11546 ( .A(n11117), .B(n11119), .Z(n11133) );
  XOR U11547 ( .A(n11159), .B(n11160), .Z(n11119) );
  AND U11548 ( .A(n518), .B(n11161), .Z(n11159) );
  XOR U11549 ( .A(n11160), .B(n11162), .Z(n11161) );
  XOR U11550 ( .A(n11163), .B(n11164), .Z(n518) );
  AND U11551 ( .A(n11165), .B(n11166), .Z(n11163) );
  XNOR U11552 ( .A(n11164), .B(n11130), .Z(n11166) );
  XNOR U11553 ( .A(n11167), .B(n11168), .Z(n11130) );
  ANDN U11554 ( .B(n11169), .A(n11170), .Z(n11167) );
  XOR U11555 ( .A(n11168), .B(n11171), .Z(n11169) );
  XOR U11556 ( .A(n11164), .B(n11132), .Z(n11165) );
  XOR U11557 ( .A(n11172), .B(n11173), .Z(n11132) );
  AND U11558 ( .A(n522), .B(n11174), .Z(n11172) );
  XOR U11559 ( .A(n11175), .B(n11173), .Z(n11174) );
  XNOR U11560 ( .A(n11176), .B(n11177), .Z(n11164) );
  NAND U11561 ( .A(n11178), .B(n11179), .Z(n11177) );
  XOR U11562 ( .A(n11180), .B(n11156), .Z(n11179) );
  XOR U11563 ( .A(n11170), .B(n11171), .Z(n11156) );
  XOR U11564 ( .A(n11181), .B(n11182), .Z(n11171) );
  ANDN U11565 ( .B(n11183), .A(n11184), .Z(n11181) );
  XOR U11566 ( .A(n11182), .B(n11185), .Z(n11183) );
  XOR U11567 ( .A(n11186), .B(n11187), .Z(n11170) );
  XOR U11568 ( .A(n11188), .B(n11189), .Z(n11187) );
  ANDN U11569 ( .B(n11190), .A(n11191), .Z(n11188) );
  XOR U11570 ( .A(n11192), .B(n11189), .Z(n11190) );
  IV U11571 ( .A(n11168), .Z(n11186) );
  XOR U11572 ( .A(n11193), .B(n11194), .Z(n11168) );
  ANDN U11573 ( .B(n11195), .A(n11196), .Z(n11193) );
  XOR U11574 ( .A(n11194), .B(n11197), .Z(n11195) );
  IV U11575 ( .A(n11176), .Z(n11180) );
  XOR U11576 ( .A(n11176), .B(n11158), .Z(n11178) );
  XOR U11577 ( .A(n11198), .B(n11199), .Z(n11158) );
  AND U11578 ( .A(n522), .B(n11200), .Z(n11198) );
  XOR U11579 ( .A(n11201), .B(n11199), .Z(n11200) );
  NANDN U11580 ( .A(n11160), .B(n11162), .Z(n11176) );
  XOR U11581 ( .A(n11202), .B(n11203), .Z(n11162) );
  AND U11582 ( .A(n522), .B(n11204), .Z(n11202) );
  XOR U11583 ( .A(n11203), .B(n11205), .Z(n11204) );
  XOR U11584 ( .A(n11206), .B(n11207), .Z(n522) );
  AND U11585 ( .A(n11208), .B(n11209), .Z(n11206) );
  XNOR U11586 ( .A(n11207), .B(n11173), .Z(n11209) );
  XNOR U11587 ( .A(n11210), .B(n11211), .Z(n11173) );
  ANDN U11588 ( .B(n11212), .A(n11213), .Z(n11210) );
  XOR U11589 ( .A(n11211), .B(n11214), .Z(n11212) );
  XOR U11590 ( .A(n11207), .B(n11175), .Z(n11208) );
  XOR U11591 ( .A(n11215), .B(n11216), .Z(n11175) );
  AND U11592 ( .A(n526), .B(n11217), .Z(n11215) );
  XOR U11593 ( .A(n11218), .B(n11216), .Z(n11217) );
  XNOR U11594 ( .A(n11219), .B(n11220), .Z(n11207) );
  NAND U11595 ( .A(n11221), .B(n11222), .Z(n11220) );
  XOR U11596 ( .A(n11223), .B(n11199), .Z(n11222) );
  XOR U11597 ( .A(n11213), .B(n11214), .Z(n11199) );
  XOR U11598 ( .A(n11224), .B(n11225), .Z(n11214) );
  ANDN U11599 ( .B(n11226), .A(n11227), .Z(n11224) );
  XOR U11600 ( .A(n11225), .B(n11228), .Z(n11226) );
  XOR U11601 ( .A(n11229), .B(n11230), .Z(n11213) );
  XOR U11602 ( .A(n11231), .B(n11232), .Z(n11230) );
  ANDN U11603 ( .B(n11233), .A(n11234), .Z(n11231) );
  XOR U11604 ( .A(n11235), .B(n11232), .Z(n11233) );
  IV U11605 ( .A(n11211), .Z(n11229) );
  XOR U11606 ( .A(n11236), .B(n11237), .Z(n11211) );
  ANDN U11607 ( .B(n11238), .A(n11239), .Z(n11236) );
  XOR U11608 ( .A(n11237), .B(n11240), .Z(n11238) );
  IV U11609 ( .A(n11219), .Z(n11223) );
  XOR U11610 ( .A(n11219), .B(n11201), .Z(n11221) );
  XOR U11611 ( .A(n11241), .B(n11242), .Z(n11201) );
  AND U11612 ( .A(n526), .B(n11243), .Z(n11241) );
  XOR U11613 ( .A(n11244), .B(n11242), .Z(n11243) );
  NANDN U11614 ( .A(n11203), .B(n11205), .Z(n11219) );
  XOR U11615 ( .A(n11245), .B(n11246), .Z(n11205) );
  AND U11616 ( .A(n526), .B(n11247), .Z(n11245) );
  XOR U11617 ( .A(n11246), .B(n11248), .Z(n11247) );
  XOR U11618 ( .A(n11249), .B(n11250), .Z(n526) );
  AND U11619 ( .A(n11251), .B(n11252), .Z(n11249) );
  XNOR U11620 ( .A(n11250), .B(n11216), .Z(n11252) );
  XNOR U11621 ( .A(n11253), .B(n11254), .Z(n11216) );
  ANDN U11622 ( .B(n11255), .A(n11256), .Z(n11253) );
  XOR U11623 ( .A(n11254), .B(n11257), .Z(n11255) );
  XOR U11624 ( .A(n11250), .B(n11218), .Z(n11251) );
  XOR U11625 ( .A(n11258), .B(n11259), .Z(n11218) );
  AND U11626 ( .A(n530), .B(n11260), .Z(n11258) );
  XOR U11627 ( .A(n11261), .B(n11259), .Z(n11260) );
  XNOR U11628 ( .A(n11262), .B(n11263), .Z(n11250) );
  NAND U11629 ( .A(n11264), .B(n11265), .Z(n11263) );
  XOR U11630 ( .A(n11266), .B(n11242), .Z(n11265) );
  XOR U11631 ( .A(n11256), .B(n11257), .Z(n11242) );
  XOR U11632 ( .A(n11267), .B(n11268), .Z(n11257) );
  ANDN U11633 ( .B(n11269), .A(n11270), .Z(n11267) );
  XOR U11634 ( .A(n11268), .B(n11271), .Z(n11269) );
  XOR U11635 ( .A(n11272), .B(n11273), .Z(n11256) );
  XOR U11636 ( .A(n11274), .B(n11275), .Z(n11273) );
  ANDN U11637 ( .B(n11276), .A(n11277), .Z(n11274) );
  XOR U11638 ( .A(n11278), .B(n11275), .Z(n11276) );
  IV U11639 ( .A(n11254), .Z(n11272) );
  XOR U11640 ( .A(n11279), .B(n11280), .Z(n11254) );
  ANDN U11641 ( .B(n11281), .A(n11282), .Z(n11279) );
  XOR U11642 ( .A(n11280), .B(n11283), .Z(n11281) );
  IV U11643 ( .A(n11262), .Z(n11266) );
  XOR U11644 ( .A(n11262), .B(n11244), .Z(n11264) );
  XOR U11645 ( .A(n11284), .B(n11285), .Z(n11244) );
  AND U11646 ( .A(n530), .B(n11286), .Z(n11284) );
  XOR U11647 ( .A(n11287), .B(n11285), .Z(n11286) );
  NANDN U11648 ( .A(n11246), .B(n11248), .Z(n11262) );
  XOR U11649 ( .A(n11288), .B(n11289), .Z(n11248) );
  AND U11650 ( .A(n530), .B(n11290), .Z(n11288) );
  XOR U11651 ( .A(n11289), .B(n11291), .Z(n11290) );
  XOR U11652 ( .A(n11292), .B(n11293), .Z(n530) );
  AND U11653 ( .A(n11294), .B(n11295), .Z(n11292) );
  XNOR U11654 ( .A(n11293), .B(n11259), .Z(n11295) );
  XNOR U11655 ( .A(n11296), .B(n11297), .Z(n11259) );
  ANDN U11656 ( .B(n11298), .A(n11299), .Z(n11296) );
  XOR U11657 ( .A(n11297), .B(n11300), .Z(n11298) );
  XOR U11658 ( .A(n11293), .B(n11261), .Z(n11294) );
  XOR U11659 ( .A(n11301), .B(n11302), .Z(n11261) );
  AND U11660 ( .A(n534), .B(n11303), .Z(n11301) );
  XOR U11661 ( .A(n11304), .B(n11302), .Z(n11303) );
  XNOR U11662 ( .A(n11305), .B(n11306), .Z(n11293) );
  NAND U11663 ( .A(n11307), .B(n11308), .Z(n11306) );
  XOR U11664 ( .A(n11309), .B(n11285), .Z(n11308) );
  XOR U11665 ( .A(n11299), .B(n11300), .Z(n11285) );
  XOR U11666 ( .A(n11310), .B(n11311), .Z(n11300) );
  ANDN U11667 ( .B(n11312), .A(n11313), .Z(n11310) );
  XOR U11668 ( .A(n11311), .B(n11314), .Z(n11312) );
  XOR U11669 ( .A(n11315), .B(n11316), .Z(n11299) );
  XOR U11670 ( .A(n11317), .B(n11318), .Z(n11316) );
  ANDN U11671 ( .B(n11319), .A(n11320), .Z(n11317) );
  XOR U11672 ( .A(n11321), .B(n11318), .Z(n11319) );
  IV U11673 ( .A(n11297), .Z(n11315) );
  XOR U11674 ( .A(n11322), .B(n11323), .Z(n11297) );
  ANDN U11675 ( .B(n11324), .A(n11325), .Z(n11322) );
  XOR U11676 ( .A(n11323), .B(n11326), .Z(n11324) );
  IV U11677 ( .A(n11305), .Z(n11309) );
  XOR U11678 ( .A(n11305), .B(n11287), .Z(n11307) );
  XOR U11679 ( .A(n11327), .B(n11328), .Z(n11287) );
  AND U11680 ( .A(n534), .B(n11329), .Z(n11327) );
  XOR U11681 ( .A(n11330), .B(n11328), .Z(n11329) );
  NANDN U11682 ( .A(n11289), .B(n11291), .Z(n11305) );
  XOR U11683 ( .A(n11331), .B(n11332), .Z(n11291) );
  AND U11684 ( .A(n534), .B(n11333), .Z(n11331) );
  XOR U11685 ( .A(n11332), .B(n11334), .Z(n11333) );
  XOR U11686 ( .A(n11335), .B(n11336), .Z(n534) );
  AND U11687 ( .A(n11337), .B(n11338), .Z(n11335) );
  XNOR U11688 ( .A(n11336), .B(n11302), .Z(n11338) );
  XNOR U11689 ( .A(n11339), .B(n11340), .Z(n11302) );
  ANDN U11690 ( .B(n11341), .A(n11342), .Z(n11339) );
  XOR U11691 ( .A(n11340), .B(n11343), .Z(n11341) );
  XOR U11692 ( .A(n11336), .B(n11304), .Z(n11337) );
  XOR U11693 ( .A(n11344), .B(n11345), .Z(n11304) );
  AND U11694 ( .A(n538), .B(n11346), .Z(n11344) );
  XOR U11695 ( .A(n11347), .B(n11345), .Z(n11346) );
  XNOR U11696 ( .A(n11348), .B(n11349), .Z(n11336) );
  NAND U11697 ( .A(n11350), .B(n11351), .Z(n11349) );
  XOR U11698 ( .A(n11352), .B(n11328), .Z(n11351) );
  XOR U11699 ( .A(n11342), .B(n11343), .Z(n11328) );
  XOR U11700 ( .A(n11353), .B(n11354), .Z(n11343) );
  ANDN U11701 ( .B(n11355), .A(n11356), .Z(n11353) );
  XOR U11702 ( .A(n11354), .B(n11357), .Z(n11355) );
  XOR U11703 ( .A(n11358), .B(n11359), .Z(n11342) );
  XOR U11704 ( .A(n11360), .B(n11361), .Z(n11359) );
  ANDN U11705 ( .B(n11362), .A(n11363), .Z(n11360) );
  XOR U11706 ( .A(n11364), .B(n11361), .Z(n11362) );
  IV U11707 ( .A(n11340), .Z(n11358) );
  XOR U11708 ( .A(n11365), .B(n11366), .Z(n11340) );
  ANDN U11709 ( .B(n11367), .A(n11368), .Z(n11365) );
  XOR U11710 ( .A(n11366), .B(n11369), .Z(n11367) );
  IV U11711 ( .A(n11348), .Z(n11352) );
  XOR U11712 ( .A(n11348), .B(n11330), .Z(n11350) );
  XOR U11713 ( .A(n11370), .B(n11371), .Z(n11330) );
  AND U11714 ( .A(n538), .B(n11372), .Z(n11370) );
  XOR U11715 ( .A(n11373), .B(n11371), .Z(n11372) );
  NANDN U11716 ( .A(n11332), .B(n11334), .Z(n11348) );
  XOR U11717 ( .A(n11374), .B(n11375), .Z(n11334) );
  AND U11718 ( .A(n538), .B(n11376), .Z(n11374) );
  XOR U11719 ( .A(n11375), .B(n11377), .Z(n11376) );
  XOR U11720 ( .A(n11378), .B(n11379), .Z(n538) );
  AND U11721 ( .A(n11380), .B(n11381), .Z(n11378) );
  XNOR U11722 ( .A(n11379), .B(n11345), .Z(n11381) );
  XNOR U11723 ( .A(n11382), .B(n11383), .Z(n11345) );
  ANDN U11724 ( .B(n11384), .A(n11385), .Z(n11382) );
  XOR U11725 ( .A(n11383), .B(n11386), .Z(n11384) );
  XOR U11726 ( .A(n11379), .B(n11347), .Z(n11380) );
  XOR U11727 ( .A(n11387), .B(n11388), .Z(n11347) );
  AND U11728 ( .A(n542), .B(n11389), .Z(n11387) );
  XOR U11729 ( .A(n11390), .B(n11388), .Z(n11389) );
  XNOR U11730 ( .A(n11391), .B(n11392), .Z(n11379) );
  NAND U11731 ( .A(n11393), .B(n11394), .Z(n11392) );
  XOR U11732 ( .A(n11395), .B(n11371), .Z(n11394) );
  XOR U11733 ( .A(n11385), .B(n11386), .Z(n11371) );
  XOR U11734 ( .A(n11396), .B(n11397), .Z(n11386) );
  ANDN U11735 ( .B(n11398), .A(n11399), .Z(n11396) );
  XOR U11736 ( .A(n11397), .B(n11400), .Z(n11398) );
  XOR U11737 ( .A(n11401), .B(n11402), .Z(n11385) );
  XOR U11738 ( .A(n11403), .B(n11404), .Z(n11402) );
  ANDN U11739 ( .B(n11405), .A(n11406), .Z(n11403) );
  XOR U11740 ( .A(n11407), .B(n11404), .Z(n11405) );
  IV U11741 ( .A(n11383), .Z(n11401) );
  XOR U11742 ( .A(n11408), .B(n11409), .Z(n11383) );
  ANDN U11743 ( .B(n11410), .A(n11411), .Z(n11408) );
  XOR U11744 ( .A(n11409), .B(n11412), .Z(n11410) );
  IV U11745 ( .A(n11391), .Z(n11395) );
  XOR U11746 ( .A(n11391), .B(n11373), .Z(n11393) );
  XOR U11747 ( .A(n11413), .B(n11414), .Z(n11373) );
  AND U11748 ( .A(n542), .B(n11415), .Z(n11413) );
  XOR U11749 ( .A(n11416), .B(n11414), .Z(n11415) );
  NANDN U11750 ( .A(n11375), .B(n11377), .Z(n11391) );
  XOR U11751 ( .A(n11417), .B(n11418), .Z(n11377) );
  AND U11752 ( .A(n542), .B(n11419), .Z(n11417) );
  XOR U11753 ( .A(n11418), .B(n11420), .Z(n11419) );
  XOR U11754 ( .A(n11421), .B(n11422), .Z(n542) );
  AND U11755 ( .A(n11423), .B(n11424), .Z(n11421) );
  XNOR U11756 ( .A(n11422), .B(n11388), .Z(n11424) );
  XNOR U11757 ( .A(n11425), .B(n11426), .Z(n11388) );
  ANDN U11758 ( .B(n11427), .A(n11428), .Z(n11425) );
  XOR U11759 ( .A(n11426), .B(n11429), .Z(n11427) );
  XOR U11760 ( .A(n11422), .B(n11390), .Z(n11423) );
  XOR U11761 ( .A(n11430), .B(n11431), .Z(n11390) );
  AND U11762 ( .A(n546), .B(n11432), .Z(n11430) );
  XOR U11763 ( .A(n11433), .B(n11431), .Z(n11432) );
  XNOR U11764 ( .A(n11434), .B(n11435), .Z(n11422) );
  NAND U11765 ( .A(n11436), .B(n11437), .Z(n11435) );
  XOR U11766 ( .A(n11438), .B(n11414), .Z(n11437) );
  XOR U11767 ( .A(n11428), .B(n11429), .Z(n11414) );
  XOR U11768 ( .A(n11439), .B(n11440), .Z(n11429) );
  ANDN U11769 ( .B(n11441), .A(n11442), .Z(n11439) );
  XOR U11770 ( .A(n11440), .B(n11443), .Z(n11441) );
  XOR U11771 ( .A(n11444), .B(n11445), .Z(n11428) );
  XOR U11772 ( .A(n11446), .B(n11447), .Z(n11445) );
  ANDN U11773 ( .B(n11448), .A(n11449), .Z(n11446) );
  XOR U11774 ( .A(n11450), .B(n11447), .Z(n11448) );
  IV U11775 ( .A(n11426), .Z(n11444) );
  XOR U11776 ( .A(n11451), .B(n11452), .Z(n11426) );
  ANDN U11777 ( .B(n11453), .A(n11454), .Z(n11451) );
  XOR U11778 ( .A(n11452), .B(n11455), .Z(n11453) );
  IV U11779 ( .A(n11434), .Z(n11438) );
  XOR U11780 ( .A(n11434), .B(n11416), .Z(n11436) );
  XOR U11781 ( .A(n11456), .B(n11457), .Z(n11416) );
  AND U11782 ( .A(n546), .B(n11458), .Z(n11456) );
  XOR U11783 ( .A(n11459), .B(n11457), .Z(n11458) );
  NANDN U11784 ( .A(n11418), .B(n11420), .Z(n11434) );
  XOR U11785 ( .A(n11460), .B(n11461), .Z(n11420) );
  AND U11786 ( .A(n546), .B(n11462), .Z(n11460) );
  XOR U11787 ( .A(n11461), .B(n11463), .Z(n11462) );
  XOR U11788 ( .A(n11464), .B(n11465), .Z(n546) );
  AND U11789 ( .A(n11466), .B(n11467), .Z(n11464) );
  XNOR U11790 ( .A(n11465), .B(n11431), .Z(n11467) );
  XNOR U11791 ( .A(n11468), .B(n11469), .Z(n11431) );
  ANDN U11792 ( .B(n11470), .A(n11471), .Z(n11468) );
  XOR U11793 ( .A(n11469), .B(n11472), .Z(n11470) );
  XOR U11794 ( .A(n11465), .B(n11433), .Z(n11466) );
  XOR U11795 ( .A(n11473), .B(n11474), .Z(n11433) );
  AND U11796 ( .A(n550), .B(n11475), .Z(n11473) );
  XOR U11797 ( .A(n11476), .B(n11474), .Z(n11475) );
  XNOR U11798 ( .A(n11477), .B(n11478), .Z(n11465) );
  NAND U11799 ( .A(n11479), .B(n11480), .Z(n11478) );
  XOR U11800 ( .A(n11481), .B(n11457), .Z(n11480) );
  XOR U11801 ( .A(n11471), .B(n11472), .Z(n11457) );
  XOR U11802 ( .A(n11482), .B(n11483), .Z(n11472) );
  ANDN U11803 ( .B(n11484), .A(n11485), .Z(n11482) );
  XOR U11804 ( .A(n11483), .B(n11486), .Z(n11484) );
  XOR U11805 ( .A(n11487), .B(n11488), .Z(n11471) );
  XOR U11806 ( .A(n11489), .B(n11490), .Z(n11488) );
  ANDN U11807 ( .B(n11491), .A(n11492), .Z(n11489) );
  XOR U11808 ( .A(n11493), .B(n11490), .Z(n11491) );
  IV U11809 ( .A(n11469), .Z(n11487) );
  XOR U11810 ( .A(n11494), .B(n11495), .Z(n11469) );
  ANDN U11811 ( .B(n11496), .A(n11497), .Z(n11494) );
  XOR U11812 ( .A(n11495), .B(n11498), .Z(n11496) );
  IV U11813 ( .A(n11477), .Z(n11481) );
  XOR U11814 ( .A(n11477), .B(n11459), .Z(n11479) );
  XOR U11815 ( .A(n11499), .B(n11500), .Z(n11459) );
  AND U11816 ( .A(n550), .B(n11501), .Z(n11499) );
  XOR U11817 ( .A(n11502), .B(n11500), .Z(n11501) );
  NANDN U11818 ( .A(n11461), .B(n11463), .Z(n11477) );
  XOR U11819 ( .A(n11503), .B(n11504), .Z(n11463) );
  AND U11820 ( .A(n550), .B(n11505), .Z(n11503) );
  XOR U11821 ( .A(n11504), .B(n11506), .Z(n11505) );
  XOR U11822 ( .A(n11507), .B(n11508), .Z(n550) );
  AND U11823 ( .A(n11509), .B(n11510), .Z(n11507) );
  XNOR U11824 ( .A(n11508), .B(n11474), .Z(n11510) );
  XNOR U11825 ( .A(n11511), .B(n11512), .Z(n11474) );
  ANDN U11826 ( .B(n11513), .A(n11514), .Z(n11511) );
  XOR U11827 ( .A(n11512), .B(n11515), .Z(n11513) );
  XOR U11828 ( .A(n11508), .B(n11476), .Z(n11509) );
  XOR U11829 ( .A(n11516), .B(n11517), .Z(n11476) );
  AND U11830 ( .A(n554), .B(n11518), .Z(n11516) );
  XOR U11831 ( .A(n11519), .B(n11517), .Z(n11518) );
  XNOR U11832 ( .A(n11520), .B(n11521), .Z(n11508) );
  NAND U11833 ( .A(n11522), .B(n11523), .Z(n11521) );
  XOR U11834 ( .A(n11524), .B(n11500), .Z(n11523) );
  XOR U11835 ( .A(n11514), .B(n11515), .Z(n11500) );
  XOR U11836 ( .A(n11525), .B(n11526), .Z(n11515) );
  ANDN U11837 ( .B(n11527), .A(n11528), .Z(n11525) );
  XOR U11838 ( .A(n11526), .B(n11529), .Z(n11527) );
  XOR U11839 ( .A(n11530), .B(n11531), .Z(n11514) );
  XOR U11840 ( .A(n11532), .B(n11533), .Z(n11531) );
  ANDN U11841 ( .B(n11534), .A(n11535), .Z(n11532) );
  XOR U11842 ( .A(n11536), .B(n11533), .Z(n11534) );
  IV U11843 ( .A(n11512), .Z(n11530) );
  XOR U11844 ( .A(n11537), .B(n11538), .Z(n11512) );
  ANDN U11845 ( .B(n11539), .A(n11540), .Z(n11537) );
  XOR U11846 ( .A(n11538), .B(n11541), .Z(n11539) );
  IV U11847 ( .A(n11520), .Z(n11524) );
  XOR U11848 ( .A(n11520), .B(n11502), .Z(n11522) );
  XOR U11849 ( .A(n11542), .B(n11543), .Z(n11502) );
  AND U11850 ( .A(n554), .B(n11544), .Z(n11542) );
  XOR U11851 ( .A(n11545), .B(n11543), .Z(n11544) );
  NANDN U11852 ( .A(n11504), .B(n11506), .Z(n11520) );
  XOR U11853 ( .A(n11546), .B(n11547), .Z(n11506) );
  AND U11854 ( .A(n554), .B(n11548), .Z(n11546) );
  XOR U11855 ( .A(n11547), .B(n11549), .Z(n11548) );
  XOR U11856 ( .A(n11550), .B(n11551), .Z(n554) );
  AND U11857 ( .A(n11552), .B(n11553), .Z(n11550) );
  XNOR U11858 ( .A(n11551), .B(n11517), .Z(n11553) );
  XNOR U11859 ( .A(n11554), .B(n11555), .Z(n11517) );
  ANDN U11860 ( .B(n11556), .A(n11557), .Z(n11554) );
  XOR U11861 ( .A(n11555), .B(n11558), .Z(n11556) );
  XOR U11862 ( .A(n11551), .B(n11519), .Z(n11552) );
  XOR U11863 ( .A(n11559), .B(n11560), .Z(n11519) );
  AND U11864 ( .A(n558), .B(n11561), .Z(n11559) );
  XOR U11865 ( .A(n11562), .B(n11560), .Z(n11561) );
  XNOR U11866 ( .A(n11563), .B(n11564), .Z(n11551) );
  NAND U11867 ( .A(n11565), .B(n11566), .Z(n11564) );
  XOR U11868 ( .A(n11567), .B(n11543), .Z(n11566) );
  XOR U11869 ( .A(n11557), .B(n11558), .Z(n11543) );
  XOR U11870 ( .A(n11568), .B(n11569), .Z(n11558) );
  ANDN U11871 ( .B(n11570), .A(n11571), .Z(n11568) );
  XOR U11872 ( .A(n11569), .B(n11572), .Z(n11570) );
  XOR U11873 ( .A(n11573), .B(n11574), .Z(n11557) );
  XOR U11874 ( .A(n11575), .B(n11576), .Z(n11574) );
  ANDN U11875 ( .B(n11577), .A(n11578), .Z(n11575) );
  XOR U11876 ( .A(n11579), .B(n11576), .Z(n11577) );
  IV U11877 ( .A(n11555), .Z(n11573) );
  XOR U11878 ( .A(n11580), .B(n11581), .Z(n11555) );
  ANDN U11879 ( .B(n11582), .A(n11583), .Z(n11580) );
  XOR U11880 ( .A(n11581), .B(n11584), .Z(n11582) );
  IV U11881 ( .A(n11563), .Z(n11567) );
  XOR U11882 ( .A(n11563), .B(n11545), .Z(n11565) );
  XOR U11883 ( .A(n11585), .B(n11586), .Z(n11545) );
  AND U11884 ( .A(n558), .B(n11587), .Z(n11585) );
  XOR U11885 ( .A(n11588), .B(n11586), .Z(n11587) );
  NANDN U11886 ( .A(n11547), .B(n11549), .Z(n11563) );
  XOR U11887 ( .A(n11589), .B(n11590), .Z(n11549) );
  AND U11888 ( .A(n558), .B(n11591), .Z(n11589) );
  XOR U11889 ( .A(n11590), .B(n11592), .Z(n11591) );
  XOR U11890 ( .A(n11593), .B(n11594), .Z(n558) );
  AND U11891 ( .A(n11595), .B(n11596), .Z(n11593) );
  XNOR U11892 ( .A(n11594), .B(n11560), .Z(n11596) );
  XNOR U11893 ( .A(n11597), .B(n11598), .Z(n11560) );
  ANDN U11894 ( .B(n11599), .A(n11600), .Z(n11597) );
  XOR U11895 ( .A(n11598), .B(n11601), .Z(n11599) );
  XOR U11896 ( .A(n11594), .B(n11562), .Z(n11595) );
  XOR U11897 ( .A(n11602), .B(n11603), .Z(n11562) );
  AND U11898 ( .A(n562), .B(n11604), .Z(n11602) );
  XOR U11899 ( .A(n11605), .B(n11603), .Z(n11604) );
  XNOR U11900 ( .A(n11606), .B(n11607), .Z(n11594) );
  NAND U11901 ( .A(n11608), .B(n11609), .Z(n11607) );
  XOR U11902 ( .A(n11610), .B(n11586), .Z(n11609) );
  XOR U11903 ( .A(n11600), .B(n11601), .Z(n11586) );
  XOR U11904 ( .A(n11611), .B(n11612), .Z(n11601) );
  ANDN U11905 ( .B(n11613), .A(n11614), .Z(n11611) );
  XOR U11906 ( .A(n11612), .B(n11615), .Z(n11613) );
  XOR U11907 ( .A(n11616), .B(n11617), .Z(n11600) );
  XOR U11908 ( .A(n11618), .B(n11619), .Z(n11617) );
  ANDN U11909 ( .B(n11620), .A(n11621), .Z(n11618) );
  XOR U11910 ( .A(n11622), .B(n11619), .Z(n11620) );
  IV U11911 ( .A(n11598), .Z(n11616) );
  XOR U11912 ( .A(n11623), .B(n11624), .Z(n11598) );
  ANDN U11913 ( .B(n11625), .A(n11626), .Z(n11623) );
  XOR U11914 ( .A(n11624), .B(n11627), .Z(n11625) );
  IV U11915 ( .A(n11606), .Z(n11610) );
  XOR U11916 ( .A(n11606), .B(n11588), .Z(n11608) );
  XOR U11917 ( .A(n11628), .B(n11629), .Z(n11588) );
  AND U11918 ( .A(n562), .B(n11630), .Z(n11628) );
  XOR U11919 ( .A(n11631), .B(n11629), .Z(n11630) );
  NANDN U11920 ( .A(n11590), .B(n11592), .Z(n11606) );
  XOR U11921 ( .A(n11632), .B(n11633), .Z(n11592) );
  AND U11922 ( .A(n562), .B(n11634), .Z(n11632) );
  XOR U11923 ( .A(n11633), .B(n11635), .Z(n11634) );
  XOR U11924 ( .A(n11636), .B(n11637), .Z(n562) );
  AND U11925 ( .A(n11638), .B(n11639), .Z(n11636) );
  XNOR U11926 ( .A(n11637), .B(n11603), .Z(n11639) );
  XNOR U11927 ( .A(n11640), .B(n11641), .Z(n11603) );
  ANDN U11928 ( .B(n11642), .A(n11643), .Z(n11640) );
  XOR U11929 ( .A(n11641), .B(n11644), .Z(n11642) );
  XOR U11930 ( .A(n11637), .B(n11605), .Z(n11638) );
  XOR U11931 ( .A(n11645), .B(n11646), .Z(n11605) );
  AND U11932 ( .A(n566), .B(n11647), .Z(n11645) );
  XOR U11933 ( .A(n11648), .B(n11646), .Z(n11647) );
  XNOR U11934 ( .A(n11649), .B(n11650), .Z(n11637) );
  NAND U11935 ( .A(n11651), .B(n11652), .Z(n11650) );
  XOR U11936 ( .A(n11653), .B(n11629), .Z(n11652) );
  XOR U11937 ( .A(n11643), .B(n11644), .Z(n11629) );
  XOR U11938 ( .A(n11654), .B(n11655), .Z(n11644) );
  ANDN U11939 ( .B(n11656), .A(n11657), .Z(n11654) );
  XOR U11940 ( .A(n11655), .B(n11658), .Z(n11656) );
  XOR U11941 ( .A(n11659), .B(n11660), .Z(n11643) );
  XOR U11942 ( .A(n11661), .B(n11662), .Z(n11660) );
  ANDN U11943 ( .B(n11663), .A(n11664), .Z(n11661) );
  XOR U11944 ( .A(n11665), .B(n11662), .Z(n11663) );
  IV U11945 ( .A(n11641), .Z(n11659) );
  XOR U11946 ( .A(n11666), .B(n11667), .Z(n11641) );
  ANDN U11947 ( .B(n11668), .A(n11669), .Z(n11666) );
  XOR U11948 ( .A(n11667), .B(n11670), .Z(n11668) );
  IV U11949 ( .A(n11649), .Z(n11653) );
  XOR U11950 ( .A(n11649), .B(n11631), .Z(n11651) );
  XOR U11951 ( .A(n11671), .B(n11672), .Z(n11631) );
  AND U11952 ( .A(n566), .B(n11673), .Z(n11671) );
  XOR U11953 ( .A(n11674), .B(n11672), .Z(n11673) );
  NANDN U11954 ( .A(n11633), .B(n11635), .Z(n11649) );
  XOR U11955 ( .A(n11675), .B(n11676), .Z(n11635) );
  AND U11956 ( .A(n566), .B(n11677), .Z(n11675) );
  XOR U11957 ( .A(n11676), .B(n11678), .Z(n11677) );
  XOR U11958 ( .A(n11679), .B(n11680), .Z(n566) );
  AND U11959 ( .A(n11681), .B(n11682), .Z(n11679) );
  XNOR U11960 ( .A(n11680), .B(n11646), .Z(n11682) );
  XNOR U11961 ( .A(n11683), .B(n11684), .Z(n11646) );
  ANDN U11962 ( .B(n11685), .A(n11686), .Z(n11683) );
  XOR U11963 ( .A(n11684), .B(n11687), .Z(n11685) );
  XOR U11964 ( .A(n11680), .B(n11648), .Z(n11681) );
  XOR U11965 ( .A(n11688), .B(n11689), .Z(n11648) );
  AND U11966 ( .A(n570), .B(n11690), .Z(n11688) );
  XOR U11967 ( .A(n11691), .B(n11689), .Z(n11690) );
  XNOR U11968 ( .A(n11692), .B(n11693), .Z(n11680) );
  NAND U11969 ( .A(n11694), .B(n11695), .Z(n11693) );
  XOR U11970 ( .A(n11696), .B(n11672), .Z(n11695) );
  XOR U11971 ( .A(n11686), .B(n11687), .Z(n11672) );
  XOR U11972 ( .A(n11697), .B(n11698), .Z(n11687) );
  ANDN U11973 ( .B(n11699), .A(n11700), .Z(n11697) );
  XOR U11974 ( .A(n11698), .B(n11701), .Z(n11699) );
  XOR U11975 ( .A(n11702), .B(n11703), .Z(n11686) );
  XOR U11976 ( .A(n11704), .B(n11705), .Z(n11703) );
  ANDN U11977 ( .B(n11706), .A(n11707), .Z(n11704) );
  XOR U11978 ( .A(n11708), .B(n11705), .Z(n11706) );
  IV U11979 ( .A(n11684), .Z(n11702) );
  XOR U11980 ( .A(n11709), .B(n11710), .Z(n11684) );
  ANDN U11981 ( .B(n11711), .A(n11712), .Z(n11709) );
  XOR U11982 ( .A(n11710), .B(n11713), .Z(n11711) );
  IV U11983 ( .A(n11692), .Z(n11696) );
  XOR U11984 ( .A(n11692), .B(n11674), .Z(n11694) );
  XOR U11985 ( .A(n11714), .B(n11715), .Z(n11674) );
  AND U11986 ( .A(n570), .B(n11716), .Z(n11714) );
  XOR U11987 ( .A(n11717), .B(n11715), .Z(n11716) );
  NANDN U11988 ( .A(n11676), .B(n11678), .Z(n11692) );
  XOR U11989 ( .A(n11718), .B(n11719), .Z(n11678) );
  AND U11990 ( .A(n570), .B(n11720), .Z(n11718) );
  XOR U11991 ( .A(n11719), .B(n11721), .Z(n11720) );
  XOR U11992 ( .A(n11722), .B(n11723), .Z(n570) );
  AND U11993 ( .A(n11724), .B(n11725), .Z(n11722) );
  XNOR U11994 ( .A(n11723), .B(n11689), .Z(n11725) );
  XNOR U11995 ( .A(n11726), .B(n11727), .Z(n11689) );
  ANDN U11996 ( .B(n11728), .A(n11729), .Z(n11726) );
  XOR U11997 ( .A(n11727), .B(n11730), .Z(n11728) );
  XOR U11998 ( .A(n11723), .B(n11691), .Z(n11724) );
  XOR U11999 ( .A(n11731), .B(n11732), .Z(n11691) );
  AND U12000 ( .A(n574), .B(n11733), .Z(n11731) );
  XOR U12001 ( .A(n11734), .B(n11732), .Z(n11733) );
  XNOR U12002 ( .A(n11735), .B(n11736), .Z(n11723) );
  NAND U12003 ( .A(n11737), .B(n11738), .Z(n11736) );
  XOR U12004 ( .A(n11739), .B(n11715), .Z(n11738) );
  XOR U12005 ( .A(n11729), .B(n11730), .Z(n11715) );
  XOR U12006 ( .A(n11740), .B(n11741), .Z(n11730) );
  ANDN U12007 ( .B(n11742), .A(n11743), .Z(n11740) );
  XOR U12008 ( .A(n11741), .B(n11744), .Z(n11742) );
  XOR U12009 ( .A(n11745), .B(n11746), .Z(n11729) );
  XOR U12010 ( .A(n11747), .B(n11748), .Z(n11746) );
  ANDN U12011 ( .B(n11749), .A(n11750), .Z(n11747) );
  XOR U12012 ( .A(n11751), .B(n11748), .Z(n11749) );
  IV U12013 ( .A(n11727), .Z(n11745) );
  XOR U12014 ( .A(n11752), .B(n11753), .Z(n11727) );
  ANDN U12015 ( .B(n11754), .A(n11755), .Z(n11752) );
  XOR U12016 ( .A(n11753), .B(n11756), .Z(n11754) );
  IV U12017 ( .A(n11735), .Z(n11739) );
  XOR U12018 ( .A(n11735), .B(n11717), .Z(n11737) );
  XOR U12019 ( .A(n11757), .B(n11758), .Z(n11717) );
  AND U12020 ( .A(n574), .B(n11759), .Z(n11757) );
  XOR U12021 ( .A(n11760), .B(n11758), .Z(n11759) );
  NANDN U12022 ( .A(n11719), .B(n11721), .Z(n11735) );
  XOR U12023 ( .A(n11761), .B(n11762), .Z(n11721) );
  AND U12024 ( .A(n574), .B(n11763), .Z(n11761) );
  XOR U12025 ( .A(n11762), .B(n11764), .Z(n11763) );
  XOR U12026 ( .A(n11765), .B(n11766), .Z(n574) );
  AND U12027 ( .A(n11767), .B(n11768), .Z(n11765) );
  XNOR U12028 ( .A(n11766), .B(n11732), .Z(n11768) );
  XNOR U12029 ( .A(n11769), .B(n11770), .Z(n11732) );
  ANDN U12030 ( .B(n11771), .A(n11772), .Z(n11769) );
  XOR U12031 ( .A(n11770), .B(n11773), .Z(n11771) );
  XOR U12032 ( .A(n11766), .B(n11734), .Z(n11767) );
  XOR U12033 ( .A(n11774), .B(n11775), .Z(n11734) );
  AND U12034 ( .A(n578), .B(n11776), .Z(n11774) );
  XOR U12035 ( .A(n11777), .B(n11775), .Z(n11776) );
  XNOR U12036 ( .A(n11778), .B(n11779), .Z(n11766) );
  NAND U12037 ( .A(n11780), .B(n11781), .Z(n11779) );
  XOR U12038 ( .A(n11782), .B(n11758), .Z(n11781) );
  XOR U12039 ( .A(n11772), .B(n11773), .Z(n11758) );
  XOR U12040 ( .A(n11783), .B(n11784), .Z(n11773) );
  ANDN U12041 ( .B(n11785), .A(n11786), .Z(n11783) );
  XOR U12042 ( .A(n11784), .B(n11787), .Z(n11785) );
  XOR U12043 ( .A(n11788), .B(n11789), .Z(n11772) );
  XOR U12044 ( .A(n11790), .B(n11791), .Z(n11789) );
  ANDN U12045 ( .B(n11792), .A(n11793), .Z(n11790) );
  XOR U12046 ( .A(n11794), .B(n11791), .Z(n11792) );
  IV U12047 ( .A(n11770), .Z(n11788) );
  XOR U12048 ( .A(n11795), .B(n11796), .Z(n11770) );
  ANDN U12049 ( .B(n11797), .A(n11798), .Z(n11795) );
  XOR U12050 ( .A(n11796), .B(n11799), .Z(n11797) );
  IV U12051 ( .A(n11778), .Z(n11782) );
  XOR U12052 ( .A(n11778), .B(n11760), .Z(n11780) );
  XOR U12053 ( .A(n11800), .B(n11801), .Z(n11760) );
  AND U12054 ( .A(n578), .B(n11802), .Z(n11800) );
  XOR U12055 ( .A(n11803), .B(n11801), .Z(n11802) );
  NANDN U12056 ( .A(n11762), .B(n11764), .Z(n11778) );
  XOR U12057 ( .A(n11804), .B(n11805), .Z(n11764) );
  AND U12058 ( .A(n578), .B(n11806), .Z(n11804) );
  XOR U12059 ( .A(n11805), .B(n11807), .Z(n11806) );
  XOR U12060 ( .A(n11808), .B(n11809), .Z(n578) );
  AND U12061 ( .A(n11810), .B(n11811), .Z(n11808) );
  XNOR U12062 ( .A(n11809), .B(n11775), .Z(n11811) );
  XNOR U12063 ( .A(n11812), .B(n11813), .Z(n11775) );
  ANDN U12064 ( .B(n11814), .A(n11815), .Z(n11812) );
  XOR U12065 ( .A(n11813), .B(n11816), .Z(n11814) );
  XOR U12066 ( .A(n11809), .B(n11777), .Z(n11810) );
  XOR U12067 ( .A(n11817), .B(n11818), .Z(n11777) );
  AND U12068 ( .A(n582), .B(n11819), .Z(n11817) );
  XOR U12069 ( .A(n11820), .B(n11818), .Z(n11819) );
  XNOR U12070 ( .A(n11821), .B(n11822), .Z(n11809) );
  NAND U12071 ( .A(n11823), .B(n11824), .Z(n11822) );
  XOR U12072 ( .A(n11825), .B(n11801), .Z(n11824) );
  XOR U12073 ( .A(n11815), .B(n11816), .Z(n11801) );
  XOR U12074 ( .A(n11826), .B(n11827), .Z(n11816) );
  ANDN U12075 ( .B(n11828), .A(n11829), .Z(n11826) );
  XOR U12076 ( .A(n11827), .B(n11830), .Z(n11828) );
  XOR U12077 ( .A(n11831), .B(n11832), .Z(n11815) );
  XOR U12078 ( .A(n11833), .B(n11834), .Z(n11832) );
  ANDN U12079 ( .B(n11835), .A(n11836), .Z(n11833) );
  XOR U12080 ( .A(n11837), .B(n11834), .Z(n11835) );
  IV U12081 ( .A(n11813), .Z(n11831) );
  XOR U12082 ( .A(n11838), .B(n11839), .Z(n11813) );
  ANDN U12083 ( .B(n11840), .A(n11841), .Z(n11838) );
  XOR U12084 ( .A(n11839), .B(n11842), .Z(n11840) );
  IV U12085 ( .A(n11821), .Z(n11825) );
  XOR U12086 ( .A(n11821), .B(n11803), .Z(n11823) );
  XOR U12087 ( .A(n11843), .B(n11844), .Z(n11803) );
  AND U12088 ( .A(n582), .B(n11845), .Z(n11843) );
  XOR U12089 ( .A(n11846), .B(n11844), .Z(n11845) );
  NANDN U12090 ( .A(n11805), .B(n11807), .Z(n11821) );
  XOR U12091 ( .A(n11847), .B(n11848), .Z(n11807) );
  AND U12092 ( .A(n582), .B(n11849), .Z(n11847) );
  XOR U12093 ( .A(n11848), .B(n11850), .Z(n11849) );
  XOR U12094 ( .A(n11851), .B(n11852), .Z(n582) );
  AND U12095 ( .A(n11853), .B(n11854), .Z(n11851) );
  XNOR U12096 ( .A(n11852), .B(n11818), .Z(n11854) );
  XNOR U12097 ( .A(n11855), .B(n11856), .Z(n11818) );
  ANDN U12098 ( .B(n11857), .A(n11858), .Z(n11855) );
  XOR U12099 ( .A(n11856), .B(n11859), .Z(n11857) );
  XOR U12100 ( .A(n11852), .B(n11820), .Z(n11853) );
  XOR U12101 ( .A(n11860), .B(n11861), .Z(n11820) );
  AND U12102 ( .A(n586), .B(n11862), .Z(n11860) );
  XOR U12103 ( .A(n11863), .B(n11861), .Z(n11862) );
  XNOR U12104 ( .A(n11864), .B(n11865), .Z(n11852) );
  NAND U12105 ( .A(n11866), .B(n11867), .Z(n11865) );
  XOR U12106 ( .A(n11868), .B(n11844), .Z(n11867) );
  XOR U12107 ( .A(n11858), .B(n11859), .Z(n11844) );
  XOR U12108 ( .A(n11869), .B(n11870), .Z(n11859) );
  ANDN U12109 ( .B(n11871), .A(n11872), .Z(n11869) );
  XOR U12110 ( .A(n11870), .B(n11873), .Z(n11871) );
  XOR U12111 ( .A(n11874), .B(n11875), .Z(n11858) );
  XOR U12112 ( .A(n11876), .B(n11877), .Z(n11875) );
  ANDN U12113 ( .B(n11878), .A(n11879), .Z(n11876) );
  XOR U12114 ( .A(n11880), .B(n11877), .Z(n11878) );
  IV U12115 ( .A(n11856), .Z(n11874) );
  XOR U12116 ( .A(n11881), .B(n11882), .Z(n11856) );
  ANDN U12117 ( .B(n11883), .A(n11884), .Z(n11881) );
  XOR U12118 ( .A(n11882), .B(n11885), .Z(n11883) );
  IV U12119 ( .A(n11864), .Z(n11868) );
  XOR U12120 ( .A(n11864), .B(n11846), .Z(n11866) );
  XOR U12121 ( .A(n11886), .B(n11887), .Z(n11846) );
  AND U12122 ( .A(n586), .B(n11888), .Z(n11886) );
  XOR U12123 ( .A(n11889), .B(n11887), .Z(n11888) );
  NANDN U12124 ( .A(n11848), .B(n11850), .Z(n11864) );
  XOR U12125 ( .A(n11890), .B(n11891), .Z(n11850) );
  AND U12126 ( .A(n586), .B(n11892), .Z(n11890) );
  XOR U12127 ( .A(n11891), .B(n11893), .Z(n11892) );
  XOR U12128 ( .A(n11894), .B(n11895), .Z(n586) );
  AND U12129 ( .A(n11896), .B(n11897), .Z(n11894) );
  XNOR U12130 ( .A(n11895), .B(n11861), .Z(n11897) );
  XNOR U12131 ( .A(n11898), .B(n11899), .Z(n11861) );
  ANDN U12132 ( .B(n11900), .A(n11901), .Z(n11898) );
  XOR U12133 ( .A(n11899), .B(n11902), .Z(n11900) );
  XOR U12134 ( .A(n11895), .B(n11863), .Z(n11896) );
  XOR U12135 ( .A(n11903), .B(n11904), .Z(n11863) );
  AND U12136 ( .A(n590), .B(n11905), .Z(n11903) );
  XOR U12137 ( .A(n11906), .B(n11904), .Z(n11905) );
  XNOR U12138 ( .A(n11907), .B(n11908), .Z(n11895) );
  NAND U12139 ( .A(n11909), .B(n11910), .Z(n11908) );
  XOR U12140 ( .A(n11911), .B(n11887), .Z(n11910) );
  XOR U12141 ( .A(n11901), .B(n11902), .Z(n11887) );
  XOR U12142 ( .A(n11912), .B(n11913), .Z(n11902) );
  ANDN U12143 ( .B(n11914), .A(n11915), .Z(n11912) );
  XOR U12144 ( .A(n11913), .B(n11916), .Z(n11914) );
  XOR U12145 ( .A(n11917), .B(n11918), .Z(n11901) );
  XOR U12146 ( .A(n11919), .B(n11920), .Z(n11918) );
  ANDN U12147 ( .B(n11921), .A(n11922), .Z(n11919) );
  XOR U12148 ( .A(n11923), .B(n11920), .Z(n11921) );
  IV U12149 ( .A(n11899), .Z(n11917) );
  XOR U12150 ( .A(n11924), .B(n11925), .Z(n11899) );
  ANDN U12151 ( .B(n11926), .A(n11927), .Z(n11924) );
  XOR U12152 ( .A(n11925), .B(n11928), .Z(n11926) );
  IV U12153 ( .A(n11907), .Z(n11911) );
  XOR U12154 ( .A(n11907), .B(n11889), .Z(n11909) );
  XOR U12155 ( .A(n11929), .B(n11930), .Z(n11889) );
  AND U12156 ( .A(n590), .B(n11931), .Z(n11929) );
  XOR U12157 ( .A(n11932), .B(n11930), .Z(n11931) );
  NANDN U12158 ( .A(n11891), .B(n11893), .Z(n11907) );
  XOR U12159 ( .A(n11933), .B(n11934), .Z(n11893) );
  AND U12160 ( .A(n590), .B(n11935), .Z(n11933) );
  XOR U12161 ( .A(n11934), .B(n11936), .Z(n11935) );
  XOR U12162 ( .A(n11937), .B(n11938), .Z(n590) );
  AND U12163 ( .A(n11939), .B(n11940), .Z(n11937) );
  XNOR U12164 ( .A(n11938), .B(n11904), .Z(n11940) );
  XNOR U12165 ( .A(n11941), .B(n11942), .Z(n11904) );
  ANDN U12166 ( .B(n11943), .A(n11944), .Z(n11941) );
  XOR U12167 ( .A(n11942), .B(n11945), .Z(n11943) );
  XOR U12168 ( .A(n11938), .B(n11906), .Z(n11939) );
  XOR U12169 ( .A(n11946), .B(n11947), .Z(n11906) );
  AND U12170 ( .A(n594), .B(n11948), .Z(n11946) );
  XOR U12171 ( .A(n11949), .B(n11947), .Z(n11948) );
  XNOR U12172 ( .A(n11950), .B(n11951), .Z(n11938) );
  NAND U12173 ( .A(n11952), .B(n11953), .Z(n11951) );
  XOR U12174 ( .A(n11954), .B(n11930), .Z(n11953) );
  XOR U12175 ( .A(n11944), .B(n11945), .Z(n11930) );
  XOR U12176 ( .A(n11955), .B(n11956), .Z(n11945) );
  ANDN U12177 ( .B(n11957), .A(n11958), .Z(n11955) );
  XOR U12178 ( .A(n11956), .B(n11959), .Z(n11957) );
  XOR U12179 ( .A(n11960), .B(n11961), .Z(n11944) );
  XOR U12180 ( .A(n11962), .B(n11963), .Z(n11961) );
  ANDN U12181 ( .B(n11964), .A(n11965), .Z(n11962) );
  XOR U12182 ( .A(n11966), .B(n11963), .Z(n11964) );
  IV U12183 ( .A(n11942), .Z(n11960) );
  XOR U12184 ( .A(n11967), .B(n11968), .Z(n11942) );
  ANDN U12185 ( .B(n11969), .A(n11970), .Z(n11967) );
  XOR U12186 ( .A(n11968), .B(n11971), .Z(n11969) );
  IV U12187 ( .A(n11950), .Z(n11954) );
  XOR U12188 ( .A(n11950), .B(n11932), .Z(n11952) );
  XOR U12189 ( .A(n11972), .B(n11973), .Z(n11932) );
  AND U12190 ( .A(n594), .B(n11974), .Z(n11972) );
  XOR U12191 ( .A(n11975), .B(n11973), .Z(n11974) );
  NANDN U12192 ( .A(n11934), .B(n11936), .Z(n11950) );
  XOR U12193 ( .A(n11976), .B(n11977), .Z(n11936) );
  AND U12194 ( .A(n594), .B(n11978), .Z(n11976) );
  XOR U12195 ( .A(n11977), .B(n11979), .Z(n11978) );
  XOR U12196 ( .A(n11980), .B(n11981), .Z(n594) );
  AND U12197 ( .A(n11982), .B(n11983), .Z(n11980) );
  XNOR U12198 ( .A(n11981), .B(n11947), .Z(n11983) );
  XNOR U12199 ( .A(n11984), .B(n11985), .Z(n11947) );
  ANDN U12200 ( .B(n11986), .A(n11987), .Z(n11984) );
  XOR U12201 ( .A(n11985), .B(n11988), .Z(n11986) );
  XOR U12202 ( .A(n11981), .B(n11949), .Z(n11982) );
  XOR U12203 ( .A(n11989), .B(n11990), .Z(n11949) );
  AND U12204 ( .A(n598), .B(n11991), .Z(n11989) );
  XOR U12205 ( .A(n11992), .B(n11990), .Z(n11991) );
  XNOR U12206 ( .A(n11993), .B(n11994), .Z(n11981) );
  NAND U12207 ( .A(n11995), .B(n11996), .Z(n11994) );
  XOR U12208 ( .A(n11997), .B(n11973), .Z(n11996) );
  XOR U12209 ( .A(n11987), .B(n11988), .Z(n11973) );
  XOR U12210 ( .A(n11998), .B(n11999), .Z(n11988) );
  ANDN U12211 ( .B(n12000), .A(n12001), .Z(n11998) );
  XOR U12212 ( .A(n11999), .B(n12002), .Z(n12000) );
  XOR U12213 ( .A(n12003), .B(n12004), .Z(n11987) );
  XOR U12214 ( .A(n12005), .B(n12006), .Z(n12004) );
  ANDN U12215 ( .B(n12007), .A(n12008), .Z(n12005) );
  XOR U12216 ( .A(n12009), .B(n12006), .Z(n12007) );
  IV U12217 ( .A(n11985), .Z(n12003) );
  XOR U12218 ( .A(n12010), .B(n12011), .Z(n11985) );
  ANDN U12219 ( .B(n12012), .A(n12013), .Z(n12010) );
  XOR U12220 ( .A(n12011), .B(n12014), .Z(n12012) );
  IV U12221 ( .A(n11993), .Z(n11997) );
  XOR U12222 ( .A(n11993), .B(n11975), .Z(n11995) );
  XOR U12223 ( .A(n12015), .B(n12016), .Z(n11975) );
  AND U12224 ( .A(n598), .B(n12017), .Z(n12015) );
  XOR U12225 ( .A(n12018), .B(n12016), .Z(n12017) );
  NANDN U12226 ( .A(n11977), .B(n11979), .Z(n11993) );
  XOR U12227 ( .A(n12019), .B(n12020), .Z(n11979) );
  AND U12228 ( .A(n598), .B(n12021), .Z(n12019) );
  XOR U12229 ( .A(n12020), .B(n12022), .Z(n12021) );
  XOR U12230 ( .A(n12023), .B(n12024), .Z(n598) );
  AND U12231 ( .A(n12025), .B(n12026), .Z(n12023) );
  XNOR U12232 ( .A(n12024), .B(n11990), .Z(n12026) );
  XNOR U12233 ( .A(n12027), .B(n12028), .Z(n11990) );
  ANDN U12234 ( .B(n12029), .A(n12030), .Z(n12027) );
  XOR U12235 ( .A(n12028), .B(n12031), .Z(n12029) );
  XOR U12236 ( .A(n12024), .B(n11992), .Z(n12025) );
  XOR U12237 ( .A(n12032), .B(n12033), .Z(n11992) );
  AND U12238 ( .A(n602), .B(n12034), .Z(n12032) );
  XOR U12239 ( .A(n12035), .B(n12033), .Z(n12034) );
  XNOR U12240 ( .A(n12036), .B(n12037), .Z(n12024) );
  NAND U12241 ( .A(n12038), .B(n12039), .Z(n12037) );
  XOR U12242 ( .A(n12040), .B(n12016), .Z(n12039) );
  XOR U12243 ( .A(n12030), .B(n12031), .Z(n12016) );
  XOR U12244 ( .A(n12041), .B(n12042), .Z(n12031) );
  ANDN U12245 ( .B(n12043), .A(n12044), .Z(n12041) );
  XOR U12246 ( .A(n12042), .B(n12045), .Z(n12043) );
  XOR U12247 ( .A(n12046), .B(n12047), .Z(n12030) );
  XOR U12248 ( .A(n12048), .B(n12049), .Z(n12047) );
  ANDN U12249 ( .B(n12050), .A(n12051), .Z(n12048) );
  XOR U12250 ( .A(n12052), .B(n12049), .Z(n12050) );
  IV U12251 ( .A(n12028), .Z(n12046) );
  XOR U12252 ( .A(n12053), .B(n12054), .Z(n12028) );
  ANDN U12253 ( .B(n12055), .A(n12056), .Z(n12053) );
  XOR U12254 ( .A(n12054), .B(n12057), .Z(n12055) );
  IV U12255 ( .A(n12036), .Z(n12040) );
  XOR U12256 ( .A(n12036), .B(n12018), .Z(n12038) );
  XOR U12257 ( .A(n12058), .B(n12059), .Z(n12018) );
  AND U12258 ( .A(n602), .B(n12060), .Z(n12058) );
  XOR U12259 ( .A(n12061), .B(n12059), .Z(n12060) );
  NANDN U12260 ( .A(n12020), .B(n12022), .Z(n12036) );
  XOR U12261 ( .A(n12062), .B(n12063), .Z(n12022) );
  AND U12262 ( .A(n602), .B(n12064), .Z(n12062) );
  XOR U12263 ( .A(n12063), .B(n12065), .Z(n12064) );
  XOR U12264 ( .A(n12066), .B(n12067), .Z(n602) );
  AND U12265 ( .A(n12068), .B(n12069), .Z(n12066) );
  XNOR U12266 ( .A(n12067), .B(n12033), .Z(n12069) );
  XNOR U12267 ( .A(n12070), .B(n12071), .Z(n12033) );
  ANDN U12268 ( .B(n12072), .A(n12073), .Z(n12070) );
  XOR U12269 ( .A(n12071), .B(n12074), .Z(n12072) );
  XOR U12270 ( .A(n12067), .B(n12035), .Z(n12068) );
  XOR U12271 ( .A(n12075), .B(n12076), .Z(n12035) );
  AND U12272 ( .A(n606), .B(n12077), .Z(n12075) );
  XOR U12273 ( .A(n12078), .B(n12076), .Z(n12077) );
  XNOR U12274 ( .A(n12079), .B(n12080), .Z(n12067) );
  NAND U12275 ( .A(n12081), .B(n12082), .Z(n12080) );
  XOR U12276 ( .A(n12083), .B(n12059), .Z(n12082) );
  XOR U12277 ( .A(n12073), .B(n12074), .Z(n12059) );
  XOR U12278 ( .A(n12084), .B(n12085), .Z(n12074) );
  ANDN U12279 ( .B(n12086), .A(n12087), .Z(n12084) );
  XOR U12280 ( .A(n12085), .B(n12088), .Z(n12086) );
  XOR U12281 ( .A(n12089), .B(n12090), .Z(n12073) );
  XOR U12282 ( .A(n12091), .B(n12092), .Z(n12090) );
  ANDN U12283 ( .B(n12093), .A(n12094), .Z(n12091) );
  XOR U12284 ( .A(n12095), .B(n12092), .Z(n12093) );
  IV U12285 ( .A(n12071), .Z(n12089) );
  XOR U12286 ( .A(n12096), .B(n12097), .Z(n12071) );
  ANDN U12287 ( .B(n12098), .A(n12099), .Z(n12096) );
  XOR U12288 ( .A(n12097), .B(n12100), .Z(n12098) );
  IV U12289 ( .A(n12079), .Z(n12083) );
  XOR U12290 ( .A(n12079), .B(n12061), .Z(n12081) );
  XOR U12291 ( .A(n12101), .B(n12102), .Z(n12061) );
  AND U12292 ( .A(n606), .B(n12103), .Z(n12101) );
  XOR U12293 ( .A(n12104), .B(n12102), .Z(n12103) );
  NANDN U12294 ( .A(n12063), .B(n12065), .Z(n12079) );
  XOR U12295 ( .A(n12105), .B(n12106), .Z(n12065) );
  AND U12296 ( .A(n606), .B(n12107), .Z(n12105) );
  XOR U12297 ( .A(n12106), .B(n12108), .Z(n12107) );
  XOR U12298 ( .A(n12109), .B(n12110), .Z(n606) );
  AND U12299 ( .A(n12111), .B(n12112), .Z(n12109) );
  XNOR U12300 ( .A(n12110), .B(n12076), .Z(n12112) );
  XNOR U12301 ( .A(n12113), .B(n12114), .Z(n12076) );
  ANDN U12302 ( .B(n12115), .A(n12116), .Z(n12113) );
  XOR U12303 ( .A(n12114), .B(n12117), .Z(n12115) );
  XOR U12304 ( .A(n12110), .B(n12078), .Z(n12111) );
  XOR U12305 ( .A(n12118), .B(n12119), .Z(n12078) );
  AND U12306 ( .A(n610), .B(n12120), .Z(n12118) );
  XOR U12307 ( .A(n12121), .B(n12119), .Z(n12120) );
  XNOR U12308 ( .A(n12122), .B(n12123), .Z(n12110) );
  NAND U12309 ( .A(n12124), .B(n12125), .Z(n12123) );
  XOR U12310 ( .A(n12126), .B(n12102), .Z(n12125) );
  XOR U12311 ( .A(n12116), .B(n12117), .Z(n12102) );
  XOR U12312 ( .A(n12127), .B(n12128), .Z(n12117) );
  ANDN U12313 ( .B(n12129), .A(n12130), .Z(n12127) );
  XOR U12314 ( .A(n12128), .B(n12131), .Z(n12129) );
  XOR U12315 ( .A(n12132), .B(n12133), .Z(n12116) );
  XOR U12316 ( .A(n12134), .B(n12135), .Z(n12133) );
  ANDN U12317 ( .B(n12136), .A(n12137), .Z(n12134) );
  XOR U12318 ( .A(n12138), .B(n12135), .Z(n12136) );
  IV U12319 ( .A(n12114), .Z(n12132) );
  XOR U12320 ( .A(n12139), .B(n12140), .Z(n12114) );
  ANDN U12321 ( .B(n12141), .A(n12142), .Z(n12139) );
  XOR U12322 ( .A(n12140), .B(n12143), .Z(n12141) );
  IV U12323 ( .A(n12122), .Z(n12126) );
  XOR U12324 ( .A(n12122), .B(n12104), .Z(n12124) );
  XOR U12325 ( .A(n12144), .B(n12145), .Z(n12104) );
  AND U12326 ( .A(n610), .B(n12146), .Z(n12144) );
  XOR U12327 ( .A(n12147), .B(n12145), .Z(n12146) );
  NANDN U12328 ( .A(n12106), .B(n12108), .Z(n12122) );
  XOR U12329 ( .A(n12148), .B(n12149), .Z(n12108) );
  AND U12330 ( .A(n610), .B(n12150), .Z(n12148) );
  XOR U12331 ( .A(n12149), .B(n12151), .Z(n12150) );
  XOR U12332 ( .A(n12152), .B(n12153), .Z(n610) );
  AND U12333 ( .A(n12154), .B(n12155), .Z(n12152) );
  XNOR U12334 ( .A(n12153), .B(n12119), .Z(n12155) );
  XNOR U12335 ( .A(n12156), .B(n12157), .Z(n12119) );
  ANDN U12336 ( .B(n12158), .A(n12159), .Z(n12156) );
  XOR U12337 ( .A(n12157), .B(n12160), .Z(n12158) );
  XOR U12338 ( .A(n12153), .B(n12121), .Z(n12154) );
  XOR U12339 ( .A(n12161), .B(n12162), .Z(n12121) );
  AND U12340 ( .A(n614), .B(n12163), .Z(n12161) );
  XOR U12341 ( .A(n12164), .B(n12162), .Z(n12163) );
  XNOR U12342 ( .A(n12165), .B(n12166), .Z(n12153) );
  NAND U12343 ( .A(n12167), .B(n12168), .Z(n12166) );
  XOR U12344 ( .A(n12169), .B(n12145), .Z(n12168) );
  XOR U12345 ( .A(n12159), .B(n12160), .Z(n12145) );
  XOR U12346 ( .A(n12170), .B(n12171), .Z(n12160) );
  ANDN U12347 ( .B(n12172), .A(n12173), .Z(n12170) );
  XOR U12348 ( .A(n12171), .B(n12174), .Z(n12172) );
  XOR U12349 ( .A(n12175), .B(n12176), .Z(n12159) );
  XOR U12350 ( .A(n12177), .B(n12178), .Z(n12176) );
  ANDN U12351 ( .B(n12179), .A(n12180), .Z(n12177) );
  XOR U12352 ( .A(n12181), .B(n12178), .Z(n12179) );
  IV U12353 ( .A(n12157), .Z(n12175) );
  XOR U12354 ( .A(n12182), .B(n12183), .Z(n12157) );
  ANDN U12355 ( .B(n12184), .A(n12185), .Z(n12182) );
  XOR U12356 ( .A(n12183), .B(n12186), .Z(n12184) );
  IV U12357 ( .A(n12165), .Z(n12169) );
  XOR U12358 ( .A(n12165), .B(n12147), .Z(n12167) );
  XOR U12359 ( .A(n12187), .B(n12188), .Z(n12147) );
  AND U12360 ( .A(n614), .B(n12189), .Z(n12187) );
  XOR U12361 ( .A(n12190), .B(n12188), .Z(n12189) );
  NANDN U12362 ( .A(n12149), .B(n12151), .Z(n12165) );
  XOR U12363 ( .A(n12191), .B(n12192), .Z(n12151) );
  AND U12364 ( .A(n614), .B(n12193), .Z(n12191) );
  XOR U12365 ( .A(n12192), .B(n12194), .Z(n12193) );
  XOR U12366 ( .A(n12195), .B(n12196), .Z(n614) );
  AND U12367 ( .A(n12197), .B(n12198), .Z(n12195) );
  XNOR U12368 ( .A(n12196), .B(n12162), .Z(n12198) );
  XNOR U12369 ( .A(n12199), .B(n12200), .Z(n12162) );
  ANDN U12370 ( .B(n12201), .A(n12202), .Z(n12199) );
  XOR U12371 ( .A(n12200), .B(n12203), .Z(n12201) );
  XOR U12372 ( .A(n12196), .B(n12164), .Z(n12197) );
  XOR U12373 ( .A(n12204), .B(n12205), .Z(n12164) );
  AND U12374 ( .A(n618), .B(n12206), .Z(n12204) );
  XOR U12375 ( .A(n12207), .B(n12205), .Z(n12206) );
  XNOR U12376 ( .A(n12208), .B(n12209), .Z(n12196) );
  NAND U12377 ( .A(n12210), .B(n12211), .Z(n12209) );
  XOR U12378 ( .A(n12212), .B(n12188), .Z(n12211) );
  XOR U12379 ( .A(n12202), .B(n12203), .Z(n12188) );
  XOR U12380 ( .A(n12213), .B(n12214), .Z(n12203) );
  ANDN U12381 ( .B(n12215), .A(n12216), .Z(n12213) );
  XOR U12382 ( .A(n12214), .B(n12217), .Z(n12215) );
  XOR U12383 ( .A(n12218), .B(n12219), .Z(n12202) );
  XOR U12384 ( .A(n12220), .B(n12221), .Z(n12219) );
  ANDN U12385 ( .B(n12222), .A(n12223), .Z(n12220) );
  XOR U12386 ( .A(n12224), .B(n12221), .Z(n12222) );
  IV U12387 ( .A(n12200), .Z(n12218) );
  XOR U12388 ( .A(n12225), .B(n12226), .Z(n12200) );
  ANDN U12389 ( .B(n12227), .A(n12228), .Z(n12225) );
  XOR U12390 ( .A(n12226), .B(n12229), .Z(n12227) );
  IV U12391 ( .A(n12208), .Z(n12212) );
  XOR U12392 ( .A(n12208), .B(n12190), .Z(n12210) );
  XOR U12393 ( .A(n12230), .B(n12231), .Z(n12190) );
  AND U12394 ( .A(n618), .B(n12232), .Z(n12230) );
  XOR U12395 ( .A(n12233), .B(n12231), .Z(n12232) );
  NANDN U12396 ( .A(n12192), .B(n12194), .Z(n12208) );
  XOR U12397 ( .A(n12234), .B(n12235), .Z(n12194) );
  AND U12398 ( .A(n618), .B(n12236), .Z(n12234) );
  XOR U12399 ( .A(n12235), .B(n12237), .Z(n12236) );
  XOR U12400 ( .A(n12238), .B(n12239), .Z(n618) );
  AND U12401 ( .A(n12240), .B(n12241), .Z(n12238) );
  XNOR U12402 ( .A(n12239), .B(n12205), .Z(n12241) );
  XNOR U12403 ( .A(n12242), .B(n12243), .Z(n12205) );
  ANDN U12404 ( .B(n12244), .A(n12245), .Z(n12242) );
  XOR U12405 ( .A(n12243), .B(n12246), .Z(n12244) );
  XOR U12406 ( .A(n12239), .B(n12207), .Z(n12240) );
  XOR U12407 ( .A(n12247), .B(n12248), .Z(n12207) );
  AND U12408 ( .A(n622), .B(n12249), .Z(n12247) );
  XOR U12409 ( .A(n12250), .B(n12248), .Z(n12249) );
  XNOR U12410 ( .A(n12251), .B(n12252), .Z(n12239) );
  NAND U12411 ( .A(n12253), .B(n12254), .Z(n12252) );
  XOR U12412 ( .A(n12255), .B(n12231), .Z(n12254) );
  XOR U12413 ( .A(n12245), .B(n12246), .Z(n12231) );
  XOR U12414 ( .A(n12256), .B(n12257), .Z(n12246) );
  ANDN U12415 ( .B(n12258), .A(n12259), .Z(n12256) );
  XOR U12416 ( .A(n12257), .B(n12260), .Z(n12258) );
  XOR U12417 ( .A(n12261), .B(n12262), .Z(n12245) );
  XOR U12418 ( .A(n12263), .B(n12264), .Z(n12262) );
  ANDN U12419 ( .B(n12265), .A(n12266), .Z(n12263) );
  XOR U12420 ( .A(n12267), .B(n12264), .Z(n12265) );
  IV U12421 ( .A(n12243), .Z(n12261) );
  XOR U12422 ( .A(n12268), .B(n12269), .Z(n12243) );
  ANDN U12423 ( .B(n12270), .A(n12271), .Z(n12268) );
  XOR U12424 ( .A(n12269), .B(n12272), .Z(n12270) );
  IV U12425 ( .A(n12251), .Z(n12255) );
  XOR U12426 ( .A(n12251), .B(n12233), .Z(n12253) );
  XOR U12427 ( .A(n12273), .B(n12274), .Z(n12233) );
  AND U12428 ( .A(n622), .B(n12275), .Z(n12273) );
  XOR U12429 ( .A(n12276), .B(n12274), .Z(n12275) );
  NANDN U12430 ( .A(n12235), .B(n12237), .Z(n12251) );
  XOR U12431 ( .A(n12277), .B(n12278), .Z(n12237) );
  AND U12432 ( .A(n622), .B(n12279), .Z(n12277) );
  XOR U12433 ( .A(n12278), .B(n12280), .Z(n12279) );
  XOR U12434 ( .A(n12281), .B(n12282), .Z(n622) );
  AND U12435 ( .A(n12283), .B(n12284), .Z(n12281) );
  XNOR U12436 ( .A(n12282), .B(n12248), .Z(n12284) );
  XNOR U12437 ( .A(n12285), .B(n12286), .Z(n12248) );
  ANDN U12438 ( .B(n12287), .A(n12288), .Z(n12285) );
  XOR U12439 ( .A(n12286), .B(n12289), .Z(n12287) );
  XOR U12440 ( .A(n12282), .B(n12250), .Z(n12283) );
  XOR U12441 ( .A(n12290), .B(n12291), .Z(n12250) );
  AND U12442 ( .A(n626), .B(n12292), .Z(n12290) );
  XOR U12443 ( .A(n12293), .B(n12291), .Z(n12292) );
  XNOR U12444 ( .A(n12294), .B(n12295), .Z(n12282) );
  NAND U12445 ( .A(n12296), .B(n12297), .Z(n12295) );
  XOR U12446 ( .A(n12298), .B(n12274), .Z(n12297) );
  XOR U12447 ( .A(n12288), .B(n12289), .Z(n12274) );
  XOR U12448 ( .A(n12299), .B(n12300), .Z(n12289) );
  ANDN U12449 ( .B(n12301), .A(n12302), .Z(n12299) );
  XOR U12450 ( .A(n12300), .B(n12303), .Z(n12301) );
  XOR U12451 ( .A(n12304), .B(n12305), .Z(n12288) );
  XOR U12452 ( .A(n12306), .B(n12307), .Z(n12305) );
  ANDN U12453 ( .B(n12308), .A(n12309), .Z(n12306) );
  XOR U12454 ( .A(n12310), .B(n12307), .Z(n12308) );
  IV U12455 ( .A(n12286), .Z(n12304) );
  XOR U12456 ( .A(n12311), .B(n12312), .Z(n12286) );
  ANDN U12457 ( .B(n12313), .A(n12314), .Z(n12311) );
  XOR U12458 ( .A(n12312), .B(n12315), .Z(n12313) );
  IV U12459 ( .A(n12294), .Z(n12298) );
  XOR U12460 ( .A(n12294), .B(n12276), .Z(n12296) );
  XOR U12461 ( .A(n12316), .B(n12317), .Z(n12276) );
  AND U12462 ( .A(n626), .B(n12318), .Z(n12316) );
  XOR U12463 ( .A(n12319), .B(n12317), .Z(n12318) );
  NANDN U12464 ( .A(n12278), .B(n12280), .Z(n12294) );
  XOR U12465 ( .A(n12320), .B(n12321), .Z(n12280) );
  AND U12466 ( .A(n626), .B(n12322), .Z(n12320) );
  XOR U12467 ( .A(n12321), .B(n12323), .Z(n12322) );
  XOR U12468 ( .A(n12324), .B(n12325), .Z(n626) );
  AND U12469 ( .A(n12326), .B(n12327), .Z(n12324) );
  XNOR U12470 ( .A(n12325), .B(n12291), .Z(n12327) );
  XNOR U12471 ( .A(n12328), .B(n12329), .Z(n12291) );
  ANDN U12472 ( .B(n12330), .A(n12331), .Z(n12328) );
  XOR U12473 ( .A(n12329), .B(n12332), .Z(n12330) );
  XOR U12474 ( .A(n12325), .B(n12293), .Z(n12326) );
  XOR U12475 ( .A(n12333), .B(n12334), .Z(n12293) );
  AND U12476 ( .A(n630), .B(n12335), .Z(n12333) );
  XOR U12477 ( .A(n12336), .B(n12334), .Z(n12335) );
  XNOR U12478 ( .A(n12337), .B(n12338), .Z(n12325) );
  NAND U12479 ( .A(n12339), .B(n12340), .Z(n12338) );
  XOR U12480 ( .A(n12341), .B(n12317), .Z(n12340) );
  XOR U12481 ( .A(n12331), .B(n12332), .Z(n12317) );
  XOR U12482 ( .A(n12342), .B(n12343), .Z(n12332) );
  ANDN U12483 ( .B(n12344), .A(n12345), .Z(n12342) );
  XOR U12484 ( .A(n12343), .B(n12346), .Z(n12344) );
  XOR U12485 ( .A(n12347), .B(n12348), .Z(n12331) );
  XOR U12486 ( .A(n12349), .B(n12350), .Z(n12348) );
  ANDN U12487 ( .B(n12351), .A(n12352), .Z(n12349) );
  XOR U12488 ( .A(n12353), .B(n12350), .Z(n12351) );
  IV U12489 ( .A(n12329), .Z(n12347) );
  XOR U12490 ( .A(n12354), .B(n12355), .Z(n12329) );
  ANDN U12491 ( .B(n12356), .A(n12357), .Z(n12354) );
  XOR U12492 ( .A(n12355), .B(n12358), .Z(n12356) );
  IV U12493 ( .A(n12337), .Z(n12341) );
  XOR U12494 ( .A(n12337), .B(n12319), .Z(n12339) );
  XOR U12495 ( .A(n12359), .B(n12360), .Z(n12319) );
  AND U12496 ( .A(n630), .B(n12361), .Z(n12359) );
  XOR U12497 ( .A(n12362), .B(n12360), .Z(n12361) );
  NANDN U12498 ( .A(n12321), .B(n12323), .Z(n12337) );
  XOR U12499 ( .A(n12363), .B(n12364), .Z(n12323) );
  AND U12500 ( .A(n630), .B(n12365), .Z(n12363) );
  XOR U12501 ( .A(n12364), .B(n12366), .Z(n12365) );
  XOR U12502 ( .A(n12367), .B(n12368), .Z(n630) );
  AND U12503 ( .A(n12369), .B(n12370), .Z(n12367) );
  XNOR U12504 ( .A(n12368), .B(n12334), .Z(n12370) );
  XNOR U12505 ( .A(n12371), .B(n12372), .Z(n12334) );
  ANDN U12506 ( .B(n12373), .A(n12374), .Z(n12371) );
  XOR U12507 ( .A(n12372), .B(n12375), .Z(n12373) );
  XOR U12508 ( .A(n12368), .B(n12336), .Z(n12369) );
  XOR U12509 ( .A(n12376), .B(n12377), .Z(n12336) );
  AND U12510 ( .A(n634), .B(n12378), .Z(n12376) );
  XOR U12511 ( .A(n12379), .B(n12377), .Z(n12378) );
  XNOR U12512 ( .A(n12380), .B(n12381), .Z(n12368) );
  NAND U12513 ( .A(n12382), .B(n12383), .Z(n12381) );
  XOR U12514 ( .A(n12384), .B(n12360), .Z(n12383) );
  XOR U12515 ( .A(n12374), .B(n12375), .Z(n12360) );
  XOR U12516 ( .A(n12385), .B(n12386), .Z(n12375) );
  ANDN U12517 ( .B(n12387), .A(n12388), .Z(n12385) );
  XOR U12518 ( .A(n12386), .B(n12389), .Z(n12387) );
  XOR U12519 ( .A(n12390), .B(n12391), .Z(n12374) );
  XOR U12520 ( .A(n12392), .B(n12393), .Z(n12391) );
  ANDN U12521 ( .B(n12394), .A(n12395), .Z(n12392) );
  XOR U12522 ( .A(n12396), .B(n12393), .Z(n12394) );
  IV U12523 ( .A(n12372), .Z(n12390) );
  XOR U12524 ( .A(n12397), .B(n12398), .Z(n12372) );
  ANDN U12525 ( .B(n12399), .A(n12400), .Z(n12397) );
  XOR U12526 ( .A(n12398), .B(n12401), .Z(n12399) );
  IV U12527 ( .A(n12380), .Z(n12384) );
  XOR U12528 ( .A(n12380), .B(n12362), .Z(n12382) );
  XOR U12529 ( .A(n12402), .B(n12403), .Z(n12362) );
  AND U12530 ( .A(n634), .B(n12404), .Z(n12402) );
  XOR U12531 ( .A(n12405), .B(n12403), .Z(n12404) );
  NANDN U12532 ( .A(n12364), .B(n12366), .Z(n12380) );
  XOR U12533 ( .A(n12406), .B(n12407), .Z(n12366) );
  AND U12534 ( .A(n634), .B(n12408), .Z(n12406) );
  XOR U12535 ( .A(n12407), .B(n12409), .Z(n12408) );
  XOR U12536 ( .A(n12410), .B(n12411), .Z(n634) );
  AND U12537 ( .A(n12412), .B(n12413), .Z(n12410) );
  XNOR U12538 ( .A(n12411), .B(n12377), .Z(n12413) );
  XNOR U12539 ( .A(n12414), .B(n12415), .Z(n12377) );
  ANDN U12540 ( .B(n12416), .A(n12417), .Z(n12414) );
  XOR U12541 ( .A(n12415), .B(n12418), .Z(n12416) );
  XOR U12542 ( .A(n12411), .B(n12379), .Z(n12412) );
  XOR U12543 ( .A(n12419), .B(n12420), .Z(n12379) );
  AND U12544 ( .A(n638), .B(n12421), .Z(n12419) );
  XOR U12545 ( .A(n12422), .B(n12420), .Z(n12421) );
  XNOR U12546 ( .A(n12423), .B(n12424), .Z(n12411) );
  NAND U12547 ( .A(n12425), .B(n12426), .Z(n12424) );
  XOR U12548 ( .A(n12427), .B(n12403), .Z(n12426) );
  XOR U12549 ( .A(n12417), .B(n12418), .Z(n12403) );
  XOR U12550 ( .A(n12428), .B(n12429), .Z(n12418) );
  ANDN U12551 ( .B(n12430), .A(n12431), .Z(n12428) );
  XOR U12552 ( .A(n12429), .B(n12432), .Z(n12430) );
  XOR U12553 ( .A(n12433), .B(n12434), .Z(n12417) );
  XOR U12554 ( .A(n12435), .B(n12436), .Z(n12434) );
  ANDN U12555 ( .B(n12437), .A(n12438), .Z(n12435) );
  XOR U12556 ( .A(n12439), .B(n12436), .Z(n12437) );
  IV U12557 ( .A(n12415), .Z(n12433) );
  XOR U12558 ( .A(n12440), .B(n12441), .Z(n12415) );
  ANDN U12559 ( .B(n12442), .A(n12443), .Z(n12440) );
  XOR U12560 ( .A(n12441), .B(n12444), .Z(n12442) );
  IV U12561 ( .A(n12423), .Z(n12427) );
  XOR U12562 ( .A(n12423), .B(n12405), .Z(n12425) );
  XOR U12563 ( .A(n12445), .B(n12446), .Z(n12405) );
  AND U12564 ( .A(n638), .B(n12447), .Z(n12445) );
  XOR U12565 ( .A(n12448), .B(n12446), .Z(n12447) );
  NANDN U12566 ( .A(n12407), .B(n12409), .Z(n12423) );
  XOR U12567 ( .A(n12449), .B(n12450), .Z(n12409) );
  AND U12568 ( .A(n638), .B(n12451), .Z(n12449) );
  XOR U12569 ( .A(n12450), .B(n12452), .Z(n12451) );
  XOR U12570 ( .A(n12453), .B(n12454), .Z(n638) );
  AND U12571 ( .A(n12455), .B(n12456), .Z(n12453) );
  XNOR U12572 ( .A(n12454), .B(n12420), .Z(n12456) );
  XNOR U12573 ( .A(n12457), .B(n12458), .Z(n12420) );
  ANDN U12574 ( .B(n12459), .A(n12460), .Z(n12457) );
  XOR U12575 ( .A(n12458), .B(n12461), .Z(n12459) );
  XOR U12576 ( .A(n12454), .B(n12422), .Z(n12455) );
  XOR U12577 ( .A(n12462), .B(n12463), .Z(n12422) );
  AND U12578 ( .A(n642), .B(n12464), .Z(n12462) );
  XOR U12579 ( .A(n12465), .B(n12463), .Z(n12464) );
  XNOR U12580 ( .A(n12466), .B(n12467), .Z(n12454) );
  NAND U12581 ( .A(n12468), .B(n12469), .Z(n12467) );
  XOR U12582 ( .A(n12470), .B(n12446), .Z(n12469) );
  XOR U12583 ( .A(n12460), .B(n12461), .Z(n12446) );
  XOR U12584 ( .A(n12471), .B(n12472), .Z(n12461) );
  ANDN U12585 ( .B(n12473), .A(n12474), .Z(n12471) );
  XOR U12586 ( .A(n12472), .B(n12475), .Z(n12473) );
  XOR U12587 ( .A(n12476), .B(n12477), .Z(n12460) );
  XOR U12588 ( .A(n12478), .B(n12479), .Z(n12477) );
  ANDN U12589 ( .B(n12480), .A(n12481), .Z(n12478) );
  XOR U12590 ( .A(n12482), .B(n12479), .Z(n12480) );
  IV U12591 ( .A(n12458), .Z(n12476) );
  XOR U12592 ( .A(n12483), .B(n12484), .Z(n12458) );
  ANDN U12593 ( .B(n12485), .A(n12486), .Z(n12483) );
  XOR U12594 ( .A(n12484), .B(n12487), .Z(n12485) );
  IV U12595 ( .A(n12466), .Z(n12470) );
  XOR U12596 ( .A(n12466), .B(n12448), .Z(n12468) );
  XOR U12597 ( .A(n12488), .B(n12489), .Z(n12448) );
  AND U12598 ( .A(n642), .B(n12490), .Z(n12488) );
  XOR U12599 ( .A(n12491), .B(n12489), .Z(n12490) );
  NANDN U12600 ( .A(n12450), .B(n12452), .Z(n12466) );
  XOR U12601 ( .A(n12492), .B(n12493), .Z(n12452) );
  AND U12602 ( .A(n642), .B(n12494), .Z(n12492) );
  XOR U12603 ( .A(n12493), .B(n12495), .Z(n12494) );
  XOR U12604 ( .A(n12496), .B(n12497), .Z(n642) );
  AND U12605 ( .A(n12498), .B(n12499), .Z(n12496) );
  XNOR U12606 ( .A(n12497), .B(n12463), .Z(n12499) );
  XNOR U12607 ( .A(n12500), .B(n12501), .Z(n12463) );
  ANDN U12608 ( .B(n12502), .A(n12503), .Z(n12500) );
  XOR U12609 ( .A(n12501), .B(n12504), .Z(n12502) );
  XOR U12610 ( .A(n12497), .B(n12465), .Z(n12498) );
  XOR U12611 ( .A(n12505), .B(n12506), .Z(n12465) );
  AND U12612 ( .A(n646), .B(n12507), .Z(n12505) );
  XOR U12613 ( .A(n12508), .B(n12506), .Z(n12507) );
  XNOR U12614 ( .A(n12509), .B(n12510), .Z(n12497) );
  NAND U12615 ( .A(n12511), .B(n12512), .Z(n12510) );
  XOR U12616 ( .A(n12513), .B(n12489), .Z(n12512) );
  XOR U12617 ( .A(n12503), .B(n12504), .Z(n12489) );
  XOR U12618 ( .A(n12514), .B(n12515), .Z(n12504) );
  ANDN U12619 ( .B(n12516), .A(n12517), .Z(n12514) );
  XOR U12620 ( .A(n12515), .B(n12518), .Z(n12516) );
  XOR U12621 ( .A(n12519), .B(n12520), .Z(n12503) );
  XOR U12622 ( .A(n12521), .B(n12522), .Z(n12520) );
  ANDN U12623 ( .B(n12523), .A(n12524), .Z(n12521) );
  XOR U12624 ( .A(n12525), .B(n12522), .Z(n12523) );
  IV U12625 ( .A(n12501), .Z(n12519) );
  XOR U12626 ( .A(n12526), .B(n12527), .Z(n12501) );
  ANDN U12627 ( .B(n12528), .A(n12529), .Z(n12526) );
  XOR U12628 ( .A(n12527), .B(n12530), .Z(n12528) );
  IV U12629 ( .A(n12509), .Z(n12513) );
  XOR U12630 ( .A(n12509), .B(n12491), .Z(n12511) );
  XOR U12631 ( .A(n12531), .B(n12532), .Z(n12491) );
  AND U12632 ( .A(n646), .B(n12533), .Z(n12531) );
  XOR U12633 ( .A(n12534), .B(n12532), .Z(n12533) );
  NANDN U12634 ( .A(n12493), .B(n12495), .Z(n12509) );
  XOR U12635 ( .A(n12535), .B(n12536), .Z(n12495) );
  AND U12636 ( .A(n646), .B(n12537), .Z(n12535) );
  XOR U12637 ( .A(n12536), .B(n12538), .Z(n12537) );
  XOR U12638 ( .A(n12539), .B(n12540), .Z(n646) );
  AND U12639 ( .A(n12541), .B(n12542), .Z(n12539) );
  XNOR U12640 ( .A(n12540), .B(n12506), .Z(n12542) );
  XNOR U12641 ( .A(n12543), .B(n12544), .Z(n12506) );
  ANDN U12642 ( .B(n12545), .A(n12546), .Z(n12543) );
  XOR U12643 ( .A(n12544), .B(n12547), .Z(n12545) );
  XOR U12644 ( .A(n12540), .B(n12508), .Z(n12541) );
  XOR U12645 ( .A(n12548), .B(n12549), .Z(n12508) );
  AND U12646 ( .A(n650), .B(n12550), .Z(n12548) );
  XOR U12647 ( .A(n12551), .B(n12549), .Z(n12550) );
  XNOR U12648 ( .A(n12552), .B(n12553), .Z(n12540) );
  NAND U12649 ( .A(n12554), .B(n12555), .Z(n12553) );
  XOR U12650 ( .A(n12556), .B(n12532), .Z(n12555) );
  XOR U12651 ( .A(n12546), .B(n12547), .Z(n12532) );
  XOR U12652 ( .A(n12557), .B(n12558), .Z(n12547) );
  ANDN U12653 ( .B(n12559), .A(n12560), .Z(n12557) );
  XOR U12654 ( .A(n12558), .B(n12561), .Z(n12559) );
  XOR U12655 ( .A(n12562), .B(n12563), .Z(n12546) );
  XOR U12656 ( .A(n12564), .B(n12565), .Z(n12563) );
  ANDN U12657 ( .B(n12566), .A(n12567), .Z(n12564) );
  XOR U12658 ( .A(n12568), .B(n12565), .Z(n12566) );
  IV U12659 ( .A(n12544), .Z(n12562) );
  XOR U12660 ( .A(n12569), .B(n12570), .Z(n12544) );
  ANDN U12661 ( .B(n12571), .A(n12572), .Z(n12569) );
  XOR U12662 ( .A(n12570), .B(n12573), .Z(n12571) );
  IV U12663 ( .A(n12552), .Z(n12556) );
  XOR U12664 ( .A(n12552), .B(n12534), .Z(n12554) );
  XOR U12665 ( .A(n12574), .B(n12575), .Z(n12534) );
  AND U12666 ( .A(n650), .B(n12576), .Z(n12574) );
  XOR U12667 ( .A(n12577), .B(n12575), .Z(n12576) );
  NANDN U12668 ( .A(n12536), .B(n12538), .Z(n12552) );
  XOR U12669 ( .A(n12578), .B(n12579), .Z(n12538) );
  AND U12670 ( .A(n650), .B(n12580), .Z(n12578) );
  XOR U12671 ( .A(n12579), .B(n12581), .Z(n12580) );
  XOR U12672 ( .A(n12582), .B(n12583), .Z(n650) );
  AND U12673 ( .A(n12584), .B(n12585), .Z(n12582) );
  XNOR U12674 ( .A(n12583), .B(n12549), .Z(n12585) );
  XNOR U12675 ( .A(n12586), .B(n12587), .Z(n12549) );
  ANDN U12676 ( .B(n12588), .A(n12589), .Z(n12586) );
  XOR U12677 ( .A(n12587), .B(n12590), .Z(n12588) );
  XOR U12678 ( .A(n12583), .B(n12551), .Z(n12584) );
  XOR U12679 ( .A(n12591), .B(n12592), .Z(n12551) );
  AND U12680 ( .A(n654), .B(n12593), .Z(n12591) );
  XOR U12681 ( .A(n12594), .B(n12592), .Z(n12593) );
  XNOR U12682 ( .A(n12595), .B(n12596), .Z(n12583) );
  NAND U12683 ( .A(n12597), .B(n12598), .Z(n12596) );
  XOR U12684 ( .A(n12599), .B(n12575), .Z(n12598) );
  XOR U12685 ( .A(n12589), .B(n12590), .Z(n12575) );
  XOR U12686 ( .A(n12600), .B(n12601), .Z(n12590) );
  ANDN U12687 ( .B(n12602), .A(n12603), .Z(n12600) );
  XOR U12688 ( .A(n12601), .B(n12604), .Z(n12602) );
  XOR U12689 ( .A(n12605), .B(n12606), .Z(n12589) );
  XOR U12690 ( .A(n12607), .B(n12608), .Z(n12606) );
  ANDN U12691 ( .B(n12609), .A(n12610), .Z(n12607) );
  XOR U12692 ( .A(n12611), .B(n12608), .Z(n12609) );
  IV U12693 ( .A(n12587), .Z(n12605) );
  XOR U12694 ( .A(n12612), .B(n12613), .Z(n12587) );
  ANDN U12695 ( .B(n12614), .A(n12615), .Z(n12612) );
  XOR U12696 ( .A(n12613), .B(n12616), .Z(n12614) );
  IV U12697 ( .A(n12595), .Z(n12599) );
  XOR U12698 ( .A(n12595), .B(n12577), .Z(n12597) );
  XOR U12699 ( .A(n12617), .B(n12618), .Z(n12577) );
  AND U12700 ( .A(n654), .B(n12619), .Z(n12617) );
  XOR U12701 ( .A(n12620), .B(n12618), .Z(n12619) );
  NANDN U12702 ( .A(n12579), .B(n12581), .Z(n12595) );
  XOR U12703 ( .A(n12621), .B(n12622), .Z(n12581) );
  AND U12704 ( .A(n654), .B(n12623), .Z(n12621) );
  XOR U12705 ( .A(n12622), .B(n12624), .Z(n12623) );
  XOR U12706 ( .A(n12625), .B(n12626), .Z(n654) );
  AND U12707 ( .A(n12627), .B(n12628), .Z(n12625) );
  XNOR U12708 ( .A(n12626), .B(n12592), .Z(n12628) );
  XNOR U12709 ( .A(n12629), .B(n12630), .Z(n12592) );
  ANDN U12710 ( .B(n12631), .A(n12632), .Z(n12629) );
  XOR U12711 ( .A(n12630), .B(n12633), .Z(n12631) );
  XOR U12712 ( .A(n12626), .B(n12594), .Z(n12627) );
  XOR U12713 ( .A(n12634), .B(n12635), .Z(n12594) );
  AND U12714 ( .A(n658), .B(n12636), .Z(n12634) );
  XOR U12715 ( .A(n12637), .B(n12635), .Z(n12636) );
  XNOR U12716 ( .A(n12638), .B(n12639), .Z(n12626) );
  NAND U12717 ( .A(n12640), .B(n12641), .Z(n12639) );
  XOR U12718 ( .A(n12642), .B(n12618), .Z(n12641) );
  XOR U12719 ( .A(n12632), .B(n12633), .Z(n12618) );
  XOR U12720 ( .A(n12643), .B(n12644), .Z(n12633) );
  ANDN U12721 ( .B(n12645), .A(n12646), .Z(n12643) );
  XOR U12722 ( .A(n12644), .B(n12647), .Z(n12645) );
  XOR U12723 ( .A(n12648), .B(n12649), .Z(n12632) );
  XOR U12724 ( .A(n12650), .B(n12651), .Z(n12649) );
  ANDN U12725 ( .B(n12652), .A(n12653), .Z(n12650) );
  XOR U12726 ( .A(n12654), .B(n12651), .Z(n12652) );
  IV U12727 ( .A(n12630), .Z(n12648) );
  XOR U12728 ( .A(n12655), .B(n12656), .Z(n12630) );
  ANDN U12729 ( .B(n12657), .A(n12658), .Z(n12655) );
  XOR U12730 ( .A(n12656), .B(n12659), .Z(n12657) );
  IV U12731 ( .A(n12638), .Z(n12642) );
  XOR U12732 ( .A(n12638), .B(n12620), .Z(n12640) );
  XOR U12733 ( .A(n12660), .B(n12661), .Z(n12620) );
  AND U12734 ( .A(n658), .B(n12662), .Z(n12660) );
  XOR U12735 ( .A(n12663), .B(n12661), .Z(n12662) );
  NANDN U12736 ( .A(n12622), .B(n12624), .Z(n12638) );
  XOR U12737 ( .A(n12664), .B(n12665), .Z(n12624) );
  AND U12738 ( .A(n658), .B(n12666), .Z(n12664) );
  XOR U12739 ( .A(n12665), .B(n12667), .Z(n12666) );
  XOR U12740 ( .A(n12668), .B(n12669), .Z(n658) );
  AND U12741 ( .A(n12670), .B(n12671), .Z(n12668) );
  XNOR U12742 ( .A(n12669), .B(n12635), .Z(n12671) );
  XNOR U12743 ( .A(n12672), .B(n12673), .Z(n12635) );
  ANDN U12744 ( .B(n12674), .A(n12675), .Z(n12672) );
  XOR U12745 ( .A(n12673), .B(n12676), .Z(n12674) );
  XOR U12746 ( .A(n12669), .B(n12637), .Z(n12670) );
  XOR U12747 ( .A(n12677), .B(n12678), .Z(n12637) );
  AND U12748 ( .A(n662), .B(n12679), .Z(n12677) );
  XOR U12749 ( .A(n12680), .B(n12678), .Z(n12679) );
  XNOR U12750 ( .A(n12681), .B(n12682), .Z(n12669) );
  NAND U12751 ( .A(n12683), .B(n12684), .Z(n12682) );
  XOR U12752 ( .A(n12685), .B(n12661), .Z(n12684) );
  XOR U12753 ( .A(n12675), .B(n12676), .Z(n12661) );
  XOR U12754 ( .A(n12686), .B(n12687), .Z(n12676) );
  ANDN U12755 ( .B(n12688), .A(n12689), .Z(n12686) );
  XOR U12756 ( .A(n12687), .B(n12690), .Z(n12688) );
  XOR U12757 ( .A(n12691), .B(n12692), .Z(n12675) );
  XOR U12758 ( .A(n12693), .B(n12694), .Z(n12692) );
  ANDN U12759 ( .B(n12695), .A(n12696), .Z(n12693) );
  XOR U12760 ( .A(n12697), .B(n12694), .Z(n12695) );
  IV U12761 ( .A(n12673), .Z(n12691) );
  XOR U12762 ( .A(n12698), .B(n12699), .Z(n12673) );
  ANDN U12763 ( .B(n12700), .A(n12701), .Z(n12698) );
  XOR U12764 ( .A(n12699), .B(n12702), .Z(n12700) );
  IV U12765 ( .A(n12681), .Z(n12685) );
  XOR U12766 ( .A(n12681), .B(n12663), .Z(n12683) );
  XOR U12767 ( .A(n12703), .B(n12704), .Z(n12663) );
  AND U12768 ( .A(n662), .B(n12705), .Z(n12703) );
  XOR U12769 ( .A(n12706), .B(n12704), .Z(n12705) );
  NANDN U12770 ( .A(n12665), .B(n12667), .Z(n12681) );
  XOR U12771 ( .A(n12707), .B(n12708), .Z(n12667) );
  AND U12772 ( .A(n662), .B(n12709), .Z(n12707) );
  XOR U12773 ( .A(n12708), .B(n12710), .Z(n12709) );
  XOR U12774 ( .A(n12711), .B(n12712), .Z(n662) );
  AND U12775 ( .A(n12713), .B(n12714), .Z(n12711) );
  XNOR U12776 ( .A(n12712), .B(n12678), .Z(n12714) );
  XNOR U12777 ( .A(n12715), .B(n12716), .Z(n12678) );
  ANDN U12778 ( .B(n12717), .A(n12718), .Z(n12715) );
  XOR U12779 ( .A(n12716), .B(n12719), .Z(n12717) );
  XOR U12780 ( .A(n12712), .B(n12680), .Z(n12713) );
  XOR U12781 ( .A(n12720), .B(n12721), .Z(n12680) );
  AND U12782 ( .A(n666), .B(n12722), .Z(n12720) );
  XOR U12783 ( .A(n12723), .B(n12721), .Z(n12722) );
  XNOR U12784 ( .A(n12724), .B(n12725), .Z(n12712) );
  NAND U12785 ( .A(n12726), .B(n12727), .Z(n12725) );
  XOR U12786 ( .A(n12728), .B(n12704), .Z(n12727) );
  XOR U12787 ( .A(n12718), .B(n12719), .Z(n12704) );
  XOR U12788 ( .A(n12729), .B(n12730), .Z(n12719) );
  ANDN U12789 ( .B(n12731), .A(n12732), .Z(n12729) );
  XOR U12790 ( .A(n12730), .B(n12733), .Z(n12731) );
  XOR U12791 ( .A(n12734), .B(n12735), .Z(n12718) );
  XOR U12792 ( .A(n12736), .B(n12737), .Z(n12735) );
  ANDN U12793 ( .B(n12738), .A(n12739), .Z(n12736) );
  XOR U12794 ( .A(n12740), .B(n12737), .Z(n12738) );
  IV U12795 ( .A(n12716), .Z(n12734) );
  XOR U12796 ( .A(n12741), .B(n12742), .Z(n12716) );
  ANDN U12797 ( .B(n12743), .A(n12744), .Z(n12741) );
  XOR U12798 ( .A(n12742), .B(n12745), .Z(n12743) );
  IV U12799 ( .A(n12724), .Z(n12728) );
  XOR U12800 ( .A(n12724), .B(n12706), .Z(n12726) );
  XOR U12801 ( .A(n12746), .B(n12747), .Z(n12706) );
  AND U12802 ( .A(n666), .B(n12748), .Z(n12746) );
  XOR U12803 ( .A(n12749), .B(n12747), .Z(n12748) );
  NANDN U12804 ( .A(n12708), .B(n12710), .Z(n12724) );
  XOR U12805 ( .A(n12750), .B(n12751), .Z(n12710) );
  AND U12806 ( .A(n666), .B(n12752), .Z(n12750) );
  XOR U12807 ( .A(n12751), .B(n12753), .Z(n12752) );
  XOR U12808 ( .A(n12754), .B(n12755), .Z(n666) );
  AND U12809 ( .A(n12756), .B(n12757), .Z(n12754) );
  XNOR U12810 ( .A(n12755), .B(n12721), .Z(n12757) );
  XNOR U12811 ( .A(n12758), .B(n12759), .Z(n12721) );
  ANDN U12812 ( .B(n12760), .A(n12761), .Z(n12758) );
  XOR U12813 ( .A(n12759), .B(n12762), .Z(n12760) );
  XOR U12814 ( .A(n12755), .B(n12723), .Z(n12756) );
  XOR U12815 ( .A(n12763), .B(n12764), .Z(n12723) );
  AND U12816 ( .A(n670), .B(n12765), .Z(n12763) );
  XOR U12817 ( .A(n12766), .B(n12764), .Z(n12765) );
  XNOR U12818 ( .A(n12767), .B(n12768), .Z(n12755) );
  NAND U12819 ( .A(n12769), .B(n12770), .Z(n12768) );
  XOR U12820 ( .A(n12771), .B(n12747), .Z(n12770) );
  XOR U12821 ( .A(n12761), .B(n12762), .Z(n12747) );
  XOR U12822 ( .A(n12772), .B(n12773), .Z(n12762) );
  ANDN U12823 ( .B(n12774), .A(n12775), .Z(n12772) );
  XOR U12824 ( .A(n12773), .B(n12776), .Z(n12774) );
  XOR U12825 ( .A(n12777), .B(n12778), .Z(n12761) );
  XOR U12826 ( .A(n12779), .B(n12780), .Z(n12778) );
  ANDN U12827 ( .B(n12781), .A(n12782), .Z(n12779) );
  XOR U12828 ( .A(n12783), .B(n12780), .Z(n12781) );
  IV U12829 ( .A(n12759), .Z(n12777) );
  XOR U12830 ( .A(n12784), .B(n12785), .Z(n12759) );
  ANDN U12831 ( .B(n12786), .A(n12787), .Z(n12784) );
  XOR U12832 ( .A(n12785), .B(n12788), .Z(n12786) );
  IV U12833 ( .A(n12767), .Z(n12771) );
  XOR U12834 ( .A(n12767), .B(n12749), .Z(n12769) );
  XOR U12835 ( .A(n12789), .B(n12790), .Z(n12749) );
  AND U12836 ( .A(n670), .B(n12791), .Z(n12789) );
  XOR U12837 ( .A(n12792), .B(n12790), .Z(n12791) );
  NANDN U12838 ( .A(n12751), .B(n12753), .Z(n12767) );
  XOR U12839 ( .A(n12793), .B(n12794), .Z(n12753) );
  AND U12840 ( .A(n670), .B(n12795), .Z(n12793) );
  XOR U12841 ( .A(n12794), .B(n12796), .Z(n12795) );
  XOR U12842 ( .A(n12797), .B(n12798), .Z(n670) );
  AND U12843 ( .A(n12799), .B(n12800), .Z(n12797) );
  XNOR U12844 ( .A(n12798), .B(n12764), .Z(n12800) );
  XNOR U12845 ( .A(n12801), .B(n12802), .Z(n12764) );
  ANDN U12846 ( .B(n12803), .A(n12804), .Z(n12801) );
  XOR U12847 ( .A(n12802), .B(n12805), .Z(n12803) );
  XOR U12848 ( .A(n12798), .B(n12766), .Z(n12799) );
  XOR U12849 ( .A(n12806), .B(n12807), .Z(n12766) );
  AND U12850 ( .A(n674), .B(n12808), .Z(n12806) );
  XOR U12851 ( .A(n12809), .B(n12807), .Z(n12808) );
  XNOR U12852 ( .A(n12810), .B(n12811), .Z(n12798) );
  NAND U12853 ( .A(n12812), .B(n12813), .Z(n12811) );
  XOR U12854 ( .A(n12814), .B(n12790), .Z(n12813) );
  XOR U12855 ( .A(n12804), .B(n12805), .Z(n12790) );
  XOR U12856 ( .A(n12815), .B(n12816), .Z(n12805) );
  ANDN U12857 ( .B(n12817), .A(n12818), .Z(n12815) );
  XOR U12858 ( .A(n12816), .B(n12819), .Z(n12817) );
  XOR U12859 ( .A(n12820), .B(n12821), .Z(n12804) );
  XOR U12860 ( .A(n12822), .B(n12823), .Z(n12821) );
  ANDN U12861 ( .B(n12824), .A(n12825), .Z(n12822) );
  XOR U12862 ( .A(n12826), .B(n12823), .Z(n12824) );
  IV U12863 ( .A(n12802), .Z(n12820) );
  XOR U12864 ( .A(n12827), .B(n12828), .Z(n12802) );
  ANDN U12865 ( .B(n12829), .A(n12830), .Z(n12827) );
  XOR U12866 ( .A(n12828), .B(n12831), .Z(n12829) );
  IV U12867 ( .A(n12810), .Z(n12814) );
  XOR U12868 ( .A(n12810), .B(n12792), .Z(n12812) );
  XOR U12869 ( .A(n12832), .B(n12833), .Z(n12792) );
  AND U12870 ( .A(n674), .B(n12834), .Z(n12832) );
  XOR U12871 ( .A(n12835), .B(n12833), .Z(n12834) );
  NANDN U12872 ( .A(n12794), .B(n12796), .Z(n12810) );
  XOR U12873 ( .A(n12836), .B(n12837), .Z(n12796) );
  AND U12874 ( .A(n674), .B(n12838), .Z(n12836) );
  XOR U12875 ( .A(n12837), .B(n12839), .Z(n12838) );
  XOR U12876 ( .A(n12840), .B(n12841), .Z(n674) );
  AND U12877 ( .A(n12842), .B(n12843), .Z(n12840) );
  XNOR U12878 ( .A(n12841), .B(n12807), .Z(n12843) );
  XNOR U12879 ( .A(n12844), .B(n12845), .Z(n12807) );
  ANDN U12880 ( .B(n12846), .A(n12847), .Z(n12844) );
  XOR U12881 ( .A(n12845), .B(n12848), .Z(n12846) );
  XOR U12882 ( .A(n12841), .B(n12809), .Z(n12842) );
  XOR U12883 ( .A(n12849), .B(n12850), .Z(n12809) );
  AND U12884 ( .A(n678), .B(n12851), .Z(n12849) );
  XOR U12885 ( .A(n12852), .B(n12850), .Z(n12851) );
  XNOR U12886 ( .A(n12853), .B(n12854), .Z(n12841) );
  NAND U12887 ( .A(n12855), .B(n12856), .Z(n12854) );
  XOR U12888 ( .A(n12857), .B(n12833), .Z(n12856) );
  XOR U12889 ( .A(n12847), .B(n12848), .Z(n12833) );
  XOR U12890 ( .A(n12858), .B(n12859), .Z(n12848) );
  ANDN U12891 ( .B(n12860), .A(n12861), .Z(n12858) );
  XOR U12892 ( .A(n12859), .B(n12862), .Z(n12860) );
  XOR U12893 ( .A(n12863), .B(n12864), .Z(n12847) );
  XOR U12894 ( .A(n12865), .B(n12866), .Z(n12864) );
  ANDN U12895 ( .B(n12867), .A(n12868), .Z(n12865) );
  XOR U12896 ( .A(n12869), .B(n12866), .Z(n12867) );
  IV U12897 ( .A(n12845), .Z(n12863) );
  XOR U12898 ( .A(n12870), .B(n12871), .Z(n12845) );
  ANDN U12899 ( .B(n12872), .A(n12873), .Z(n12870) );
  XOR U12900 ( .A(n12871), .B(n12874), .Z(n12872) );
  IV U12901 ( .A(n12853), .Z(n12857) );
  XOR U12902 ( .A(n12853), .B(n12835), .Z(n12855) );
  XOR U12903 ( .A(n12875), .B(n12876), .Z(n12835) );
  AND U12904 ( .A(n678), .B(n12877), .Z(n12875) );
  XOR U12905 ( .A(n12878), .B(n12876), .Z(n12877) );
  NANDN U12906 ( .A(n12837), .B(n12839), .Z(n12853) );
  XOR U12907 ( .A(n12879), .B(n12880), .Z(n12839) );
  AND U12908 ( .A(n678), .B(n12881), .Z(n12879) );
  XOR U12909 ( .A(n12880), .B(n12882), .Z(n12881) );
  XOR U12910 ( .A(n12883), .B(n12884), .Z(n678) );
  AND U12911 ( .A(n12885), .B(n12886), .Z(n12883) );
  XNOR U12912 ( .A(n12884), .B(n12850), .Z(n12886) );
  XNOR U12913 ( .A(n12887), .B(n12888), .Z(n12850) );
  ANDN U12914 ( .B(n12889), .A(n12890), .Z(n12887) );
  XOR U12915 ( .A(n12888), .B(n12891), .Z(n12889) );
  XOR U12916 ( .A(n12884), .B(n12852), .Z(n12885) );
  XOR U12917 ( .A(n12892), .B(n12893), .Z(n12852) );
  AND U12918 ( .A(n682), .B(n12894), .Z(n12892) );
  XOR U12919 ( .A(n12895), .B(n12893), .Z(n12894) );
  XNOR U12920 ( .A(n12896), .B(n12897), .Z(n12884) );
  NAND U12921 ( .A(n12898), .B(n12899), .Z(n12897) );
  XOR U12922 ( .A(n12900), .B(n12876), .Z(n12899) );
  XOR U12923 ( .A(n12890), .B(n12891), .Z(n12876) );
  XOR U12924 ( .A(n12901), .B(n12902), .Z(n12891) );
  ANDN U12925 ( .B(n12903), .A(n12904), .Z(n12901) );
  XOR U12926 ( .A(n12902), .B(n12905), .Z(n12903) );
  XOR U12927 ( .A(n12906), .B(n12907), .Z(n12890) );
  XOR U12928 ( .A(n12908), .B(n12909), .Z(n12907) );
  ANDN U12929 ( .B(n12910), .A(n12911), .Z(n12908) );
  XOR U12930 ( .A(n12912), .B(n12909), .Z(n12910) );
  IV U12931 ( .A(n12888), .Z(n12906) );
  XOR U12932 ( .A(n12913), .B(n12914), .Z(n12888) );
  ANDN U12933 ( .B(n12915), .A(n12916), .Z(n12913) );
  XOR U12934 ( .A(n12914), .B(n12917), .Z(n12915) );
  IV U12935 ( .A(n12896), .Z(n12900) );
  XOR U12936 ( .A(n12896), .B(n12878), .Z(n12898) );
  XOR U12937 ( .A(n12918), .B(n12919), .Z(n12878) );
  AND U12938 ( .A(n682), .B(n12920), .Z(n12918) );
  XOR U12939 ( .A(n12921), .B(n12919), .Z(n12920) );
  NANDN U12940 ( .A(n12880), .B(n12882), .Z(n12896) );
  XOR U12941 ( .A(n12922), .B(n12923), .Z(n12882) );
  AND U12942 ( .A(n682), .B(n12924), .Z(n12922) );
  XOR U12943 ( .A(n12923), .B(n12925), .Z(n12924) );
  XOR U12944 ( .A(n12926), .B(n12927), .Z(n682) );
  AND U12945 ( .A(n12928), .B(n12929), .Z(n12926) );
  XNOR U12946 ( .A(n12927), .B(n12893), .Z(n12929) );
  XNOR U12947 ( .A(n12930), .B(n12931), .Z(n12893) );
  ANDN U12948 ( .B(n12932), .A(n12933), .Z(n12930) );
  XOR U12949 ( .A(n12931), .B(n12934), .Z(n12932) );
  XOR U12950 ( .A(n12927), .B(n12895), .Z(n12928) );
  XOR U12951 ( .A(n12935), .B(n12936), .Z(n12895) );
  AND U12952 ( .A(n686), .B(n12937), .Z(n12935) );
  XOR U12953 ( .A(n12938), .B(n12936), .Z(n12937) );
  XNOR U12954 ( .A(n12939), .B(n12940), .Z(n12927) );
  NAND U12955 ( .A(n12941), .B(n12942), .Z(n12940) );
  XOR U12956 ( .A(n12943), .B(n12919), .Z(n12942) );
  XOR U12957 ( .A(n12933), .B(n12934), .Z(n12919) );
  XOR U12958 ( .A(n12944), .B(n12945), .Z(n12934) );
  ANDN U12959 ( .B(n12946), .A(n12947), .Z(n12944) );
  XOR U12960 ( .A(n12945), .B(n12948), .Z(n12946) );
  XOR U12961 ( .A(n12949), .B(n12950), .Z(n12933) );
  XOR U12962 ( .A(n12951), .B(n12952), .Z(n12950) );
  ANDN U12963 ( .B(n12953), .A(n12954), .Z(n12951) );
  XOR U12964 ( .A(n12955), .B(n12952), .Z(n12953) );
  IV U12965 ( .A(n12931), .Z(n12949) );
  XOR U12966 ( .A(n12956), .B(n12957), .Z(n12931) );
  ANDN U12967 ( .B(n12958), .A(n12959), .Z(n12956) );
  XOR U12968 ( .A(n12957), .B(n12960), .Z(n12958) );
  IV U12969 ( .A(n12939), .Z(n12943) );
  XOR U12970 ( .A(n12939), .B(n12921), .Z(n12941) );
  XOR U12971 ( .A(n12961), .B(n12962), .Z(n12921) );
  AND U12972 ( .A(n686), .B(n12963), .Z(n12961) );
  XOR U12973 ( .A(n12964), .B(n12962), .Z(n12963) );
  NANDN U12974 ( .A(n12923), .B(n12925), .Z(n12939) );
  XOR U12975 ( .A(n12965), .B(n12966), .Z(n12925) );
  AND U12976 ( .A(n686), .B(n12967), .Z(n12965) );
  XOR U12977 ( .A(n12966), .B(n12968), .Z(n12967) );
  XOR U12978 ( .A(n12969), .B(n12970), .Z(n686) );
  AND U12979 ( .A(n12971), .B(n12972), .Z(n12969) );
  XNOR U12980 ( .A(n12970), .B(n12936), .Z(n12972) );
  XNOR U12981 ( .A(n12973), .B(n12974), .Z(n12936) );
  ANDN U12982 ( .B(n12975), .A(n12976), .Z(n12973) );
  XOR U12983 ( .A(n12974), .B(n12977), .Z(n12975) );
  XOR U12984 ( .A(n12970), .B(n12938), .Z(n12971) );
  XOR U12985 ( .A(n12978), .B(n12979), .Z(n12938) );
  AND U12986 ( .A(n690), .B(n12980), .Z(n12978) );
  XOR U12987 ( .A(n12981), .B(n12979), .Z(n12980) );
  XNOR U12988 ( .A(n12982), .B(n12983), .Z(n12970) );
  NAND U12989 ( .A(n12984), .B(n12985), .Z(n12983) );
  XOR U12990 ( .A(n12986), .B(n12962), .Z(n12985) );
  XOR U12991 ( .A(n12976), .B(n12977), .Z(n12962) );
  XOR U12992 ( .A(n12987), .B(n12988), .Z(n12977) );
  ANDN U12993 ( .B(n12989), .A(n12990), .Z(n12987) );
  XOR U12994 ( .A(n12988), .B(n12991), .Z(n12989) );
  XOR U12995 ( .A(n12992), .B(n12993), .Z(n12976) );
  XOR U12996 ( .A(n12994), .B(n12995), .Z(n12993) );
  ANDN U12997 ( .B(n12996), .A(n12997), .Z(n12994) );
  XOR U12998 ( .A(n12998), .B(n12995), .Z(n12996) );
  IV U12999 ( .A(n12974), .Z(n12992) );
  XOR U13000 ( .A(n12999), .B(n13000), .Z(n12974) );
  ANDN U13001 ( .B(n13001), .A(n13002), .Z(n12999) );
  XOR U13002 ( .A(n13000), .B(n13003), .Z(n13001) );
  IV U13003 ( .A(n12982), .Z(n12986) );
  XOR U13004 ( .A(n12982), .B(n12964), .Z(n12984) );
  XOR U13005 ( .A(n13004), .B(n13005), .Z(n12964) );
  AND U13006 ( .A(n690), .B(n13006), .Z(n13004) );
  XOR U13007 ( .A(n13007), .B(n13005), .Z(n13006) );
  NANDN U13008 ( .A(n12966), .B(n12968), .Z(n12982) );
  XOR U13009 ( .A(n13008), .B(n13009), .Z(n12968) );
  AND U13010 ( .A(n690), .B(n13010), .Z(n13008) );
  XOR U13011 ( .A(n13009), .B(n13011), .Z(n13010) );
  XOR U13012 ( .A(n13012), .B(n13013), .Z(n690) );
  AND U13013 ( .A(n13014), .B(n13015), .Z(n13012) );
  XNOR U13014 ( .A(n13013), .B(n12979), .Z(n13015) );
  XNOR U13015 ( .A(n13016), .B(n13017), .Z(n12979) );
  ANDN U13016 ( .B(n13018), .A(n13019), .Z(n13016) );
  XOR U13017 ( .A(n13017), .B(n13020), .Z(n13018) );
  XOR U13018 ( .A(n13013), .B(n12981), .Z(n13014) );
  XOR U13019 ( .A(n13021), .B(n13022), .Z(n12981) );
  AND U13020 ( .A(n694), .B(n13023), .Z(n13021) );
  XOR U13021 ( .A(n13024), .B(n13022), .Z(n13023) );
  XNOR U13022 ( .A(n13025), .B(n13026), .Z(n13013) );
  NAND U13023 ( .A(n13027), .B(n13028), .Z(n13026) );
  XOR U13024 ( .A(n13029), .B(n13005), .Z(n13028) );
  XOR U13025 ( .A(n13019), .B(n13020), .Z(n13005) );
  XOR U13026 ( .A(n13030), .B(n13031), .Z(n13020) );
  ANDN U13027 ( .B(n13032), .A(n13033), .Z(n13030) );
  XOR U13028 ( .A(n13031), .B(n13034), .Z(n13032) );
  XOR U13029 ( .A(n13035), .B(n13036), .Z(n13019) );
  XOR U13030 ( .A(n13037), .B(n13038), .Z(n13036) );
  ANDN U13031 ( .B(n13039), .A(n13040), .Z(n13037) );
  XOR U13032 ( .A(n13041), .B(n13038), .Z(n13039) );
  IV U13033 ( .A(n13017), .Z(n13035) );
  XOR U13034 ( .A(n13042), .B(n13043), .Z(n13017) );
  ANDN U13035 ( .B(n13044), .A(n13045), .Z(n13042) );
  XOR U13036 ( .A(n13043), .B(n13046), .Z(n13044) );
  IV U13037 ( .A(n13025), .Z(n13029) );
  XOR U13038 ( .A(n13025), .B(n13007), .Z(n13027) );
  XOR U13039 ( .A(n13047), .B(n13048), .Z(n13007) );
  AND U13040 ( .A(n694), .B(n13049), .Z(n13047) );
  XOR U13041 ( .A(n13050), .B(n13048), .Z(n13049) );
  NANDN U13042 ( .A(n13009), .B(n13011), .Z(n13025) );
  XOR U13043 ( .A(n13051), .B(n13052), .Z(n13011) );
  AND U13044 ( .A(n694), .B(n13053), .Z(n13051) );
  XOR U13045 ( .A(n13052), .B(n13054), .Z(n13053) );
  XOR U13046 ( .A(n13055), .B(n13056), .Z(n694) );
  AND U13047 ( .A(n13057), .B(n13058), .Z(n13055) );
  XNOR U13048 ( .A(n13056), .B(n13022), .Z(n13058) );
  XNOR U13049 ( .A(n13059), .B(n13060), .Z(n13022) );
  ANDN U13050 ( .B(n13061), .A(n13062), .Z(n13059) );
  XOR U13051 ( .A(n13060), .B(n13063), .Z(n13061) );
  XOR U13052 ( .A(n13056), .B(n13024), .Z(n13057) );
  XOR U13053 ( .A(n13064), .B(n13065), .Z(n13024) );
  AND U13054 ( .A(n698), .B(n13066), .Z(n13064) );
  XOR U13055 ( .A(n13067), .B(n13065), .Z(n13066) );
  XNOR U13056 ( .A(n13068), .B(n13069), .Z(n13056) );
  NAND U13057 ( .A(n13070), .B(n13071), .Z(n13069) );
  XOR U13058 ( .A(n13072), .B(n13048), .Z(n13071) );
  XOR U13059 ( .A(n13062), .B(n13063), .Z(n13048) );
  XOR U13060 ( .A(n13073), .B(n13074), .Z(n13063) );
  ANDN U13061 ( .B(n13075), .A(n13076), .Z(n13073) );
  XOR U13062 ( .A(n13074), .B(n13077), .Z(n13075) );
  XOR U13063 ( .A(n13078), .B(n13079), .Z(n13062) );
  XOR U13064 ( .A(n13080), .B(n13081), .Z(n13079) );
  ANDN U13065 ( .B(n13082), .A(n13083), .Z(n13080) );
  XOR U13066 ( .A(n13084), .B(n13081), .Z(n13082) );
  IV U13067 ( .A(n13060), .Z(n13078) );
  XOR U13068 ( .A(n13085), .B(n13086), .Z(n13060) );
  ANDN U13069 ( .B(n13087), .A(n13088), .Z(n13085) );
  XOR U13070 ( .A(n13086), .B(n13089), .Z(n13087) );
  IV U13071 ( .A(n13068), .Z(n13072) );
  XOR U13072 ( .A(n13068), .B(n13050), .Z(n13070) );
  XOR U13073 ( .A(n13090), .B(n13091), .Z(n13050) );
  AND U13074 ( .A(n698), .B(n13092), .Z(n13090) );
  XOR U13075 ( .A(n13093), .B(n13091), .Z(n13092) );
  NANDN U13076 ( .A(n13052), .B(n13054), .Z(n13068) );
  XOR U13077 ( .A(n13094), .B(n13095), .Z(n13054) );
  AND U13078 ( .A(n698), .B(n13096), .Z(n13094) );
  XOR U13079 ( .A(n13095), .B(n13097), .Z(n13096) );
  XOR U13080 ( .A(n13098), .B(n13099), .Z(n698) );
  AND U13081 ( .A(n13100), .B(n13101), .Z(n13098) );
  XNOR U13082 ( .A(n13099), .B(n13065), .Z(n13101) );
  XNOR U13083 ( .A(n13102), .B(n13103), .Z(n13065) );
  ANDN U13084 ( .B(n13104), .A(n13105), .Z(n13102) );
  XOR U13085 ( .A(n13103), .B(n13106), .Z(n13104) );
  XOR U13086 ( .A(n13099), .B(n13067), .Z(n13100) );
  XOR U13087 ( .A(n13107), .B(n13108), .Z(n13067) );
  AND U13088 ( .A(n702), .B(n13109), .Z(n13107) );
  XOR U13089 ( .A(n13110), .B(n13108), .Z(n13109) );
  XNOR U13090 ( .A(n13111), .B(n13112), .Z(n13099) );
  NAND U13091 ( .A(n13113), .B(n13114), .Z(n13112) );
  XOR U13092 ( .A(n13115), .B(n13091), .Z(n13114) );
  XOR U13093 ( .A(n13105), .B(n13106), .Z(n13091) );
  XOR U13094 ( .A(n13116), .B(n13117), .Z(n13106) );
  ANDN U13095 ( .B(n13118), .A(n13119), .Z(n13116) );
  XOR U13096 ( .A(n13117), .B(n13120), .Z(n13118) );
  XOR U13097 ( .A(n13121), .B(n13122), .Z(n13105) );
  XOR U13098 ( .A(n13123), .B(n13124), .Z(n13122) );
  ANDN U13099 ( .B(n13125), .A(n13126), .Z(n13123) );
  XOR U13100 ( .A(n13127), .B(n13124), .Z(n13125) );
  IV U13101 ( .A(n13103), .Z(n13121) );
  XOR U13102 ( .A(n13128), .B(n13129), .Z(n13103) );
  ANDN U13103 ( .B(n13130), .A(n13131), .Z(n13128) );
  XOR U13104 ( .A(n13129), .B(n13132), .Z(n13130) );
  IV U13105 ( .A(n13111), .Z(n13115) );
  XOR U13106 ( .A(n13111), .B(n13093), .Z(n13113) );
  XOR U13107 ( .A(n13133), .B(n13134), .Z(n13093) );
  AND U13108 ( .A(n702), .B(n13135), .Z(n13133) );
  XOR U13109 ( .A(n13136), .B(n13134), .Z(n13135) );
  NANDN U13110 ( .A(n13095), .B(n13097), .Z(n13111) );
  XOR U13111 ( .A(n13137), .B(n13138), .Z(n13097) );
  AND U13112 ( .A(n702), .B(n13139), .Z(n13137) );
  XOR U13113 ( .A(n13138), .B(n13140), .Z(n13139) );
  XOR U13114 ( .A(n13141), .B(n13142), .Z(n702) );
  AND U13115 ( .A(n13143), .B(n13144), .Z(n13141) );
  XNOR U13116 ( .A(n13142), .B(n13108), .Z(n13144) );
  XNOR U13117 ( .A(n13145), .B(n13146), .Z(n13108) );
  ANDN U13118 ( .B(n13147), .A(n13148), .Z(n13145) );
  XOR U13119 ( .A(n13146), .B(n13149), .Z(n13147) );
  XOR U13120 ( .A(n13142), .B(n13110), .Z(n13143) );
  XOR U13121 ( .A(n13150), .B(n13151), .Z(n13110) );
  AND U13122 ( .A(n706), .B(n13152), .Z(n13150) );
  XOR U13123 ( .A(n13153), .B(n13151), .Z(n13152) );
  XNOR U13124 ( .A(n13154), .B(n13155), .Z(n13142) );
  NAND U13125 ( .A(n13156), .B(n13157), .Z(n13155) );
  XOR U13126 ( .A(n13158), .B(n13134), .Z(n13157) );
  XOR U13127 ( .A(n13148), .B(n13149), .Z(n13134) );
  XOR U13128 ( .A(n13159), .B(n13160), .Z(n13149) );
  ANDN U13129 ( .B(n13161), .A(n13162), .Z(n13159) );
  XOR U13130 ( .A(n13160), .B(n13163), .Z(n13161) );
  XOR U13131 ( .A(n13164), .B(n13165), .Z(n13148) );
  XOR U13132 ( .A(n13166), .B(n13167), .Z(n13165) );
  ANDN U13133 ( .B(n13168), .A(n13169), .Z(n13166) );
  XOR U13134 ( .A(n13170), .B(n13167), .Z(n13168) );
  IV U13135 ( .A(n13146), .Z(n13164) );
  XOR U13136 ( .A(n13171), .B(n13172), .Z(n13146) );
  ANDN U13137 ( .B(n13173), .A(n13174), .Z(n13171) );
  XOR U13138 ( .A(n13172), .B(n13175), .Z(n13173) );
  IV U13139 ( .A(n13154), .Z(n13158) );
  XOR U13140 ( .A(n13154), .B(n13136), .Z(n13156) );
  XOR U13141 ( .A(n13176), .B(n13177), .Z(n13136) );
  AND U13142 ( .A(n706), .B(n13178), .Z(n13176) );
  XOR U13143 ( .A(n13179), .B(n13177), .Z(n13178) );
  NANDN U13144 ( .A(n13138), .B(n13140), .Z(n13154) );
  XOR U13145 ( .A(n13180), .B(n13181), .Z(n13140) );
  AND U13146 ( .A(n706), .B(n13182), .Z(n13180) );
  XOR U13147 ( .A(n13181), .B(n13183), .Z(n13182) );
  XOR U13148 ( .A(n13184), .B(n13185), .Z(n706) );
  AND U13149 ( .A(n13186), .B(n13187), .Z(n13184) );
  XNOR U13150 ( .A(n13185), .B(n13151), .Z(n13187) );
  XNOR U13151 ( .A(n13188), .B(n13189), .Z(n13151) );
  ANDN U13152 ( .B(n13190), .A(n13191), .Z(n13188) );
  XOR U13153 ( .A(n13189), .B(n13192), .Z(n13190) );
  XOR U13154 ( .A(n13185), .B(n13153), .Z(n13186) );
  XOR U13155 ( .A(n13193), .B(n13194), .Z(n13153) );
  AND U13156 ( .A(n710), .B(n13195), .Z(n13193) );
  XOR U13157 ( .A(n13196), .B(n13194), .Z(n13195) );
  XNOR U13158 ( .A(n13197), .B(n13198), .Z(n13185) );
  NAND U13159 ( .A(n13199), .B(n13200), .Z(n13198) );
  XOR U13160 ( .A(n13201), .B(n13177), .Z(n13200) );
  XOR U13161 ( .A(n13191), .B(n13192), .Z(n13177) );
  XOR U13162 ( .A(n13202), .B(n13203), .Z(n13192) );
  ANDN U13163 ( .B(n13204), .A(n13205), .Z(n13202) );
  XOR U13164 ( .A(n13203), .B(n13206), .Z(n13204) );
  XOR U13165 ( .A(n13207), .B(n13208), .Z(n13191) );
  XOR U13166 ( .A(n13209), .B(n13210), .Z(n13208) );
  ANDN U13167 ( .B(n13211), .A(n13212), .Z(n13209) );
  XOR U13168 ( .A(n13213), .B(n13210), .Z(n13211) );
  IV U13169 ( .A(n13189), .Z(n13207) );
  XOR U13170 ( .A(n13214), .B(n13215), .Z(n13189) );
  ANDN U13171 ( .B(n13216), .A(n13217), .Z(n13214) );
  XOR U13172 ( .A(n13215), .B(n13218), .Z(n13216) );
  IV U13173 ( .A(n13197), .Z(n13201) );
  XOR U13174 ( .A(n13197), .B(n13179), .Z(n13199) );
  XOR U13175 ( .A(n13219), .B(n13220), .Z(n13179) );
  AND U13176 ( .A(n710), .B(n13221), .Z(n13219) );
  XOR U13177 ( .A(n13222), .B(n13220), .Z(n13221) );
  NANDN U13178 ( .A(n13181), .B(n13183), .Z(n13197) );
  XOR U13179 ( .A(n13223), .B(n13224), .Z(n13183) );
  AND U13180 ( .A(n710), .B(n13225), .Z(n13223) );
  XOR U13181 ( .A(n13224), .B(n13226), .Z(n13225) );
  XOR U13182 ( .A(n13227), .B(n13228), .Z(n710) );
  AND U13183 ( .A(n13229), .B(n13230), .Z(n13227) );
  XNOR U13184 ( .A(n13228), .B(n13194), .Z(n13230) );
  XNOR U13185 ( .A(n13231), .B(n13232), .Z(n13194) );
  ANDN U13186 ( .B(n13233), .A(n13234), .Z(n13231) );
  XOR U13187 ( .A(n13232), .B(n13235), .Z(n13233) );
  XOR U13188 ( .A(n13228), .B(n13196), .Z(n13229) );
  XOR U13189 ( .A(n13236), .B(n13237), .Z(n13196) );
  AND U13190 ( .A(n714), .B(n13238), .Z(n13236) );
  XOR U13191 ( .A(n13239), .B(n13237), .Z(n13238) );
  XNOR U13192 ( .A(n13240), .B(n13241), .Z(n13228) );
  NAND U13193 ( .A(n13242), .B(n13243), .Z(n13241) );
  XOR U13194 ( .A(n13244), .B(n13220), .Z(n13243) );
  XOR U13195 ( .A(n13234), .B(n13235), .Z(n13220) );
  XOR U13196 ( .A(n13245), .B(n13246), .Z(n13235) );
  ANDN U13197 ( .B(n13247), .A(n13248), .Z(n13245) );
  XOR U13198 ( .A(n13246), .B(n13249), .Z(n13247) );
  XOR U13199 ( .A(n13250), .B(n13251), .Z(n13234) );
  XOR U13200 ( .A(n13252), .B(n13253), .Z(n13251) );
  ANDN U13201 ( .B(n13254), .A(n13255), .Z(n13252) );
  XOR U13202 ( .A(n13256), .B(n13253), .Z(n13254) );
  IV U13203 ( .A(n13232), .Z(n13250) );
  XOR U13204 ( .A(n13257), .B(n13258), .Z(n13232) );
  ANDN U13205 ( .B(n13259), .A(n13260), .Z(n13257) );
  XOR U13206 ( .A(n13258), .B(n13261), .Z(n13259) );
  IV U13207 ( .A(n13240), .Z(n13244) );
  XOR U13208 ( .A(n13240), .B(n13222), .Z(n13242) );
  XOR U13209 ( .A(n13262), .B(n13263), .Z(n13222) );
  AND U13210 ( .A(n714), .B(n13264), .Z(n13262) );
  XOR U13211 ( .A(n13265), .B(n13263), .Z(n13264) );
  NANDN U13212 ( .A(n13224), .B(n13226), .Z(n13240) );
  XOR U13213 ( .A(n13266), .B(n13267), .Z(n13226) );
  AND U13214 ( .A(n714), .B(n13268), .Z(n13266) );
  XOR U13215 ( .A(n13267), .B(n13269), .Z(n13268) );
  XOR U13216 ( .A(n13270), .B(n13271), .Z(n714) );
  AND U13217 ( .A(n13272), .B(n13273), .Z(n13270) );
  XNOR U13218 ( .A(n13271), .B(n13237), .Z(n13273) );
  XNOR U13219 ( .A(n13274), .B(n13275), .Z(n13237) );
  ANDN U13220 ( .B(n13276), .A(n13277), .Z(n13274) );
  XOR U13221 ( .A(n13275), .B(n13278), .Z(n13276) );
  XOR U13222 ( .A(n13271), .B(n13239), .Z(n13272) );
  XOR U13223 ( .A(n13279), .B(n13280), .Z(n13239) );
  AND U13224 ( .A(n718), .B(n13281), .Z(n13279) );
  XOR U13225 ( .A(n13282), .B(n13280), .Z(n13281) );
  XNOR U13226 ( .A(n13283), .B(n13284), .Z(n13271) );
  NAND U13227 ( .A(n13285), .B(n13286), .Z(n13284) );
  XOR U13228 ( .A(n13287), .B(n13263), .Z(n13286) );
  XOR U13229 ( .A(n13277), .B(n13278), .Z(n13263) );
  XOR U13230 ( .A(n13288), .B(n13289), .Z(n13278) );
  ANDN U13231 ( .B(n13290), .A(n13291), .Z(n13288) );
  XOR U13232 ( .A(n13289), .B(n13292), .Z(n13290) );
  XOR U13233 ( .A(n13293), .B(n13294), .Z(n13277) );
  XOR U13234 ( .A(n13295), .B(n13296), .Z(n13294) );
  ANDN U13235 ( .B(n13297), .A(n13298), .Z(n13295) );
  XOR U13236 ( .A(n13299), .B(n13296), .Z(n13297) );
  IV U13237 ( .A(n13275), .Z(n13293) );
  XOR U13238 ( .A(n13300), .B(n13301), .Z(n13275) );
  ANDN U13239 ( .B(n13302), .A(n13303), .Z(n13300) );
  XOR U13240 ( .A(n13301), .B(n13304), .Z(n13302) );
  IV U13241 ( .A(n13283), .Z(n13287) );
  XOR U13242 ( .A(n13283), .B(n13265), .Z(n13285) );
  XOR U13243 ( .A(n13305), .B(n13306), .Z(n13265) );
  AND U13244 ( .A(n718), .B(n13307), .Z(n13305) );
  XOR U13245 ( .A(n13308), .B(n13306), .Z(n13307) );
  NANDN U13246 ( .A(n13267), .B(n13269), .Z(n13283) );
  XOR U13247 ( .A(n13309), .B(n13310), .Z(n13269) );
  AND U13248 ( .A(n718), .B(n13311), .Z(n13309) );
  XOR U13249 ( .A(n13310), .B(n13312), .Z(n13311) );
  XOR U13250 ( .A(n13313), .B(n13314), .Z(n718) );
  AND U13251 ( .A(n13315), .B(n13316), .Z(n13313) );
  XNOR U13252 ( .A(n13314), .B(n13280), .Z(n13316) );
  XNOR U13253 ( .A(n13317), .B(n13318), .Z(n13280) );
  ANDN U13254 ( .B(n13319), .A(n13320), .Z(n13317) );
  XOR U13255 ( .A(n13318), .B(n13321), .Z(n13319) );
  XOR U13256 ( .A(n13314), .B(n13282), .Z(n13315) );
  XOR U13257 ( .A(n13322), .B(n13323), .Z(n13282) );
  AND U13258 ( .A(n722), .B(n13324), .Z(n13322) );
  XOR U13259 ( .A(n13325), .B(n13323), .Z(n13324) );
  XNOR U13260 ( .A(n13326), .B(n13327), .Z(n13314) );
  NAND U13261 ( .A(n13328), .B(n13329), .Z(n13327) );
  XOR U13262 ( .A(n13330), .B(n13306), .Z(n13329) );
  XOR U13263 ( .A(n13320), .B(n13321), .Z(n13306) );
  XOR U13264 ( .A(n13331), .B(n13332), .Z(n13321) );
  ANDN U13265 ( .B(n13333), .A(n13334), .Z(n13331) );
  XOR U13266 ( .A(n13332), .B(n13335), .Z(n13333) );
  XOR U13267 ( .A(n13336), .B(n13337), .Z(n13320) );
  XOR U13268 ( .A(n13338), .B(n13339), .Z(n13337) );
  ANDN U13269 ( .B(n13340), .A(n13341), .Z(n13338) );
  XOR U13270 ( .A(n13342), .B(n13339), .Z(n13340) );
  IV U13271 ( .A(n13318), .Z(n13336) );
  XOR U13272 ( .A(n13343), .B(n13344), .Z(n13318) );
  ANDN U13273 ( .B(n13345), .A(n13346), .Z(n13343) );
  XOR U13274 ( .A(n13344), .B(n13347), .Z(n13345) );
  IV U13275 ( .A(n13326), .Z(n13330) );
  XOR U13276 ( .A(n13326), .B(n13308), .Z(n13328) );
  XOR U13277 ( .A(n13348), .B(n13349), .Z(n13308) );
  AND U13278 ( .A(n722), .B(n13350), .Z(n13348) );
  XOR U13279 ( .A(n13351), .B(n13349), .Z(n13350) );
  NANDN U13280 ( .A(n13310), .B(n13312), .Z(n13326) );
  XOR U13281 ( .A(n13352), .B(n13353), .Z(n13312) );
  AND U13282 ( .A(n722), .B(n13354), .Z(n13352) );
  XOR U13283 ( .A(n13353), .B(n13355), .Z(n13354) );
  XOR U13284 ( .A(n13356), .B(n13357), .Z(n722) );
  AND U13285 ( .A(n13358), .B(n13359), .Z(n13356) );
  XNOR U13286 ( .A(n13357), .B(n13323), .Z(n13359) );
  XNOR U13287 ( .A(n13360), .B(n13361), .Z(n13323) );
  ANDN U13288 ( .B(n13362), .A(n13363), .Z(n13360) );
  XOR U13289 ( .A(n13361), .B(n13364), .Z(n13362) );
  XOR U13290 ( .A(n13357), .B(n13325), .Z(n13358) );
  XOR U13291 ( .A(n13365), .B(n13366), .Z(n13325) );
  AND U13292 ( .A(n726), .B(n13367), .Z(n13365) );
  XOR U13293 ( .A(n13368), .B(n13366), .Z(n13367) );
  XNOR U13294 ( .A(n13369), .B(n13370), .Z(n13357) );
  NAND U13295 ( .A(n13371), .B(n13372), .Z(n13370) );
  XOR U13296 ( .A(n13373), .B(n13349), .Z(n13372) );
  XOR U13297 ( .A(n13363), .B(n13364), .Z(n13349) );
  XOR U13298 ( .A(n13374), .B(n13375), .Z(n13364) );
  ANDN U13299 ( .B(n13376), .A(n13377), .Z(n13374) );
  XOR U13300 ( .A(n13375), .B(n13378), .Z(n13376) );
  XOR U13301 ( .A(n13379), .B(n13380), .Z(n13363) );
  XOR U13302 ( .A(n13381), .B(n13382), .Z(n13380) );
  ANDN U13303 ( .B(n13383), .A(n13384), .Z(n13381) );
  XOR U13304 ( .A(n13385), .B(n13382), .Z(n13383) );
  IV U13305 ( .A(n13361), .Z(n13379) );
  XOR U13306 ( .A(n13386), .B(n13387), .Z(n13361) );
  ANDN U13307 ( .B(n13388), .A(n13389), .Z(n13386) );
  XOR U13308 ( .A(n13387), .B(n13390), .Z(n13388) );
  IV U13309 ( .A(n13369), .Z(n13373) );
  XOR U13310 ( .A(n13369), .B(n13351), .Z(n13371) );
  XOR U13311 ( .A(n13391), .B(n13392), .Z(n13351) );
  AND U13312 ( .A(n726), .B(n13393), .Z(n13391) );
  XOR U13313 ( .A(n13394), .B(n13392), .Z(n13393) );
  NANDN U13314 ( .A(n13353), .B(n13355), .Z(n13369) );
  XOR U13315 ( .A(n13395), .B(n13396), .Z(n13355) );
  AND U13316 ( .A(n726), .B(n13397), .Z(n13395) );
  XOR U13317 ( .A(n13396), .B(n13398), .Z(n13397) );
  XOR U13318 ( .A(n13399), .B(n13400), .Z(n726) );
  AND U13319 ( .A(n13401), .B(n13402), .Z(n13399) );
  XNOR U13320 ( .A(n13400), .B(n13366), .Z(n13402) );
  XNOR U13321 ( .A(n13403), .B(n13404), .Z(n13366) );
  ANDN U13322 ( .B(n13405), .A(n13406), .Z(n13403) );
  XOR U13323 ( .A(n13404), .B(n13407), .Z(n13405) );
  XOR U13324 ( .A(n13400), .B(n13368), .Z(n13401) );
  XOR U13325 ( .A(n13408), .B(n13409), .Z(n13368) );
  AND U13326 ( .A(n730), .B(n13410), .Z(n13408) );
  XOR U13327 ( .A(n13411), .B(n13409), .Z(n13410) );
  XNOR U13328 ( .A(n13412), .B(n13413), .Z(n13400) );
  NAND U13329 ( .A(n13414), .B(n13415), .Z(n13413) );
  XOR U13330 ( .A(n13416), .B(n13392), .Z(n13415) );
  XOR U13331 ( .A(n13406), .B(n13407), .Z(n13392) );
  XOR U13332 ( .A(n13417), .B(n13418), .Z(n13407) );
  ANDN U13333 ( .B(n13419), .A(n13420), .Z(n13417) );
  XOR U13334 ( .A(n13418), .B(n13421), .Z(n13419) );
  XOR U13335 ( .A(n13422), .B(n13423), .Z(n13406) );
  XOR U13336 ( .A(n13424), .B(n13425), .Z(n13423) );
  ANDN U13337 ( .B(n13426), .A(n13427), .Z(n13424) );
  XOR U13338 ( .A(n13428), .B(n13425), .Z(n13426) );
  IV U13339 ( .A(n13404), .Z(n13422) );
  XOR U13340 ( .A(n13429), .B(n13430), .Z(n13404) );
  ANDN U13341 ( .B(n13431), .A(n13432), .Z(n13429) );
  XOR U13342 ( .A(n13430), .B(n13433), .Z(n13431) );
  IV U13343 ( .A(n13412), .Z(n13416) );
  XOR U13344 ( .A(n13412), .B(n13394), .Z(n13414) );
  XOR U13345 ( .A(n13434), .B(n13435), .Z(n13394) );
  AND U13346 ( .A(n730), .B(n13436), .Z(n13434) );
  XOR U13347 ( .A(n13437), .B(n13435), .Z(n13436) );
  NANDN U13348 ( .A(n13396), .B(n13398), .Z(n13412) );
  XOR U13349 ( .A(n13438), .B(n13439), .Z(n13398) );
  AND U13350 ( .A(n730), .B(n13440), .Z(n13438) );
  XOR U13351 ( .A(n13439), .B(n13441), .Z(n13440) );
  XOR U13352 ( .A(n13442), .B(n13443), .Z(n730) );
  AND U13353 ( .A(n13444), .B(n13445), .Z(n13442) );
  XNOR U13354 ( .A(n13443), .B(n13409), .Z(n13445) );
  XNOR U13355 ( .A(n13446), .B(n13447), .Z(n13409) );
  ANDN U13356 ( .B(n13448), .A(n13449), .Z(n13446) );
  XOR U13357 ( .A(n13447), .B(n13450), .Z(n13448) );
  XOR U13358 ( .A(n13443), .B(n13411), .Z(n13444) );
  XOR U13359 ( .A(n13451), .B(n13452), .Z(n13411) );
  AND U13360 ( .A(n734), .B(n13453), .Z(n13451) );
  XOR U13361 ( .A(n13454), .B(n13452), .Z(n13453) );
  XNOR U13362 ( .A(n13455), .B(n13456), .Z(n13443) );
  NAND U13363 ( .A(n13457), .B(n13458), .Z(n13456) );
  XOR U13364 ( .A(n13459), .B(n13435), .Z(n13458) );
  XOR U13365 ( .A(n13449), .B(n13450), .Z(n13435) );
  XOR U13366 ( .A(n13460), .B(n13461), .Z(n13450) );
  ANDN U13367 ( .B(n13462), .A(n13463), .Z(n13460) );
  XOR U13368 ( .A(n13461), .B(n13464), .Z(n13462) );
  XOR U13369 ( .A(n13465), .B(n13466), .Z(n13449) );
  XOR U13370 ( .A(n13467), .B(n13468), .Z(n13466) );
  ANDN U13371 ( .B(n13469), .A(n13470), .Z(n13467) );
  XOR U13372 ( .A(n13471), .B(n13468), .Z(n13469) );
  IV U13373 ( .A(n13447), .Z(n13465) );
  XOR U13374 ( .A(n13472), .B(n13473), .Z(n13447) );
  ANDN U13375 ( .B(n13474), .A(n13475), .Z(n13472) );
  XOR U13376 ( .A(n13473), .B(n13476), .Z(n13474) );
  IV U13377 ( .A(n13455), .Z(n13459) );
  XOR U13378 ( .A(n13455), .B(n13437), .Z(n13457) );
  XOR U13379 ( .A(n13477), .B(n13478), .Z(n13437) );
  AND U13380 ( .A(n734), .B(n13479), .Z(n13477) );
  XOR U13381 ( .A(n13480), .B(n13478), .Z(n13479) );
  NANDN U13382 ( .A(n13439), .B(n13441), .Z(n13455) );
  XOR U13383 ( .A(n13481), .B(n13482), .Z(n13441) );
  AND U13384 ( .A(n734), .B(n13483), .Z(n13481) );
  XOR U13385 ( .A(n13482), .B(n13484), .Z(n13483) );
  XOR U13386 ( .A(n13485), .B(n13486), .Z(n734) );
  AND U13387 ( .A(n13487), .B(n13488), .Z(n13485) );
  XNOR U13388 ( .A(n13486), .B(n13452), .Z(n13488) );
  XNOR U13389 ( .A(n13489), .B(n13490), .Z(n13452) );
  ANDN U13390 ( .B(n13491), .A(n13492), .Z(n13489) );
  XOR U13391 ( .A(n13490), .B(n13493), .Z(n13491) );
  XOR U13392 ( .A(n13486), .B(n13454), .Z(n13487) );
  XOR U13393 ( .A(n13494), .B(n13495), .Z(n13454) );
  AND U13394 ( .A(n738), .B(n13496), .Z(n13494) );
  XOR U13395 ( .A(n13497), .B(n13495), .Z(n13496) );
  XNOR U13396 ( .A(n13498), .B(n13499), .Z(n13486) );
  NAND U13397 ( .A(n13500), .B(n13501), .Z(n13499) );
  XOR U13398 ( .A(n13502), .B(n13478), .Z(n13501) );
  XOR U13399 ( .A(n13492), .B(n13493), .Z(n13478) );
  XOR U13400 ( .A(n13503), .B(n13504), .Z(n13493) );
  ANDN U13401 ( .B(n13505), .A(n13506), .Z(n13503) );
  XOR U13402 ( .A(n13504), .B(n13507), .Z(n13505) );
  XOR U13403 ( .A(n13508), .B(n13509), .Z(n13492) );
  XOR U13404 ( .A(n13510), .B(n13511), .Z(n13509) );
  ANDN U13405 ( .B(n13512), .A(n13513), .Z(n13510) );
  XOR U13406 ( .A(n13514), .B(n13511), .Z(n13512) );
  IV U13407 ( .A(n13490), .Z(n13508) );
  XOR U13408 ( .A(n13515), .B(n13516), .Z(n13490) );
  ANDN U13409 ( .B(n13517), .A(n13518), .Z(n13515) );
  XOR U13410 ( .A(n13516), .B(n13519), .Z(n13517) );
  IV U13411 ( .A(n13498), .Z(n13502) );
  XOR U13412 ( .A(n13498), .B(n13480), .Z(n13500) );
  XOR U13413 ( .A(n13520), .B(n13521), .Z(n13480) );
  AND U13414 ( .A(n738), .B(n13522), .Z(n13520) );
  XOR U13415 ( .A(n13523), .B(n13521), .Z(n13522) );
  NANDN U13416 ( .A(n13482), .B(n13484), .Z(n13498) );
  XOR U13417 ( .A(n13524), .B(n13525), .Z(n13484) );
  AND U13418 ( .A(n738), .B(n13526), .Z(n13524) );
  XOR U13419 ( .A(n13525), .B(n13527), .Z(n13526) );
  XOR U13420 ( .A(n13528), .B(n13529), .Z(n738) );
  AND U13421 ( .A(n13530), .B(n13531), .Z(n13528) );
  XNOR U13422 ( .A(n13529), .B(n13495), .Z(n13531) );
  XNOR U13423 ( .A(n13532), .B(n13533), .Z(n13495) );
  ANDN U13424 ( .B(n13534), .A(n13535), .Z(n13532) );
  XOR U13425 ( .A(n13533), .B(n13536), .Z(n13534) );
  XOR U13426 ( .A(n13529), .B(n13497), .Z(n13530) );
  XOR U13427 ( .A(n13537), .B(n13538), .Z(n13497) );
  AND U13428 ( .A(n742), .B(n13539), .Z(n13537) );
  XOR U13429 ( .A(n13540), .B(n13538), .Z(n13539) );
  XNOR U13430 ( .A(n13541), .B(n13542), .Z(n13529) );
  NAND U13431 ( .A(n13543), .B(n13544), .Z(n13542) );
  XOR U13432 ( .A(n13545), .B(n13521), .Z(n13544) );
  XOR U13433 ( .A(n13535), .B(n13536), .Z(n13521) );
  XOR U13434 ( .A(n13546), .B(n13547), .Z(n13536) );
  ANDN U13435 ( .B(n13548), .A(n13549), .Z(n13546) );
  XOR U13436 ( .A(n13547), .B(n13550), .Z(n13548) );
  XOR U13437 ( .A(n13551), .B(n13552), .Z(n13535) );
  XOR U13438 ( .A(n13553), .B(n13554), .Z(n13552) );
  ANDN U13439 ( .B(n13555), .A(n13556), .Z(n13553) );
  XOR U13440 ( .A(n13557), .B(n13554), .Z(n13555) );
  IV U13441 ( .A(n13533), .Z(n13551) );
  XOR U13442 ( .A(n13558), .B(n13559), .Z(n13533) );
  ANDN U13443 ( .B(n13560), .A(n13561), .Z(n13558) );
  XOR U13444 ( .A(n13559), .B(n13562), .Z(n13560) );
  IV U13445 ( .A(n13541), .Z(n13545) );
  XOR U13446 ( .A(n13541), .B(n13523), .Z(n13543) );
  XOR U13447 ( .A(n13563), .B(n13564), .Z(n13523) );
  AND U13448 ( .A(n742), .B(n13565), .Z(n13563) );
  XOR U13449 ( .A(n13566), .B(n13564), .Z(n13565) );
  NANDN U13450 ( .A(n13525), .B(n13527), .Z(n13541) );
  XOR U13451 ( .A(n13567), .B(n13568), .Z(n13527) );
  AND U13452 ( .A(n742), .B(n13569), .Z(n13567) );
  XOR U13453 ( .A(n13568), .B(n13570), .Z(n13569) );
  XOR U13454 ( .A(n13571), .B(n13572), .Z(n742) );
  AND U13455 ( .A(n13573), .B(n13574), .Z(n13571) );
  XNOR U13456 ( .A(n13572), .B(n13538), .Z(n13574) );
  XNOR U13457 ( .A(n13575), .B(n13576), .Z(n13538) );
  ANDN U13458 ( .B(n13577), .A(n13578), .Z(n13575) );
  XOR U13459 ( .A(n13576), .B(n13579), .Z(n13577) );
  XOR U13460 ( .A(n13572), .B(n13540), .Z(n13573) );
  XOR U13461 ( .A(n13580), .B(n13581), .Z(n13540) );
  AND U13462 ( .A(n746), .B(n13582), .Z(n13580) );
  XOR U13463 ( .A(n13583), .B(n13581), .Z(n13582) );
  XNOR U13464 ( .A(n13584), .B(n13585), .Z(n13572) );
  NAND U13465 ( .A(n13586), .B(n13587), .Z(n13585) );
  XOR U13466 ( .A(n13588), .B(n13564), .Z(n13587) );
  XOR U13467 ( .A(n13578), .B(n13579), .Z(n13564) );
  XOR U13468 ( .A(n13589), .B(n13590), .Z(n13579) );
  ANDN U13469 ( .B(n13591), .A(n13592), .Z(n13589) );
  XOR U13470 ( .A(n13590), .B(n13593), .Z(n13591) );
  XOR U13471 ( .A(n13594), .B(n13595), .Z(n13578) );
  XOR U13472 ( .A(n13596), .B(n13597), .Z(n13595) );
  ANDN U13473 ( .B(n13598), .A(n13599), .Z(n13596) );
  XOR U13474 ( .A(n13600), .B(n13597), .Z(n13598) );
  IV U13475 ( .A(n13576), .Z(n13594) );
  XOR U13476 ( .A(n13601), .B(n13602), .Z(n13576) );
  ANDN U13477 ( .B(n13603), .A(n13604), .Z(n13601) );
  XOR U13478 ( .A(n13602), .B(n13605), .Z(n13603) );
  IV U13479 ( .A(n13584), .Z(n13588) );
  XOR U13480 ( .A(n13584), .B(n13566), .Z(n13586) );
  XOR U13481 ( .A(n13606), .B(n13607), .Z(n13566) );
  AND U13482 ( .A(n746), .B(n13608), .Z(n13606) );
  XOR U13483 ( .A(n13609), .B(n13607), .Z(n13608) );
  NANDN U13484 ( .A(n13568), .B(n13570), .Z(n13584) );
  XOR U13485 ( .A(n13610), .B(n13611), .Z(n13570) );
  AND U13486 ( .A(n746), .B(n13612), .Z(n13610) );
  XOR U13487 ( .A(n13611), .B(n13613), .Z(n13612) );
  XOR U13488 ( .A(n13614), .B(n13615), .Z(n746) );
  AND U13489 ( .A(n13616), .B(n13617), .Z(n13614) );
  XNOR U13490 ( .A(n13615), .B(n13581), .Z(n13617) );
  XNOR U13491 ( .A(n13618), .B(n13619), .Z(n13581) );
  ANDN U13492 ( .B(n13620), .A(n13621), .Z(n13618) );
  XOR U13493 ( .A(n13619), .B(n13622), .Z(n13620) );
  XOR U13494 ( .A(n13615), .B(n13583), .Z(n13616) );
  XOR U13495 ( .A(n13623), .B(n13624), .Z(n13583) );
  AND U13496 ( .A(n750), .B(n13625), .Z(n13623) );
  XOR U13497 ( .A(n13626), .B(n13624), .Z(n13625) );
  XNOR U13498 ( .A(n13627), .B(n13628), .Z(n13615) );
  NAND U13499 ( .A(n13629), .B(n13630), .Z(n13628) );
  XOR U13500 ( .A(n13631), .B(n13607), .Z(n13630) );
  XOR U13501 ( .A(n13621), .B(n13622), .Z(n13607) );
  XOR U13502 ( .A(n13632), .B(n13633), .Z(n13622) );
  ANDN U13503 ( .B(n13634), .A(n13635), .Z(n13632) );
  XOR U13504 ( .A(n13633), .B(n13636), .Z(n13634) );
  XOR U13505 ( .A(n13637), .B(n13638), .Z(n13621) );
  XOR U13506 ( .A(n13639), .B(n13640), .Z(n13638) );
  ANDN U13507 ( .B(n13641), .A(n13642), .Z(n13639) );
  XOR U13508 ( .A(n13643), .B(n13640), .Z(n13641) );
  IV U13509 ( .A(n13619), .Z(n13637) );
  XOR U13510 ( .A(n13644), .B(n13645), .Z(n13619) );
  ANDN U13511 ( .B(n13646), .A(n13647), .Z(n13644) );
  XOR U13512 ( .A(n13645), .B(n13648), .Z(n13646) );
  IV U13513 ( .A(n13627), .Z(n13631) );
  XOR U13514 ( .A(n13627), .B(n13609), .Z(n13629) );
  XOR U13515 ( .A(n13649), .B(n13650), .Z(n13609) );
  AND U13516 ( .A(n750), .B(n13651), .Z(n13649) );
  XOR U13517 ( .A(n13652), .B(n13650), .Z(n13651) );
  NANDN U13518 ( .A(n13611), .B(n13613), .Z(n13627) );
  XOR U13519 ( .A(n13653), .B(n13654), .Z(n13613) );
  AND U13520 ( .A(n750), .B(n13655), .Z(n13653) );
  XOR U13521 ( .A(n13654), .B(n13656), .Z(n13655) );
  XOR U13522 ( .A(n13657), .B(n13658), .Z(n750) );
  AND U13523 ( .A(n13659), .B(n13660), .Z(n13657) );
  XNOR U13524 ( .A(n13658), .B(n13624), .Z(n13660) );
  XNOR U13525 ( .A(n13661), .B(n13662), .Z(n13624) );
  ANDN U13526 ( .B(n13663), .A(n13664), .Z(n13661) );
  XOR U13527 ( .A(n13662), .B(n13665), .Z(n13663) );
  XOR U13528 ( .A(n13658), .B(n13626), .Z(n13659) );
  XOR U13529 ( .A(n13666), .B(n13667), .Z(n13626) );
  AND U13530 ( .A(n754), .B(n13668), .Z(n13666) );
  XOR U13531 ( .A(n13669), .B(n13667), .Z(n13668) );
  XNOR U13532 ( .A(n13670), .B(n13671), .Z(n13658) );
  NAND U13533 ( .A(n13672), .B(n13673), .Z(n13671) );
  XOR U13534 ( .A(n13674), .B(n13650), .Z(n13673) );
  XOR U13535 ( .A(n13664), .B(n13665), .Z(n13650) );
  XOR U13536 ( .A(n13675), .B(n13676), .Z(n13665) );
  ANDN U13537 ( .B(n13677), .A(n13678), .Z(n13675) );
  XOR U13538 ( .A(n13676), .B(n13679), .Z(n13677) );
  XOR U13539 ( .A(n13680), .B(n13681), .Z(n13664) );
  XOR U13540 ( .A(n13682), .B(n13683), .Z(n13681) );
  ANDN U13541 ( .B(n13684), .A(n13685), .Z(n13682) );
  XOR U13542 ( .A(n13686), .B(n13683), .Z(n13684) );
  IV U13543 ( .A(n13662), .Z(n13680) );
  XOR U13544 ( .A(n13687), .B(n13688), .Z(n13662) );
  ANDN U13545 ( .B(n13689), .A(n13690), .Z(n13687) );
  XOR U13546 ( .A(n13688), .B(n13691), .Z(n13689) );
  IV U13547 ( .A(n13670), .Z(n13674) );
  XOR U13548 ( .A(n13670), .B(n13652), .Z(n13672) );
  XOR U13549 ( .A(n13692), .B(n13693), .Z(n13652) );
  AND U13550 ( .A(n754), .B(n13694), .Z(n13692) );
  XOR U13551 ( .A(n13695), .B(n13693), .Z(n13694) );
  NANDN U13552 ( .A(n13654), .B(n13656), .Z(n13670) );
  XOR U13553 ( .A(n13696), .B(n13697), .Z(n13656) );
  AND U13554 ( .A(n754), .B(n13698), .Z(n13696) );
  XOR U13555 ( .A(n13697), .B(n13699), .Z(n13698) );
  XOR U13556 ( .A(n13700), .B(n13701), .Z(n754) );
  AND U13557 ( .A(n13702), .B(n13703), .Z(n13700) );
  XNOR U13558 ( .A(n13701), .B(n13667), .Z(n13703) );
  XNOR U13559 ( .A(n13704), .B(n13705), .Z(n13667) );
  ANDN U13560 ( .B(n13706), .A(n13707), .Z(n13704) );
  XOR U13561 ( .A(n13705), .B(n13708), .Z(n13706) );
  XOR U13562 ( .A(n13701), .B(n13669), .Z(n13702) );
  XOR U13563 ( .A(n13709), .B(n13710), .Z(n13669) );
  AND U13564 ( .A(n758), .B(n13711), .Z(n13709) );
  XOR U13565 ( .A(n13712), .B(n13710), .Z(n13711) );
  XNOR U13566 ( .A(n13713), .B(n13714), .Z(n13701) );
  NAND U13567 ( .A(n13715), .B(n13716), .Z(n13714) );
  XOR U13568 ( .A(n13717), .B(n13693), .Z(n13716) );
  XOR U13569 ( .A(n13707), .B(n13708), .Z(n13693) );
  XOR U13570 ( .A(n13718), .B(n13719), .Z(n13708) );
  ANDN U13571 ( .B(n13720), .A(n13721), .Z(n13718) );
  XOR U13572 ( .A(n13719), .B(n13722), .Z(n13720) );
  XOR U13573 ( .A(n13723), .B(n13724), .Z(n13707) );
  XOR U13574 ( .A(n13725), .B(n13726), .Z(n13724) );
  ANDN U13575 ( .B(n13727), .A(n13728), .Z(n13725) );
  XOR U13576 ( .A(n13729), .B(n13726), .Z(n13727) );
  IV U13577 ( .A(n13705), .Z(n13723) );
  XOR U13578 ( .A(n13730), .B(n13731), .Z(n13705) );
  ANDN U13579 ( .B(n13732), .A(n13733), .Z(n13730) );
  XOR U13580 ( .A(n13731), .B(n13734), .Z(n13732) );
  IV U13581 ( .A(n13713), .Z(n13717) );
  XOR U13582 ( .A(n13713), .B(n13695), .Z(n13715) );
  XOR U13583 ( .A(n13735), .B(n13736), .Z(n13695) );
  AND U13584 ( .A(n758), .B(n13737), .Z(n13735) );
  XOR U13585 ( .A(n13738), .B(n13736), .Z(n13737) );
  NANDN U13586 ( .A(n13697), .B(n13699), .Z(n13713) );
  XOR U13587 ( .A(n13739), .B(n13740), .Z(n13699) );
  AND U13588 ( .A(n758), .B(n13741), .Z(n13739) );
  XOR U13589 ( .A(n13740), .B(n13742), .Z(n13741) );
  XOR U13590 ( .A(n13743), .B(n13744), .Z(n758) );
  AND U13591 ( .A(n13745), .B(n13746), .Z(n13743) );
  XNOR U13592 ( .A(n13744), .B(n13710), .Z(n13746) );
  XNOR U13593 ( .A(n13747), .B(n13748), .Z(n13710) );
  ANDN U13594 ( .B(n13749), .A(n13750), .Z(n13747) );
  XOR U13595 ( .A(n13748), .B(n13751), .Z(n13749) );
  XOR U13596 ( .A(n13744), .B(n13712), .Z(n13745) );
  XOR U13597 ( .A(n13752), .B(n13753), .Z(n13712) );
  AND U13598 ( .A(n762), .B(n13754), .Z(n13752) );
  XOR U13599 ( .A(n13755), .B(n13753), .Z(n13754) );
  XNOR U13600 ( .A(n13756), .B(n13757), .Z(n13744) );
  NAND U13601 ( .A(n13758), .B(n13759), .Z(n13757) );
  XOR U13602 ( .A(n13760), .B(n13736), .Z(n13759) );
  XOR U13603 ( .A(n13750), .B(n13751), .Z(n13736) );
  XOR U13604 ( .A(n13761), .B(n13762), .Z(n13751) );
  ANDN U13605 ( .B(n13763), .A(n13764), .Z(n13761) );
  XOR U13606 ( .A(n13762), .B(n13765), .Z(n13763) );
  XOR U13607 ( .A(n13766), .B(n13767), .Z(n13750) );
  XOR U13608 ( .A(n13768), .B(n13769), .Z(n13767) );
  ANDN U13609 ( .B(n13770), .A(n13771), .Z(n13768) );
  XOR U13610 ( .A(n13772), .B(n13769), .Z(n13770) );
  IV U13611 ( .A(n13748), .Z(n13766) );
  XOR U13612 ( .A(n13773), .B(n13774), .Z(n13748) );
  ANDN U13613 ( .B(n13775), .A(n13776), .Z(n13773) );
  XOR U13614 ( .A(n13774), .B(n13777), .Z(n13775) );
  IV U13615 ( .A(n13756), .Z(n13760) );
  XOR U13616 ( .A(n13756), .B(n13738), .Z(n13758) );
  XOR U13617 ( .A(n13778), .B(n13779), .Z(n13738) );
  AND U13618 ( .A(n762), .B(n13780), .Z(n13778) );
  XOR U13619 ( .A(n13781), .B(n13779), .Z(n13780) );
  NANDN U13620 ( .A(n13740), .B(n13742), .Z(n13756) );
  XOR U13621 ( .A(n13782), .B(n13783), .Z(n13742) );
  AND U13622 ( .A(n762), .B(n13784), .Z(n13782) );
  XOR U13623 ( .A(n13783), .B(n13785), .Z(n13784) );
  XOR U13624 ( .A(n13786), .B(n13787), .Z(n762) );
  AND U13625 ( .A(n13788), .B(n13789), .Z(n13786) );
  XNOR U13626 ( .A(n13787), .B(n13753), .Z(n13789) );
  XNOR U13627 ( .A(n13790), .B(n13791), .Z(n13753) );
  ANDN U13628 ( .B(n13792), .A(n13793), .Z(n13790) );
  XOR U13629 ( .A(n13791), .B(n13794), .Z(n13792) );
  XOR U13630 ( .A(n13787), .B(n13755), .Z(n13788) );
  XOR U13631 ( .A(n13795), .B(n13796), .Z(n13755) );
  AND U13632 ( .A(n766), .B(n13797), .Z(n13795) );
  XOR U13633 ( .A(n13798), .B(n13796), .Z(n13797) );
  XNOR U13634 ( .A(n13799), .B(n13800), .Z(n13787) );
  NAND U13635 ( .A(n13801), .B(n13802), .Z(n13800) );
  XOR U13636 ( .A(n13803), .B(n13779), .Z(n13802) );
  XOR U13637 ( .A(n13793), .B(n13794), .Z(n13779) );
  XOR U13638 ( .A(n13804), .B(n13805), .Z(n13794) );
  ANDN U13639 ( .B(n13806), .A(n13807), .Z(n13804) );
  XOR U13640 ( .A(n13805), .B(n13808), .Z(n13806) );
  XOR U13641 ( .A(n13809), .B(n13810), .Z(n13793) );
  XOR U13642 ( .A(n13811), .B(n13812), .Z(n13810) );
  ANDN U13643 ( .B(n13813), .A(n13814), .Z(n13811) );
  XOR U13644 ( .A(n13815), .B(n13812), .Z(n13813) );
  IV U13645 ( .A(n13791), .Z(n13809) );
  XOR U13646 ( .A(n13816), .B(n13817), .Z(n13791) );
  ANDN U13647 ( .B(n13818), .A(n13819), .Z(n13816) );
  XOR U13648 ( .A(n13817), .B(n13820), .Z(n13818) );
  IV U13649 ( .A(n13799), .Z(n13803) );
  XOR U13650 ( .A(n13799), .B(n13781), .Z(n13801) );
  XOR U13651 ( .A(n13821), .B(n13822), .Z(n13781) );
  AND U13652 ( .A(n766), .B(n13823), .Z(n13821) );
  XOR U13653 ( .A(n13824), .B(n13822), .Z(n13823) );
  NANDN U13654 ( .A(n13783), .B(n13785), .Z(n13799) );
  XOR U13655 ( .A(n13825), .B(n13826), .Z(n13785) );
  AND U13656 ( .A(n766), .B(n13827), .Z(n13825) );
  XOR U13657 ( .A(n13826), .B(n13828), .Z(n13827) );
  XOR U13658 ( .A(n13829), .B(n13830), .Z(n766) );
  AND U13659 ( .A(n13831), .B(n13832), .Z(n13829) );
  XNOR U13660 ( .A(n13830), .B(n13796), .Z(n13832) );
  XNOR U13661 ( .A(n13833), .B(n13834), .Z(n13796) );
  ANDN U13662 ( .B(n13835), .A(n13836), .Z(n13833) );
  XOR U13663 ( .A(n13834), .B(n13837), .Z(n13835) );
  XOR U13664 ( .A(n13830), .B(n13798), .Z(n13831) );
  XOR U13665 ( .A(n13838), .B(n13839), .Z(n13798) );
  AND U13666 ( .A(n770), .B(n13840), .Z(n13838) );
  XOR U13667 ( .A(n13841), .B(n13839), .Z(n13840) );
  XNOR U13668 ( .A(n13842), .B(n13843), .Z(n13830) );
  NAND U13669 ( .A(n13844), .B(n13845), .Z(n13843) );
  XOR U13670 ( .A(n13846), .B(n13822), .Z(n13845) );
  XOR U13671 ( .A(n13836), .B(n13837), .Z(n13822) );
  XOR U13672 ( .A(n13847), .B(n13848), .Z(n13837) );
  ANDN U13673 ( .B(n13849), .A(n13850), .Z(n13847) );
  XOR U13674 ( .A(n13848), .B(n13851), .Z(n13849) );
  XOR U13675 ( .A(n13852), .B(n13853), .Z(n13836) );
  XOR U13676 ( .A(n13854), .B(n13855), .Z(n13853) );
  ANDN U13677 ( .B(n13856), .A(n13857), .Z(n13854) );
  XOR U13678 ( .A(n13858), .B(n13855), .Z(n13856) );
  IV U13679 ( .A(n13834), .Z(n13852) );
  XOR U13680 ( .A(n13859), .B(n13860), .Z(n13834) );
  ANDN U13681 ( .B(n13861), .A(n13862), .Z(n13859) );
  XOR U13682 ( .A(n13860), .B(n13863), .Z(n13861) );
  IV U13683 ( .A(n13842), .Z(n13846) );
  XOR U13684 ( .A(n13842), .B(n13824), .Z(n13844) );
  XOR U13685 ( .A(n13864), .B(n13865), .Z(n13824) );
  AND U13686 ( .A(n770), .B(n13866), .Z(n13864) );
  XOR U13687 ( .A(n13867), .B(n13865), .Z(n13866) );
  NANDN U13688 ( .A(n13826), .B(n13828), .Z(n13842) );
  XOR U13689 ( .A(n13868), .B(n13869), .Z(n13828) );
  AND U13690 ( .A(n770), .B(n13870), .Z(n13868) );
  XOR U13691 ( .A(n13869), .B(n13871), .Z(n13870) );
  XOR U13692 ( .A(n13872), .B(n13873), .Z(n770) );
  AND U13693 ( .A(n13874), .B(n13875), .Z(n13872) );
  XNOR U13694 ( .A(n13873), .B(n13839), .Z(n13875) );
  XNOR U13695 ( .A(n13876), .B(n13877), .Z(n13839) );
  ANDN U13696 ( .B(n13878), .A(n13879), .Z(n13876) );
  XOR U13697 ( .A(n13877), .B(n13880), .Z(n13878) );
  XOR U13698 ( .A(n13873), .B(n13841), .Z(n13874) );
  XOR U13699 ( .A(n13881), .B(n13882), .Z(n13841) );
  AND U13700 ( .A(n774), .B(n13883), .Z(n13881) );
  XOR U13701 ( .A(n13884), .B(n13882), .Z(n13883) );
  XNOR U13702 ( .A(n13885), .B(n13886), .Z(n13873) );
  NAND U13703 ( .A(n13887), .B(n13888), .Z(n13886) );
  XOR U13704 ( .A(n13889), .B(n13865), .Z(n13888) );
  XOR U13705 ( .A(n13879), .B(n13880), .Z(n13865) );
  XOR U13706 ( .A(n13890), .B(n13891), .Z(n13880) );
  ANDN U13707 ( .B(n13892), .A(n13893), .Z(n13890) );
  XOR U13708 ( .A(n13891), .B(n13894), .Z(n13892) );
  XOR U13709 ( .A(n13895), .B(n13896), .Z(n13879) );
  XOR U13710 ( .A(n13897), .B(n13898), .Z(n13896) );
  ANDN U13711 ( .B(n13899), .A(n13900), .Z(n13897) );
  XOR U13712 ( .A(n13901), .B(n13898), .Z(n13899) );
  IV U13713 ( .A(n13877), .Z(n13895) );
  XOR U13714 ( .A(n13902), .B(n13903), .Z(n13877) );
  ANDN U13715 ( .B(n13904), .A(n13905), .Z(n13902) );
  XOR U13716 ( .A(n13903), .B(n13906), .Z(n13904) );
  IV U13717 ( .A(n13885), .Z(n13889) );
  XOR U13718 ( .A(n13885), .B(n13867), .Z(n13887) );
  XOR U13719 ( .A(n13907), .B(n13908), .Z(n13867) );
  AND U13720 ( .A(n774), .B(n13909), .Z(n13907) );
  XOR U13721 ( .A(n13910), .B(n13908), .Z(n13909) );
  NANDN U13722 ( .A(n13869), .B(n13871), .Z(n13885) );
  XOR U13723 ( .A(n13911), .B(n13912), .Z(n13871) );
  AND U13724 ( .A(n774), .B(n13913), .Z(n13911) );
  XOR U13725 ( .A(n13912), .B(n13914), .Z(n13913) );
  XOR U13726 ( .A(n13915), .B(n13916), .Z(n774) );
  AND U13727 ( .A(n13917), .B(n13918), .Z(n13915) );
  XNOR U13728 ( .A(n13916), .B(n13882), .Z(n13918) );
  XNOR U13729 ( .A(n13919), .B(n13920), .Z(n13882) );
  ANDN U13730 ( .B(n13921), .A(n13922), .Z(n13919) );
  XOR U13731 ( .A(n13920), .B(n13923), .Z(n13921) );
  XOR U13732 ( .A(n13916), .B(n13884), .Z(n13917) );
  XOR U13733 ( .A(n13924), .B(n13925), .Z(n13884) );
  AND U13734 ( .A(n778), .B(n13926), .Z(n13924) );
  XOR U13735 ( .A(n13927), .B(n13925), .Z(n13926) );
  XNOR U13736 ( .A(n13928), .B(n13929), .Z(n13916) );
  NAND U13737 ( .A(n13930), .B(n13931), .Z(n13929) );
  XOR U13738 ( .A(n13932), .B(n13908), .Z(n13931) );
  XOR U13739 ( .A(n13922), .B(n13923), .Z(n13908) );
  XOR U13740 ( .A(n13933), .B(n13934), .Z(n13923) );
  ANDN U13741 ( .B(n13935), .A(n13936), .Z(n13933) );
  XOR U13742 ( .A(n13934), .B(n13937), .Z(n13935) );
  XOR U13743 ( .A(n13938), .B(n13939), .Z(n13922) );
  XOR U13744 ( .A(n13940), .B(n13941), .Z(n13939) );
  ANDN U13745 ( .B(n13942), .A(n13943), .Z(n13940) );
  XOR U13746 ( .A(n13944), .B(n13941), .Z(n13942) );
  IV U13747 ( .A(n13920), .Z(n13938) );
  XOR U13748 ( .A(n13945), .B(n13946), .Z(n13920) );
  ANDN U13749 ( .B(n13947), .A(n13948), .Z(n13945) );
  XOR U13750 ( .A(n13946), .B(n13949), .Z(n13947) );
  IV U13751 ( .A(n13928), .Z(n13932) );
  XOR U13752 ( .A(n13928), .B(n13910), .Z(n13930) );
  XOR U13753 ( .A(n13950), .B(n13951), .Z(n13910) );
  AND U13754 ( .A(n778), .B(n13952), .Z(n13950) );
  XOR U13755 ( .A(n13953), .B(n13951), .Z(n13952) );
  NANDN U13756 ( .A(n13912), .B(n13914), .Z(n13928) );
  XOR U13757 ( .A(n13954), .B(n13955), .Z(n13914) );
  AND U13758 ( .A(n778), .B(n13956), .Z(n13954) );
  XOR U13759 ( .A(n13955), .B(n13957), .Z(n13956) );
  XOR U13760 ( .A(n13958), .B(n13959), .Z(n778) );
  AND U13761 ( .A(n13960), .B(n13961), .Z(n13958) );
  XNOR U13762 ( .A(n13959), .B(n13925), .Z(n13961) );
  XNOR U13763 ( .A(n13962), .B(n13963), .Z(n13925) );
  ANDN U13764 ( .B(n13964), .A(n13965), .Z(n13962) );
  XOR U13765 ( .A(n13963), .B(n13966), .Z(n13964) );
  XOR U13766 ( .A(n13959), .B(n13927), .Z(n13960) );
  XOR U13767 ( .A(n13967), .B(n13968), .Z(n13927) );
  AND U13768 ( .A(n782), .B(n13969), .Z(n13967) );
  XOR U13769 ( .A(n13970), .B(n13968), .Z(n13969) );
  XNOR U13770 ( .A(n13971), .B(n13972), .Z(n13959) );
  NAND U13771 ( .A(n13973), .B(n13974), .Z(n13972) );
  XOR U13772 ( .A(n13975), .B(n13951), .Z(n13974) );
  XOR U13773 ( .A(n13965), .B(n13966), .Z(n13951) );
  XOR U13774 ( .A(n13976), .B(n13977), .Z(n13966) );
  ANDN U13775 ( .B(n13978), .A(n13979), .Z(n13976) );
  XOR U13776 ( .A(n13977), .B(n13980), .Z(n13978) );
  XOR U13777 ( .A(n13981), .B(n13982), .Z(n13965) );
  XOR U13778 ( .A(n13983), .B(n13984), .Z(n13982) );
  ANDN U13779 ( .B(n13985), .A(n13986), .Z(n13983) );
  XOR U13780 ( .A(n13987), .B(n13984), .Z(n13985) );
  IV U13781 ( .A(n13963), .Z(n13981) );
  XOR U13782 ( .A(n13988), .B(n13989), .Z(n13963) );
  ANDN U13783 ( .B(n13990), .A(n13991), .Z(n13988) );
  XOR U13784 ( .A(n13989), .B(n13992), .Z(n13990) );
  IV U13785 ( .A(n13971), .Z(n13975) );
  XOR U13786 ( .A(n13971), .B(n13953), .Z(n13973) );
  XOR U13787 ( .A(n13993), .B(n13994), .Z(n13953) );
  AND U13788 ( .A(n782), .B(n13995), .Z(n13993) );
  XOR U13789 ( .A(n13996), .B(n13994), .Z(n13995) );
  NANDN U13790 ( .A(n13955), .B(n13957), .Z(n13971) );
  XOR U13791 ( .A(n13997), .B(n13998), .Z(n13957) );
  AND U13792 ( .A(n782), .B(n13999), .Z(n13997) );
  XOR U13793 ( .A(n13998), .B(n14000), .Z(n13999) );
  XOR U13794 ( .A(n14001), .B(n14002), .Z(n782) );
  AND U13795 ( .A(n14003), .B(n14004), .Z(n14001) );
  XNOR U13796 ( .A(n14002), .B(n13968), .Z(n14004) );
  XNOR U13797 ( .A(n14005), .B(n14006), .Z(n13968) );
  ANDN U13798 ( .B(n14007), .A(n14008), .Z(n14005) );
  XOR U13799 ( .A(n14006), .B(n14009), .Z(n14007) );
  XOR U13800 ( .A(n14002), .B(n13970), .Z(n14003) );
  XOR U13801 ( .A(n14010), .B(n14011), .Z(n13970) );
  AND U13802 ( .A(n786), .B(n14012), .Z(n14010) );
  XOR U13803 ( .A(n14013), .B(n14011), .Z(n14012) );
  XNOR U13804 ( .A(n14014), .B(n14015), .Z(n14002) );
  NAND U13805 ( .A(n14016), .B(n14017), .Z(n14015) );
  XOR U13806 ( .A(n14018), .B(n13994), .Z(n14017) );
  XOR U13807 ( .A(n14008), .B(n14009), .Z(n13994) );
  XOR U13808 ( .A(n14019), .B(n14020), .Z(n14009) );
  ANDN U13809 ( .B(n14021), .A(n14022), .Z(n14019) );
  XOR U13810 ( .A(n14020), .B(n14023), .Z(n14021) );
  XOR U13811 ( .A(n14024), .B(n14025), .Z(n14008) );
  XOR U13812 ( .A(n14026), .B(n14027), .Z(n14025) );
  ANDN U13813 ( .B(n14028), .A(n14029), .Z(n14026) );
  XOR U13814 ( .A(n14030), .B(n14027), .Z(n14028) );
  IV U13815 ( .A(n14006), .Z(n14024) );
  XOR U13816 ( .A(n14031), .B(n14032), .Z(n14006) );
  ANDN U13817 ( .B(n14033), .A(n14034), .Z(n14031) );
  XOR U13818 ( .A(n14032), .B(n14035), .Z(n14033) );
  IV U13819 ( .A(n14014), .Z(n14018) );
  XOR U13820 ( .A(n14014), .B(n13996), .Z(n14016) );
  XOR U13821 ( .A(n14036), .B(n14037), .Z(n13996) );
  AND U13822 ( .A(n786), .B(n14038), .Z(n14036) );
  XOR U13823 ( .A(n14039), .B(n14037), .Z(n14038) );
  NANDN U13824 ( .A(n13998), .B(n14000), .Z(n14014) );
  XOR U13825 ( .A(n14040), .B(n14041), .Z(n14000) );
  AND U13826 ( .A(n786), .B(n14042), .Z(n14040) );
  XOR U13827 ( .A(n14041), .B(n14043), .Z(n14042) );
  XOR U13828 ( .A(n14044), .B(n14045), .Z(n786) );
  AND U13829 ( .A(n14046), .B(n14047), .Z(n14044) );
  XNOR U13830 ( .A(n14045), .B(n14011), .Z(n14047) );
  XNOR U13831 ( .A(n14048), .B(n14049), .Z(n14011) );
  ANDN U13832 ( .B(n14050), .A(n14051), .Z(n14048) );
  XOR U13833 ( .A(n14049), .B(n14052), .Z(n14050) );
  XOR U13834 ( .A(n14045), .B(n14013), .Z(n14046) );
  XOR U13835 ( .A(n14053), .B(n14054), .Z(n14013) );
  AND U13836 ( .A(n790), .B(n14055), .Z(n14053) );
  XOR U13837 ( .A(n14056), .B(n14054), .Z(n14055) );
  XNOR U13838 ( .A(n14057), .B(n14058), .Z(n14045) );
  NAND U13839 ( .A(n14059), .B(n14060), .Z(n14058) );
  XOR U13840 ( .A(n14061), .B(n14037), .Z(n14060) );
  XOR U13841 ( .A(n14051), .B(n14052), .Z(n14037) );
  XOR U13842 ( .A(n14062), .B(n14063), .Z(n14052) );
  ANDN U13843 ( .B(n14064), .A(n14065), .Z(n14062) );
  XOR U13844 ( .A(n14063), .B(n14066), .Z(n14064) );
  XOR U13845 ( .A(n14067), .B(n14068), .Z(n14051) );
  XOR U13846 ( .A(n14069), .B(n14070), .Z(n14068) );
  ANDN U13847 ( .B(n14071), .A(n14072), .Z(n14069) );
  XOR U13848 ( .A(n14073), .B(n14070), .Z(n14071) );
  IV U13849 ( .A(n14049), .Z(n14067) );
  XOR U13850 ( .A(n14074), .B(n14075), .Z(n14049) );
  ANDN U13851 ( .B(n14076), .A(n14077), .Z(n14074) );
  XOR U13852 ( .A(n14075), .B(n14078), .Z(n14076) );
  IV U13853 ( .A(n14057), .Z(n14061) );
  XOR U13854 ( .A(n14057), .B(n14039), .Z(n14059) );
  XOR U13855 ( .A(n14079), .B(n14080), .Z(n14039) );
  AND U13856 ( .A(n790), .B(n14081), .Z(n14079) );
  XOR U13857 ( .A(n14082), .B(n14080), .Z(n14081) );
  NANDN U13858 ( .A(n14041), .B(n14043), .Z(n14057) );
  XOR U13859 ( .A(n14083), .B(n14084), .Z(n14043) );
  AND U13860 ( .A(n790), .B(n14085), .Z(n14083) );
  XOR U13861 ( .A(n14084), .B(n14086), .Z(n14085) );
  XOR U13862 ( .A(n14087), .B(n14088), .Z(n790) );
  AND U13863 ( .A(n14089), .B(n14090), .Z(n14087) );
  XNOR U13864 ( .A(n14088), .B(n14054), .Z(n14090) );
  XNOR U13865 ( .A(n14091), .B(n14092), .Z(n14054) );
  ANDN U13866 ( .B(n14093), .A(n14094), .Z(n14091) );
  XOR U13867 ( .A(n14092), .B(n14095), .Z(n14093) );
  XOR U13868 ( .A(n14088), .B(n14056), .Z(n14089) );
  XOR U13869 ( .A(n14096), .B(n14097), .Z(n14056) );
  AND U13870 ( .A(n794), .B(n14098), .Z(n14096) );
  XOR U13871 ( .A(n14099), .B(n14097), .Z(n14098) );
  XNOR U13872 ( .A(n14100), .B(n14101), .Z(n14088) );
  NAND U13873 ( .A(n14102), .B(n14103), .Z(n14101) );
  XOR U13874 ( .A(n14104), .B(n14080), .Z(n14103) );
  XOR U13875 ( .A(n14094), .B(n14095), .Z(n14080) );
  XOR U13876 ( .A(n14105), .B(n14106), .Z(n14095) );
  ANDN U13877 ( .B(n14107), .A(n14108), .Z(n14105) );
  XOR U13878 ( .A(n14106), .B(n14109), .Z(n14107) );
  XOR U13879 ( .A(n14110), .B(n14111), .Z(n14094) );
  XOR U13880 ( .A(n14112), .B(n14113), .Z(n14111) );
  ANDN U13881 ( .B(n14114), .A(n14115), .Z(n14112) );
  XOR U13882 ( .A(n14116), .B(n14113), .Z(n14114) );
  IV U13883 ( .A(n14092), .Z(n14110) );
  XOR U13884 ( .A(n14117), .B(n14118), .Z(n14092) );
  ANDN U13885 ( .B(n14119), .A(n14120), .Z(n14117) );
  XOR U13886 ( .A(n14118), .B(n14121), .Z(n14119) );
  IV U13887 ( .A(n14100), .Z(n14104) );
  XOR U13888 ( .A(n14100), .B(n14082), .Z(n14102) );
  XOR U13889 ( .A(n14122), .B(n14123), .Z(n14082) );
  AND U13890 ( .A(n794), .B(n14124), .Z(n14122) );
  XOR U13891 ( .A(n14125), .B(n14123), .Z(n14124) );
  NANDN U13892 ( .A(n14084), .B(n14086), .Z(n14100) );
  XOR U13893 ( .A(n14126), .B(n14127), .Z(n14086) );
  AND U13894 ( .A(n794), .B(n14128), .Z(n14126) );
  XOR U13895 ( .A(n14127), .B(n14129), .Z(n14128) );
  XOR U13896 ( .A(n14130), .B(n14131), .Z(n794) );
  AND U13897 ( .A(n14132), .B(n14133), .Z(n14130) );
  XNOR U13898 ( .A(n14131), .B(n14097), .Z(n14133) );
  XNOR U13899 ( .A(n14134), .B(n14135), .Z(n14097) );
  ANDN U13900 ( .B(n14136), .A(n14137), .Z(n14134) );
  XOR U13901 ( .A(n14135), .B(n14138), .Z(n14136) );
  XOR U13902 ( .A(n14131), .B(n14099), .Z(n14132) );
  XOR U13903 ( .A(n14139), .B(n14140), .Z(n14099) );
  AND U13904 ( .A(n798), .B(n14141), .Z(n14139) );
  XOR U13905 ( .A(n14142), .B(n14140), .Z(n14141) );
  XNOR U13906 ( .A(n14143), .B(n14144), .Z(n14131) );
  NAND U13907 ( .A(n14145), .B(n14146), .Z(n14144) );
  XOR U13908 ( .A(n14147), .B(n14123), .Z(n14146) );
  XOR U13909 ( .A(n14137), .B(n14138), .Z(n14123) );
  XOR U13910 ( .A(n14148), .B(n14149), .Z(n14138) );
  ANDN U13911 ( .B(n14150), .A(n14151), .Z(n14148) );
  XOR U13912 ( .A(n14149), .B(n14152), .Z(n14150) );
  XOR U13913 ( .A(n14153), .B(n14154), .Z(n14137) );
  XOR U13914 ( .A(n14155), .B(n14156), .Z(n14154) );
  ANDN U13915 ( .B(n14157), .A(n14158), .Z(n14155) );
  XOR U13916 ( .A(n14159), .B(n14156), .Z(n14157) );
  IV U13917 ( .A(n14135), .Z(n14153) );
  XOR U13918 ( .A(n14160), .B(n14161), .Z(n14135) );
  ANDN U13919 ( .B(n14162), .A(n14163), .Z(n14160) );
  XOR U13920 ( .A(n14161), .B(n14164), .Z(n14162) );
  IV U13921 ( .A(n14143), .Z(n14147) );
  XOR U13922 ( .A(n14143), .B(n14125), .Z(n14145) );
  XOR U13923 ( .A(n14165), .B(n14166), .Z(n14125) );
  AND U13924 ( .A(n798), .B(n14167), .Z(n14165) );
  XOR U13925 ( .A(n14168), .B(n14166), .Z(n14167) );
  NANDN U13926 ( .A(n14127), .B(n14129), .Z(n14143) );
  XOR U13927 ( .A(n14169), .B(n14170), .Z(n14129) );
  AND U13928 ( .A(n798), .B(n14171), .Z(n14169) );
  XOR U13929 ( .A(n14170), .B(n14172), .Z(n14171) );
  XOR U13930 ( .A(n14173), .B(n14174), .Z(n798) );
  AND U13931 ( .A(n14175), .B(n14176), .Z(n14173) );
  XNOR U13932 ( .A(n14174), .B(n14140), .Z(n14176) );
  XNOR U13933 ( .A(n14177), .B(n14178), .Z(n14140) );
  ANDN U13934 ( .B(n14179), .A(n14180), .Z(n14177) );
  XOR U13935 ( .A(n14178), .B(n14181), .Z(n14179) );
  XOR U13936 ( .A(n14174), .B(n14142), .Z(n14175) );
  XOR U13937 ( .A(n14182), .B(n14183), .Z(n14142) );
  AND U13938 ( .A(n802), .B(n14184), .Z(n14182) );
  XOR U13939 ( .A(n14185), .B(n14183), .Z(n14184) );
  XNOR U13940 ( .A(n14186), .B(n14187), .Z(n14174) );
  NAND U13941 ( .A(n14188), .B(n14189), .Z(n14187) );
  XOR U13942 ( .A(n14190), .B(n14166), .Z(n14189) );
  XOR U13943 ( .A(n14180), .B(n14181), .Z(n14166) );
  XOR U13944 ( .A(n14191), .B(n14192), .Z(n14181) );
  ANDN U13945 ( .B(n14193), .A(n14194), .Z(n14191) );
  XOR U13946 ( .A(n14192), .B(n14195), .Z(n14193) );
  XOR U13947 ( .A(n14196), .B(n14197), .Z(n14180) );
  XOR U13948 ( .A(n14198), .B(n14199), .Z(n14197) );
  ANDN U13949 ( .B(n14200), .A(n14201), .Z(n14198) );
  XOR U13950 ( .A(n14202), .B(n14199), .Z(n14200) );
  IV U13951 ( .A(n14178), .Z(n14196) );
  XOR U13952 ( .A(n14203), .B(n14204), .Z(n14178) );
  ANDN U13953 ( .B(n14205), .A(n14206), .Z(n14203) );
  XOR U13954 ( .A(n14204), .B(n14207), .Z(n14205) );
  IV U13955 ( .A(n14186), .Z(n14190) );
  XOR U13956 ( .A(n14186), .B(n14168), .Z(n14188) );
  XOR U13957 ( .A(n14208), .B(n14209), .Z(n14168) );
  AND U13958 ( .A(n802), .B(n14210), .Z(n14208) );
  XOR U13959 ( .A(n14211), .B(n14209), .Z(n14210) );
  NANDN U13960 ( .A(n14170), .B(n14172), .Z(n14186) );
  XOR U13961 ( .A(n14212), .B(n14213), .Z(n14172) );
  AND U13962 ( .A(n802), .B(n14214), .Z(n14212) );
  XOR U13963 ( .A(n14213), .B(n14215), .Z(n14214) );
  XOR U13964 ( .A(n14216), .B(n14217), .Z(n802) );
  AND U13965 ( .A(n14218), .B(n14219), .Z(n14216) );
  XNOR U13966 ( .A(n14217), .B(n14183), .Z(n14219) );
  XNOR U13967 ( .A(n14220), .B(n14221), .Z(n14183) );
  ANDN U13968 ( .B(n14222), .A(n14223), .Z(n14220) );
  XOR U13969 ( .A(n14221), .B(n14224), .Z(n14222) );
  XOR U13970 ( .A(n14217), .B(n14185), .Z(n14218) );
  XOR U13971 ( .A(n14225), .B(n14226), .Z(n14185) );
  AND U13972 ( .A(n806), .B(n14227), .Z(n14225) );
  XOR U13973 ( .A(n14228), .B(n14226), .Z(n14227) );
  XNOR U13974 ( .A(n14229), .B(n14230), .Z(n14217) );
  NAND U13975 ( .A(n14231), .B(n14232), .Z(n14230) );
  XOR U13976 ( .A(n14233), .B(n14209), .Z(n14232) );
  XOR U13977 ( .A(n14223), .B(n14224), .Z(n14209) );
  XOR U13978 ( .A(n14234), .B(n14235), .Z(n14224) );
  ANDN U13979 ( .B(n14236), .A(n14237), .Z(n14234) );
  XOR U13980 ( .A(n14235), .B(n14238), .Z(n14236) );
  XOR U13981 ( .A(n14239), .B(n14240), .Z(n14223) );
  XOR U13982 ( .A(n14241), .B(n14242), .Z(n14240) );
  ANDN U13983 ( .B(n14243), .A(n14244), .Z(n14241) );
  XOR U13984 ( .A(n14245), .B(n14242), .Z(n14243) );
  IV U13985 ( .A(n14221), .Z(n14239) );
  XOR U13986 ( .A(n14246), .B(n14247), .Z(n14221) );
  ANDN U13987 ( .B(n14248), .A(n14249), .Z(n14246) );
  XOR U13988 ( .A(n14247), .B(n14250), .Z(n14248) );
  IV U13989 ( .A(n14229), .Z(n14233) );
  XOR U13990 ( .A(n14229), .B(n14211), .Z(n14231) );
  XOR U13991 ( .A(n14251), .B(n14252), .Z(n14211) );
  AND U13992 ( .A(n806), .B(n14253), .Z(n14251) );
  XOR U13993 ( .A(n14254), .B(n14252), .Z(n14253) );
  NANDN U13994 ( .A(n14213), .B(n14215), .Z(n14229) );
  XOR U13995 ( .A(n14255), .B(n14256), .Z(n14215) );
  AND U13996 ( .A(n806), .B(n14257), .Z(n14255) );
  XOR U13997 ( .A(n14256), .B(n14258), .Z(n14257) );
  XOR U13998 ( .A(n14259), .B(n14260), .Z(n806) );
  AND U13999 ( .A(n14261), .B(n14262), .Z(n14259) );
  XNOR U14000 ( .A(n14260), .B(n14226), .Z(n14262) );
  XNOR U14001 ( .A(n14263), .B(n14264), .Z(n14226) );
  ANDN U14002 ( .B(n14265), .A(n14266), .Z(n14263) );
  XOR U14003 ( .A(n14264), .B(n14267), .Z(n14265) );
  XOR U14004 ( .A(n14260), .B(n14228), .Z(n14261) );
  XOR U14005 ( .A(n14268), .B(n14269), .Z(n14228) );
  AND U14006 ( .A(n810), .B(n14270), .Z(n14268) );
  XOR U14007 ( .A(n14271), .B(n14269), .Z(n14270) );
  XNOR U14008 ( .A(n14272), .B(n14273), .Z(n14260) );
  NAND U14009 ( .A(n14274), .B(n14275), .Z(n14273) );
  XOR U14010 ( .A(n14276), .B(n14252), .Z(n14275) );
  XOR U14011 ( .A(n14266), .B(n14267), .Z(n14252) );
  XOR U14012 ( .A(n14277), .B(n14278), .Z(n14267) );
  ANDN U14013 ( .B(n14279), .A(n14280), .Z(n14277) );
  XOR U14014 ( .A(n14278), .B(n14281), .Z(n14279) );
  XOR U14015 ( .A(n14282), .B(n14283), .Z(n14266) );
  XOR U14016 ( .A(n14284), .B(n14285), .Z(n14283) );
  ANDN U14017 ( .B(n14286), .A(n14287), .Z(n14284) );
  XOR U14018 ( .A(n14288), .B(n14285), .Z(n14286) );
  IV U14019 ( .A(n14264), .Z(n14282) );
  XOR U14020 ( .A(n14289), .B(n14290), .Z(n14264) );
  ANDN U14021 ( .B(n14291), .A(n14292), .Z(n14289) );
  XOR U14022 ( .A(n14290), .B(n14293), .Z(n14291) );
  IV U14023 ( .A(n14272), .Z(n14276) );
  XOR U14024 ( .A(n14272), .B(n14254), .Z(n14274) );
  XOR U14025 ( .A(n14294), .B(n14295), .Z(n14254) );
  AND U14026 ( .A(n810), .B(n14296), .Z(n14294) );
  XOR U14027 ( .A(n14297), .B(n14295), .Z(n14296) );
  NANDN U14028 ( .A(n14256), .B(n14258), .Z(n14272) );
  XOR U14029 ( .A(n14298), .B(n14299), .Z(n14258) );
  AND U14030 ( .A(n810), .B(n14300), .Z(n14298) );
  XOR U14031 ( .A(n14299), .B(n14301), .Z(n14300) );
  XOR U14032 ( .A(n14302), .B(n14303), .Z(n810) );
  AND U14033 ( .A(n14304), .B(n14305), .Z(n14302) );
  XNOR U14034 ( .A(n14303), .B(n14269), .Z(n14305) );
  XNOR U14035 ( .A(n14306), .B(n14307), .Z(n14269) );
  ANDN U14036 ( .B(n14308), .A(n14309), .Z(n14306) );
  XOR U14037 ( .A(n14307), .B(n14310), .Z(n14308) );
  XOR U14038 ( .A(n14303), .B(n14271), .Z(n14304) );
  XOR U14039 ( .A(n14311), .B(n14312), .Z(n14271) );
  AND U14040 ( .A(n814), .B(n14313), .Z(n14311) );
  XOR U14041 ( .A(n14314), .B(n14312), .Z(n14313) );
  XNOR U14042 ( .A(n14315), .B(n14316), .Z(n14303) );
  NAND U14043 ( .A(n14317), .B(n14318), .Z(n14316) );
  XOR U14044 ( .A(n14319), .B(n14295), .Z(n14318) );
  XOR U14045 ( .A(n14309), .B(n14310), .Z(n14295) );
  XOR U14046 ( .A(n14320), .B(n14321), .Z(n14310) );
  ANDN U14047 ( .B(n14322), .A(n14323), .Z(n14320) );
  XOR U14048 ( .A(n14321), .B(n14324), .Z(n14322) );
  XOR U14049 ( .A(n14325), .B(n14326), .Z(n14309) );
  XOR U14050 ( .A(n14327), .B(n14328), .Z(n14326) );
  ANDN U14051 ( .B(n14329), .A(n14330), .Z(n14327) );
  XOR U14052 ( .A(n14331), .B(n14328), .Z(n14329) );
  IV U14053 ( .A(n14307), .Z(n14325) );
  XOR U14054 ( .A(n14332), .B(n14333), .Z(n14307) );
  ANDN U14055 ( .B(n14334), .A(n14335), .Z(n14332) );
  XOR U14056 ( .A(n14333), .B(n14336), .Z(n14334) );
  IV U14057 ( .A(n14315), .Z(n14319) );
  XOR U14058 ( .A(n14315), .B(n14297), .Z(n14317) );
  XOR U14059 ( .A(n14337), .B(n14338), .Z(n14297) );
  AND U14060 ( .A(n814), .B(n14339), .Z(n14337) );
  XOR U14061 ( .A(n14340), .B(n14338), .Z(n14339) );
  NANDN U14062 ( .A(n14299), .B(n14301), .Z(n14315) );
  XOR U14063 ( .A(n14341), .B(n14342), .Z(n14301) );
  AND U14064 ( .A(n814), .B(n14343), .Z(n14341) );
  XOR U14065 ( .A(n14342), .B(n14344), .Z(n14343) );
  XOR U14066 ( .A(n14345), .B(n14346), .Z(n814) );
  AND U14067 ( .A(n14347), .B(n14348), .Z(n14345) );
  XNOR U14068 ( .A(n14346), .B(n14312), .Z(n14348) );
  XNOR U14069 ( .A(n14349), .B(n14350), .Z(n14312) );
  ANDN U14070 ( .B(n14351), .A(n14352), .Z(n14349) );
  XOR U14071 ( .A(n14350), .B(n14353), .Z(n14351) );
  XOR U14072 ( .A(n14346), .B(n14314), .Z(n14347) );
  XOR U14073 ( .A(n14354), .B(n14355), .Z(n14314) );
  AND U14074 ( .A(n818), .B(n14356), .Z(n14354) );
  XOR U14075 ( .A(n14357), .B(n14355), .Z(n14356) );
  XNOR U14076 ( .A(n14358), .B(n14359), .Z(n14346) );
  NAND U14077 ( .A(n14360), .B(n14361), .Z(n14359) );
  XOR U14078 ( .A(n14362), .B(n14338), .Z(n14361) );
  XOR U14079 ( .A(n14352), .B(n14353), .Z(n14338) );
  XOR U14080 ( .A(n14363), .B(n14364), .Z(n14353) );
  ANDN U14081 ( .B(n14365), .A(n14366), .Z(n14363) );
  XOR U14082 ( .A(n14364), .B(n14367), .Z(n14365) );
  XOR U14083 ( .A(n14368), .B(n14369), .Z(n14352) );
  XOR U14084 ( .A(n14370), .B(n14371), .Z(n14369) );
  ANDN U14085 ( .B(n14372), .A(n14373), .Z(n14370) );
  XOR U14086 ( .A(n14374), .B(n14371), .Z(n14372) );
  IV U14087 ( .A(n14350), .Z(n14368) );
  XOR U14088 ( .A(n14375), .B(n14376), .Z(n14350) );
  ANDN U14089 ( .B(n14377), .A(n14378), .Z(n14375) );
  XOR U14090 ( .A(n14376), .B(n14379), .Z(n14377) );
  IV U14091 ( .A(n14358), .Z(n14362) );
  XOR U14092 ( .A(n14358), .B(n14340), .Z(n14360) );
  XOR U14093 ( .A(n14380), .B(n14381), .Z(n14340) );
  AND U14094 ( .A(n818), .B(n14382), .Z(n14380) );
  XOR U14095 ( .A(n14383), .B(n14381), .Z(n14382) );
  NANDN U14096 ( .A(n14342), .B(n14344), .Z(n14358) );
  XOR U14097 ( .A(n14384), .B(n14385), .Z(n14344) );
  AND U14098 ( .A(n818), .B(n14386), .Z(n14384) );
  XOR U14099 ( .A(n14385), .B(n14387), .Z(n14386) );
  XOR U14100 ( .A(n14388), .B(n14389), .Z(n818) );
  AND U14101 ( .A(n14390), .B(n14391), .Z(n14388) );
  XNOR U14102 ( .A(n14389), .B(n14355), .Z(n14391) );
  XNOR U14103 ( .A(n14392), .B(n14393), .Z(n14355) );
  ANDN U14104 ( .B(n14394), .A(n14395), .Z(n14392) );
  XOR U14105 ( .A(n14393), .B(n14396), .Z(n14394) );
  XOR U14106 ( .A(n14389), .B(n14357), .Z(n14390) );
  XOR U14107 ( .A(n14397), .B(n14398), .Z(n14357) );
  AND U14108 ( .A(n822), .B(n14399), .Z(n14397) );
  XOR U14109 ( .A(n14400), .B(n14398), .Z(n14399) );
  XNOR U14110 ( .A(n14401), .B(n14402), .Z(n14389) );
  NAND U14111 ( .A(n14403), .B(n14404), .Z(n14402) );
  XOR U14112 ( .A(n14405), .B(n14381), .Z(n14404) );
  XOR U14113 ( .A(n14395), .B(n14396), .Z(n14381) );
  XOR U14114 ( .A(n14406), .B(n14407), .Z(n14396) );
  ANDN U14115 ( .B(n14408), .A(n14409), .Z(n14406) );
  XOR U14116 ( .A(n14407), .B(n14410), .Z(n14408) );
  XOR U14117 ( .A(n14411), .B(n14412), .Z(n14395) );
  XOR U14118 ( .A(n14413), .B(n14414), .Z(n14412) );
  ANDN U14119 ( .B(n14415), .A(n14416), .Z(n14413) );
  XOR U14120 ( .A(n14417), .B(n14414), .Z(n14415) );
  IV U14121 ( .A(n14393), .Z(n14411) );
  XOR U14122 ( .A(n14418), .B(n14419), .Z(n14393) );
  ANDN U14123 ( .B(n14420), .A(n14421), .Z(n14418) );
  XOR U14124 ( .A(n14419), .B(n14422), .Z(n14420) );
  IV U14125 ( .A(n14401), .Z(n14405) );
  XOR U14126 ( .A(n14401), .B(n14383), .Z(n14403) );
  XOR U14127 ( .A(n14423), .B(n14424), .Z(n14383) );
  AND U14128 ( .A(n822), .B(n14425), .Z(n14423) );
  XOR U14129 ( .A(n14426), .B(n14424), .Z(n14425) );
  NANDN U14130 ( .A(n14385), .B(n14387), .Z(n14401) );
  XOR U14131 ( .A(n14427), .B(n14428), .Z(n14387) );
  AND U14132 ( .A(n822), .B(n14429), .Z(n14427) );
  XOR U14133 ( .A(n14428), .B(n14430), .Z(n14429) );
  XOR U14134 ( .A(n14431), .B(n14432), .Z(n822) );
  AND U14135 ( .A(n14433), .B(n14434), .Z(n14431) );
  XNOR U14136 ( .A(n14432), .B(n14398), .Z(n14434) );
  XNOR U14137 ( .A(n14435), .B(n14436), .Z(n14398) );
  ANDN U14138 ( .B(n14437), .A(n14438), .Z(n14435) );
  XOR U14139 ( .A(n14436), .B(n14439), .Z(n14437) );
  XOR U14140 ( .A(n14432), .B(n14400), .Z(n14433) );
  XOR U14141 ( .A(n14440), .B(n14441), .Z(n14400) );
  AND U14142 ( .A(n826), .B(n14442), .Z(n14440) );
  XOR U14143 ( .A(n14443), .B(n14441), .Z(n14442) );
  XNOR U14144 ( .A(n14444), .B(n14445), .Z(n14432) );
  NAND U14145 ( .A(n14446), .B(n14447), .Z(n14445) );
  XOR U14146 ( .A(n14448), .B(n14424), .Z(n14447) );
  XOR U14147 ( .A(n14438), .B(n14439), .Z(n14424) );
  XOR U14148 ( .A(n14449), .B(n14450), .Z(n14439) );
  ANDN U14149 ( .B(n14451), .A(n14452), .Z(n14449) );
  XOR U14150 ( .A(n14450), .B(n14453), .Z(n14451) );
  XOR U14151 ( .A(n14454), .B(n14455), .Z(n14438) );
  XOR U14152 ( .A(n14456), .B(n14457), .Z(n14455) );
  ANDN U14153 ( .B(n14458), .A(n14459), .Z(n14456) );
  XOR U14154 ( .A(n14460), .B(n14457), .Z(n14458) );
  IV U14155 ( .A(n14436), .Z(n14454) );
  XOR U14156 ( .A(n14461), .B(n14462), .Z(n14436) );
  ANDN U14157 ( .B(n14463), .A(n14464), .Z(n14461) );
  XOR U14158 ( .A(n14462), .B(n14465), .Z(n14463) );
  IV U14159 ( .A(n14444), .Z(n14448) );
  XOR U14160 ( .A(n14444), .B(n14426), .Z(n14446) );
  XOR U14161 ( .A(n14466), .B(n14467), .Z(n14426) );
  AND U14162 ( .A(n826), .B(n14468), .Z(n14466) );
  XOR U14163 ( .A(n14469), .B(n14467), .Z(n14468) );
  NANDN U14164 ( .A(n14428), .B(n14430), .Z(n14444) );
  XOR U14165 ( .A(n14470), .B(n14471), .Z(n14430) );
  AND U14166 ( .A(n826), .B(n14472), .Z(n14470) );
  XOR U14167 ( .A(n14471), .B(n14473), .Z(n14472) );
  XOR U14168 ( .A(n14474), .B(n14475), .Z(n826) );
  AND U14169 ( .A(n14476), .B(n14477), .Z(n14474) );
  XNOR U14170 ( .A(n14475), .B(n14441), .Z(n14477) );
  XNOR U14171 ( .A(n14478), .B(n14479), .Z(n14441) );
  ANDN U14172 ( .B(n14480), .A(n14481), .Z(n14478) );
  XOR U14173 ( .A(n14479), .B(n14482), .Z(n14480) );
  XOR U14174 ( .A(n14475), .B(n14443), .Z(n14476) );
  XOR U14175 ( .A(n14483), .B(n14484), .Z(n14443) );
  AND U14176 ( .A(n830), .B(n14485), .Z(n14483) );
  XOR U14177 ( .A(n14486), .B(n14484), .Z(n14485) );
  XNOR U14178 ( .A(n14487), .B(n14488), .Z(n14475) );
  NAND U14179 ( .A(n14489), .B(n14490), .Z(n14488) );
  XOR U14180 ( .A(n14491), .B(n14467), .Z(n14490) );
  XOR U14181 ( .A(n14481), .B(n14482), .Z(n14467) );
  XOR U14182 ( .A(n14492), .B(n14493), .Z(n14482) );
  ANDN U14183 ( .B(n14494), .A(n14495), .Z(n14492) );
  XOR U14184 ( .A(n14493), .B(n14496), .Z(n14494) );
  XOR U14185 ( .A(n14497), .B(n14498), .Z(n14481) );
  XOR U14186 ( .A(n14499), .B(n14500), .Z(n14498) );
  ANDN U14187 ( .B(n14501), .A(n14502), .Z(n14499) );
  XOR U14188 ( .A(n14503), .B(n14500), .Z(n14501) );
  IV U14189 ( .A(n14479), .Z(n14497) );
  XOR U14190 ( .A(n14504), .B(n14505), .Z(n14479) );
  ANDN U14191 ( .B(n14506), .A(n14507), .Z(n14504) );
  XOR U14192 ( .A(n14505), .B(n14508), .Z(n14506) );
  IV U14193 ( .A(n14487), .Z(n14491) );
  XOR U14194 ( .A(n14487), .B(n14469), .Z(n14489) );
  XOR U14195 ( .A(n14509), .B(n14510), .Z(n14469) );
  AND U14196 ( .A(n830), .B(n14511), .Z(n14509) );
  XOR U14197 ( .A(n14512), .B(n14510), .Z(n14511) );
  NANDN U14198 ( .A(n14471), .B(n14473), .Z(n14487) );
  XOR U14199 ( .A(n14513), .B(n14514), .Z(n14473) );
  AND U14200 ( .A(n830), .B(n14515), .Z(n14513) );
  XOR U14201 ( .A(n14514), .B(n14516), .Z(n14515) );
  XOR U14202 ( .A(n14517), .B(n14518), .Z(n830) );
  AND U14203 ( .A(n14519), .B(n14520), .Z(n14517) );
  XNOR U14204 ( .A(n14518), .B(n14484), .Z(n14520) );
  XNOR U14205 ( .A(n14521), .B(n14522), .Z(n14484) );
  ANDN U14206 ( .B(n14523), .A(n14524), .Z(n14521) );
  XOR U14207 ( .A(n14522), .B(n14525), .Z(n14523) );
  XOR U14208 ( .A(n14518), .B(n14486), .Z(n14519) );
  XOR U14209 ( .A(n14526), .B(n14527), .Z(n14486) );
  AND U14210 ( .A(n834), .B(n14528), .Z(n14526) );
  XOR U14211 ( .A(n14529), .B(n14527), .Z(n14528) );
  XNOR U14212 ( .A(n14530), .B(n14531), .Z(n14518) );
  NAND U14213 ( .A(n14532), .B(n14533), .Z(n14531) );
  XOR U14214 ( .A(n14534), .B(n14510), .Z(n14533) );
  XOR U14215 ( .A(n14524), .B(n14525), .Z(n14510) );
  XOR U14216 ( .A(n14535), .B(n14536), .Z(n14525) );
  ANDN U14217 ( .B(n14537), .A(n14538), .Z(n14535) );
  XOR U14218 ( .A(n14536), .B(n14539), .Z(n14537) );
  XOR U14219 ( .A(n14540), .B(n14541), .Z(n14524) );
  XOR U14220 ( .A(n14542), .B(n14543), .Z(n14541) );
  ANDN U14221 ( .B(n14544), .A(n14545), .Z(n14542) );
  XOR U14222 ( .A(n14546), .B(n14543), .Z(n14544) );
  IV U14223 ( .A(n14522), .Z(n14540) );
  XOR U14224 ( .A(n14547), .B(n14548), .Z(n14522) );
  ANDN U14225 ( .B(n14549), .A(n14550), .Z(n14547) );
  XOR U14226 ( .A(n14548), .B(n14551), .Z(n14549) );
  IV U14227 ( .A(n14530), .Z(n14534) );
  XOR U14228 ( .A(n14530), .B(n14512), .Z(n14532) );
  XOR U14229 ( .A(n14552), .B(n14553), .Z(n14512) );
  AND U14230 ( .A(n834), .B(n14554), .Z(n14552) );
  XOR U14231 ( .A(n14555), .B(n14553), .Z(n14554) );
  NANDN U14232 ( .A(n14514), .B(n14516), .Z(n14530) );
  XOR U14233 ( .A(n14556), .B(n14557), .Z(n14516) );
  AND U14234 ( .A(n834), .B(n14558), .Z(n14556) );
  XOR U14235 ( .A(n14557), .B(n14559), .Z(n14558) );
  XOR U14236 ( .A(n14560), .B(n14561), .Z(n834) );
  AND U14237 ( .A(n14562), .B(n14563), .Z(n14560) );
  XNOR U14238 ( .A(n14561), .B(n14527), .Z(n14563) );
  XNOR U14239 ( .A(n14564), .B(n14565), .Z(n14527) );
  ANDN U14240 ( .B(n14566), .A(n14567), .Z(n14564) );
  XOR U14241 ( .A(n14565), .B(n14568), .Z(n14566) );
  XOR U14242 ( .A(n14561), .B(n14529), .Z(n14562) );
  XOR U14243 ( .A(n14569), .B(n14570), .Z(n14529) );
  AND U14244 ( .A(n838), .B(n14571), .Z(n14569) );
  XOR U14245 ( .A(n14572), .B(n14570), .Z(n14571) );
  XNOR U14246 ( .A(n14573), .B(n14574), .Z(n14561) );
  NAND U14247 ( .A(n14575), .B(n14576), .Z(n14574) );
  XOR U14248 ( .A(n14577), .B(n14553), .Z(n14576) );
  XOR U14249 ( .A(n14567), .B(n14568), .Z(n14553) );
  XOR U14250 ( .A(n14578), .B(n14579), .Z(n14568) );
  ANDN U14251 ( .B(n14580), .A(n14581), .Z(n14578) );
  XOR U14252 ( .A(n14579), .B(n14582), .Z(n14580) );
  XOR U14253 ( .A(n14583), .B(n14584), .Z(n14567) );
  XOR U14254 ( .A(n14585), .B(n14586), .Z(n14584) );
  ANDN U14255 ( .B(n14587), .A(n14588), .Z(n14585) );
  XOR U14256 ( .A(n14589), .B(n14586), .Z(n14587) );
  IV U14257 ( .A(n14565), .Z(n14583) );
  XOR U14258 ( .A(n14590), .B(n14591), .Z(n14565) );
  ANDN U14259 ( .B(n14592), .A(n14593), .Z(n14590) );
  XOR U14260 ( .A(n14591), .B(n14594), .Z(n14592) );
  IV U14261 ( .A(n14573), .Z(n14577) );
  XOR U14262 ( .A(n14573), .B(n14555), .Z(n14575) );
  XOR U14263 ( .A(n14595), .B(n14596), .Z(n14555) );
  AND U14264 ( .A(n838), .B(n14597), .Z(n14595) );
  XOR U14265 ( .A(n14598), .B(n14596), .Z(n14597) );
  NANDN U14266 ( .A(n14557), .B(n14559), .Z(n14573) );
  XOR U14267 ( .A(n14599), .B(n14600), .Z(n14559) );
  AND U14268 ( .A(n838), .B(n14601), .Z(n14599) );
  XOR U14269 ( .A(n14600), .B(n14602), .Z(n14601) );
  XOR U14270 ( .A(n14603), .B(n14604), .Z(n838) );
  AND U14271 ( .A(n14605), .B(n14606), .Z(n14603) );
  XNOR U14272 ( .A(n14604), .B(n14570), .Z(n14606) );
  XNOR U14273 ( .A(n14607), .B(n14608), .Z(n14570) );
  ANDN U14274 ( .B(n14609), .A(n14610), .Z(n14607) );
  XOR U14275 ( .A(n14608), .B(n14611), .Z(n14609) );
  XOR U14276 ( .A(n14604), .B(n14572), .Z(n14605) );
  XOR U14277 ( .A(n14612), .B(n14613), .Z(n14572) );
  AND U14278 ( .A(n842), .B(n14614), .Z(n14612) );
  XOR U14279 ( .A(n14615), .B(n14613), .Z(n14614) );
  XNOR U14280 ( .A(n14616), .B(n14617), .Z(n14604) );
  NAND U14281 ( .A(n14618), .B(n14619), .Z(n14617) );
  XOR U14282 ( .A(n14620), .B(n14596), .Z(n14619) );
  XOR U14283 ( .A(n14610), .B(n14611), .Z(n14596) );
  XOR U14284 ( .A(n14621), .B(n14622), .Z(n14611) );
  ANDN U14285 ( .B(n14623), .A(n14624), .Z(n14621) );
  XOR U14286 ( .A(n14622), .B(n14625), .Z(n14623) );
  XOR U14287 ( .A(n14626), .B(n14627), .Z(n14610) );
  XOR U14288 ( .A(n14628), .B(n14629), .Z(n14627) );
  ANDN U14289 ( .B(n14630), .A(n14631), .Z(n14628) );
  XOR U14290 ( .A(n14632), .B(n14629), .Z(n14630) );
  IV U14291 ( .A(n14608), .Z(n14626) );
  XOR U14292 ( .A(n14633), .B(n14634), .Z(n14608) );
  ANDN U14293 ( .B(n14635), .A(n14636), .Z(n14633) );
  XOR U14294 ( .A(n14634), .B(n14637), .Z(n14635) );
  IV U14295 ( .A(n14616), .Z(n14620) );
  XOR U14296 ( .A(n14616), .B(n14598), .Z(n14618) );
  XOR U14297 ( .A(n14638), .B(n14639), .Z(n14598) );
  AND U14298 ( .A(n842), .B(n14640), .Z(n14638) );
  XOR U14299 ( .A(n14641), .B(n14639), .Z(n14640) );
  NANDN U14300 ( .A(n14600), .B(n14602), .Z(n14616) );
  XOR U14301 ( .A(n14642), .B(n14643), .Z(n14602) );
  AND U14302 ( .A(n842), .B(n14644), .Z(n14642) );
  XOR U14303 ( .A(n14643), .B(n14645), .Z(n14644) );
  XOR U14304 ( .A(n14646), .B(n14647), .Z(n842) );
  AND U14305 ( .A(n14648), .B(n14649), .Z(n14646) );
  XNOR U14306 ( .A(n14647), .B(n14613), .Z(n14649) );
  XNOR U14307 ( .A(n14650), .B(n14651), .Z(n14613) );
  ANDN U14308 ( .B(n14652), .A(n14653), .Z(n14650) );
  XOR U14309 ( .A(n14651), .B(n14654), .Z(n14652) );
  XOR U14310 ( .A(n14647), .B(n14615), .Z(n14648) );
  XOR U14311 ( .A(n14655), .B(n14656), .Z(n14615) );
  AND U14312 ( .A(n846), .B(n14657), .Z(n14655) );
  XOR U14313 ( .A(n14658), .B(n14656), .Z(n14657) );
  XNOR U14314 ( .A(n14659), .B(n14660), .Z(n14647) );
  NAND U14315 ( .A(n14661), .B(n14662), .Z(n14660) );
  XOR U14316 ( .A(n14663), .B(n14639), .Z(n14662) );
  XOR U14317 ( .A(n14653), .B(n14654), .Z(n14639) );
  XOR U14318 ( .A(n14664), .B(n14665), .Z(n14654) );
  ANDN U14319 ( .B(n14666), .A(n14667), .Z(n14664) );
  XOR U14320 ( .A(n14665), .B(n14668), .Z(n14666) );
  XOR U14321 ( .A(n14669), .B(n14670), .Z(n14653) );
  XOR U14322 ( .A(n14671), .B(n14672), .Z(n14670) );
  ANDN U14323 ( .B(n14673), .A(n14674), .Z(n14671) );
  XOR U14324 ( .A(n14675), .B(n14672), .Z(n14673) );
  IV U14325 ( .A(n14651), .Z(n14669) );
  XOR U14326 ( .A(n14676), .B(n14677), .Z(n14651) );
  ANDN U14327 ( .B(n14678), .A(n14679), .Z(n14676) );
  XOR U14328 ( .A(n14677), .B(n14680), .Z(n14678) );
  IV U14329 ( .A(n14659), .Z(n14663) );
  XOR U14330 ( .A(n14659), .B(n14641), .Z(n14661) );
  XOR U14331 ( .A(n14681), .B(n14682), .Z(n14641) );
  AND U14332 ( .A(n846), .B(n14683), .Z(n14681) );
  XOR U14333 ( .A(n14684), .B(n14682), .Z(n14683) );
  NANDN U14334 ( .A(n14643), .B(n14645), .Z(n14659) );
  XOR U14335 ( .A(n14685), .B(n14686), .Z(n14645) );
  AND U14336 ( .A(n846), .B(n14687), .Z(n14685) );
  XOR U14337 ( .A(n14686), .B(n14688), .Z(n14687) );
  XOR U14338 ( .A(n14689), .B(n14690), .Z(n846) );
  AND U14339 ( .A(n14691), .B(n14692), .Z(n14689) );
  XNOR U14340 ( .A(n14690), .B(n14656), .Z(n14692) );
  XNOR U14341 ( .A(n14693), .B(n14694), .Z(n14656) );
  ANDN U14342 ( .B(n14695), .A(n14696), .Z(n14693) );
  XOR U14343 ( .A(n14694), .B(n14697), .Z(n14695) );
  XOR U14344 ( .A(n14690), .B(n14658), .Z(n14691) );
  XOR U14345 ( .A(n14698), .B(n14699), .Z(n14658) );
  AND U14346 ( .A(n850), .B(n14700), .Z(n14698) );
  XOR U14347 ( .A(n14701), .B(n14699), .Z(n14700) );
  XNOR U14348 ( .A(n14702), .B(n14703), .Z(n14690) );
  NAND U14349 ( .A(n14704), .B(n14705), .Z(n14703) );
  XOR U14350 ( .A(n14706), .B(n14682), .Z(n14705) );
  XOR U14351 ( .A(n14696), .B(n14697), .Z(n14682) );
  XOR U14352 ( .A(n14707), .B(n14708), .Z(n14697) );
  ANDN U14353 ( .B(n14709), .A(n14710), .Z(n14707) );
  XOR U14354 ( .A(n14708), .B(n14711), .Z(n14709) );
  XOR U14355 ( .A(n14712), .B(n14713), .Z(n14696) );
  XOR U14356 ( .A(n14714), .B(n14715), .Z(n14713) );
  ANDN U14357 ( .B(n14716), .A(n14717), .Z(n14714) );
  XOR U14358 ( .A(n14718), .B(n14715), .Z(n14716) );
  IV U14359 ( .A(n14694), .Z(n14712) );
  XOR U14360 ( .A(n14719), .B(n14720), .Z(n14694) );
  ANDN U14361 ( .B(n14721), .A(n14722), .Z(n14719) );
  XOR U14362 ( .A(n14720), .B(n14723), .Z(n14721) );
  IV U14363 ( .A(n14702), .Z(n14706) );
  XOR U14364 ( .A(n14702), .B(n14684), .Z(n14704) );
  XOR U14365 ( .A(n14724), .B(n14725), .Z(n14684) );
  AND U14366 ( .A(n850), .B(n14726), .Z(n14724) );
  XOR U14367 ( .A(n14727), .B(n14725), .Z(n14726) );
  NANDN U14368 ( .A(n14686), .B(n14688), .Z(n14702) );
  XOR U14369 ( .A(n14728), .B(n14729), .Z(n14688) );
  AND U14370 ( .A(n850), .B(n14730), .Z(n14728) );
  XOR U14371 ( .A(n14729), .B(n14731), .Z(n14730) );
  XOR U14372 ( .A(n14732), .B(n14733), .Z(n850) );
  AND U14373 ( .A(n14734), .B(n14735), .Z(n14732) );
  XNOR U14374 ( .A(n14733), .B(n14699), .Z(n14735) );
  XNOR U14375 ( .A(n14736), .B(n14737), .Z(n14699) );
  ANDN U14376 ( .B(n14738), .A(n14739), .Z(n14736) );
  XOR U14377 ( .A(n14737), .B(n14740), .Z(n14738) );
  XOR U14378 ( .A(n14733), .B(n14701), .Z(n14734) );
  XOR U14379 ( .A(n14741), .B(n14742), .Z(n14701) );
  AND U14380 ( .A(n854), .B(n14743), .Z(n14741) );
  XOR U14381 ( .A(n14744), .B(n14742), .Z(n14743) );
  XNOR U14382 ( .A(n14745), .B(n14746), .Z(n14733) );
  NAND U14383 ( .A(n14747), .B(n14748), .Z(n14746) );
  XOR U14384 ( .A(n14749), .B(n14725), .Z(n14748) );
  XOR U14385 ( .A(n14739), .B(n14740), .Z(n14725) );
  XOR U14386 ( .A(n14750), .B(n14751), .Z(n14740) );
  ANDN U14387 ( .B(n14752), .A(n14753), .Z(n14750) );
  XOR U14388 ( .A(n14751), .B(n14754), .Z(n14752) );
  XOR U14389 ( .A(n14755), .B(n14756), .Z(n14739) );
  XOR U14390 ( .A(n14757), .B(n14758), .Z(n14756) );
  ANDN U14391 ( .B(n14759), .A(n14760), .Z(n14757) );
  XOR U14392 ( .A(n14761), .B(n14758), .Z(n14759) );
  IV U14393 ( .A(n14737), .Z(n14755) );
  XOR U14394 ( .A(n14762), .B(n14763), .Z(n14737) );
  ANDN U14395 ( .B(n14764), .A(n14765), .Z(n14762) );
  XOR U14396 ( .A(n14763), .B(n14766), .Z(n14764) );
  IV U14397 ( .A(n14745), .Z(n14749) );
  XOR U14398 ( .A(n14745), .B(n14727), .Z(n14747) );
  XOR U14399 ( .A(n14767), .B(n14768), .Z(n14727) );
  AND U14400 ( .A(n854), .B(n14769), .Z(n14767) );
  XOR U14401 ( .A(n14770), .B(n14768), .Z(n14769) );
  NANDN U14402 ( .A(n14729), .B(n14731), .Z(n14745) );
  XOR U14403 ( .A(n14771), .B(n14772), .Z(n14731) );
  AND U14404 ( .A(n854), .B(n14773), .Z(n14771) );
  XOR U14405 ( .A(n14772), .B(n14774), .Z(n14773) );
  XOR U14406 ( .A(n14775), .B(n14776), .Z(n854) );
  AND U14407 ( .A(n14777), .B(n14778), .Z(n14775) );
  XNOR U14408 ( .A(n14776), .B(n14742), .Z(n14778) );
  XNOR U14409 ( .A(n14779), .B(n14780), .Z(n14742) );
  ANDN U14410 ( .B(n14781), .A(n14782), .Z(n14779) );
  XOR U14411 ( .A(n14780), .B(n14783), .Z(n14781) );
  XOR U14412 ( .A(n14776), .B(n14744), .Z(n14777) );
  XOR U14413 ( .A(n14784), .B(n14785), .Z(n14744) );
  AND U14414 ( .A(n858), .B(n14786), .Z(n14784) );
  XOR U14415 ( .A(n14787), .B(n14785), .Z(n14786) );
  XNOR U14416 ( .A(n14788), .B(n14789), .Z(n14776) );
  NAND U14417 ( .A(n14790), .B(n14791), .Z(n14789) );
  XOR U14418 ( .A(n14792), .B(n14768), .Z(n14791) );
  XOR U14419 ( .A(n14782), .B(n14783), .Z(n14768) );
  XOR U14420 ( .A(n14793), .B(n14794), .Z(n14783) );
  ANDN U14421 ( .B(n14795), .A(n14796), .Z(n14793) );
  XOR U14422 ( .A(n14794), .B(n14797), .Z(n14795) );
  XOR U14423 ( .A(n14798), .B(n14799), .Z(n14782) );
  XOR U14424 ( .A(n14800), .B(n14801), .Z(n14799) );
  ANDN U14425 ( .B(n14802), .A(n14803), .Z(n14800) );
  XOR U14426 ( .A(n14804), .B(n14801), .Z(n14802) );
  IV U14427 ( .A(n14780), .Z(n14798) );
  XOR U14428 ( .A(n14805), .B(n14806), .Z(n14780) );
  ANDN U14429 ( .B(n14807), .A(n14808), .Z(n14805) );
  XOR U14430 ( .A(n14806), .B(n14809), .Z(n14807) );
  IV U14431 ( .A(n14788), .Z(n14792) );
  XOR U14432 ( .A(n14788), .B(n14770), .Z(n14790) );
  XOR U14433 ( .A(n14810), .B(n14811), .Z(n14770) );
  AND U14434 ( .A(n858), .B(n14812), .Z(n14810) );
  XOR U14435 ( .A(n14813), .B(n14811), .Z(n14812) );
  NANDN U14436 ( .A(n14772), .B(n14774), .Z(n14788) );
  XOR U14437 ( .A(n14814), .B(n14815), .Z(n14774) );
  AND U14438 ( .A(n858), .B(n14816), .Z(n14814) );
  XOR U14439 ( .A(n14815), .B(n14817), .Z(n14816) );
  XOR U14440 ( .A(n14818), .B(n14819), .Z(n858) );
  AND U14441 ( .A(n14820), .B(n14821), .Z(n14818) );
  XNOR U14442 ( .A(n14819), .B(n14785), .Z(n14821) );
  XNOR U14443 ( .A(n14822), .B(n14823), .Z(n14785) );
  ANDN U14444 ( .B(n14824), .A(n14825), .Z(n14822) );
  XOR U14445 ( .A(n14823), .B(n14826), .Z(n14824) );
  XOR U14446 ( .A(n14819), .B(n14787), .Z(n14820) );
  XOR U14447 ( .A(n14827), .B(n14828), .Z(n14787) );
  AND U14448 ( .A(n862), .B(n14829), .Z(n14827) );
  XOR U14449 ( .A(n14830), .B(n14828), .Z(n14829) );
  XNOR U14450 ( .A(n14831), .B(n14832), .Z(n14819) );
  NAND U14451 ( .A(n14833), .B(n14834), .Z(n14832) );
  XOR U14452 ( .A(n14835), .B(n14811), .Z(n14834) );
  XOR U14453 ( .A(n14825), .B(n14826), .Z(n14811) );
  XOR U14454 ( .A(n14836), .B(n14837), .Z(n14826) );
  ANDN U14455 ( .B(n14838), .A(n14839), .Z(n14836) );
  XOR U14456 ( .A(n14837), .B(n14840), .Z(n14838) );
  XOR U14457 ( .A(n14841), .B(n14842), .Z(n14825) );
  XOR U14458 ( .A(n14843), .B(n14844), .Z(n14842) );
  ANDN U14459 ( .B(n14845), .A(n14846), .Z(n14843) );
  XOR U14460 ( .A(n14847), .B(n14844), .Z(n14845) );
  IV U14461 ( .A(n14823), .Z(n14841) );
  XOR U14462 ( .A(n14848), .B(n14849), .Z(n14823) );
  ANDN U14463 ( .B(n14850), .A(n14851), .Z(n14848) );
  XOR U14464 ( .A(n14849), .B(n14852), .Z(n14850) );
  IV U14465 ( .A(n14831), .Z(n14835) );
  XOR U14466 ( .A(n14831), .B(n14813), .Z(n14833) );
  XOR U14467 ( .A(n14853), .B(n14854), .Z(n14813) );
  AND U14468 ( .A(n862), .B(n14855), .Z(n14853) );
  XOR U14469 ( .A(n14856), .B(n14854), .Z(n14855) );
  NANDN U14470 ( .A(n14815), .B(n14817), .Z(n14831) );
  XOR U14471 ( .A(n14857), .B(n14858), .Z(n14817) );
  AND U14472 ( .A(n862), .B(n14859), .Z(n14857) );
  XOR U14473 ( .A(n14858), .B(n14860), .Z(n14859) );
  XOR U14474 ( .A(n14861), .B(n14862), .Z(n862) );
  AND U14475 ( .A(n14863), .B(n14864), .Z(n14861) );
  XNOR U14476 ( .A(n14862), .B(n14828), .Z(n14864) );
  XNOR U14477 ( .A(n14865), .B(n14866), .Z(n14828) );
  ANDN U14478 ( .B(n14867), .A(n14868), .Z(n14865) );
  XOR U14479 ( .A(n14866), .B(n14869), .Z(n14867) );
  XOR U14480 ( .A(n14862), .B(n14830), .Z(n14863) );
  XOR U14481 ( .A(n14870), .B(n14871), .Z(n14830) );
  AND U14482 ( .A(n866), .B(n14872), .Z(n14870) );
  XOR U14483 ( .A(n14873), .B(n14871), .Z(n14872) );
  XNOR U14484 ( .A(n14874), .B(n14875), .Z(n14862) );
  NAND U14485 ( .A(n14876), .B(n14877), .Z(n14875) );
  XOR U14486 ( .A(n14878), .B(n14854), .Z(n14877) );
  XOR U14487 ( .A(n14868), .B(n14869), .Z(n14854) );
  XOR U14488 ( .A(n14879), .B(n14880), .Z(n14869) );
  ANDN U14489 ( .B(n14881), .A(n14882), .Z(n14879) );
  XOR U14490 ( .A(n14880), .B(n14883), .Z(n14881) );
  XOR U14491 ( .A(n14884), .B(n14885), .Z(n14868) );
  XOR U14492 ( .A(n14886), .B(n14887), .Z(n14885) );
  ANDN U14493 ( .B(n14888), .A(n14889), .Z(n14886) );
  XOR U14494 ( .A(n14890), .B(n14887), .Z(n14888) );
  IV U14495 ( .A(n14866), .Z(n14884) );
  XOR U14496 ( .A(n14891), .B(n14892), .Z(n14866) );
  ANDN U14497 ( .B(n14893), .A(n14894), .Z(n14891) );
  XOR U14498 ( .A(n14892), .B(n14895), .Z(n14893) );
  IV U14499 ( .A(n14874), .Z(n14878) );
  XOR U14500 ( .A(n14874), .B(n14856), .Z(n14876) );
  XOR U14501 ( .A(n14896), .B(n14897), .Z(n14856) );
  AND U14502 ( .A(n866), .B(n14898), .Z(n14896) );
  XOR U14503 ( .A(n14899), .B(n14897), .Z(n14898) );
  NANDN U14504 ( .A(n14858), .B(n14860), .Z(n14874) );
  XOR U14505 ( .A(n14900), .B(n14901), .Z(n14860) );
  AND U14506 ( .A(n866), .B(n14902), .Z(n14900) );
  XOR U14507 ( .A(n14901), .B(n14903), .Z(n14902) );
  XOR U14508 ( .A(n14904), .B(n14905), .Z(n866) );
  AND U14509 ( .A(n14906), .B(n14907), .Z(n14904) );
  XNOR U14510 ( .A(n14905), .B(n14871), .Z(n14907) );
  XNOR U14511 ( .A(n14908), .B(n14909), .Z(n14871) );
  ANDN U14512 ( .B(n14910), .A(n14911), .Z(n14908) );
  XOR U14513 ( .A(n14909), .B(n14912), .Z(n14910) );
  XOR U14514 ( .A(n14905), .B(n14873), .Z(n14906) );
  XOR U14515 ( .A(n14913), .B(n14914), .Z(n14873) );
  AND U14516 ( .A(n870), .B(n14915), .Z(n14913) );
  XOR U14517 ( .A(n14916), .B(n14914), .Z(n14915) );
  XNOR U14518 ( .A(n14917), .B(n14918), .Z(n14905) );
  NAND U14519 ( .A(n14919), .B(n14920), .Z(n14918) );
  XOR U14520 ( .A(n14921), .B(n14897), .Z(n14920) );
  XOR U14521 ( .A(n14911), .B(n14912), .Z(n14897) );
  XOR U14522 ( .A(n14922), .B(n14923), .Z(n14912) );
  ANDN U14523 ( .B(n14924), .A(n14925), .Z(n14922) );
  XOR U14524 ( .A(n14923), .B(n14926), .Z(n14924) );
  XOR U14525 ( .A(n14927), .B(n14928), .Z(n14911) );
  XOR U14526 ( .A(n14929), .B(n14930), .Z(n14928) );
  ANDN U14527 ( .B(n14931), .A(n14932), .Z(n14929) );
  XOR U14528 ( .A(n14933), .B(n14930), .Z(n14931) );
  IV U14529 ( .A(n14909), .Z(n14927) );
  XOR U14530 ( .A(n14934), .B(n14935), .Z(n14909) );
  ANDN U14531 ( .B(n14936), .A(n14937), .Z(n14934) );
  XOR U14532 ( .A(n14935), .B(n14938), .Z(n14936) );
  IV U14533 ( .A(n14917), .Z(n14921) );
  XOR U14534 ( .A(n14917), .B(n14899), .Z(n14919) );
  XOR U14535 ( .A(n14939), .B(n14940), .Z(n14899) );
  AND U14536 ( .A(n870), .B(n14941), .Z(n14939) );
  XOR U14537 ( .A(n14942), .B(n14940), .Z(n14941) );
  NANDN U14538 ( .A(n14901), .B(n14903), .Z(n14917) );
  XOR U14539 ( .A(n14943), .B(n14944), .Z(n14903) );
  AND U14540 ( .A(n870), .B(n14945), .Z(n14943) );
  XOR U14541 ( .A(n14944), .B(n14946), .Z(n14945) );
  XOR U14542 ( .A(n14947), .B(n14948), .Z(n870) );
  AND U14543 ( .A(n14949), .B(n14950), .Z(n14947) );
  XNOR U14544 ( .A(n14948), .B(n14914), .Z(n14950) );
  XNOR U14545 ( .A(n14951), .B(n14952), .Z(n14914) );
  ANDN U14546 ( .B(n14953), .A(n14954), .Z(n14951) );
  XOR U14547 ( .A(n14952), .B(n14955), .Z(n14953) );
  XOR U14548 ( .A(n14948), .B(n14916), .Z(n14949) );
  XOR U14549 ( .A(n14956), .B(n14957), .Z(n14916) );
  AND U14550 ( .A(n874), .B(n14958), .Z(n14956) );
  XOR U14551 ( .A(n14959), .B(n14957), .Z(n14958) );
  XNOR U14552 ( .A(n14960), .B(n14961), .Z(n14948) );
  NAND U14553 ( .A(n14962), .B(n14963), .Z(n14961) );
  XOR U14554 ( .A(n14964), .B(n14940), .Z(n14963) );
  XOR U14555 ( .A(n14954), .B(n14955), .Z(n14940) );
  XOR U14556 ( .A(n14965), .B(n14966), .Z(n14955) );
  ANDN U14557 ( .B(n14967), .A(n14968), .Z(n14965) );
  XOR U14558 ( .A(n14966), .B(n14969), .Z(n14967) );
  XOR U14559 ( .A(n14970), .B(n14971), .Z(n14954) );
  XOR U14560 ( .A(n14972), .B(n14973), .Z(n14971) );
  ANDN U14561 ( .B(n14974), .A(n14975), .Z(n14972) );
  XOR U14562 ( .A(n14976), .B(n14973), .Z(n14974) );
  IV U14563 ( .A(n14952), .Z(n14970) );
  XOR U14564 ( .A(n14977), .B(n14978), .Z(n14952) );
  ANDN U14565 ( .B(n14979), .A(n14980), .Z(n14977) );
  XOR U14566 ( .A(n14978), .B(n14981), .Z(n14979) );
  IV U14567 ( .A(n14960), .Z(n14964) );
  XOR U14568 ( .A(n14960), .B(n14942), .Z(n14962) );
  XOR U14569 ( .A(n14982), .B(n14983), .Z(n14942) );
  AND U14570 ( .A(n874), .B(n14984), .Z(n14982) );
  XOR U14571 ( .A(n14985), .B(n14983), .Z(n14984) );
  NANDN U14572 ( .A(n14944), .B(n14946), .Z(n14960) );
  XOR U14573 ( .A(n14986), .B(n14987), .Z(n14946) );
  AND U14574 ( .A(n874), .B(n14988), .Z(n14986) );
  XOR U14575 ( .A(n14987), .B(n14989), .Z(n14988) );
  XOR U14576 ( .A(n14990), .B(n14991), .Z(n874) );
  AND U14577 ( .A(n14992), .B(n14993), .Z(n14990) );
  XNOR U14578 ( .A(n14991), .B(n14957), .Z(n14993) );
  XNOR U14579 ( .A(n14994), .B(n14995), .Z(n14957) );
  ANDN U14580 ( .B(n14996), .A(n14997), .Z(n14994) );
  XOR U14581 ( .A(n14995), .B(n14998), .Z(n14996) );
  XOR U14582 ( .A(n14991), .B(n14959), .Z(n14992) );
  XOR U14583 ( .A(n14999), .B(n15000), .Z(n14959) );
  AND U14584 ( .A(n878), .B(n15001), .Z(n14999) );
  XOR U14585 ( .A(n15002), .B(n15000), .Z(n15001) );
  XNOR U14586 ( .A(n15003), .B(n15004), .Z(n14991) );
  NAND U14587 ( .A(n15005), .B(n15006), .Z(n15004) );
  XOR U14588 ( .A(n15007), .B(n14983), .Z(n15006) );
  XOR U14589 ( .A(n14997), .B(n14998), .Z(n14983) );
  XOR U14590 ( .A(n15008), .B(n15009), .Z(n14998) );
  ANDN U14591 ( .B(n15010), .A(n15011), .Z(n15008) );
  XOR U14592 ( .A(n15009), .B(n15012), .Z(n15010) );
  XOR U14593 ( .A(n15013), .B(n15014), .Z(n14997) );
  XOR U14594 ( .A(n15015), .B(n15016), .Z(n15014) );
  ANDN U14595 ( .B(n15017), .A(n15018), .Z(n15015) );
  XOR U14596 ( .A(n15019), .B(n15016), .Z(n15017) );
  IV U14597 ( .A(n14995), .Z(n15013) );
  XOR U14598 ( .A(n15020), .B(n15021), .Z(n14995) );
  ANDN U14599 ( .B(n15022), .A(n15023), .Z(n15020) );
  XOR U14600 ( .A(n15021), .B(n15024), .Z(n15022) );
  IV U14601 ( .A(n15003), .Z(n15007) );
  XOR U14602 ( .A(n15003), .B(n14985), .Z(n15005) );
  XOR U14603 ( .A(n15025), .B(n15026), .Z(n14985) );
  AND U14604 ( .A(n878), .B(n15027), .Z(n15025) );
  XOR U14605 ( .A(n15028), .B(n15026), .Z(n15027) );
  NANDN U14606 ( .A(n14987), .B(n14989), .Z(n15003) );
  XOR U14607 ( .A(n15029), .B(n15030), .Z(n14989) );
  AND U14608 ( .A(n878), .B(n15031), .Z(n15029) );
  XOR U14609 ( .A(n15030), .B(n15032), .Z(n15031) );
  XOR U14610 ( .A(n15033), .B(n15034), .Z(n878) );
  AND U14611 ( .A(n15035), .B(n15036), .Z(n15033) );
  XNOR U14612 ( .A(n15034), .B(n15000), .Z(n15036) );
  XNOR U14613 ( .A(n15037), .B(n15038), .Z(n15000) );
  ANDN U14614 ( .B(n15039), .A(n15040), .Z(n15037) );
  XOR U14615 ( .A(n15038), .B(n15041), .Z(n15039) );
  XOR U14616 ( .A(n15034), .B(n15002), .Z(n15035) );
  XOR U14617 ( .A(n15042), .B(n15043), .Z(n15002) );
  AND U14618 ( .A(n882), .B(n15044), .Z(n15042) );
  XOR U14619 ( .A(n15045), .B(n15043), .Z(n15044) );
  XNOR U14620 ( .A(n15046), .B(n15047), .Z(n15034) );
  NAND U14621 ( .A(n15048), .B(n15049), .Z(n15047) );
  XOR U14622 ( .A(n15050), .B(n15026), .Z(n15049) );
  XOR U14623 ( .A(n15040), .B(n15041), .Z(n15026) );
  XOR U14624 ( .A(n15051), .B(n15052), .Z(n15041) );
  ANDN U14625 ( .B(n15053), .A(n15054), .Z(n15051) );
  XOR U14626 ( .A(n15052), .B(n15055), .Z(n15053) );
  XOR U14627 ( .A(n15056), .B(n15057), .Z(n15040) );
  XOR U14628 ( .A(n15058), .B(n15059), .Z(n15057) );
  ANDN U14629 ( .B(n15060), .A(n15061), .Z(n15058) );
  XOR U14630 ( .A(n15062), .B(n15059), .Z(n15060) );
  IV U14631 ( .A(n15038), .Z(n15056) );
  XOR U14632 ( .A(n15063), .B(n15064), .Z(n15038) );
  ANDN U14633 ( .B(n15065), .A(n15066), .Z(n15063) );
  XOR U14634 ( .A(n15064), .B(n15067), .Z(n15065) );
  IV U14635 ( .A(n15046), .Z(n15050) );
  XOR U14636 ( .A(n15046), .B(n15028), .Z(n15048) );
  XOR U14637 ( .A(n15068), .B(n15069), .Z(n15028) );
  AND U14638 ( .A(n882), .B(n15070), .Z(n15068) );
  XOR U14639 ( .A(n15071), .B(n15069), .Z(n15070) );
  NANDN U14640 ( .A(n15030), .B(n15032), .Z(n15046) );
  XOR U14641 ( .A(n15072), .B(n15073), .Z(n15032) );
  AND U14642 ( .A(n882), .B(n15074), .Z(n15072) );
  XOR U14643 ( .A(n15073), .B(n15075), .Z(n15074) );
  XOR U14644 ( .A(n15076), .B(n15077), .Z(n882) );
  AND U14645 ( .A(n15078), .B(n15079), .Z(n15076) );
  XNOR U14646 ( .A(n15077), .B(n15043), .Z(n15079) );
  XNOR U14647 ( .A(n15080), .B(n15081), .Z(n15043) );
  ANDN U14648 ( .B(n15082), .A(n15083), .Z(n15080) );
  XOR U14649 ( .A(n15081), .B(n15084), .Z(n15082) );
  XOR U14650 ( .A(n15077), .B(n15045), .Z(n15078) );
  XOR U14651 ( .A(n15085), .B(n15086), .Z(n15045) );
  AND U14652 ( .A(n886), .B(n15087), .Z(n15085) );
  XOR U14653 ( .A(n15088), .B(n15086), .Z(n15087) );
  XNOR U14654 ( .A(n15089), .B(n15090), .Z(n15077) );
  NAND U14655 ( .A(n15091), .B(n15092), .Z(n15090) );
  XOR U14656 ( .A(n15093), .B(n15069), .Z(n15092) );
  XOR U14657 ( .A(n15083), .B(n15084), .Z(n15069) );
  XOR U14658 ( .A(n15094), .B(n15095), .Z(n15084) );
  ANDN U14659 ( .B(n15096), .A(n15097), .Z(n15094) );
  XOR U14660 ( .A(n15095), .B(n15098), .Z(n15096) );
  XOR U14661 ( .A(n15099), .B(n15100), .Z(n15083) );
  XOR U14662 ( .A(n15101), .B(n15102), .Z(n15100) );
  ANDN U14663 ( .B(n15103), .A(n15104), .Z(n15101) );
  XOR U14664 ( .A(n15105), .B(n15102), .Z(n15103) );
  IV U14665 ( .A(n15081), .Z(n15099) );
  XOR U14666 ( .A(n15106), .B(n15107), .Z(n15081) );
  ANDN U14667 ( .B(n15108), .A(n15109), .Z(n15106) );
  XOR U14668 ( .A(n15107), .B(n15110), .Z(n15108) );
  IV U14669 ( .A(n15089), .Z(n15093) );
  XOR U14670 ( .A(n15089), .B(n15071), .Z(n15091) );
  XOR U14671 ( .A(n15111), .B(n15112), .Z(n15071) );
  AND U14672 ( .A(n886), .B(n15113), .Z(n15111) );
  XOR U14673 ( .A(n15114), .B(n15112), .Z(n15113) );
  NANDN U14674 ( .A(n15073), .B(n15075), .Z(n15089) );
  XOR U14675 ( .A(n15115), .B(n15116), .Z(n15075) );
  AND U14676 ( .A(n886), .B(n15117), .Z(n15115) );
  XOR U14677 ( .A(n15116), .B(n15118), .Z(n15117) );
  XOR U14678 ( .A(n15119), .B(n15120), .Z(n886) );
  AND U14679 ( .A(n15121), .B(n15122), .Z(n15119) );
  XNOR U14680 ( .A(n15120), .B(n15086), .Z(n15122) );
  XNOR U14681 ( .A(n15123), .B(n15124), .Z(n15086) );
  ANDN U14682 ( .B(n15125), .A(n15126), .Z(n15123) );
  XOR U14683 ( .A(n15124), .B(n15127), .Z(n15125) );
  XOR U14684 ( .A(n15120), .B(n15088), .Z(n15121) );
  XOR U14685 ( .A(n15128), .B(n15129), .Z(n15088) );
  AND U14686 ( .A(n890), .B(n15130), .Z(n15128) );
  XOR U14687 ( .A(n15131), .B(n15129), .Z(n15130) );
  XNOR U14688 ( .A(n15132), .B(n15133), .Z(n15120) );
  NAND U14689 ( .A(n15134), .B(n15135), .Z(n15133) );
  XOR U14690 ( .A(n15136), .B(n15112), .Z(n15135) );
  XOR U14691 ( .A(n15126), .B(n15127), .Z(n15112) );
  XOR U14692 ( .A(n15137), .B(n15138), .Z(n15127) );
  ANDN U14693 ( .B(n15139), .A(n15140), .Z(n15137) );
  XOR U14694 ( .A(n15138), .B(n15141), .Z(n15139) );
  XOR U14695 ( .A(n15142), .B(n15143), .Z(n15126) );
  XOR U14696 ( .A(n15144), .B(n15145), .Z(n15143) );
  ANDN U14697 ( .B(n15146), .A(n15147), .Z(n15144) );
  XOR U14698 ( .A(n15148), .B(n15145), .Z(n15146) );
  IV U14699 ( .A(n15124), .Z(n15142) );
  XOR U14700 ( .A(n15149), .B(n15150), .Z(n15124) );
  ANDN U14701 ( .B(n15151), .A(n15152), .Z(n15149) );
  XOR U14702 ( .A(n15150), .B(n15153), .Z(n15151) );
  IV U14703 ( .A(n15132), .Z(n15136) );
  XOR U14704 ( .A(n15132), .B(n15114), .Z(n15134) );
  XOR U14705 ( .A(n15154), .B(n15155), .Z(n15114) );
  AND U14706 ( .A(n890), .B(n15156), .Z(n15154) );
  XOR U14707 ( .A(n15157), .B(n15155), .Z(n15156) );
  NANDN U14708 ( .A(n15116), .B(n15118), .Z(n15132) );
  XOR U14709 ( .A(n15158), .B(n15159), .Z(n15118) );
  AND U14710 ( .A(n890), .B(n15160), .Z(n15158) );
  XOR U14711 ( .A(n15159), .B(n15161), .Z(n15160) );
  XOR U14712 ( .A(n15162), .B(n15163), .Z(n890) );
  AND U14713 ( .A(n15164), .B(n15165), .Z(n15162) );
  XNOR U14714 ( .A(n15163), .B(n15129), .Z(n15165) );
  XNOR U14715 ( .A(n15166), .B(n15167), .Z(n15129) );
  ANDN U14716 ( .B(n15168), .A(n15169), .Z(n15166) );
  XOR U14717 ( .A(n15167), .B(n15170), .Z(n15168) );
  XOR U14718 ( .A(n15163), .B(n15131), .Z(n15164) );
  XOR U14719 ( .A(n15171), .B(n15172), .Z(n15131) );
  AND U14720 ( .A(n894), .B(n15173), .Z(n15171) );
  XOR U14721 ( .A(n15174), .B(n15172), .Z(n15173) );
  XNOR U14722 ( .A(n15175), .B(n15176), .Z(n15163) );
  NAND U14723 ( .A(n15177), .B(n15178), .Z(n15176) );
  XOR U14724 ( .A(n15179), .B(n15155), .Z(n15178) );
  XOR U14725 ( .A(n15169), .B(n15170), .Z(n15155) );
  XOR U14726 ( .A(n15180), .B(n15181), .Z(n15170) );
  ANDN U14727 ( .B(n15182), .A(n15183), .Z(n15180) );
  XOR U14728 ( .A(n15181), .B(n15184), .Z(n15182) );
  XOR U14729 ( .A(n15185), .B(n15186), .Z(n15169) );
  XOR U14730 ( .A(n15187), .B(n15188), .Z(n15186) );
  ANDN U14731 ( .B(n15189), .A(n15190), .Z(n15187) );
  XOR U14732 ( .A(n15191), .B(n15188), .Z(n15189) );
  IV U14733 ( .A(n15167), .Z(n15185) );
  XOR U14734 ( .A(n15192), .B(n15193), .Z(n15167) );
  ANDN U14735 ( .B(n15194), .A(n15195), .Z(n15192) );
  XOR U14736 ( .A(n15193), .B(n15196), .Z(n15194) );
  IV U14737 ( .A(n15175), .Z(n15179) );
  XOR U14738 ( .A(n15175), .B(n15157), .Z(n15177) );
  XOR U14739 ( .A(n15197), .B(n15198), .Z(n15157) );
  AND U14740 ( .A(n894), .B(n15199), .Z(n15197) );
  XOR U14741 ( .A(n15200), .B(n15198), .Z(n15199) );
  NANDN U14742 ( .A(n15159), .B(n15161), .Z(n15175) );
  XOR U14743 ( .A(n15201), .B(n15202), .Z(n15161) );
  AND U14744 ( .A(n894), .B(n15203), .Z(n15201) );
  XOR U14745 ( .A(n15202), .B(n15204), .Z(n15203) );
  XOR U14746 ( .A(n15205), .B(n15206), .Z(n894) );
  AND U14747 ( .A(n15207), .B(n15208), .Z(n15205) );
  XNOR U14748 ( .A(n15206), .B(n15172), .Z(n15208) );
  XNOR U14749 ( .A(n15209), .B(n15210), .Z(n15172) );
  ANDN U14750 ( .B(n15211), .A(n15212), .Z(n15209) );
  XOR U14751 ( .A(n15210), .B(n15213), .Z(n15211) );
  XOR U14752 ( .A(n15206), .B(n15174), .Z(n15207) );
  XOR U14753 ( .A(n15214), .B(n15215), .Z(n15174) );
  AND U14754 ( .A(n898), .B(n15216), .Z(n15214) );
  XOR U14755 ( .A(n15217), .B(n15215), .Z(n15216) );
  XNOR U14756 ( .A(n15218), .B(n15219), .Z(n15206) );
  NAND U14757 ( .A(n15220), .B(n15221), .Z(n15219) );
  XOR U14758 ( .A(n15222), .B(n15198), .Z(n15221) );
  XOR U14759 ( .A(n15212), .B(n15213), .Z(n15198) );
  XOR U14760 ( .A(n15223), .B(n15224), .Z(n15213) );
  ANDN U14761 ( .B(n15225), .A(n15226), .Z(n15223) );
  XOR U14762 ( .A(n15224), .B(n15227), .Z(n15225) );
  XOR U14763 ( .A(n15228), .B(n15229), .Z(n15212) );
  XOR U14764 ( .A(n15230), .B(n15231), .Z(n15229) );
  ANDN U14765 ( .B(n15232), .A(n15233), .Z(n15230) );
  XOR U14766 ( .A(n15234), .B(n15231), .Z(n15232) );
  IV U14767 ( .A(n15210), .Z(n15228) );
  XOR U14768 ( .A(n15235), .B(n15236), .Z(n15210) );
  ANDN U14769 ( .B(n15237), .A(n15238), .Z(n15235) );
  XOR U14770 ( .A(n15236), .B(n15239), .Z(n15237) );
  IV U14771 ( .A(n15218), .Z(n15222) );
  XOR U14772 ( .A(n15218), .B(n15200), .Z(n15220) );
  XOR U14773 ( .A(n15240), .B(n15241), .Z(n15200) );
  AND U14774 ( .A(n898), .B(n15242), .Z(n15240) );
  XOR U14775 ( .A(n15243), .B(n15241), .Z(n15242) );
  NANDN U14776 ( .A(n15202), .B(n15204), .Z(n15218) );
  XOR U14777 ( .A(n15244), .B(n15245), .Z(n15204) );
  AND U14778 ( .A(n898), .B(n15246), .Z(n15244) );
  XOR U14779 ( .A(n15245), .B(n15247), .Z(n15246) );
  XOR U14780 ( .A(n15248), .B(n15249), .Z(n898) );
  AND U14781 ( .A(n15250), .B(n15251), .Z(n15248) );
  XNOR U14782 ( .A(n15249), .B(n15215), .Z(n15251) );
  XNOR U14783 ( .A(n15252), .B(n15253), .Z(n15215) );
  ANDN U14784 ( .B(n15254), .A(n15255), .Z(n15252) );
  XOR U14785 ( .A(n15253), .B(n15256), .Z(n15254) );
  XOR U14786 ( .A(n15249), .B(n15217), .Z(n15250) );
  XOR U14787 ( .A(n15257), .B(n15258), .Z(n15217) );
  AND U14788 ( .A(n902), .B(n15259), .Z(n15257) );
  XOR U14789 ( .A(n15260), .B(n15258), .Z(n15259) );
  XNOR U14790 ( .A(n15261), .B(n15262), .Z(n15249) );
  NAND U14791 ( .A(n15263), .B(n15264), .Z(n15262) );
  XOR U14792 ( .A(n15265), .B(n15241), .Z(n15264) );
  XOR U14793 ( .A(n15255), .B(n15256), .Z(n15241) );
  XOR U14794 ( .A(n15266), .B(n15267), .Z(n15256) );
  ANDN U14795 ( .B(n15268), .A(n15269), .Z(n15266) );
  XOR U14796 ( .A(n15267), .B(n15270), .Z(n15268) );
  XOR U14797 ( .A(n15271), .B(n15272), .Z(n15255) );
  XOR U14798 ( .A(n15273), .B(n15274), .Z(n15272) );
  ANDN U14799 ( .B(n15275), .A(n15276), .Z(n15273) );
  XOR U14800 ( .A(n15277), .B(n15274), .Z(n15275) );
  IV U14801 ( .A(n15253), .Z(n15271) );
  XOR U14802 ( .A(n15278), .B(n15279), .Z(n15253) );
  ANDN U14803 ( .B(n15280), .A(n15281), .Z(n15278) );
  XOR U14804 ( .A(n15279), .B(n15282), .Z(n15280) );
  IV U14805 ( .A(n15261), .Z(n15265) );
  XOR U14806 ( .A(n15261), .B(n15243), .Z(n15263) );
  XOR U14807 ( .A(n15283), .B(n15284), .Z(n15243) );
  AND U14808 ( .A(n902), .B(n15285), .Z(n15283) );
  XOR U14809 ( .A(n15286), .B(n15284), .Z(n15285) );
  NANDN U14810 ( .A(n15245), .B(n15247), .Z(n15261) );
  XOR U14811 ( .A(n15287), .B(n15288), .Z(n15247) );
  AND U14812 ( .A(n902), .B(n15289), .Z(n15287) );
  XOR U14813 ( .A(n15288), .B(n15290), .Z(n15289) );
  XOR U14814 ( .A(n15291), .B(n15292), .Z(n902) );
  AND U14815 ( .A(n15293), .B(n15294), .Z(n15291) );
  XNOR U14816 ( .A(n15292), .B(n15258), .Z(n15294) );
  XNOR U14817 ( .A(n15295), .B(n15296), .Z(n15258) );
  ANDN U14818 ( .B(n15297), .A(n15298), .Z(n15295) );
  XOR U14819 ( .A(n15296), .B(n15299), .Z(n15297) );
  XOR U14820 ( .A(n15292), .B(n15260), .Z(n15293) );
  XOR U14821 ( .A(n15300), .B(n15301), .Z(n15260) );
  AND U14822 ( .A(n906), .B(n15302), .Z(n15300) );
  XOR U14823 ( .A(n15303), .B(n15301), .Z(n15302) );
  XNOR U14824 ( .A(n15304), .B(n15305), .Z(n15292) );
  NAND U14825 ( .A(n15306), .B(n15307), .Z(n15305) );
  XOR U14826 ( .A(n15308), .B(n15284), .Z(n15307) );
  XOR U14827 ( .A(n15298), .B(n15299), .Z(n15284) );
  XOR U14828 ( .A(n15309), .B(n15310), .Z(n15299) );
  ANDN U14829 ( .B(n15311), .A(n15312), .Z(n15309) );
  XOR U14830 ( .A(n15310), .B(n15313), .Z(n15311) );
  XOR U14831 ( .A(n15314), .B(n15315), .Z(n15298) );
  XOR U14832 ( .A(n15316), .B(n15317), .Z(n15315) );
  ANDN U14833 ( .B(n15318), .A(n15319), .Z(n15316) );
  XOR U14834 ( .A(n15320), .B(n15317), .Z(n15318) );
  IV U14835 ( .A(n15296), .Z(n15314) );
  XOR U14836 ( .A(n15321), .B(n15322), .Z(n15296) );
  ANDN U14837 ( .B(n15323), .A(n15324), .Z(n15321) );
  XOR U14838 ( .A(n15322), .B(n15325), .Z(n15323) );
  IV U14839 ( .A(n15304), .Z(n15308) );
  XOR U14840 ( .A(n15304), .B(n15286), .Z(n15306) );
  XOR U14841 ( .A(n15326), .B(n15327), .Z(n15286) );
  AND U14842 ( .A(n906), .B(n15328), .Z(n15326) );
  XOR U14843 ( .A(n15329), .B(n15327), .Z(n15328) );
  NANDN U14844 ( .A(n15288), .B(n15290), .Z(n15304) );
  XOR U14845 ( .A(n15330), .B(n15331), .Z(n15290) );
  AND U14846 ( .A(n906), .B(n15332), .Z(n15330) );
  XOR U14847 ( .A(n15331), .B(n15333), .Z(n15332) );
  XOR U14848 ( .A(n15334), .B(n15335), .Z(n906) );
  AND U14849 ( .A(n15336), .B(n15337), .Z(n15334) );
  XNOR U14850 ( .A(n15335), .B(n15301), .Z(n15337) );
  XNOR U14851 ( .A(n15338), .B(n15339), .Z(n15301) );
  ANDN U14852 ( .B(n15340), .A(n15341), .Z(n15338) );
  XOR U14853 ( .A(n15339), .B(n15342), .Z(n15340) );
  XOR U14854 ( .A(n15335), .B(n15303), .Z(n15336) );
  XOR U14855 ( .A(n15343), .B(n15344), .Z(n15303) );
  AND U14856 ( .A(n910), .B(n15345), .Z(n15343) );
  XOR U14857 ( .A(n15346), .B(n15344), .Z(n15345) );
  XNOR U14858 ( .A(n15347), .B(n15348), .Z(n15335) );
  NAND U14859 ( .A(n15349), .B(n15350), .Z(n15348) );
  XOR U14860 ( .A(n15351), .B(n15327), .Z(n15350) );
  XOR U14861 ( .A(n15341), .B(n15342), .Z(n15327) );
  XOR U14862 ( .A(n15352), .B(n15353), .Z(n15342) );
  ANDN U14863 ( .B(n15354), .A(n15355), .Z(n15352) );
  XOR U14864 ( .A(n15353), .B(n15356), .Z(n15354) );
  XOR U14865 ( .A(n15357), .B(n15358), .Z(n15341) );
  XOR U14866 ( .A(n15359), .B(n15360), .Z(n15358) );
  ANDN U14867 ( .B(n15361), .A(n15362), .Z(n15359) );
  XOR U14868 ( .A(n15363), .B(n15360), .Z(n15361) );
  IV U14869 ( .A(n15339), .Z(n15357) );
  XOR U14870 ( .A(n15364), .B(n15365), .Z(n15339) );
  ANDN U14871 ( .B(n15366), .A(n15367), .Z(n15364) );
  XOR U14872 ( .A(n15365), .B(n15368), .Z(n15366) );
  IV U14873 ( .A(n15347), .Z(n15351) );
  XOR U14874 ( .A(n15347), .B(n15329), .Z(n15349) );
  XOR U14875 ( .A(n15369), .B(n15370), .Z(n15329) );
  AND U14876 ( .A(n910), .B(n15371), .Z(n15369) );
  XOR U14877 ( .A(n15372), .B(n15370), .Z(n15371) );
  NANDN U14878 ( .A(n15331), .B(n15333), .Z(n15347) );
  XOR U14879 ( .A(n15373), .B(n15374), .Z(n15333) );
  AND U14880 ( .A(n910), .B(n15375), .Z(n15373) );
  XOR U14881 ( .A(n15374), .B(n15376), .Z(n15375) );
  XOR U14882 ( .A(n15377), .B(n15378), .Z(n910) );
  AND U14883 ( .A(n15379), .B(n15380), .Z(n15377) );
  XNOR U14884 ( .A(n15378), .B(n15344), .Z(n15380) );
  XNOR U14885 ( .A(n15381), .B(n15382), .Z(n15344) );
  ANDN U14886 ( .B(n15383), .A(n15384), .Z(n15381) );
  XOR U14887 ( .A(n15382), .B(n15385), .Z(n15383) );
  XOR U14888 ( .A(n15378), .B(n15346), .Z(n15379) );
  XOR U14889 ( .A(n15386), .B(n15387), .Z(n15346) );
  AND U14890 ( .A(n914), .B(n15388), .Z(n15386) );
  XOR U14891 ( .A(n15389), .B(n15387), .Z(n15388) );
  XNOR U14892 ( .A(n15390), .B(n15391), .Z(n15378) );
  NAND U14893 ( .A(n15392), .B(n15393), .Z(n15391) );
  XOR U14894 ( .A(n15394), .B(n15370), .Z(n15393) );
  XOR U14895 ( .A(n15384), .B(n15385), .Z(n15370) );
  XOR U14896 ( .A(n15395), .B(n15396), .Z(n15385) );
  ANDN U14897 ( .B(n15397), .A(n15398), .Z(n15395) );
  XOR U14898 ( .A(n15396), .B(n15399), .Z(n15397) );
  XOR U14899 ( .A(n15400), .B(n15401), .Z(n15384) );
  XOR U14900 ( .A(n15402), .B(n15403), .Z(n15401) );
  ANDN U14901 ( .B(n15404), .A(n15405), .Z(n15402) );
  XOR U14902 ( .A(n15406), .B(n15403), .Z(n15404) );
  IV U14903 ( .A(n15382), .Z(n15400) );
  XOR U14904 ( .A(n15407), .B(n15408), .Z(n15382) );
  ANDN U14905 ( .B(n15409), .A(n15410), .Z(n15407) );
  XOR U14906 ( .A(n15408), .B(n15411), .Z(n15409) );
  IV U14907 ( .A(n15390), .Z(n15394) );
  XOR U14908 ( .A(n15390), .B(n15372), .Z(n15392) );
  XOR U14909 ( .A(n15412), .B(n15413), .Z(n15372) );
  AND U14910 ( .A(n914), .B(n15414), .Z(n15412) );
  XOR U14911 ( .A(n15415), .B(n15413), .Z(n15414) );
  NANDN U14912 ( .A(n15374), .B(n15376), .Z(n15390) );
  XOR U14913 ( .A(n15416), .B(n15417), .Z(n15376) );
  AND U14914 ( .A(n914), .B(n15418), .Z(n15416) );
  XOR U14915 ( .A(n15417), .B(n15419), .Z(n15418) );
  XOR U14916 ( .A(n15420), .B(n15421), .Z(n914) );
  AND U14917 ( .A(n15422), .B(n15423), .Z(n15420) );
  XNOR U14918 ( .A(n15421), .B(n15387), .Z(n15423) );
  XNOR U14919 ( .A(n15424), .B(n15425), .Z(n15387) );
  ANDN U14920 ( .B(n15426), .A(n15427), .Z(n15424) );
  XOR U14921 ( .A(n15425), .B(n15428), .Z(n15426) );
  XOR U14922 ( .A(n15421), .B(n15389), .Z(n15422) );
  XOR U14923 ( .A(n15429), .B(n15430), .Z(n15389) );
  AND U14924 ( .A(n918), .B(n15431), .Z(n15429) );
  XOR U14925 ( .A(n15432), .B(n15430), .Z(n15431) );
  XNOR U14926 ( .A(n15433), .B(n15434), .Z(n15421) );
  NAND U14927 ( .A(n15435), .B(n15436), .Z(n15434) );
  XOR U14928 ( .A(n15437), .B(n15413), .Z(n15436) );
  XOR U14929 ( .A(n15427), .B(n15428), .Z(n15413) );
  XOR U14930 ( .A(n15438), .B(n15439), .Z(n15428) );
  ANDN U14931 ( .B(n15440), .A(n15441), .Z(n15438) );
  XOR U14932 ( .A(n15439), .B(n15442), .Z(n15440) );
  XOR U14933 ( .A(n15443), .B(n15444), .Z(n15427) );
  XOR U14934 ( .A(n15445), .B(n15446), .Z(n15444) );
  ANDN U14935 ( .B(n15447), .A(n15448), .Z(n15445) );
  XOR U14936 ( .A(n15449), .B(n15446), .Z(n15447) );
  IV U14937 ( .A(n15425), .Z(n15443) );
  XOR U14938 ( .A(n15450), .B(n15451), .Z(n15425) );
  ANDN U14939 ( .B(n15452), .A(n15453), .Z(n15450) );
  XOR U14940 ( .A(n15451), .B(n15454), .Z(n15452) );
  IV U14941 ( .A(n15433), .Z(n15437) );
  XOR U14942 ( .A(n15433), .B(n15415), .Z(n15435) );
  XOR U14943 ( .A(n15455), .B(n15456), .Z(n15415) );
  AND U14944 ( .A(n918), .B(n15457), .Z(n15455) );
  XOR U14945 ( .A(n15458), .B(n15456), .Z(n15457) );
  NANDN U14946 ( .A(n15417), .B(n15419), .Z(n15433) );
  XOR U14947 ( .A(n15459), .B(n15460), .Z(n15419) );
  AND U14948 ( .A(n918), .B(n15461), .Z(n15459) );
  XOR U14949 ( .A(n15460), .B(n15462), .Z(n15461) );
  XOR U14950 ( .A(n15463), .B(n15464), .Z(n918) );
  AND U14951 ( .A(n15465), .B(n15466), .Z(n15463) );
  XNOR U14952 ( .A(n15464), .B(n15430), .Z(n15466) );
  XNOR U14953 ( .A(n15467), .B(n15468), .Z(n15430) );
  ANDN U14954 ( .B(n15469), .A(n15470), .Z(n15467) );
  XOR U14955 ( .A(n15468), .B(n15471), .Z(n15469) );
  XOR U14956 ( .A(n15464), .B(n15432), .Z(n15465) );
  XOR U14957 ( .A(n15472), .B(n15473), .Z(n15432) );
  AND U14958 ( .A(n922), .B(n15474), .Z(n15472) );
  XOR U14959 ( .A(n15475), .B(n15473), .Z(n15474) );
  XNOR U14960 ( .A(n15476), .B(n15477), .Z(n15464) );
  NAND U14961 ( .A(n15478), .B(n15479), .Z(n15477) );
  XOR U14962 ( .A(n15480), .B(n15456), .Z(n15479) );
  XOR U14963 ( .A(n15470), .B(n15471), .Z(n15456) );
  XOR U14964 ( .A(n15481), .B(n15482), .Z(n15471) );
  ANDN U14965 ( .B(n15483), .A(n15484), .Z(n15481) );
  XOR U14966 ( .A(n15482), .B(n15485), .Z(n15483) );
  XOR U14967 ( .A(n15486), .B(n15487), .Z(n15470) );
  XOR U14968 ( .A(n15488), .B(n15489), .Z(n15487) );
  ANDN U14969 ( .B(n15490), .A(n15491), .Z(n15488) );
  XOR U14970 ( .A(n15492), .B(n15489), .Z(n15490) );
  IV U14971 ( .A(n15468), .Z(n15486) );
  XOR U14972 ( .A(n15493), .B(n15494), .Z(n15468) );
  ANDN U14973 ( .B(n15495), .A(n15496), .Z(n15493) );
  XOR U14974 ( .A(n15494), .B(n15497), .Z(n15495) );
  IV U14975 ( .A(n15476), .Z(n15480) );
  XOR U14976 ( .A(n15476), .B(n15458), .Z(n15478) );
  XOR U14977 ( .A(n15498), .B(n15499), .Z(n15458) );
  AND U14978 ( .A(n922), .B(n15500), .Z(n15498) );
  XOR U14979 ( .A(n15501), .B(n15499), .Z(n15500) );
  NANDN U14980 ( .A(n15460), .B(n15462), .Z(n15476) );
  XOR U14981 ( .A(n15502), .B(n15503), .Z(n15462) );
  AND U14982 ( .A(n922), .B(n15504), .Z(n15502) );
  XOR U14983 ( .A(n15503), .B(n15505), .Z(n15504) );
  XOR U14984 ( .A(n15506), .B(n15507), .Z(n922) );
  AND U14985 ( .A(n15508), .B(n15509), .Z(n15506) );
  XNOR U14986 ( .A(n15507), .B(n15473), .Z(n15509) );
  XNOR U14987 ( .A(n15510), .B(n15511), .Z(n15473) );
  ANDN U14988 ( .B(n15512), .A(n15513), .Z(n15510) );
  XOR U14989 ( .A(n15511), .B(n15514), .Z(n15512) );
  XOR U14990 ( .A(n15507), .B(n15475), .Z(n15508) );
  XOR U14991 ( .A(n15515), .B(n15516), .Z(n15475) );
  AND U14992 ( .A(n926), .B(n15517), .Z(n15515) );
  XOR U14993 ( .A(n15518), .B(n15516), .Z(n15517) );
  XNOR U14994 ( .A(n15519), .B(n15520), .Z(n15507) );
  NAND U14995 ( .A(n15521), .B(n15522), .Z(n15520) );
  XOR U14996 ( .A(n15523), .B(n15499), .Z(n15522) );
  XOR U14997 ( .A(n15513), .B(n15514), .Z(n15499) );
  XOR U14998 ( .A(n15524), .B(n15525), .Z(n15514) );
  ANDN U14999 ( .B(n15526), .A(n15527), .Z(n15524) );
  XOR U15000 ( .A(n15525), .B(n15528), .Z(n15526) );
  XOR U15001 ( .A(n15529), .B(n15530), .Z(n15513) );
  XOR U15002 ( .A(n15531), .B(n15532), .Z(n15530) );
  ANDN U15003 ( .B(n15533), .A(n15534), .Z(n15531) );
  XOR U15004 ( .A(n15535), .B(n15532), .Z(n15533) );
  IV U15005 ( .A(n15511), .Z(n15529) );
  XOR U15006 ( .A(n15536), .B(n15537), .Z(n15511) );
  ANDN U15007 ( .B(n15538), .A(n15539), .Z(n15536) );
  XOR U15008 ( .A(n15537), .B(n15540), .Z(n15538) );
  IV U15009 ( .A(n15519), .Z(n15523) );
  XOR U15010 ( .A(n15519), .B(n15501), .Z(n15521) );
  XOR U15011 ( .A(n15541), .B(n15542), .Z(n15501) );
  AND U15012 ( .A(n926), .B(n15543), .Z(n15541) );
  XOR U15013 ( .A(n15544), .B(n15542), .Z(n15543) );
  NANDN U15014 ( .A(n15503), .B(n15505), .Z(n15519) );
  XOR U15015 ( .A(n15545), .B(n15546), .Z(n15505) );
  AND U15016 ( .A(n926), .B(n15547), .Z(n15545) );
  XOR U15017 ( .A(n15546), .B(n15548), .Z(n15547) );
  XOR U15018 ( .A(n15549), .B(n15550), .Z(n926) );
  AND U15019 ( .A(n15551), .B(n15552), .Z(n15549) );
  XNOR U15020 ( .A(n15550), .B(n15516), .Z(n15552) );
  XNOR U15021 ( .A(n15553), .B(n15554), .Z(n15516) );
  ANDN U15022 ( .B(n15555), .A(n15556), .Z(n15553) );
  XOR U15023 ( .A(n15554), .B(n15557), .Z(n15555) );
  XOR U15024 ( .A(n15550), .B(n15518), .Z(n15551) );
  XOR U15025 ( .A(n15558), .B(n15559), .Z(n15518) );
  AND U15026 ( .A(n930), .B(n15560), .Z(n15558) );
  XOR U15027 ( .A(n15561), .B(n15559), .Z(n15560) );
  XNOR U15028 ( .A(n15562), .B(n15563), .Z(n15550) );
  NAND U15029 ( .A(n15564), .B(n15565), .Z(n15563) );
  XOR U15030 ( .A(n15566), .B(n15542), .Z(n15565) );
  XOR U15031 ( .A(n15556), .B(n15557), .Z(n15542) );
  XOR U15032 ( .A(n15567), .B(n15568), .Z(n15557) );
  ANDN U15033 ( .B(n15569), .A(n15570), .Z(n15567) );
  XOR U15034 ( .A(n15568), .B(n15571), .Z(n15569) );
  XOR U15035 ( .A(n15572), .B(n15573), .Z(n15556) );
  XOR U15036 ( .A(n15574), .B(n15575), .Z(n15573) );
  ANDN U15037 ( .B(n15576), .A(n15577), .Z(n15574) );
  XOR U15038 ( .A(n15578), .B(n15575), .Z(n15576) );
  IV U15039 ( .A(n15554), .Z(n15572) );
  XOR U15040 ( .A(n15579), .B(n15580), .Z(n15554) );
  ANDN U15041 ( .B(n15581), .A(n15582), .Z(n15579) );
  XOR U15042 ( .A(n15580), .B(n15583), .Z(n15581) );
  IV U15043 ( .A(n15562), .Z(n15566) );
  XOR U15044 ( .A(n15562), .B(n15544), .Z(n15564) );
  XOR U15045 ( .A(n15584), .B(n15585), .Z(n15544) );
  AND U15046 ( .A(n930), .B(n15586), .Z(n15584) );
  XOR U15047 ( .A(n15587), .B(n15585), .Z(n15586) );
  NANDN U15048 ( .A(n15546), .B(n15548), .Z(n15562) );
  XOR U15049 ( .A(n15588), .B(n15589), .Z(n15548) );
  AND U15050 ( .A(n930), .B(n15590), .Z(n15588) );
  XOR U15051 ( .A(n15589), .B(n15591), .Z(n15590) );
  XOR U15052 ( .A(n15592), .B(n15593), .Z(n930) );
  AND U15053 ( .A(n15594), .B(n15595), .Z(n15592) );
  XNOR U15054 ( .A(n15593), .B(n15559), .Z(n15595) );
  XNOR U15055 ( .A(n15596), .B(n15597), .Z(n15559) );
  ANDN U15056 ( .B(n15598), .A(n15599), .Z(n15596) );
  XOR U15057 ( .A(n15597), .B(n15600), .Z(n15598) );
  XOR U15058 ( .A(n15593), .B(n15561), .Z(n15594) );
  XOR U15059 ( .A(n15601), .B(n15602), .Z(n15561) );
  AND U15060 ( .A(n934), .B(n15603), .Z(n15601) );
  XOR U15061 ( .A(n15604), .B(n15602), .Z(n15603) );
  XNOR U15062 ( .A(n15605), .B(n15606), .Z(n15593) );
  NAND U15063 ( .A(n15607), .B(n15608), .Z(n15606) );
  XOR U15064 ( .A(n15609), .B(n15585), .Z(n15608) );
  XOR U15065 ( .A(n15599), .B(n15600), .Z(n15585) );
  XOR U15066 ( .A(n15610), .B(n15611), .Z(n15600) );
  ANDN U15067 ( .B(n15612), .A(n15613), .Z(n15610) );
  XOR U15068 ( .A(n15611), .B(n15614), .Z(n15612) );
  XOR U15069 ( .A(n15615), .B(n15616), .Z(n15599) );
  XOR U15070 ( .A(n15617), .B(n15618), .Z(n15616) );
  ANDN U15071 ( .B(n15619), .A(n15620), .Z(n15617) );
  XOR U15072 ( .A(n15621), .B(n15618), .Z(n15619) );
  IV U15073 ( .A(n15597), .Z(n15615) );
  XOR U15074 ( .A(n15622), .B(n15623), .Z(n15597) );
  ANDN U15075 ( .B(n15624), .A(n15625), .Z(n15622) );
  XOR U15076 ( .A(n15623), .B(n15626), .Z(n15624) );
  IV U15077 ( .A(n15605), .Z(n15609) );
  XOR U15078 ( .A(n15605), .B(n15587), .Z(n15607) );
  XOR U15079 ( .A(n15627), .B(n15628), .Z(n15587) );
  AND U15080 ( .A(n934), .B(n15629), .Z(n15627) );
  XOR U15081 ( .A(n15630), .B(n15628), .Z(n15629) );
  NANDN U15082 ( .A(n15589), .B(n15591), .Z(n15605) );
  XOR U15083 ( .A(n15631), .B(n15632), .Z(n15591) );
  AND U15084 ( .A(n934), .B(n15633), .Z(n15631) );
  XOR U15085 ( .A(n15632), .B(n15634), .Z(n15633) );
  XOR U15086 ( .A(n15635), .B(n15636), .Z(n934) );
  AND U15087 ( .A(n15637), .B(n15638), .Z(n15635) );
  XNOR U15088 ( .A(n15636), .B(n15602), .Z(n15638) );
  XNOR U15089 ( .A(n15639), .B(n15640), .Z(n15602) );
  ANDN U15090 ( .B(n15641), .A(n15642), .Z(n15639) );
  XOR U15091 ( .A(n15640), .B(n15643), .Z(n15641) );
  XOR U15092 ( .A(n15636), .B(n15604), .Z(n15637) );
  XOR U15093 ( .A(n15644), .B(n15645), .Z(n15604) );
  AND U15094 ( .A(n938), .B(n15646), .Z(n15644) );
  XOR U15095 ( .A(n15647), .B(n15645), .Z(n15646) );
  XNOR U15096 ( .A(n15648), .B(n15649), .Z(n15636) );
  NAND U15097 ( .A(n15650), .B(n15651), .Z(n15649) );
  XOR U15098 ( .A(n15652), .B(n15628), .Z(n15651) );
  XOR U15099 ( .A(n15642), .B(n15643), .Z(n15628) );
  XOR U15100 ( .A(n15653), .B(n15654), .Z(n15643) );
  ANDN U15101 ( .B(n15655), .A(n15656), .Z(n15653) );
  XOR U15102 ( .A(n15654), .B(n15657), .Z(n15655) );
  XOR U15103 ( .A(n15658), .B(n15659), .Z(n15642) );
  XOR U15104 ( .A(n15660), .B(n15661), .Z(n15659) );
  ANDN U15105 ( .B(n15662), .A(n15663), .Z(n15660) );
  XOR U15106 ( .A(n15664), .B(n15661), .Z(n15662) );
  IV U15107 ( .A(n15640), .Z(n15658) );
  XOR U15108 ( .A(n15665), .B(n15666), .Z(n15640) );
  ANDN U15109 ( .B(n15667), .A(n15668), .Z(n15665) );
  XOR U15110 ( .A(n15666), .B(n15669), .Z(n15667) );
  IV U15111 ( .A(n15648), .Z(n15652) );
  XOR U15112 ( .A(n15648), .B(n15630), .Z(n15650) );
  XOR U15113 ( .A(n15670), .B(n15671), .Z(n15630) );
  AND U15114 ( .A(n938), .B(n15672), .Z(n15670) );
  XOR U15115 ( .A(n15673), .B(n15671), .Z(n15672) );
  NANDN U15116 ( .A(n15632), .B(n15634), .Z(n15648) );
  XOR U15117 ( .A(n15674), .B(n15675), .Z(n15634) );
  AND U15118 ( .A(n938), .B(n15676), .Z(n15674) );
  XOR U15119 ( .A(n15675), .B(n15677), .Z(n15676) );
  XOR U15120 ( .A(n15678), .B(n15679), .Z(n938) );
  AND U15121 ( .A(n15680), .B(n15681), .Z(n15678) );
  XNOR U15122 ( .A(n15679), .B(n15645), .Z(n15681) );
  XNOR U15123 ( .A(n15682), .B(n15683), .Z(n15645) );
  ANDN U15124 ( .B(n15684), .A(n15685), .Z(n15682) );
  XOR U15125 ( .A(n15683), .B(n15686), .Z(n15684) );
  XOR U15126 ( .A(n15679), .B(n15647), .Z(n15680) );
  XOR U15127 ( .A(n15687), .B(n15688), .Z(n15647) );
  AND U15128 ( .A(n942), .B(n15689), .Z(n15687) );
  XOR U15129 ( .A(n15690), .B(n15688), .Z(n15689) );
  XNOR U15130 ( .A(n15691), .B(n15692), .Z(n15679) );
  NAND U15131 ( .A(n15693), .B(n15694), .Z(n15692) );
  XOR U15132 ( .A(n15695), .B(n15671), .Z(n15694) );
  XOR U15133 ( .A(n15685), .B(n15686), .Z(n15671) );
  XOR U15134 ( .A(n15696), .B(n15697), .Z(n15686) );
  ANDN U15135 ( .B(n15698), .A(n15699), .Z(n15696) );
  XOR U15136 ( .A(n15697), .B(n15700), .Z(n15698) );
  XOR U15137 ( .A(n15701), .B(n15702), .Z(n15685) );
  XOR U15138 ( .A(n15703), .B(n15704), .Z(n15702) );
  ANDN U15139 ( .B(n15705), .A(n15706), .Z(n15703) );
  XOR U15140 ( .A(n15707), .B(n15704), .Z(n15705) );
  IV U15141 ( .A(n15683), .Z(n15701) );
  XOR U15142 ( .A(n15708), .B(n15709), .Z(n15683) );
  ANDN U15143 ( .B(n15710), .A(n15711), .Z(n15708) );
  XOR U15144 ( .A(n15709), .B(n15712), .Z(n15710) );
  IV U15145 ( .A(n15691), .Z(n15695) );
  XOR U15146 ( .A(n15691), .B(n15673), .Z(n15693) );
  XOR U15147 ( .A(n15713), .B(n15714), .Z(n15673) );
  AND U15148 ( .A(n942), .B(n15715), .Z(n15713) );
  XOR U15149 ( .A(n15716), .B(n15714), .Z(n15715) );
  NANDN U15150 ( .A(n15675), .B(n15677), .Z(n15691) );
  XOR U15151 ( .A(n15717), .B(n15718), .Z(n15677) );
  AND U15152 ( .A(n942), .B(n15719), .Z(n15717) );
  XOR U15153 ( .A(n15718), .B(n15720), .Z(n15719) );
  XOR U15154 ( .A(n15721), .B(n15722), .Z(n942) );
  AND U15155 ( .A(n15723), .B(n15724), .Z(n15721) );
  XNOR U15156 ( .A(n15722), .B(n15688), .Z(n15724) );
  XNOR U15157 ( .A(n15725), .B(n15726), .Z(n15688) );
  ANDN U15158 ( .B(n15727), .A(n15728), .Z(n15725) );
  XOR U15159 ( .A(n15726), .B(n15729), .Z(n15727) );
  XOR U15160 ( .A(n15722), .B(n15690), .Z(n15723) );
  XOR U15161 ( .A(n15730), .B(n15731), .Z(n15690) );
  AND U15162 ( .A(n946), .B(n15732), .Z(n15730) );
  XOR U15163 ( .A(n15733), .B(n15731), .Z(n15732) );
  XNOR U15164 ( .A(n15734), .B(n15735), .Z(n15722) );
  NAND U15165 ( .A(n15736), .B(n15737), .Z(n15735) );
  XOR U15166 ( .A(n15738), .B(n15714), .Z(n15737) );
  XOR U15167 ( .A(n15728), .B(n15729), .Z(n15714) );
  XOR U15168 ( .A(n15739), .B(n15740), .Z(n15729) );
  ANDN U15169 ( .B(n15741), .A(n15742), .Z(n15739) );
  XOR U15170 ( .A(n15740), .B(n15743), .Z(n15741) );
  XOR U15171 ( .A(n15744), .B(n15745), .Z(n15728) );
  XOR U15172 ( .A(n15746), .B(n15747), .Z(n15745) );
  ANDN U15173 ( .B(n15748), .A(n15749), .Z(n15746) );
  XOR U15174 ( .A(n15750), .B(n15747), .Z(n15748) );
  IV U15175 ( .A(n15726), .Z(n15744) );
  XOR U15176 ( .A(n15751), .B(n15752), .Z(n15726) );
  ANDN U15177 ( .B(n15753), .A(n15754), .Z(n15751) );
  XOR U15178 ( .A(n15752), .B(n15755), .Z(n15753) );
  IV U15179 ( .A(n15734), .Z(n15738) );
  XOR U15180 ( .A(n15734), .B(n15716), .Z(n15736) );
  XOR U15181 ( .A(n15756), .B(n15757), .Z(n15716) );
  AND U15182 ( .A(n946), .B(n15758), .Z(n15756) );
  XOR U15183 ( .A(n15759), .B(n15757), .Z(n15758) );
  NANDN U15184 ( .A(n15718), .B(n15720), .Z(n15734) );
  XOR U15185 ( .A(n15760), .B(n15761), .Z(n15720) );
  AND U15186 ( .A(n946), .B(n15762), .Z(n15760) );
  XOR U15187 ( .A(n15761), .B(n15763), .Z(n15762) );
  XOR U15188 ( .A(n15764), .B(n15765), .Z(n946) );
  AND U15189 ( .A(n15766), .B(n15767), .Z(n15764) );
  XNOR U15190 ( .A(n15765), .B(n15731), .Z(n15767) );
  XNOR U15191 ( .A(n15768), .B(n15769), .Z(n15731) );
  ANDN U15192 ( .B(n15770), .A(n15771), .Z(n15768) );
  XOR U15193 ( .A(n15769), .B(n15772), .Z(n15770) );
  XOR U15194 ( .A(n15765), .B(n15733), .Z(n15766) );
  XOR U15195 ( .A(n15773), .B(n15774), .Z(n15733) );
  AND U15196 ( .A(n950), .B(n15775), .Z(n15773) );
  XOR U15197 ( .A(n15776), .B(n15774), .Z(n15775) );
  XNOR U15198 ( .A(n15777), .B(n15778), .Z(n15765) );
  NAND U15199 ( .A(n15779), .B(n15780), .Z(n15778) );
  XOR U15200 ( .A(n15781), .B(n15757), .Z(n15780) );
  XOR U15201 ( .A(n15771), .B(n15772), .Z(n15757) );
  XOR U15202 ( .A(n15782), .B(n15783), .Z(n15772) );
  ANDN U15203 ( .B(n15784), .A(n15785), .Z(n15782) );
  XOR U15204 ( .A(n15783), .B(n15786), .Z(n15784) );
  XOR U15205 ( .A(n15787), .B(n15788), .Z(n15771) );
  XOR U15206 ( .A(n15789), .B(n15790), .Z(n15788) );
  ANDN U15207 ( .B(n15791), .A(n15792), .Z(n15789) );
  XOR U15208 ( .A(n15793), .B(n15790), .Z(n15791) );
  IV U15209 ( .A(n15769), .Z(n15787) );
  XOR U15210 ( .A(n15794), .B(n15795), .Z(n15769) );
  ANDN U15211 ( .B(n15796), .A(n15797), .Z(n15794) );
  XOR U15212 ( .A(n15795), .B(n15798), .Z(n15796) );
  IV U15213 ( .A(n15777), .Z(n15781) );
  XOR U15214 ( .A(n15777), .B(n15759), .Z(n15779) );
  XOR U15215 ( .A(n15799), .B(n15800), .Z(n15759) );
  AND U15216 ( .A(n950), .B(n15801), .Z(n15799) );
  XOR U15217 ( .A(n15802), .B(n15800), .Z(n15801) );
  NANDN U15218 ( .A(n15761), .B(n15763), .Z(n15777) );
  XOR U15219 ( .A(n15803), .B(n15804), .Z(n15763) );
  AND U15220 ( .A(n950), .B(n15805), .Z(n15803) );
  XOR U15221 ( .A(n15804), .B(n15806), .Z(n15805) );
  XOR U15222 ( .A(n15807), .B(n15808), .Z(n950) );
  AND U15223 ( .A(n15809), .B(n15810), .Z(n15807) );
  XNOR U15224 ( .A(n15808), .B(n15774), .Z(n15810) );
  XNOR U15225 ( .A(n15811), .B(n15812), .Z(n15774) );
  ANDN U15226 ( .B(n15813), .A(n15814), .Z(n15811) );
  XOR U15227 ( .A(n15812), .B(n15815), .Z(n15813) );
  XOR U15228 ( .A(n15808), .B(n15776), .Z(n15809) );
  XOR U15229 ( .A(n15816), .B(n15817), .Z(n15776) );
  AND U15230 ( .A(n954), .B(n15818), .Z(n15816) );
  XOR U15231 ( .A(n15819), .B(n15817), .Z(n15818) );
  XNOR U15232 ( .A(n15820), .B(n15821), .Z(n15808) );
  NAND U15233 ( .A(n15822), .B(n15823), .Z(n15821) );
  XOR U15234 ( .A(n15824), .B(n15800), .Z(n15823) );
  XOR U15235 ( .A(n15814), .B(n15815), .Z(n15800) );
  XOR U15236 ( .A(n15825), .B(n15826), .Z(n15815) );
  ANDN U15237 ( .B(n15827), .A(n15828), .Z(n15825) );
  XOR U15238 ( .A(n15826), .B(n15829), .Z(n15827) );
  XOR U15239 ( .A(n15830), .B(n15831), .Z(n15814) );
  XOR U15240 ( .A(n15832), .B(n15833), .Z(n15831) );
  ANDN U15241 ( .B(n15834), .A(n15835), .Z(n15832) );
  XOR U15242 ( .A(n15836), .B(n15833), .Z(n15834) );
  IV U15243 ( .A(n15812), .Z(n15830) );
  XOR U15244 ( .A(n15837), .B(n15838), .Z(n15812) );
  ANDN U15245 ( .B(n15839), .A(n15840), .Z(n15837) );
  XOR U15246 ( .A(n15838), .B(n15841), .Z(n15839) );
  IV U15247 ( .A(n15820), .Z(n15824) );
  XOR U15248 ( .A(n15820), .B(n15802), .Z(n15822) );
  XOR U15249 ( .A(n15842), .B(n15843), .Z(n15802) );
  AND U15250 ( .A(n954), .B(n15844), .Z(n15842) );
  XOR U15251 ( .A(n15845), .B(n15843), .Z(n15844) );
  NANDN U15252 ( .A(n15804), .B(n15806), .Z(n15820) );
  XOR U15253 ( .A(n15846), .B(n15847), .Z(n15806) );
  AND U15254 ( .A(n954), .B(n15848), .Z(n15846) );
  XOR U15255 ( .A(n15847), .B(n15849), .Z(n15848) );
  XOR U15256 ( .A(n15850), .B(n15851), .Z(n954) );
  AND U15257 ( .A(n15852), .B(n15853), .Z(n15850) );
  XNOR U15258 ( .A(n15851), .B(n15817), .Z(n15853) );
  XNOR U15259 ( .A(n15854), .B(n15855), .Z(n15817) );
  ANDN U15260 ( .B(n15856), .A(n15857), .Z(n15854) );
  XOR U15261 ( .A(n15855), .B(n15858), .Z(n15856) );
  XOR U15262 ( .A(n15851), .B(n15819), .Z(n15852) );
  XOR U15263 ( .A(n15859), .B(n15860), .Z(n15819) );
  AND U15264 ( .A(n958), .B(n15861), .Z(n15859) );
  XOR U15265 ( .A(n15862), .B(n15860), .Z(n15861) );
  XNOR U15266 ( .A(n15863), .B(n15864), .Z(n15851) );
  NAND U15267 ( .A(n15865), .B(n15866), .Z(n15864) );
  XOR U15268 ( .A(n15867), .B(n15843), .Z(n15866) );
  XOR U15269 ( .A(n15857), .B(n15858), .Z(n15843) );
  XOR U15270 ( .A(n15868), .B(n15869), .Z(n15858) );
  ANDN U15271 ( .B(n15870), .A(n15871), .Z(n15868) );
  XOR U15272 ( .A(n15869), .B(n15872), .Z(n15870) );
  XOR U15273 ( .A(n15873), .B(n15874), .Z(n15857) );
  XOR U15274 ( .A(n15875), .B(n15876), .Z(n15874) );
  ANDN U15275 ( .B(n15877), .A(n15878), .Z(n15875) );
  XOR U15276 ( .A(n15879), .B(n15876), .Z(n15877) );
  IV U15277 ( .A(n15855), .Z(n15873) );
  XOR U15278 ( .A(n15880), .B(n15881), .Z(n15855) );
  ANDN U15279 ( .B(n15882), .A(n15883), .Z(n15880) );
  XOR U15280 ( .A(n15881), .B(n15884), .Z(n15882) );
  IV U15281 ( .A(n15863), .Z(n15867) );
  XOR U15282 ( .A(n15863), .B(n15845), .Z(n15865) );
  XOR U15283 ( .A(n15885), .B(n15886), .Z(n15845) );
  AND U15284 ( .A(n958), .B(n15887), .Z(n15885) );
  XOR U15285 ( .A(n15888), .B(n15886), .Z(n15887) );
  NANDN U15286 ( .A(n15847), .B(n15849), .Z(n15863) );
  XOR U15287 ( .A(n15889), .B(n15890), .Z(n15849) );
  AND U15288 ( .A(n958), .B(n15891), .Z(n15889) );
  XOR U15289 ( .A(n15890), .B(n15892), .Z(n15891) );
  XOR U15290 ( .A(n15893), .B(n15894), .Z(n958) );
  AND U15291 ( .A(n15895), .B(n15896), .Z(n15893) );
  XNOR U15292 ( .A(n15894), .B(n15860), .Z(n15896) );
  XNOR U15293 ( .A(n15897), .B(n15898), .Z(n15860) );
  ANDN U15294 ( .B(n15899), .A(n15900), .Z(n15897) );
  XOR U15295 ( .A(n15898), .B(n15901), .Z(n15899) );
  XOR U15296 ( .A(n15894), .B(n15862), .Z(n15895) );
  XOR U15297 ( .A(n15902), .B(n15903), .Z(n15862) );
  AND U15298 ( .A(n962), .B(n15904), .Z(n15902) );
  XOR U15299 ( .A(n15905), .B(n15903), .Z(n15904) );
  XNOR U15300 ( .A(n15906), .B(n15907), .Z(n15894) );
  NAND U15301 ( .A(n15908), .B(n15909), .Z(n15907) );
  XOR U15302 ( .A(n15910), .B(n15886), .Z(n15909) );
  XOR U15303 ( .A(n15900), .B(n15901), .Z(n15886) );
  XOR U15304 ( .A(n15911), .B(n15912), .Z(n15901) );
  ANDN U15305 ( .B(n15913), .A(n15914), .Z(n15911) );
  XOR U15306 ( .A(n15912), .B(n15915), .Z(n15913) );
  XOR U15307 ( .A(n15916), .B(n15917), .Z(n15900) );
  XOR U15308 ( .A(n15918), .B(n15919), .Z(n15917) );
  ANDN U15309 ( .B(n15920), .A(n15921), .Z(n15918) );
  XOR U15310 ( .A(n15922), .B(n15919), .Z(n15920) );
  IV U15311 ( .A(n15898), .Z(n15916) );
  XOR U15312 ( .A(n15923), .B(n15924), .Z(n15898) );
  ANDN U15313 ( .B(n15925), .A(n15926), .Z(n15923) );
  XOR U15314 ( .A(n15924), .B(n15927), .Z(n15925) );
  IV U15315 ( .A(n15906), .Z(n15910) );
  XOR U15316 ( .A(n15906), .B(n15888), .Z(n15908) );
  XOR U15317 ( .A(n15928), .B(n15929), .Z(n15888) );
  AND U15318 ( .A(n962), .B(n15930), .Z(n15928) );
  XOR U15319 ( .A(n15931), .B(n15929), .Z(n15930) );
  NANDN U15320 ( .A(n15890), .B(n15892), .Z(n15906) );
  XOR U15321 ( .A(n15932), .B(n15933), .Z(n15892) );
  AND U15322 ( .A(n962), .B(n15934), .Z(n15932) );
  XOR U15323 ( .A(n15933), .B(n15935), .Z(n15934) );
  XOR U15324 ( .A(n15936), .B(n15937), .Z(n962) );
  AND U15325 ( .A(n15938), .B(n15939), .Z(n15936) );
  XNOR U15326 ( .A(n15937), .B(n15903), .Z(n15939) );
  XNOR U15327 ( .A(n15940), .B(n15941), .Z(n15903) );
  ANDN U15328 ( .B(n15942), .A(n15943), .Z(n15940) );
  XOR U15329 ( .A(n15941), .B(n15944), .Z(n15942) );
  XOR U15330 ( .A(n15937), .B(n15905), .Z(n15938) );
  XOR U15331 ( .A(n15945), .B(n15946), .Z(n15905) );
  AND U15332 ( .A(n966), .B(n15947), .Z(n15945) );
  XOR U15333 ( .A(n15948), .B(n15946), .Z(n15947) );
  XNOR U15334 ( .A(n15949), .B(n15950), .Z(n15937) );
  NAND U15335 ( .A(n15951), .B(n15952), .Z(n15950) );
  XOR U15336 ( .A(n15953), .B(n15929), .Z(n15952) );
  XOR U15337 ( .A(n15943), .B(n15944), .Z(n15929) );
  XOR U15338 ( .A(n15954), .B(n15955), .Z(n15944) );
  ANDN U15339 ( .B(n15956), .A(n15957), .Z(n15954) );
  XOR U15340 ( .A(n15955), .B(n15958), .Z(n15956) );
  XOR U15341 ( .A(n15959), .B(n15960), .Z(n15943) );
  XOR U15342 ( .A(n15961), .B(n15962), .Z(n15960) );
  ANDN U15343 ( .B(n15963), .A(n15964), .Z(n15961) );
  XOR U15344 ( .A(n15965), .B(n15962), .Z(n15963) );
  IV U15345 ( .A(n15941), .Z(n15959) );
  XOR U15346 ( .A(n15966), .B(n15967), .Z(n15941) );
  ANDN U15347 ( .B(n15968), .A(n15969), .Z(n15966) );
  XOR U15348 ( .A(n15967), .B(n15970), .Z(n15968) );
  IV U15349 ( .A(n15949), .Z(n15953) );
  XOR U15350 ( .A(n15949), .B(n15931), .Z(n15951) );
  XOR U15351 ( .A(n15971), .B(n15972), .Z(n15931) );
  AND U15352 ( .A(n966), .B(n15973), .Z(n15971) );
  XOR U15353 ( .A(n15974), .B(n15972), .Z(n15973) );
  NANDN U15354 ( .A(n15933), .B(n15935), .Z(n15949) );
  XOR U15355 ( .A(n15975), .B(n15976), .Z(n15935) );
  AND U15356 ( .A(n966), .B(n15977), .Z(n15975) );
  XOR U15357 ( .A(n15976), .B(n15978), .Z(n15977) );
  XOR U15358 ( .A(n15979), .B(n15980), .Z(n966) );
  AND U15359 ( .A(n15981), .B(n15982), .Z(n15979) );
  XNOR U15360 ( .A(n15980), .B(n15946), .Z(n15982) );
  XNOR U15361 ( .A(n15983), .B(n15984), .Z(n15946) );
  ANDN U15362 ( .B(n15985), .A(n15986), .Z(n15983) );
  XOR U15363 ( .A(n15984), .B(n15987), .Z(n15985) );
  XOR U15364 ( .A(n15980), .B(n15948), .Z(n15981) );
  XOR U15365 ( .A(n15988), .B(n15989), .Z(n15948) );
  AND U15366 ( .A(n970), .B(n15990), .Z(n15988) );
  XOR U15367 ( .A(n15991), .B(n15989), .Z(n15990) );
  XNOR U15368 ( .A(n15992), .B(n15993), .Z(n15980) );
  NAND U15369 ( .A(n15994), .B(n15995), .Z(n15993) );
  XOR U15370 ( .A(n15996), .B(n15972), .Z(n15995) );
  XOR U15371 ( .A(n15986), .B(n15987), .Z(n15972) );
  XOR U15372 ( .A(n15997), .B(n15998), .Z(n15987) );
  ANDN U15373 ( .B(n15999), .A(n16000), .Z(n15997) );
  XOR U15374 ( .A(n15998), .B(n16001), .Z(n15999) );
  XOR U15375 ( .A(n16002), .B(n16003), .Z(n15986) );
  XOR U15376 ( .A(n16004), .B(n16005), .Z(n16003) );
  ANDN U15377 ( .B(n16006), .A(n16007), .Z(n16004) );
  XOR U15378 ( .A(n16008), .B(n16005), .Z(n16006) );
  IV U15379 ( .A(n15984), .Z(n16002) );
  XOR U15380 ( .A(n16009), .B(n16010), .Z(n15984) );
  ANDN U15381 ( .B(n16011), .A(n16012), .Z(n16009) );
  XOR U15382 ( .A(n16010), .B(n16013), .Z(n16011) );
  IV U15383 ( .A(n15992), .Z(n15996) );
  XOR U15384 ( .A(n15992), .B(n15974), .Z(n15994) );
  XOR U15385 ( .A(n16014), .B(n16015), .Z(n15974) );
  AND U15386 ( .A(n970), .B(n16016), .Z(n16014) );
  XOR U15387 ( .A(n16017), .B(n16015), .Z(n16016) );
  NANDN U15388 ( .A(n15976), .B(n15978), .Z(n15992) );
  XOR U15389 ( .A(n16018), .B(n16019), .Z(n15978) );
  AND U15390 ( .A(n970), .B(n16020), .Z(n16018) );
  XOR U15391 ( .A(n16019), .B(n16021), .Z(n16020) );
  XOR U15392 ( .A(n16022), .B(n16023), .Z(n970) );
  AND U15393 ( .A(n16024), .B(n16025), .Z(n16022) );
  XNOR U15394 ( .A(n16023), .B(n15989), .Z(n16025) );
  XNOR U15395 ( .A(n16026), .B(n16027), .Z(n15989) );
  ANDN U15396 ( .B(n16028), .A(n16029), .Z(n16026) );
  XOR U15397 ( .A(n16027), .B(n16030), .Z(n16028) );
  XOR U15398 ( .A(n16023), .B(n15991), .Z(n16024) );
  XOR U15399 ( .A(n16031), .B(n16032), .Z(n15991) );
  AND U15400 ( .A(n974), .B(n16033), .Z(n16031) );
  XOR U15401 ( .A(n16034), .B(n16032), .Z(n16033) );
  XNOR U15402 ( .A(n16035), .B(n16036), .Z(n16023) );
  NAND U15403 ( .A(n16037), .B(n16038), .Z(n16036) );
  XOR U15404 ( .A(n16039), .B(n16015), .Z(n16038) );
  XOR U15405 ( .A(n16029), .B(n16030), .Z(n16015) );
  XOR U15406 ( .A(n16040), .B(n16041), .Z(n16030) );
  ANDN U15407 ( .B(n16042), .A(n16043), .Z(n16040) );
  XOR U15408 ( .A(n16041), .B(n16044), .Z(n16042) );
  XOR U15409 ( .A(n16045), .B(n16046), .Z(n16029) );
  XOR U15410 ( .A(n16047), .B(n16048), .Z(n16046) );
  ANDN U15411 ( .B(n16049), .A(n16050), .Z(n16047) );
  XOR U15412 ( .A(n16051), .B(n16048), .Z(n16049) );
  IV U15413 ( .A(n16027), .Z(n16045) );
  XOR U15414 ( .A(n16052), .B(n16053), .Z(n16027) );
  ANDN U15415 ( .B(n16054), .A(n16055), .Z(n16052) );
  XOR U15416 ( .A(n16053), .B(n16056), .Z(n16054) );
  IV U15417 ( .A(n16035), .Z(n16039) );
  XOR U15418 ( .A(n16035), .B(n16017), .Z(n16037) );
  XOR U15419 ( .A(n16057), .B(n16058), .Z(n16017) );
  AND U15420 ( .A(n974), .B(n16059), .Z(n16057) );
  XOR U15421 ( .A(n16060), .B(n16058), .Z(n16059) );
  NANDN U15422 ( .A(n16019), .B(n16021), .Z(n16035) );
  XOR U15423 ( .A(n16061), .B(n16062), .Z(n16021) );
  AND U15424 ( .A(n974), .B(n16063), .Z(n16061) );
  XOR U15425 ( .A(n16062), .B(n16064), .Z(n16063) );
  XOR U15426 ( .A(n16065), .B(n16066), .Z(n974) );
  AND U15427 ( .A(n16067), .B(n16068), .Z(n16065) );
  XNOR U15428 ( .A(n16066), .B(n16032), .Z(n16068) );
  XNOR U15429 ( .A(n16069), .B(n16070), .Z(n16032) );
  ANDN U15430 ( .B(n16071), .A(n16072), .Z(n16069) );
  XOR U15431 ( .A(n16070), .B(n16073), .Z(n16071) );
  XOR U15432 ( .A(n16066), .B(n16034), .Z(n16067) );
  XOR U15433 ( .A(n16074), .B(n16075), .Z(n16034) );
  AND U15434 ( .A(n978), .B(n16076), .Z(n16074) );
  XOR U15435 ( .A(n16077), .B(n16075), .Z(n16076) );
  XNOR U15436 ( .A(n16078), .B(n16079), .Z(n16066) );
  NAND U15437 ( .A(n16080), .B(n16081), .Z(n16079) );
  XOR U15438 ( .A(n16082), .B(n16058), .Z(n16081) );
  XOR U15439 ( .A(n16072), .B(n16073), .Z(n16058) );
  XOR U15440 ( .A(n16083), .B(n16084), .Z(n16073) );
  ANDN U15441 ( .B(n16085), .A(n16086), .Z(n16083) );
  XOR U15442 ( .A(n16084), .B(n16087), .Z(n16085) );
  XOR U15443 ( .A(n16088), .B(n16089), .Z(n16072) );
  XOR U15444 ( .A(n16090), .B(n16091), .Z(n16089) );
  ANDN U15445 ( .B(n16092), .A(n16093), .Z(n16090) );
  XOR U15446 ( .A(n16094), .B(n16091), .Z(n16092) );
  IV U15447 ( .A(n16070), .Z(n16088) );
  XOR U15448 ( .A(n16095), .B(n16096), .Z(n16070) );
  ANDN U15449 ( .B(n16097), .A(n16098), .Z(n16095) );
  XOR U15450 ( .A(n16096), .B(n16099), .Z(n16097) );
  IV U15451 ( .A(n16078), .Z(n16082) );
  XOR U15452 ( .A(n16078), .B(n16060), .Z(n16080) );
  XOR U15453 ( .A(n16100), .B(n16101), .Z(n16060) );
  AND U15454 ( .A(n978), .B(n16102), .Z(n16100) );
  XOR U15455 ( .A(n16103), .B(n16101), .Z(n16102) );
  NANDN U15456 ( .A(n16062), .B(n16064), .Z(n16078) );
  XOR U15457 ( .A(n16104), .B(n16105), .Z(n16064) );
  AND U15458 ( .A(n978), .B(n16106), .Z(n16104) );
  XOR U15459 ( .A(n16105), .B(n16107), .Z(n16106) );
  XOR U15460 ( .A(n16108), .B(n16109), .Z(n978) );
  AND U15461 ( .A(n16110), .B(n16111), .Z(n16108) );
  XNOR U15462 ( .A(n16109), .B(n16075), .Z(n16111) );
  XNOR U15463 ( .A(n16112), .B(n16113), .Z(n16075) );
  ANDN U15464 ( .B(n16114), .A(n16115), .Z(n16112) );
  XOR U15465 ( .A(n16113), .B(n16116), .Z(n16114) );
  XOR U15466 ( .A(n16109), .B(n16077), .Z(n16110) );
  XOR U15467 ( .A(n16117), .B(n16118), .Z(n16077) );
  AND U15468 ( .A(n982), .B(n16119), .Z(n16117) );
  XOR U15469 ( .A(n16120), .B(n16118), .Z(n16119) );
  XNOR U15470 ( .A(n16121), .B(n16122), .Z(n16109) );
  NAND U15471 ( .A(n16123), .B(n16124), .Z(n16122) );
  XOR U15472 ( .A(n16125), .B(n16101), .Z(n16124) );
  XOR U15473 ( .A(n16115), .B(n16116), .Z(n16101) );
  XOR U15474 ( .A(n16126), .B(n16127), .Z(n16116) );
  ANDN U15475 ( .B(n16128), .A(n16129), .Z(n16126) );
  XOR U15476 ( .A(n16127), .B(n16130), .Z(n16128) );
  XOR U15477 ( .A(n16131), .B(n16132), .Z(n16115) );
  XOR U15478 ( .A(n16133), .B(n16134), .Z(n16132) );
  ANDN U15479 ( .B(n16135), .A(n16136), .Z(n16133) );
  XOR U15480 ( .A(n16137), .B(n16134), .Z(n16135) );
  IV U15481 ( .A(n16113), .Z(n16131) );
  XOR U15482 ( .A(n16138), .B(n16139), .Z(n16113) );
  ANDN U15483 ( .B(n16140), .A(n16141), .Z(n16138) );
  XOR U15484 ( .A(n16139), .B(n16142), .Z(n16140) );
  IV U15485 ( .A(n16121), .Z(n16125) );
  XOR U15486 ( .A(n16121), .B(n16103), .Z(n16123) );
  XOR U15487 ( .A(n16143), .B(n16144), .Z(n16103) );
  AND U15488 ( .A(n982), .B(n16145), .Z(n16143) );
  XOR U15489 ( .A(n16146), .B(n16144), .Z(n16145) );
  NANDN U15490 ( .A(n16105), .B(n16107), .Z(n16121) );
  XOR U15491 ( .A(n16147), .B(n16148), .Z(n16107) );
  AND U15492 ( .A(n982), .B(n16149), .Z(n16147) );
  XOR U15493 ( .A(n16148), .B(n16150), .Z(n16149) );
  XOR U15494 ( .A(n16151), .B(n16152), .Z(n982) );
  AND U15495 ( .A(n16153), .B(n16154), .Z(n16151) );
  XNOR U15496 ( .A(n16152), .B(n16118), .Z(n16154) );
  XNOR U15497 ( .A(n16155), .B(n16156), .Z(n16118) );
  ANDN U15498 ( .B(n16157), .A(n16158), .Z(n16155) );
  XOR U15499 ( .A(n16156), .B(n16159), .Z(n16157) );
  XOR U15500 ( .A(n16152), .B(n16120), .Z(n16153) );
  XOR U15501 ( .A(n16160), .B(n16161), .Z(n16120) );
  AND U15502 ( .A(n986), .B(n16162), .Z(n16160) );
  XOR U15503 ( .A(n16163), .B(n16161), .Z(n16162) );
  XNOR U15504 ( .A(n16164), .B(n16165), .Z(n16152) );
  NAND U15505 ( .A(n16166), .B(n16167), .Z(n16165) );
  XOR U15506 ( .A(n16168), .B(n16144), .Z(n16167) );
  XOR U15507 ( .A(n16158), .B(n16159), .Z(n16144) );
  XOR U15508 ( .A(n16169), .B(n16170), .Z(n16159) );
  ANDN U15509 ( .B(n16171), .A(n16172), .Z(n16169) );
  XOR U15510 ( .A(n16170), .B(n16173), .Z(n16171) );
  XOR U15511 ( .A(n16174), .B(n16175), .Z(n16158) );
  XOR U15512 ( .A(n16176), .B(n16177), .Z(n16175) );
  ANDN U15513 ( .B(n16178), .A(n16179), .Z(n16176) );
  XOR U15514 ( .A(n16180), .B(n16177), .Z(n16178) );
  IV U15515 ( .A(n16156), .Z(n16174) );
  XOR U15516 ( .A(n16181), .B(n16182), .Z(n16156) );
  ANDN U15517 ( .B(n16183), .A(n16184), .Z(n16181) );
  XOR U15518 ( .A(n16182), .B(n16185), .Z(n16183) );
  IV U15519 ( .A(n16164), .Z(n16168) );
  XOR U15520 ( .A(n16164), .B(n16146), .Z(n16166) );
  XOR U15521 ( .A(n16186), .B(n16187), .Z(n16146) );
  AND U15522 ( .A(n986), .B(n16188), .Z(n16186) );
  XOR U15523 ( .A(n16189), .B(n16187), .Z(n16188) );
  NANDN U15524 ( .A(n16148), .B(n16150), .Z(n16164) );
  XOR U15525 ( .A(n16190), .B(n16191), .Z(n16150) );
  AND U15526 ( .A(n986), .B(n16192), .Z(n16190) );
  XOR U15527 ( .A(n16191), .B(n16193), .Z(n16192) );
  XOR U15528 ( .A(n16194), .B(n16195), .Z(n986) );
  AND U15529 ( .A(n16196), .B(n16197), .Z(n16194) );
  XNOR U15530 ( .A(n16195), .B(n16161), .Z(n16197) );
  XNOR U15531 ( .A(n16198), .B(n16199), .Z(n16161) );
  ANDN U15532 ( .B(n16200), .A(n16201), .Z(n16198) );
  XOR U15533 ( .A(n16199), .B(n16202), .Z(n16200) );
  XOR U15534 ( .A(n16195), .B(n16163), .Z(n16196) );
  XOR U15535 ( .A(n16203), .B(n16204), .Z(n16163) );
  AND U15536 ( .A(n990), .B(n16205), .Z(n16203) );
  XOR U15537 ( .A(n16206), .B(n16204), .Z(n16205) );
  XNOR U15538 ( .A(n16207), .B(n16208), .Z(n16195) );
  NAND U15539 ( .A(n16209), .B(n16210), .Z(n16208) );
  XOR U15540 ( .A(n16211), .B(n16187), .Z(n16210) );
  XOR U15541 ( .A(n16201), .B(n16202), .Z(n16187) );
  XOR U15542 ( .A(n16212), .B(n16213), .Z(n16202) );
  ANDN U15543 ( .B(n16214), .A(n16215), .Z(n16212) );
  XOR U15544 ( .A(n16213), .B(n16216), .Z(n16214) );
  XOR U15545 ( .A(n16217), .B(n16218), .Z(n16201) );
  XOR U15546 ( .A(n16219), .B(n16220), .Z(n16218) );
  ANDN U15547 ( .B(n16221), .A(n16222), .Z(n16219) );
  XOR U15548 ( .A(n16223), .B(n16220), .Z(n16221) );
  IV U15549 ( .A(n16199), .Z(n16217) );
  XOR U15550 ( .A(n16224), .B(n16225), .Z(n16199) );
  ANDN U15551 ( .B(n16226), .A(n16227), .Z(n16224) );
  XOR U15552 ( .A(n16225), .B(n16228), .Z(n16226) );
  IV U15553 ( .A(n16207), .Z(n16211) );
  XOR U15554 ( .A(n16207), .B(n16189), .Z(n16209) );
  XOR U15555 ( .A(n16229), .B(n16230), .Z(n16189) );
  AND U15556 ( .A(n990), .B(n16231), .Z(n16229) );
  XOR U15557 ( .A(n16232), .B(n16230), .Z(n16231) );
  NANDN U15558 ( .A(n16191), .B(n16193), .Z(n16207) );
  XOR U15559 ( .A(n16233), .B(n16234), .Z(n16193) );
  AND U15560 ( .A(n990), .B(n16235), .Z(n16233) );
  XOR U15561 ( .A(n16234), .B(n16236), .Z(n16235) );
  XOR U15562 ( .A(n16237), .B(n16238), .Z(n990) );
  AND U15563 ( .A(n16239), .B(n16240), .Z(n16237) );
  XNOR U15564 ( .A(n16238), .B(n16204), .Z(n16240) );
  XNOR U15565 ( .A(n16241), .B(n16242), .Z(n16204) );
  ANDN U15566 ( .B(n16243), .A(n16244), .Z(n16241) );
  XOR U15567 ( .A(n16242), .B(n16245), .Z(n16243) );
  XOR U15568 ( .A(n16238), .B(n16206), .Z(n16239) );
  XOR U15569 ( .A(n16246), .B(n16247), .Z(n16206) );
  AND U15570 ( .A(n994), .B(n16248), .Z(n16246) );
  XOR U15571 ( .A(n16249), .B(n16247), .Z(n16248) );
  XNOR U15572 ( .A(n16250), .B(n16251), .Z(n16238) );
  NAND U15573 ( .A(n16252), .B(n16253), .Z(n16251) );
  XOR U15574 ( .A(n16254), .B(n16230), .Z(n16253) );
  XOR U15575 ( .A(n16244), .B(n16245), .Z(n16230) );
  XOR U15576 ( .A(n16255), .B(n16256), .Z(n16245) );
  ANDN U15577 ( .B(n16257), .A(n16258), .Z(n16255) );
  XOR U15578 ( .A(n16256), .B(n16259), .Z(n16257) );
  XOR U15579 ( .A(n16260), .B(n16261), .Z(n16244) );
  XOR U15580 ( .A(n16262), .B(n16263), .Z(n16261) );
  ANDN U15581 ( .B(n16264), .A(n16265), .Z(n16262) );
  XOR U15582 ( .A(n16266), .B(n16263), .Z(n16264) );
  IV U15583 ( .A(n16242), .Z(n16260) );
  XOR U15584 ( .A(n16267), .B(n16268), .Z(n16242) );
  ANDN U15585 ( .B(n16269), .A(n16270), .Z(n16267) );
  XOR U15586 ( .A(n16268), .B(n16271), .Z(n16269) );
  IV U15587 ( .A(n16250), .Z(n16254) );
  XOR U15588 ( .A(n16250), .B(n16232), .Z(n16252) );
  XOR U15589 ( .A(n16272), .B(n16273), .Z(n16232) );
  AND U15590 ( .A(n994), .B(n16274), .Z(n16272) );
  XOR U15591 ( .A(n16275), .B(n16273), .Z(n16274) );
  NANDN U15592 ( .A(n16234), .B(n16236), .Z(n16250) );
  XOR U15593 ( .A(n16276), .B(n16277), .Z(n16236) );
  AND U15594 ( .A(n994), .B(n16278), .Z(n16276) );
  XOR U15595 ( .A(n16277), .B(n16279), .Z(n16278) );
  XOR U15596 ( .A(n16280), .B(n16281), .Z(n994) );
  AND U15597 ( .A(n16282), .B(n16283), .Z(n16280) );
  XNOR U15598 ( .A(n16281), .B(n16247), .Z(n16283) );
  XNOR U15599 ( .A(n16284), .B(n16285), .Z(n16247) );
  ANDN U15600 ( .B(n16286), .A(n16287), .Z(n16284) );
  XOR U15601 ( .A(n16285), .B(n16288), .Z(n16286) );
  XOR U15602 ( .A(n16281), .B(n16249), .Z(n16282) );
  XOR U15603 ( .A(n16289), .B(n16290), .Z(n16249) );
  AND U15604 ( .A(n998), .B(n16291), .Z(n16289) );
  XOR U15605 ( .A(n16292), .B(n16290), .Z(n16291) );
  XNOR U15606 ( .A(n16293), .B(n16294), .Z(n16281) );
  NAND U15607 ( .A(n16295), .B(n16296), .Z(n16294) );
  XOR U15608 ( .A(n16297), .B(n16273), .Z(n16296) );
  XOR U15609 ( .A(n16287), .B(n16288), .Z(n16273) );
  XOR U15610 ( .A(n16298), .B(n16299), .Z(n16288) );
  ANDN U15611 ( .B(n16300), .A(n16301), .Z(n16298) );
  XOR U15612 ( .A(n16299), .B(n16302), .Z(n16300) );
  XOR U15613 ( .A(n16303), .B(n16304), .Z(n16287) );
  XOR U15614 ( .A(n16305), .B(n16306), .Z(n16304) );
  ANDN U15615 ( .B(n16307), .A(n16308), .Z(n16305) );
  XOR U15616 ( .A(n16309), .B(n16306), .Z(n16307) );
  IV U15617 ( .A(n16285), .Z(n16303) );
  XOR U15618 ( .A(n16310), .B(n16311), .Z(n16285) );
  ANDN U15619 ( .B(n16312), .A(n16313), .Z(n16310) );
  XOR U15620 ( .A(n16311), .B(n16314), .Z(n16312) );
  IV U15621 ( .A(n16293), .Z(n16297) );
  XOR U15622 ( .A(n16293), .B(n16275), .Z(n16295) );
  XOR U15623 ( .A(n16315), .B(n16316), .Z(n16275) );
  AND U15624 ( .A(n998), .B(n16317), .Z(n16315) );
  XOR U15625 ( .A(n16318), .B(n16316), .Z(n16317) );
  NANDN U15626 ( .A(n16277), .B(n16279), .Z(n16293) );
  XOR U15627 ( .A(n16319), .B(n16320), .Z(n16279) );
  AND U15628 ( .A(n998), .B(n16321), .Z(n16319) );
  XOR U15629 ( .A(n16320), .B(n16322), .Z(n16321) );
  XOR U15630 ( .A(n16323), .B(n16324), .Z(n998) );
  AND U15631 ( .A(n16325), .B(n16326), .Z(n16323) );
  XNOR U15632 ( .A(n16324), .B(n16290), .Z(n16326) );
  XNOR U15633 ( .A(n16327), .B(n16328), .Z(n16290) );
  ANDN U15634 ( .B(n16329), .A(n16330), .Z(n16327) );
  XOR U15635 ( .A(n16328), .B(n16331), .Z(n16329) );
  XOR U15636 ( .A(n16324), .B(n16292), .Z(n16325) );
  XOR U15637 ( .A(n16332), .B(n16333), .Z(n16292) );
  AND U15638 ( .A(n1002), .B(n16334), .Z(n16332) );
  XOR U15639 ( .A(n16335), .B(n16333), .Z(n16334) );
  XNOR U15640 ( .A(n16336), .B(n16337), .Z(n16324) );
  NAND U15641 ( .A(n16338), .B(n16339), .Z(n16337) );
  XOR U15642 ( .A(n16340), .B(n16316), .Z(n16339) );
  XOR U15643 ( .A(n16330), .B(n16331), .Z(n16316) );
  XOR U15644 ( .A(n16341), .B(n16342), .Z(n16331) );
  ANDN U15645 ( .B(n16343), .A(n16344), .Z(n16341) );
  XOR U15646 ( .A(n16342), .B(n16345), .Z(n16343) );
  XOR U15647 ( .A(n16346), .B(n16347), .Z(n16330) );
  XOR U15648 ( .A(n16348), .B(n16349), .Z(n16347) );
  ANDN U15649 ( .B(n16350), .A(n16351), .Z(n16348) );
  XOR U15650 ( .A(n16352), .B(n16349), .Z(n16350) );
  IV U15651 ( .A(n16328), .Z(n16346) );
  XOR U15652 ( .A(n16353), .B(n16354), .Z(n16328) );
  ANDN U15653 ( .B(n16355), .A(n16356), .Z(n16353) );
  XOR U15654 ( .A(n16354), .B(n16357), .Z(n16355) );
  IV U15655 ( .A(n16336), .Z(n16340) );
  XOR U15656 ( .A(n16336), .B(n16318), .Z(n16338) );
  XOR U15657 ( .A(n16358), .B(n16359), .Z(n16318) );
  AND U15658 ( .A(n1002), .B(n16360), .Z(n16358) );
  XOR U15659 ( .A(n16361), .B(n16359), .Z(n16360) );
  NANDN U15660 ( .A(n16320), .B(n16322), .Z(n16336) );
  XOR U15661 ( .A(n16362), .B(n16363), .Z(n16322) );
  AND U15662 ( .A(n1002), .B(n16364), .Z(n16362) );
  XOR U15663 ( .A(n16363), .B(n16365), .Z(n16364) );
  XOR U15664 ( .A(n16366), .B(n16367), .Z(n1002) );
  AND U15665 ( .A(n16368), .B(n16369), .Z(n16366) );
  XNOR U15666 ( .A(n16367), .B(n16333), .Z(n16369) );
  XNOR U15667 ( .A(n16370), .B(n16371), .Z(n16333) );
  ANDN U15668 ( .B(n16372), .A(n16373), .Z(n16370) );
  XOR U15669 ( .A(n16371), .B(n16374), .Z(n16372) );
  XOR U15670 ( .A(n16367), .B(n16335), .Z(n16368) );
  XOR U15671 ( .A(n16375), .B(n16376), .Z(n16335) );
  AND U15672 ( .A(n1006), .B(n16377), .Z(n16375) );
  XOR U15673 ( .A(n16378), .B(n16376), .Z(n16377) );
  XNOR U15674 ( .A(n16379), .B(n16380), .Z(n16367) );
  NAND U15675 ( .A(n16381), .B(n16382), .Z(n16380) );
  XOR U15676 ( .A(n16383), .B(n16359), .Z(n16382) );
  XOR U15677 ( .A(n16373), .B(n16374), .Z(n16359) );
  XOR U15678 ( .A(n16384), .B(n16385), .Z(n16374) );
  ANDN U15679 ( .B(n16386), .A(n16387), .Z(n16384) );
  XOR U15680 ( .A(n16385), .B(n16388), .Z(n16386) );
  XOR U15681 ( .A(n16389), .B(n16390), .Z(n16373) );
  XOR U15682 ( .A(n16391), .B(n16392), .Z(n16390) );
  ANDN U15683 ( .B(n16393), .A(n16394), .Z(n16391) );
  XOR U15684 ( .A(n16395), .B(n16392), .Z(n16393) );
  IV U15685 ( .A(n16371), .Z(n16389) );
  XOR U15686 ( .A(n16396), .B(n16397), .Z(n16371) );
  ANDN U15687 ( .B(n16398), .A(n16399), .Z(n16396) );
  XOR U15688 ( .A(n16397), .B(n16400), .Z(n16398) );
  IV U15689 ( .A(n16379), .Z(n16383) );
  XOR U15690 ( .A(n16379), .B(n16361), .Z(n16381) );
  XOR U15691 ( .A(n16401), .B(n16402), .Z(n16361) );
  AND U15692 ( .A(n1006), .B(n16403), .Z(n16401) );
  XOR U15693 ( .A(n16404), .B(n16402), .Z(n16403) );
  NANDN U15694 ( .A(n16363), .B(n16365), .Z(n16379) );
  XOR U15695 ( .A(n16405), .B(n16406), .Z(n16365) );
  AND U15696 ( .A(n1006), .B(n16407), .Z(n16405) );
  XOR U15697 ( .A(n16406), .B(n16408), .Z(n16407) );
  XOR U15698 ( .A(n16409), .B(n16410), .Z(n1006) );
  AND U15699 ( .A(n16411), .B(n16412), .Z(n16409) );
  XNOR U15700 ( .A(n16410), .B(n16376), .Z(n16412) );
  XNOR U15701 ( .A(n16413), .B(n16414), .Z(n16376) );
  ANDN U15702 ( .B(n16415), .A(n16416), .Z(n16413) );
  XOR U15703 ( .A(n16414), .B(n16417), .Z(n16415) );
  XOR U15704 ( .A(n16410), .B(n16378), .Z(n16411) );
  XOR U15705 ( .A(n16418), .B(n16419), .Z(n16378) );
  AND U15706 ( .A(n1010), .B(n16420), .Z(n16418) );
  XOR U15707 ( .A(n16421), .B(n16419), .Z(n16420) );
  XNOR U15708 ( .A(n16422), .B(n16423), .Z(n16410) );
  NAND U15709 ( .A(n16424), .B(n16425), .Z(n16423) );
  XOR U15710 ( .A(n16426), .B(n16402), .Z(n16425) );
  XOR U15711 ( .A(n16416), .B(n16417), .Z(n16402) );
  XOR U15712 ( .A(n16427), .B(n16428), .Z(n16417) );
  ANDN U15713 ( .B(n16429), .A(n16430), .Z(n16427) );
  XOR U15714 ( .A(n16428), .B(n16431), .Z(n16429) );
  XOR U15715 ( .A(n16432), .B(n16433), .Z(n16416) );
  XOR U15716 ( .A(n16434), .B(n16435), .Z(n16433) );
  ANDN U15717 ( .B(n16436), .A(n16437), .Z(n16434) );
  XOR U15718 ( .A(n16438), .B(n16435), .Z(n16436) );
  IV U15719 ( .A(n16414), .Z(n16432) );
  XOR U15720 ( .A(n16439), .B(n16440), .Z(n16414) );
  ANDN U15721 ( .B(n16441), .A(n16442), .Z(n16439) );
  XOR U15722 ( .A(n16440), .B(n16443), .Z(n16441) );
  IV U15723 ( .A(n16422), .Z(n16426) );
  XOR U15724 ( .A(n16422), .B(n16404), .Z(n16424) );
  XOR U15725 ( .A(n16444), .B(n16445), .Z(n16404) );
  AND U15726 ( .A(n1010), .B(n16446), .Z(n16444) );
  XOR U15727 ( .A(n16447), .B(n16445), .Z(n16446) );
  NANDN U15728 ( .A(n16406), .B(n16408), .Z(n16422) );
  XOR U15729 ( .A(n16448), .B(n16449), .Z(n16408) );
  AND U15730 ( .A(n1010), .B(n16450), .Z(n16448) );
  XOR U15731 ( .A(n16449), .B(n16451), .Z(n16450) );
  XOR U15732 ( .A(n16452), .B(n16453), .Z(n1010) );
  AND U15733 ( .A(n16454), .B(n16455), .Z(n16452) );
  XNOR U15734 ( .A(n16453), .B(n16419), .Z(n16455) );
  XNOR U15735 ( .A(n16456), .B(n16457), .Z(n16419) );
  ANDN U15736 ( .B(n16458), .A(n16459), .Z(n16456) );
  XOR U15737 ( .A(n16457), .B(n16460), .Z(n16458) );
  XOR U15738 ( .A(n16453), .B(n16421), .Z(n16454) );
  XOR U15739 ( .A(n16461), .B(n16462), .Z(n16421) );
  AND U15740 ( .A(n1014), .B(n16463), .Z(n16461) );
  XOR U15741 ( .A(n16464), .B(n16462), .Z(n16463) );
  XNOR U15742 ( .A(n16465), .B(n16466), .Z(n16453) );
  NAND U15743 ( .A(n16467), .B(n16468), .Z(n16466) );
  XOR U15744 ( .A(n16469), .B(n16445), .Z(n16468) );
  XOR U15745 ( .A(n16459), .B(n16460), .Z(n16445) );
  XOR U15746 ( .A(n16470), .B(n16471), .Z(n16460) );
  ANDN U15747 ( .B(n16472), .A(n16473), .Z(n16470) );
  XOR U15748 ( .A(n16471), .B(n16474), .Z(n16472) );
  XOR U15749 ( .A(n16475), .B(n16476), .Z(n16459) );
  XOR U15750 ( .A(n16477), .B(n16478), .Z(n16476) );
  ANDN U15751 ( .B(n16479), .A(n16480), .Z(n16477) );
  XOR U15752 ( .A(n16481), .B(n16478), .Z(n16479) );
  IV U15753 ( .A(n16457), .Z(n16475) );
  XOR U15754 ( .A(n16482), .B(n16483), .Z(n16457) );
  ANDN U15755 ( .B(n16484), .A(n16485), .Z(n16482) );
  XOR U15756 ( .A(n16483), .B(n16486), .Z(n16484) );
  IV U15757 ( .A(n16465), .Z(n16469) );
  XOR U15758 ( .A(n16465), .B(n16447), .Z(n16467) );
  XOR U15759 ( .A(n16487), .B(n16488), .Z(n16447) );
  AND U15760 ( .A(n1014), .B(n16489), .Z(n16487) );
  XOR U15761 ( .A(n16490), .B(n16488), .Z(n16489) );
  NANDN U15762 ( .A(n16449), .B(n16451), .Z(n16465) );
  XOR U15763 ( .A(n16491), .B(n16492), .Z(n16451) );
  AND U15764 ( .A(n1014), .B(n16493), .Z(n16491) );
  XOR U15765 ( .A(n16492), .B(n16494), .Z(n16493) );
  XOR U15766 ( .A(n16495), .B(n16496), .Z(n1014) );
  AND U15767 ( .A(n16497), .B(n16498), .Z(n16495) );
  XNOR U15768 ( .A(n16496), .B(n16462), .Z(n16498) );
  XNOR U15769 ( .A(n16499), .B(n16500), .Z(n16462) );
  ANDN U15770 ( .B(n16501), .A(n16502), .Z(n16499) );
  XOR U15771 ( .A(n16500), .B(n16503), .Z(n16501) );
  XOR U15772 ( .A(n16496), .B(n16464), .Z(n16497) );
  XOR U15773 ( .A(n16504), .B(n16505), .Z(n16464) );
  AND U15774 ( .A(n1018), .B(n16506), .Z(n16504) );
  XOR U15775 ( .A(n16507), .B(n16505), .Z(n16506) );
  XNOR U15776 ( .A(n16508), .B(n16509), .Z(n16496) );
  NAND U15777 ( .A(n16510), .B(n16511), .Z(n16509) );
  XOR U15778 ( .A(n16512), .B(n16488), .Z(n16511) );
  XOR U15779 ( .A(n16502), .B(n16503), .Z(n16488) );
  XOR U15780 ( .A(n16513), .B(n16514), .Z(n16503) );
  ANDN U15781 ( .B(n16515), .A(n16516), .Z(n16513) );
  XOR U15782 ( .A(n16514), .B(n16517), .Z(n16515) );
  XOR U15783 ( .A(n16518), .B(n16519), .Z(n16502) );
  XOR U15784 ( .A(n16520), .B(n16521), .Z(n16519) );
  ANDN U15785 ( .B(n16522), .A(n16523), .Z(n16520) );
  XOR U15786 ( .A(n16524), .B(n16521), .Z(n16522) );
  IV U15787 ( .A(n16500), .Z(n16518) );
  XOR U15788 ( .A(n16525), .B(n16526), .Z(n16500) );
  ANDN U15789 ( .B(n16527), .A(n16528), .Z(n16525) );
  XOR U15790 ( .A(n16526), .B(n16529), .Z(n16527) );
  IV U15791 ( .A(n16508), .Z(n16512) );
  XOR U15792 ( .A(n16508), .B(n16490), .Z(n16510) );
  XOR U15793 ( .A(n16530), .B(n16531), .Z(n16490) );
  AND U15794 ( .A(n1018), .B(n16532), .Z(n16530) );
  XNOR U15795 ( .A(n16533), .B(n16531), .Z(n16532) );
  NANDN U15796 ( .A(n16492), .B(n16494), .Z(n16508) );
  XOR U15797 ( .A(n16534), .B(n16535), .Z(n16494) );
  AND U15798 ( .A(n1018), .B(n16536), .Z(n16534) );
  XOR U15799 ( .A(n16535), .B(n16537), .Z(n16536) );
  XOR U15800 ( .A(n16538), .B(n16539), .Z(n1018) );
  AND U15801 ( .A(n16540), .B(n16541), .Z(n16538) );
  XNOR U15802 ( .A(n16539), .B(n16505), .Z(n16541) );
  XNOR U15803 ( .A(n16542), .B(n16543), .Z(n16505) );
  ANDN U15804 ( .B(n16544), .A(n16545), .Z(n16542) );
  XOR U15805 ( .A(n16543), .B(n16546), .Z(n16544) );
  XOR U15806 ( .A(n16539), .B(n16507), .Z(n16540) );
  XNOR U15807 ( .A(n16547), .B(n16548), .Z(n16507) );
  ANDN U15808 ( .B(n16549), .A(n16550), .Z(n16547) );
  XOR U15809 ( .A(n16548), .B(n16551), .Z(n16549) );
  XNOR U15810 ( .A(n16552), .B(n16553), .Z(n16539) );
  NAND U15811 ( .A(n16554), .B(n16555), .Z(n16553) );
  XOR U15812 ( .A(n16556), .B(n16531), .Z(n16555) );
  XOR U15813 ( .A(n16545), .B(n16546), .Z(n16531) );
  XOR U15814 ( .A(n16557), .B(n16558), .Z(n16546) );
  ANDN U15815 ( .B(n16559), .A(n16560), .Z(n16557) );
  XOR U15816 ( .A(n16558), .B(n16561), .Z(n16559) );
  XOR U15817 ( .A(n16562), .B(n16563), .Z(n16545) );
  XOR U15818 ( .A(n16564), .B(n16565), .Z(n16563) );
  ANDN U15819 ( .B(n16566), .A(n16567), .Z(n16564) );
  XOR U15820 ( .A(n16568), .B(n16565), .Z(n16566) );
  IV U15821 ( .A(n16543), .Z(n16562) );
  XOR U15822 ( .A(n16569), .B(n16570), .Z(n16543) );
  ANDN U15823 ( .B(n16571), .A(n16572), .Z(n16569) );
  XOR U15824 ( .A(n16570), .B(n16573), .Z(n16571) );
  IV U15825 ( .A(n16552), .Z(n16556) );
  XNOR U15826 ( .A(n16552), .B(n16533), .Z(n16554) );
  XOR U15827 ( .A(n16574), .B(n16551), .Z(n16533) );
  XOR U15828 ( .A(n16575), .B(n16576), .Z(n16551) );
  ANDN U15829 ( .B(n16577), .A(n16578), .Z(n16575) );
  XOR U15830 ( .A(n16576), .B(n16579), .Z(n16577) );
  IV U15831 ( .A(n16550), .Z(n16574) );
  XOR U15832 ( .A(n16580), .B(n16581), .Z(n16550) );
  XOR U15833 ( .A(n16582), .B(n16583), .Z(n16581) );
  ANDN U15834 ( .B(n16584), .A(n16585), .Z(n16582) );
  XOR U15835 ( .A(n16586), .B(n16583), .Z(n16584) );
  IV U15836 ( .A(n16548), .Z(n16580) );
  XNOR U15837 ( .A(n16587), .B(n16588), .Z(n16548) );
  ANDN U15838 ( .B(n16589), .A(n16590), .Z(n16587) );
  XNOR U15839 ( .A(n16588), .B(n16591), .Z(n16589) );
  NANDN U15840 ( .A(n16535), .B(n16537), .Z(n16552) );
  XOR U15841 ( .A(n16592), .B(n16591), .Z(n16537) );
  XOR U15842 ( .A(n16593), .B(n16579), .Z(n16591) );
  XNOR U15843 ( .A(q[6]), .B(DB[6]), .Z(n16579) );
  IV U15844 ( .A(n16578), .Z(n16593) );
  XNOR U15845 ( .A(n16576), .B(n16594), .Z(n16578) );
  XNOR U15846 ( .A(q[5]), .B(DB[5]), .Z(n16594) );
  XNOR U15847 ( .A(q[4]), .B(DB[4]), .Z(n16576) );
  IV U15848 ( .A(n16590), .Z(n16592) );
  XOR U15849 ( .A(n16595), .B(n16596), .Z(n16590) );
  XOR U15850 ( .A(n16588), .B(n16586), .Z(n16596) );
  XNOR U15851 ( .A(q[3]), .B(DB[3]), .Z(n16586) );
  XOR U15852 ( .A(q[0]), .B(DB[0]), .Z(n16588) );
  IV U15853 ( .A(n16585), .Z(n16595) );
  XNOR U15854 ( .A(n16583), .B(n16597), .Z(n16585) );
  XNOR U15855 ( .A(q[2]), .B(DB[2]), .Z(n16597) );
  XNOR U15856 ( .A(q[1]), .B(DB[1]), .Z(n16583) );
  XOR U15857 ( .A(n16598), .B(n16573), .Z(n16535) );
  XOR U15858 ( .A(n16599), .B(n16561), .Z(n16573) );
  XNOR U15859 ( .A(q[6]), .B(DB[13]), .Z(n16561) );
  IV U15860 ( .A(n16560), .Z(n16599) );
  XNOR U15861 ( .A(n16558), .B(n16600), .Z(n16560) );
  XNOR U15862 ( .A(q[5]), .B(DB[12]), .Z(n16600) );
  XNOR U15863 ( .A(q[4]), .B(DB[11]), .Z(n16558) );
  IV U15864 ( .A(n16572), .Z(n16598) );
  XOR U15865 ( .A(n16601), .B(n16602), .Z(n16572) );
  XNOR U15866 ( .A(n16568), .B(n16570), .Z(n16602) );
  XNOR U15867 ( .A(q[0]), .B(DB[7]), .Z(n16570) );
  XNOR U15868 ( .A(q[3]), .B(DB[10]), .Z(n16568) );
  IV U15869 ( .A(n16567), .Z(n16601) );
  XNOR U15870 ( .A(n16565), .B(n16603), .Z(n16567) );
  XNOR U15871 ( .A(q[2]), .B(DB[9]), .Z(n16603) );
  XNOR U15872 ( .A(q[1]), .B(DB[8]), .Z(n16565) );
  XOR U15873 ( .A(n16604), .B(n16529), .Z(n16492) );
  XOR U15874 ( .A(n16605), .B(n16517), .Z(n16529) );
  XNOR U15875 ( .A(q[6]), .B(DB[20]), .Z(n16517) );
  IV U15876 ( .A(n16516), .Z(n16605) );
  XNOR U15877 ( .A(n16514), .B(n16606), .Z(n16516) );
  XNOR U15878 ( .A(q[5]), .B(DB[19]), .Z(n16606) );
  XNOR U15879 ( .A(q[4]), .B(DB[18]), .Z(n16514) );
  IV U15880 ( .A(n16528), .Z(n16604) );
  XOR U15881 ( .A(n16607), .B(n16608), .Z(n16528) );
  XNOR U15882 ( .A(n16524), .B(n16526), .Z(n16608) );
  XNOR U15883 ( .A(q[0]), .B(DB[14]), .Z(n16526) );
  XNOR U15884 ( .A(q[3]), .B(DB[17]), .Z(n16524) );
  IV U15885 ( .A(n16523), .Z(n16607) );
  XNOR U15886 ( .A(n16521), .B(n16609), .Z(n16523) );
  XNOR U15887 ( .A(q[2]), .B(DB[16]), .Z(n16609) );
  XNOR U15888 ( .A(q[1]), .B(DB[15]), .Z(n16521) );
  XOR U15889 ( .A(n16610), .B(n16486), .Z(n16449) );
  XOR U15890 ( .A(n16611), .B(n16474), .Z(n16486) );
  XNOR U15891 ( .A(q[6]), .B(DB[27]), .Z(n16474) );
  IV U15892 ( .A(n16473), .Z(n16611) );
  XNOR U15893 ( .A(n16471), .B(n16612), .Z(n16473) );
  XNOR U15894 ( .A(q[5]), .B(DB[26]), .Z(n16612) );
  XNOR U15895 ( .A(q[4]), .B(DB[25]), .Z(n16471) );
  IV U15896 ( .A(n16485), .Z(n16610) );
  XOR U15897 ( .A(n16613), .B(n16614), .Z(n16485) );
  XNOR U15898 ( .A(n16481), .B(n16483), .Z(n16614) );
  XNOR U15899 ( .A(q[0]), .B(DB[21]), .Z(n16483) );
  XNOR U15900 ( .A(q[3]), .B(DB[24]), .Z(n16481) );
  IV U15901 ( .A(n16480), .Z(n16613) );
  XNOR U15902 ( .A(n16478), .B(n16615), .Z(n16480) );
  XNOR U15903 ( .A(q[2]), .B(DB[23]), .Z(n16615) );
  XNOR U15904 ( .A(q[1]), .B(DB[22]), .Z(n16478) );
  XOR U15905 ( .A(n16616), .B(n16443), .Z(n16406) );
  XOR U15906 ( .A(n16617), .B(n16431), .Z(n16443) );
  XNOR U15907 ( .A(q[6]), .B(DB[34]), .Z(n16431) );
  IV U15908 ( .A(n16430), .Z(n16617) );
  XNOR U15909 ( .A(n16428), .B(n16618), .Z(n16430) );
  XNOR U15910 ( .A(q[5]), .B(DB[33]), .Z(n16618) );
  XNOR U15911 ( .A(q[4]), .B(DB[32]), .Z(n16428) );
  IV U15912 ( .A(n16442), .Z(n16616) );
  XOR U15913 ( .A(n16619), .B(n16620), .Z(n16442) );
  XNOR U15914 ( .A(n16438), .B(n16440), .Z(n16620) );
  XNOR U15915 ( .A(q[0]), .B(DB[28]), .Z(n16440) );
  XNOR U15916 ( .A(q[3]), .B(DB[31]), .Z(n16438) );
  IV U15917 ( .A(n16437), .Z(n16619) );
  XNOR U15918 ( .A(n16435), .B(n16621), .Z(n16437) );
  XNOR U15919 ( .A(q[2]), .B(DB[30]), .Z(n16621) );
  XNOR U15920 ( .A(q[1]), .B(DB[29]), .Z(n16435) );
  XOR U15921 ( .A(n16622), .B(n16400), .Z(n16363) );
  XOR U15922 ( .A(n16623), .B(n16388), .Z(n16400) );
  XNOR U15923 ( .A(q[6]), .B(DB[41]), .Z(n16388) );
  IV U15924 ( .A(n16387), .Z(n16623) );
  XNOR U15925 ( .A(n16385), .B(n16624), .Z(n16387) );
  XNOR U15926 ( .A(q[5]), .B(DB[40]), .Z(n16624) );
  XNOR U15927 ( .A(q[4]), .B(DB[39]), .Z(n16385) );
  IV U15928 ( .A(n16399), .Z(n16622) );
  XOR U15929 ( .A(n16625), .B(n16626), .Z(n16399) );
  XNOR U15930 ( .A(n16395), .B(n16397), .Z(n16626) );
  XNOR U15931 ( .A(q[0]), .B(DB[35]), .Z(n16397) );
  XNOR U15932 ( .A(q[3]), .B(DB[38]), .Z(n16395) );
  IV U15933 ( .A(n16394), .Z(n16625) );
  XNOR U15934 ( .A(n16392), .B(n16627), .Z(n16394) );
  XNOR U15935 ( .A(q[2]), .B(DB[37]), .Z(n16627) );
  XNOR U15936 ( .A(q[1]), .B(DB[36]), .Z(n16392) );
  XOR U15937 ( .A(n16628), .B(n16357), .Z(n16320) );
  XOR U15938 ( .A(n16629), .B(n16345), .Z(n16357) );
  XNOR U15939 ( .A(q[6]), .B(DB[48]), .Z(n16345) );
  IV U15940 ( .A(n16344), .Z(n16629) );
  XNOR U15941 ( .A(n16342), .B(n16630), .Z(n16344) );
  XNOR U15942 ( .A(q[5]), .B(DB[47]), .Z(n16630) );
  XNOR U15943 ( .A(q[4]), .B(DB[46]), .Z(n16342) );
  IV U15944 ( .A(n16356), .Z(n16628) );
  XOR U15945 ( .A(n16631), .B(n16632), .Z(n16356) );
  XNOR U15946 ( .A(n16352), .B(n16354), .Z(n16632) );
  XNOR U15947 ( .A(q[0]), .B(DB[42]), .Z(n16354) );
  XNOR U15948 ( .A(q[3]), .B(DB[45]), .Z(n16352) );
  IV U15949 ( .A(n16351), .Z(n16631) );
  XNOR U15950 ( .A(n16349), .B(n16633), .Z(n16351) );
  XNOR U15951 ( .A(q[2]), .B(DB[44]), .Z(n16633) );
  XNOR U15952 ( .A(q[1]), .B(DB[43]), .Z(n16349) );
  XOR U15953 ( .A(n16634), .B(n16314), .Z(n16277) );
  XOR U15954 ( .A(n16635), .B(n16302), .Z(n16314) );
  XNOR U15955 ( .A(q[6]), .B(DB[55]), .Z(n16302) );
  IV U15956 ( .A(n16301), .Z(n16635) );
  XNOR U15957 ( .A(n16299), .B(n16636), .Z(n16301) );
  XNOR U15958 ( .A(q[5]), .B(DB[54]), .Z(n16636) );
  XNOR U15959 ( .A(q[4]), .B(DB[53]), .Z(n16299) );
  IV U15960 ( .A(n16313), .Z(n16634) );
  XOR U15961 ( .A(n16637), .B(n16638), .Z(n16313) );
  XNOR U15962 ( .A(n16309), .B(n16311), .Z(n16638) );
  XNOR U15963 ( .A(q[0]), .B(DB[49]), .Z(n16311) );
  XNOR U15964 ( .A(q[3]), .B(DB[52]), .Z(n16309) );
  IV U15965 ( .A(n16308), .Z(n16637) );
  XNOR U15966 ( .A(n16306), .B(n16639), .Z(n16308) );
  XNOR U15967 ( .A(q[2]), .B(DB[51]), .Z(n16639) );
  XNOR U15968 ( .A(q[1]), .B(DB[50]), .Z(n16306) );
  XOR U15969 ( .A(n16640), .B(n16271), .Z(n16234) );
  XOR U15970 ( .A(n16641), .B(n16259), .Z(n16271) );
  XNOR U15971 ( .A(q[6]), .B(DB[62]), .Z(n16259) );
  IV U15972 ( .A(n16258), .Z(n16641) );
  XNOR U15973 ( .A(n16256), .B(n16642), .Z(n16258) );
  XNOR U15974 ( .A(q[5]), .B(DB[61]), .Z(n16642) );
  XNOR U15975 ( .A(q[4]), .B(DB[60]), .Z(n16256) );
  IV U15976 ( .A(n16270), .Z(n16640) );
  XOR U15977 ( .A(n16643), .B(n16644), .Z(n16270) );
  XNOR U15978 ( .A(n16266), .B(n16268), .Z(n16644) );
  XNOR U15979 ( .A(q[0]), .B(DB[56]), .Z(n16268) );
  XNOR U15980 ( .A(q[3]), .B(DB[59]), .Z(n16266) );
  IV U15981 ( .A(n16265), .Z(n16643) );
  XNOR U15982 ( .A(n16263), .B(n16645), .Z(n16265) );
  XNOR U15983 ( .A(q[2]), .B(DB[58]), .Z(n16645) );
  XNOR U15984 ( .A(q[1]), .B(DB[57]), .Z(n16263) );
  XOR U15985 ( .A(n16646), .B(n16228), .Z(n16191) );
  XOR U15986 ( .A(n16647), .B(n16216), .Z(n16228) );
  XNOR U15987 ( .A(q[6]), .B(DB[69]), .Z(n16216) );
  IV U15988 ( .A(n16215), .Z(n16647) );
  XNOR U15989 ( .A(n16213), .B(n16648), .Z(n16215) );
  XNOR U15990 ( .A(q[5]), .B(DB[68]), .Z(n16648) );
  XNOR U15991 ( .A(q[4]), .B(DB[67]), .Z(n16213) );
  IV U15992 ( .A(n16227), .Z(n16646) );
  XOR U15993 ( .A(n16649), .B(n16650), .Z(n16227) );
  XNOR U15994 ( .A(n16223), .B(n16225), .Z(n16650) );
  XNOR U15995 ( .A(q[0]), .B(DB[63]), .Z(n16225) );
  XNOR U15996 ( .A(q[3]), .B(DB[66]), .Z(n16223) );
  IV U15997 ( .A(n16222), .Z(n16649) );
  XNOR U15998 ( .A(n16220), .B(n16651), .Z(n16222) );
  XNOR U15999 ( .A(q[2]), .B(DB[65]), .Z(n16651) );
  XNOR U16000 ( .A(q[1]), .B(DB[64]), .Z(n16220) );
  XOR U16001 ( .A(n16652), .B(n16185), .Z(n16148) );
  XOR U16002 ( .A(n16653), .B(n16173), .Z(n16185) );
  XNOR U16003 ( .A(q[6]), .B(DB[76]), .Z(n16173) );
  IV U16004 ( .A(n16172), .Z(n16653) );
  XNOR U16005 ( .A(n16170), .B(n16654), .Z(n16172) );
  XNOR U16006 ( .A(q[5]), .B(DB[75]), .Z(n16654) );
  XNOR U16007 ( .A(q[4]), .B(DB[74]), .Z(n16170) );
  IV U16008 ( .A(n16184), .Z(n16652) );
  XOR U16009 ( .A(n16655), .B(n16656), .Z(n16184) );
  XNOR U16010 ( .A(n16180), .B(n16182), .Z(n16656) );
  XNOR U16011 ( .A(q[0]), .B(DB[70]), .Z(n16182) );
  XNOR U16012 ( .A(q[3]), .B(DB[73]), .Z(n16180) );
  IV U16013 ( .A(n16179), .Z(n16655) );
  XNOR U16014 ( .A(n16177), .B(n16657), .Z(n16179) );
  XNOR U16015 ( .A(q[2]), .B(DB[72]), .Z(n16657) );
  XNOR U16016 ( .A(q[1]), .B(DB[71]), .Z(n16177) );
  XOR U16017 ( .A(n16658), .B(n16142), .Z(n16105) );
  XOR U16018 ( .A(n16659), .B(n16130), .Z(n16142) );
  XNOR U16019 ( .A(q[6]), .B(DB[83]), .Z(n16130) );
  IV U16020 ( .A(n16129), .Z(n16659) );
  XNOR U16021 ( .A(n16127), .B(n16660), .Z(n16129) );
  XNOR U16022 ( .A(q[5]), .B(DB[82]), .Z(n16660) );
  XNOR U16023 ( .A(q[4]), .B(DB[81]), .Z(n16127) );
  IV U16024 ( .A(n16141), .Z(n16658) );
  XOR U16025 ( .A(n16661), .B(n16662), .Z(n16141) );
  XNOR U16026 ( .A(n16137), .B(n16139), .Z(n16662) );
  XNOR U16027 ( .A(q[0]), .B(DB[77]), .Z(n16139) );
  XNOR U16028 ( .A(q[3]), .B(DB[80]), .Z(n16137) );
  IV U16029 ( .A(n16136), .Z(n16661) );
  XNOR U16030 ( .A(n16134), .B(n16663), .Z(n16136) );
  XNOR U16031 ( .A(q[2]), .B(DB[79]), .Z(n16663) );
  XNOR U16032 ( .A(q[1]), .B(DB[78]), .Z(n16134) );
  XOR U16033 ( .A(n16664), .B(n16099), .Z(n16062) );
  XOR U16034 ( .A(n16665), .B(n16087), .Z(n16099) );
  XNOR U16035 ( .A(q[6]), .B(DB[90]), .Z(n16087) );
  IV U16036 ( .A(n16086), .Z(n16665) );
  XNOR U16037 ( .A(n16084), .B(n16666), .Z(n16086) );
  XNOR U16038 ( .A(q[5]), .B(DB[89]), .Z(n16666) );
  XNOR U16039 ( .A(q[4]), .B(DB[88]), .Z(n16084) );
  IV U16040 ( .A(n16098), .Z(n16664) );
  XOR U16041 ( .A(n16667), .B(n16668), .Z(n16098) );
  XNOR U16042 ( .A(n16094), .B(n16096), .Z(n16668) );
  XNOR U16043 ( .A(q[0]), .B(DB[84]), .Z(n16096) );
  XNOR U16044 ( .A(q[3]), .B(DB[87]), .Z(n16094) );
  IV U16045 ( .A(n16093), .Z(n16667) );
  XNOR U16046 ( .A(n16091), .B(n16669), .Z(n16093) );
  XNOR U16047 ( .A(q[2]), .B(DB[86]), .Z(n16669) );
  XNOR U16048 ( .A(q[1]), .B(DB[85]), .Z(n16091) );
  XOR U16049 ( .A(n16670), .B(n16056), .Z(n16019) );
  XOR U16050 ( .A(n16671), .B(n16044), .Z(n16056) );
  XNOR U16051 ( .A(q[6]), .B(DB[97]), .Z(n16044) );
  IV U16052 ( .A(n16043), .Z(n16671) );
  XNOR U16053 ( .A(n16041), .B(n16672), .Z(n16043) );
  XNOR U16054 ( .A(q[5]), .B(DB[96]), .Z(n16672) );
  XNOR U16055 ( .A(q[4]), .B(DB[95]), .Z(n16041) );
  IV U16056 ( .A(n16055), .Z(n16670) );
  XOR U16057 ( .A(n16673), .B(n16674), .Z(n16055) );
  XNOR U16058 ( .A(n16051), .B(n16053), .Z(n16674) );
  XNOR U16059 ( .A(q[0]), .B(DB[91]), .Z(n16053) );
  XNOR U16060 ( .A(q[3]), .B(DB[94]), .Z(n16051) );
  IV U16061 ( .A(n16050), .Z(n16673) );
  XNOR U16062 ( .A(n16048), .B(n16675), .Z(n16050) );
  XNOR U16063 ( .A(q[2]), .B(DB[93]), .Z(n16675) );
  XNOR U16064 ( .A(q[1]), .B(DB[92]), .Z(n16048) );
  XOR U16065 ( .A(n16676), .B(n16013), .Z(n15976) );
  XOR U16066 ( .A(n16677), .B(n16001), .Z(n16013) );
  XNOR U16067 ( .A(q[6]), .B(DB[104]), .Z(n16001) );
  IV U16068 ( .A(n16000), .Z(n16677) );
  XNOR U16069 ( .A(n15998), .B(n16678), .Z(n16000) );
  XNOR U16070 ( .A(q[5]), .B(DB[103]), .Z(n16678) );
  XNOR U16071 ( .A(q[4]), .B(DB[102]), .Z(n15998) );
  IV U16072 ( .A(n16012), .Z(n16676) );
  XOR U16073 ( .A(n16679), .B(n16680), .Z(n16012) );
  XNOR U16074 ( .A(n16008), .B(n16010), .Z(n16680) );
  XNOR U16075 ( .A(q[0]), .B(DB[98]), .Z(n16010) );
  XNOR U16076 ( .A(q[3]), .B(DB[101]), .Z(n16008) );
  IV U16077 ( .A(n16007), .Z(n16679) );
  XNOR U16078 ( .A(n16005), .B(n16681), .Z(n16007) );
  XNOR U16079 ( .A(q[2]), .B(DB[100]), .Z(n16681) );
  XNOR U16080 ( .A(q[1]), .B(DB[99]), .Z(n16005) );
  XOR U16081 ( .A(n16682), .B(n15970), .Z(n15933) );
  XOR U16082 ( .A(n16683), .B(n15958), .Z(n15970) );
  XNOR U16083 ( .A(q[6]), .B(DB[111]), .Z(n15958) );
  IV U16084 ( .A(n15957), .Z(n16683) );
  XNOR U16085 ( .A(n15955), .B(n16684), .Z(n15957) );
  XNOR U16086 ( .A(q[5]), .B(DB[110]), .Z(n16684) );
  XNOR U16087 ( .A(q[4]), .B(DB[109]), .Z(n15955) );
  IV U16088 ( .A(n15969), .Z(n16682) );
  XOR U16089 ( .A(n16685), .B(n16686), .Z(n15969) );
  XNOR U16090 ( .A(n15965), .B(n15967), .Z(n16686) );
  XNOR U16091 ( .A(q[0]), .B(DB[105]), .Z(n15967) );
  XNOR U16092 ( .A(q[3]), .B(DB[108]), .Z(n15965) );
  IV U16093 ( .A(n15964), .Z(n16685) );
  XNOR U16094 ( .A(n15962), .B(n16687), .Z(n15964) );
  XNOR U16095 ( .A(q[2]), .B(DB[107]), .Z(n16687) );
  XNOR U16096 ( .A(q[1]), .B(DB[106]), .Z(n15962) );
  XOR U16097 ( .A(n16688), .B(n15927), .Z(n15890) );
  XOR U16098 ( .A(n16689), .B(n15915), .Z(n15927) );
  XNOR U16099 ( .A(q[6]), .B(DB[118]), .Z(n15915) );
  IV U16100 ( .A(n15914), .Z(n16689) );
  XNOR U16101 ( .A(n15912), .B(n16690), .Z(n15914) );
  XNOR U16102 ( .A(q[5]), .B(DB[117]), .Z(n16690) );
  XNOR U16103 ( .A(q[4]), .B(DB[116]), .Z(n15912) );
  IV U16104 ( .A(n15926), .Z(n16688) );
  XOR U16105 ( .A(n16691), .B(n16692), .Z(n15926) );
  XNOR U16106 ( .A(n15922), .B(n15924), .Z(n16692) );
  XNOR U16107 ( .A(q[0]), .B(DB[112]), .Z(n15924) );
  XNOR U16108 ( .A(q[3]), .B(DB[115]), .Z(n15922) );
  IV U16109 ( .A(n15921), .Z(n16691) );
  XNOR U16110 ( .A(n15919), .B(n16693), .Z(n15921) );
  XNOR U16111 ( .A(q[2]), .B(DB[114]), .Z(n16693) );
  XNOR U16112 ( .A(q[1]), .B(DB[113]), .Z(n15919) );
  XOR U16113 ( .A(n16694), .B(n15884), .Z(n15847) );
  XOR U16114 ( .A(n16695), .B(n15872), .Z(n15884) );
  XNOR U16115 ( .A(q[6]), .B(DB[125]), .Z(n15872) );
  IV U16116 ( .A(n15871), .Z(n16695) );
  XNOR U16117 ( .A(n15869), .B(n16696), .Z(n15871) );
  XNOR U16118 ( .A(q[5]), .B(DB[124]), .Z(n16696) );
  XNOR U16119 ( .A(q[4]), .B(DB[123]), .Z(n15869) );
  IV U16120 ( .A(n15883), .Z(n16694) );
  XOR U16121 ( .A(n16697), .B(n16698), .Z(n15883) );
  XNOR U16122 ( .A(n15879), .B(n15881), .Z(n16698) );
  XNOR U16123 ( .A(q[0]), .B(DB[119]), .Z(n15881) );
  XNOR U16124 ( .A(q[3]), .B(DB[122]), .Z(n15879) );
  IV U16125 ( .A(n15878), .Z(n16697) );
  XNOR U16126 ( .A(n15876), .B(n16699), .Z(n15878) );
  XNOR U16127 ( .A(q[2]), .B(DB[121]), .Z(n16699) );
  XNOR U16128 ( .A(q[1]), .B(DB[120]), .Z(n15876) );
  XOR U16129 ( .A(n16700), .B(n15841), .Z(n15804) );
  XOR U16130 ( .A(n16701), .B(n15829), .Z(n15841) );
  XNOR U16131 ( .A(q[6]), .B(DB[132]), .Z(n15829) );
  IV U16132 ( .A(n15828), .Z(n16701) );
  XNOR U16133 ( .A(n15826), .B(n16702), .Z(n15828) );
  XNOR U16134 ( .A(q[5]), .B(DB[131]), .Z(n16702) );
  XNOR U16135 ( .A(q[4]), .B(DB[130]), .Z(n15826) );
  IV U16136 ( .A(n15840), .Z(n16700) );
  XOR U16137 ( .A(n16703), .B(n16704), .Z(n15840) );
  XNOR U16138 ( .A(n15836), .B(n15838), .Z(n16704) );
  XNOR U16139 ( .A(q[0]), .B(DB[126]), .Z(n15838) );
  XNOR U16140 ( .A(q[3]), .B(DB[129]), .Z(n15836) );
  IV U16141 ( .A(n15835), .Z(n16703) );
  XNOR U16142 ( .A(n15833), .B(n16705), .Z(n15835) );
  XNOR U16143 ( .A(q[2]), .B(DB[128]), .Z(n16705) );
  XNOR U16144 ( .A(q[1]), .B(DB[127]), .Z(n15833) );
  XOR U16145 ( .A(n16706), .B(n15798), .Z(n15761) );
  XOR U16146 ( .A(n16707), .B(n15786), .Z(n15798) );
  XNOR U16147 ( .A(q[6]), .B(DB[139]), .Z(n15786) );
  IV U16148 ( .A(n15785), .Z(n16707) );
  XNOR U16149 ( .A(n15783), .B(n16708), .Z(n15785) );
  XNOR U16150 ( .A(q[5]), .B(DB[138]), .Z(n16708) );
  XNOR U16151 ( .A(q[4]), .B(DB[137]), .Z(n15783) );
  IV U16152 ( .A(n15797), .Z(n16706) );
  XOR U16153 ( .A(n16709), .B(n16710), .Z(n15797) );
  XNOR U16154 ( .A(n15793), .B(n15795), .Z(n16710) );
  XNOR U16155 ( .A(q[0]), .B(DB[133]), .Z(n15795) );
  XNOR U16156 ( .A(q[3]), .B(DB[136]), .Z(n15793) );
  IV U16157 ( .A(n15792), .Z(n16709) );
  XNOR U16158 ( .A(n15790), .B(n16711), .Z(n15792) );
  XNOR U16159 ( .A(q[2]), .B(DB[135]), .Z(n16711) );
  XNOR U16160 ( .A(q[1]), .B(DB[134]), .Z(n15790) );
  XOR U16161 ( .A(n16712), .B(n15755), .Z(n15718) );
  XOR U16162 ( .A(n16713), .B(n15743), .Z(n15755) );
  XNOR U16163 ( .A(q[6]), .B(DB[146]), .Z(n15743) );
  IV U16164 ( .A(n15742), .Z(n16713) );
  XNOR U16165 ( .A(n15740), .B(n16714), .Z(n15742) );
  XNOR U16166 ( .A(q[5]), .B(DB[145]), .Z(n16714) );
  XNOR U16167 ( .A(q[4]), .B(DB[144]), .Z(n15740) );
  IV U16168 ( .A(n15754), .Z(n16712) );
  XOR U16169 ( .A(n16715), .B(n16716), .Z(n15754) );
  XNOR U16170 ( .A(n15750), .B(n15752), .Z(n16716) );
  XNOR U16171 ( .A(q[0]), .B(DB[140]), .Z(n15752) );
  XNOR U16172 ( .A(q[3]), .B(DB[143]), .Z(n15750) );
  IV U16173 ( .A(n15749), .Z(n16715) );
  XNOR U16174 ( .A(n15747), .B(n16717), .Z(n15749) );
  XNOR U16175 ( .A(q[2]), .B(DB[142]), .Z(n16717) );
  XNOR U16176 ( .A(q[1]), .B(DB[141]), .Z(n15747) );
  XOR U16177 ( .A(n16718), .B(n15712), .Z(n15675) );
  XOR U16178 ( .A(n16719), .B(n15700), .Z(n15712) );
  XNOR U16179 ( .A(q[6]), .B(DB[153]), .Z(n15700) );
  IV U16180 ( .A(n15699), .Z(n16719) );
  XNOR U16181 ( .A(n15697), .B(n16720), .Z(n15699) );
  XNOR U16182 ( .A(q[5]), .B(DB[152]), .Z(n16720) );
  XNOR U16183 ( .A(q[4]), .B(DB[151]), .Z(n15697) );
  IV U16184 ( .A(n15711), .Z(n16718) );
  XOR U16185 ( .A(n16721), .B(n16722), .Z(n15711) );
  XNOR U16186 ( .A(n15707), .B(n15709), .Z(n16722) );
  XNOR U16187 ( .A(q[0]), .B(DB[147]), .Z(n15709) );
  XNOR U16188 ( .A(q[3]), .B(DB[150]), .Z(n15707) );
  IV U16189 ( .A(n15706), .Z(n16721) );
  XNOR U16190 ( .A(n15704), .B(n16723), .Z(n15706) );
  XNOR U16191 ( .A(q[2]), .B(DB[149]), .Z(n16723) );
  XNOR U16192 ( .A(q[1]), .B(DB[148]), .Z(n15704) );
  XOR U16193 ( .A(n16724), .B(n15669), .Z(n15632) );
  XOR U16194 ( .A(n16725), .B(n15657), .Z(n15669) );
  XNOR U16195 ( .A(q[6]), .B(DB[160]), .Z(n15657) );
  IV U16196 ( .A(n15656), .Z(n16725) );
  XNOR U16197 ( .A(n15654), .B(n16726), .Z(n15656) );
  XNOR U16198 ( .A(q[5]), .B(DB[159]), .Z(n16726) );
  XNOR U16199 ( .A(q[4]), .B(DB[158]), .Z(n15654) );
  IV U16200 ( .A(n15668), .Z(n16724) );
  XOR U16201 ( .A(n16727), .B(n16728), .Z(n15668) );
  XNOR U16202 ( .A(n15664), .B(n15666), .Z(n16728) );
  XNOR U16203 ( .A(q[0]), .B(DB[154]), .Z(n15666) );
  XNOR U16204 ( .A(q[3]), .B(DB[157]), .Z(n15664) );
  IV U16205 ( .A(n15663), .Z(n16727) );
  XNOR U16206 ( .A(n15661), .B(n16729), .Z(n15663) );
  XNOR U16207 ( .A(q[2]), .B(DB[156]), .Z(n16729) );
  XNOR U16208 ( .A(q[1]), .B(DB[155]), .Z(n15661) );
  XOR U16209 ( .A(n16730), .B(n15626), .Z(n15589) );
  XOR U16210 ( .A(n16731), .B(n15614), .Z(n15626) );
  XNOR U16211 ( .A(q[6]), .B(DB[167]), .Z(n15614) );
  IV U16212 ( .A(n15613), .Z(n16731) );
  XNOR U16213 ( .A(n15611), .B(n16732), .Z(n15613) );
  XNOR U16214 ( .A(q[5]), .B(DB[166]), .Z(n16732) );
  XNOR U16215 ( .A(q[4]), .B(DB[165]), .Z(n15611) );
  IV U16216 ( .A(n15625), .Z(n16730) );
  XOR U16217 ( .A(n16733), .B(n16734), .Z(n15625) );
  XNOR U16218 ( .A(n15621), .B(n15623), .Z(n16734) );
  XNOR U16219 ( .A(q[0]), .B(DB[161]), .Z(n15623) );
  XNOR U16220 ( .A(q[3]), .B(DB[164]), .Z(n15621) );
  IV U16221 ( .A(n15620), .Z(n16733) );
  XNOR U16222 ( .A(n15618), .B(n16735), .Z(n15620) );
  XNOR U16223 ( .A(q[2]), .B(DB[163]), .Z(n16735) );
  XNOR U16224 ( .A(q[1]), .B(DB[162]), .Z(n15618) );
  XOR U16225 ( .A(n16736), .B(n15583), .Z(n15546) );
  XOR U16226 ( .A(n16737), .B(n15571), .Z(n15583) );
  XNOR U16227 ( .A(q[6]), .B(DB[174]), .Z(n15571) );
  IV U16228 ( .A(n15570), .Z(n16737) );
  XNOR U16229 ( .A(n15568), .B(n16738), .Z(n15570) );
  XNOR U16230 ( .A(q[5]), .B(DB[173]), .Z(n16738) );
  XNOR U16231 ( .A(q[4]), .B(DB[172]), .Z(n15568) );
  IV U16232 ( .A(n15582), .Z(n16736) );
  XOR U16233 ( .A(n16739), .B(n16740), .Z(n15582) );
  XNOR U16234 ( .A(n15578), .B(n15580), .Z(n16740) );
  XNOR U16235 ( .A(q[0]), .B(DB[168]), .Z(n15580) );
  XNOR U16236 ( .A(q[3]), .B(DB[171]), .Z(n15578) );
  IV U16237 ( .A(n15577), .Z(n16739) );
  XNOR U16238 ( .A(n15575), .B(n16741), .Z(n15577) );
  XNOR U16239 ( .A(q[2]), .B(DB[170]), .Z(n16741) );
  XNOR U16240 ( .A(q[1]), .B(DB[169]), .Z(n15575) );
  XOR U16241 ( .A(n16742), .B(n15540), .Z(n15503) );
  XOR U16242 ( .A(n16743), .B(n15528), .Z(n15540) );
  XNOR U16243 ( .A(q[6]), .B(DB[181]), .Z(n15528) );
  IV U16244 ( .A(n15527), .Z(n16743) );
  XNOR U16245 ( .A(n15525), .B(n16744), .Z(n15527) );
  XNOR U16246 ( .A(q[5]), .B(DB[180]), .Z(n16744) );
  XNOR U16247 ( .A(q[4]), .B(DB[179]), .Z(n15525) );
  IV U16248 ( .A(n15539), .Z(n16742) );
  XOR U16249 ( .A(n16745), .B(n16746), .Z(n15539) );
  XNOR U16250 ( .A(n15535), .B(n15537), .Z(n16746) );
  XNOR U16251 ( .A(q[0]), .B(DB[175]), .Z(n15537) );
  XNOR U16252 ( .A(q[3]), .B(DB[178]), .Z(n15535) );
  IV U16253 ( .A(n15534), .Z(n16745) );
  XNOR U16254 ( .A(n15532), .B(n16747), .Z(n15534) );
  XNOR U16255 ( .A(q[2]), .B(DB[177]), .Z(n16747) );
  XNOR U16256 ( .A(q[1]), .B(DB[176]), .Z(n15532) );
  XOR U16257 ( .A(n16748), .B(n15497), .Z(n15460) );
  XOR U16258 ( .A(n16749), .B(n15485), .Z(n15497) );
  XNOR U16259 ( .A(q[6]), .B(DB[188]), .Z(n15485) );
  IV U16260 ( .A(n15484), .Z(n16749) );
  XNOR U16261 ( .A(n15482), .B(n16750), .Z(n15484) );
  XNOR U16262 ( .A(q[5]), .B(DB[187]), .Z(n16750) );
  XNOR U16263 ( .A(q[4]), .B(DB[186]), .Z(n15482) );
  IV U16264 ( .A(n15496), .Z(n16748) );
  XOR U16265 ( .A(n16751), .B(n16752), .Z(n15496) );
  XNOR U16266 ( .A(n15492), .B(n15494), .Z(n16752) );
  XNOR U16267 ( .A(q[0]), .B(DB[182]), .Z(n15494) );
  XNOR U16268 ( .A(q[3]), .B(DB[185]), .Z(n15492) );
  IV U16269 ( .A(n15491), .Z(n16751) );
  XNOR U16270 ( .A(n15489), .B(n16753), .Z(n15491) );
  XNOR U16271 ( .A(q[2]), .B(DB[184]), .Z(n16753) );
  XNOR U16272 ( .A(q[1]), .B(DB[183]), .Z(n15489) );
  XOR U16273 ( .A(n16754), .B(n15454), .Z(n15417) );
  XOR U16274 ( .A(n16755), .B(n15442), .Z(n15454) );
  XNOR U16275 ( .A(q[6]), .B(DB[195]), .Z(n15442) );
  IV U16276 ( .A(n15441), .Z(n16755) );
  XNOR U16277 ( .A(n15439), .B(n16756), .Z(n15441) );
  XNOR U16278 ( .A(q[5]), .B(DB[194]), .Z(n16756) );
  XNOR U16279 ( .A(q[4]), .B(DB[193]), .Z(n15439) );
  IV U16280 ( .A(n15453), .Z(n16754) );
  XOR U16281 ( .A(n16757), .B(n16758), .Z(n15453) );
  XNOR U16282 ( .A(n15449), .B(n15451), .Z(n16758) );
  XNOR U16283 ( .A(q[0]), .B(DB[189]), .Z(n15451) );
  XNOR U16284 ( .A(q[3]), .B(DB[192]), .Z(n15449) );
  IV U16285 ( .A(n15448), .Z(n16757) );
  XNOR U16286 ( .A(n15446), .B(n16759), .Z(n15448) );
  XNOR U16287 ( .A(q[2]), .B(DB[191]), .Z(n16759) );
  XNOR U16288 ( .A(q[1]), .B(DB[190]), .Z(n15446) );
  XOR U16289 ( .A(n16760), .B(n15411), .Z(n15374) );
  XOR U16290 ( .A(n16761), .B(n15399), .Z(n15411) );
  XNOR U16291 ( .A(q[6]), .B(DB[202]), .Z(n15399) );
  IV U16292 ( .A(n15398), .Z(n16761) );
  XNOR U16293 ( .A(n15396), .B(n16762), .Z(n15398) );
  XNOR U16294 ( .A(q[5]), .B(DB[201]), .Z(n16762) );
  XNOR U16295 ( .A(q[4]), .B(DB[200]), .Z(n15396) );
  IV U16296 ( .A(n15410), .Z(n16760) );
  XOR U16297 ( .A(n16763), .B(n16764), .Z(n15410) );
  XNOR U16298 ( .A(n15406), .B(n15408), .Z(n16764) );
  XNOR U16299 ( .A(q[0]), .B(DB[196]), .Z(n15408) );
  XNOR U16300 ( .A(q[3]), .B(DB[199]), .Z(n15406) );
  IV U16301 ( .A(n15405), .Z(n16763) );
  XNOR U16302 ( .A(n15403), .B(n16765), .Z(n15405) );
  XNOR U16303 ( .A(q[2]), .B(DB[198]), .Z(n16765) );
  XNOR U16304 ( .A(q[1]), .B(DB[197]), .Z(n15403) );
  XOR U16305 ( .A(n16766), .B(n15368), .Z(n15331) );
  XOR U16306 ( .A(n16767), .B(n15356), .Z(n15368) );
  XNOR U16307 ( .A(q[6]), .B(DB[209]), .Z(n15356) );
  IV U16308 ( .A(n15355), .Z(n16767) );
  XNOR U16309 ( .A(n15353), .B(n16768), .Z(n15355) );
  XNOR U16310 ( .A(q[5]), .B(DB[208]), .Z(n16768) );
  XNOR U16311 ( .A(q[4]), .B(DB[207]), .Z(n15353) );
  IV U16312 ( .A(n15367), .Z(n16766) );
  XOR U16313 ( .A(n16769), .B(n16770), .Z(n15367) );
  XNOR U16314 ( .A(n15363), .B(n15365), .Z(n16770) );
  XNOR U16315 ( .A(q[0]), .B(DB[203]), .Z(n15365) );
  XNOR U16316 ( .A(q[3]), .B(DB[206]), .Z(n15363) );
  IV U16317 ( .A(n15362), .Z(n16769) );
  XNOR U16318 ( .A(n15360), .B(n16771), .Z(n15362) );
  XNOR U16319 ( .A(q[2]), .B(DB[205]), .Z(n16771) );
  XNOR U16320 ( .A(q[1]), .B(DB[204]), .Z(n15360) );
  XOR U16321 ( .A(n16772), .B(n15325), .Z(n15288) );
  XOR U16322 ( .A(n16773), .B(n15313), .Z(n15325) );
  XNOR U16323 ( .A(q[6]), .B(DB[216]), .Z(n15313) );
  IV U16324 ( .A(n15312), .Z(n16773) );
  XNOR U16325 ( .A(n15310), .B(n16774), .Z(n15312) );
  XNOR U16326 ( .A(q[5]), .B(DB[215]), .Z(n16774) );
  XNOR U16327 ( .A(q[4]), .B(DB[214]), .Z(n15310) );
  IV U16328 ( .A(n15324), .Z(n16772) );
  XOR U16329 ( .A(n16775), .B(n16776), .Z(n15324) );
  XNOR U16330 ( .A(n15320), .B(n15322), .Z(n16776) );
  XNOR U16331 ( .A(q[0]), .B(DB[210]), .Z(n15322) );
  XNOR U16332 ( .A(q[3]), .B(DB[213]), .Z(n15320) );
  IV U16333 ( .A(n15319), .Z(n16775) );
  XNOR U16334 ( .A(n15317), .B(n16777), .Z(n15319) );
  XNOR U16335 ( .A(q[2]), .B(DB[212]), .Z(n16777) );
  XNOR U16336 ( .A(q[1]), .B(DB[211]), .Z(n15317) );
  XOR U16337 ( .A(n16778), .B(n15282), .Z(n15245) );
  XOR U16338 ( .A(n16779), .B(n15270), .Z(n15282) );
  XNOR U16339 ( .A(q[6]), .B(DB[223]), .Z(n15270) );
  IV U16340 ( .A(n15269), .Z(n16779) );
  XNOR U16341 ( .A(n15267), .B(n16780), .Z(n15269) );
  XNOR U16342 ( .A(q[5]), .B(DB[222]), .Z(n16780) );
  XNOR U16343 ( .A(q[4]), .B(DB[221]), .Z(n15267) );
  IV U16344 ( .A(n15281), .Z(n16778) );
  XOR U16345 ( .A(n16781), .B(n16782), .Z(n15281) );
  XNOR U16346 ( .A(n15277), .B(n15279), .Z(n16782) );
  XNOR U16347 ( .A(q[0]), .B(DB[217]), .Z(n15279) );
  XNOR U16348 ( .A(q[3]), .B(DB[220]), .Z(n15277) );
  IV U16349 ( .A(n15276), .Z(n16781) );
  XNOR U16350 ( .A(n15274), .B(n16783), .Z(n15276) );
  XNOR U16351 ( .A(q[2]), .B(DB[219]), .Z(n16783) );
  XNOR U16352 ( .A(q[1]), .B(DB[218]), .Z(n15274) );
  XOR U16353 ( .A(n16784), .B(n15239), .Z(n15202) );
  XOR U16354 ( .A(n16785), .B(n15227), .Z(n15239) );
  XNOR U16355 ( .A(q[6]), .B(DB[230]), .Z(n15227) );
  IV U16356 ( .A(n15226), .Z(n16785) );
  XNOR U16357 ( .A(n15224), .B(n16786), .Z(n15226) );
  XNOR U16358 ( .A(q[5]), .B(DB[229]), .Z(n16786) );
  XNOR U16359 ( .A(q[4]), .B(DB[228]), .Z(n15224) );
  IV U16360 ( .A(n15238), .Z(n16784) );
  XOR U16361 ( .A(n16787), .B(n16788), .Z(n15238) );
  XNOR U16362 ( .A(n15234), .B(n15236), .Z(n16788) );
  XNOR U16363 ( .A(q[0]), .B(DB[224]), .Z(n15236) );
  XNOR U16364 ( .A(q[3]), .B(DB[227]), .Z(n15234) );
  IV U16365 ( .A(n15233), .Z(n16787) );
  XNOR U16366 ( .A(n15231), .B(n16789), .Z(n15233) );
  XNOR U16367 ( .A(q[2]), .B(DB[226]), .Z(n16789) );
  XNOR U16368 ( .A(q[1]), .B(DB[225]), .Z(n15231) );
  XOR U16369 ( .A(n16790), .B(n15196), .Z(n15159) );
  XOR U16370 ( .A(n16791), .B(n15184), .Z(n15196) );
  XNOR U16371 ( .A(q[6]), .B(DB[237]), .Z(n15184) );
  IV U16372 ( .A(n15183), .Z(n16791) );
  XNOR U16373 ( .A(n15181), .B(n16792), .Z(n15183) );
  XNOR U16374 ( .A(q[5]), .B(DB[236]), .Z(n16792) );
  XNOR U16375 ( .A(q[4]), .B(DB[235]), .Z(n15181) );
  IV U16376 ( .A(n15195), .Z(n16790) );
  XOR U16377 ( .A(n16793), .B(n16794), .Z(n15195) );
  XNOR U16378 ( .A(n15191), .B(n15193), .Z(n16794) );
  XNOR U16379 ( .A(q[0]), .B(DB[231]), .Z(n15193) );
  XNOR U16380 ( .A(q[3]), .B(DB[234]), .Z(n15191) );
  IV U16381 ( .A(n15190), .Z(n16793) );
  XNOR U16382 ( .A(n15188), .B(n16795), .Z(n15190) );
  XNOR U16383 ( .A(q[2]), .B(DB[233]), .Z(n16795) );
  XNOR U16384 ( .A(q[1]), .B(DB[232]), .Z(n15188) );
  XOR U16385 ( .A(n16796), .B(n15153), .Z(n15116) );
  XOR U16386 ( .A(n16797), .B(n15141), .Z(n15153) );
  XNOR U16387 ( .A(q[6]), .B(DB[244]), .Z(n15141) );
  IV U16388 ( .A(n15140), .Z(n16797) );
  XNOR U16389 ( .A(n15138), .B(n16798), .Z(n15140) );
  XNOR U16390 ( .A(q[5]), .B(DB[243]), .Z(n16798) );
  XNOR U16391 ( .A(q[4]), .B(DB[242]), .Z(n15138) );
  IV U16392 ( .A(n15152), .Z(n16796) );
  XOR U16393 ( .A(n16799), .B(n16800), .Z(n15152) );
  XNOR U16394 ( .A(n15148), .B(n15150), .Z(n16800) );
  XNOR U16395 ( .A(q[0]), .B(DB[238]), .Z(n15150) );
  XNOR U16396 ( .A(q[3]), .B(DB[241]), .Z(n15148) );
  IV U16397 ( .A(n15147), .Z(n16799) );
  XNOR U16398 ( .A(n15145), .B(n16801), .Z(n15147) );
  XNOR U16399 ( .A(q[2]), .B(DB[240]), .Z(n16801) );
  XNOR U16400 ( .A(q[1]), .B(DB[239]), .Z(n15145) );
  XOR U16401 ( .A(n16802), .B(n15110), .Z(n15073) );
  XOR U16402 ( .A(n16803), .B(n15098), .Z(n15110) );
  XNOR U16403 ( .A(q[6]), .B(DB[251]), .Z(n15098) );
  IV U16404 ( .A(n15097), .Z(n16803) );
  XNOR U16405 ( .A(n15095), .B(n16804), .Z(n15097) );
  XNOR U16406 ( .A(q[5]), .B(DB[250]), .Z(n16804) );
  XNOR U16407 ( .A(q[4]), .B(DB[249]), .Z(n15095) );
  IV U16408 ( .A(n15109), .Z(n16802) );
  XOR U16409 ( .A(n16805), .B(n16806), .Z(n15109) );
  XNOR U16410 ( .A(n15105), .B(n15107), .Z(n16806) );
  XNOR U16411 ( .A(q[0]), .B(DB[245]), .Z(n15107) );
  XNOR U16412 ( .A(q[3]), .B(DB[248]), .Z(n15105) );
  IV U16413 ( .A(n15104), .Z(n16805) );
  XNOR U16414 ( .A(n15102), .B(n16807), .Z(n15104) );
  XNOR U16415 ( .A(q[2]), .B(DB[247]), .Z(n16807) );
  XNOR U16416 ( .A(q[1]), .B(DB[246]), .Z(n15102) );
  XOR U16417 ( .A(n16808), .B(n15067), .Z(n15030) );
  XOR U16418 ( .A(n16809), .B(n15055), .Z(n15067) );
  XNOR U16419 ( .A(q[6]), .B(DB[258]), .Z(n15055) );
  IV U16420 ( .A(n15054), .Z(n16809) );
  XNOR U16421 ( .A(n15052), .B(n16810), .Z(n15054) );
  XNOR U16422 ( .A(q[5]), .B(DB[257]), .Z(n16810) );
  XNOR U16423 ( .A(q[4]), .B(DB[256]), .Z(n15052) );
  IV U16424 ( .A(n15066), .Z(n16808) );
  XOR U16425 ( .A(n16811), .B(n16812), .Z(n15066) );
  XNOR U16426 ( .A(n15062), .B(n15064), .Z(n16812) );
  XNOR U16427 ( .A(q[0]), .B(DB[252]), .Z(n15064) );
  XNOR U16428 ( .A(q[3]), .B(DB[255]), .Z(n15062) );
  IV U16429 ( .A(n15061), .Z(n16811) );
  XNOR U16430 ( .A(n15059), .B(n16813), .Z(n15061) );
  XNOR U16431 ( .A(q[2]), .B(DB[254]), .Z(n16813) );
  XNOR U16432 ( .A(q[1]), .B(DB[253]), .Z(n15059) );
  XOR U16433 ( .A(n16814), .B(n15024), .Z(n14987) );
  XOR U16434 ( .A(n16815), .B(n15012), .Z(n15024) );
  XNOR U16435 ( .A(q[6]), .B(DB[265]), .Z(n15012) );
  IV U16436 ( .A(n15011), .Z(n16815) );
  XNOR U16437 ( .A(n15009), .B(n16816), .Z(n15011) );
  XNOR U16438 ( .A(q[5]), .B(DB[264]), .Z(n16816) );
  XNOR U16439 ( .A(q[4]), .B(DB[263]), .Z(n15009) );
  IV U16440 ( .A(n15023), .Z(n16814) );
  XOR U16441 ( .A(n16817), .B(n16818), .Z(n15023) );
  XNOR U16442 ( .A(n15019), .B(n15021), .Z(n16818) );
  XNOR U16443 ( .A(q[0]), .B(DB[259]), .Z(n15021) );
  XNOR U16444 ( .A(q[3]), .B(DB[262]), .Z(n15019) );
  IV U16445 ( .A(n15018), .Z(n16817) );
  XNOR U16446 ( .A(n15016), .B(n16819), .Z(n15018) );
  XNOR U16447 ( .A(q[2]), .B(DB[261]), .Z(n16819) );
  XNOR U16448 ( .A(q[1]), .B(DB[260]), .Z(n15016) );
  XOR U16449 ( .A(n16820), .B(n14981), .Z(n14944) );
  XOR U16450 ( .A(n16821), .B(n14969), .Z(n14981) );
  XNOR U16451 ( .A(q[6]), .B(DB[272]), .Z(n14969) );
  IV U16452 ( .A(n14968), .Z(n16821) );
  XNOR U16453 ( .A(n14966), .B(n16822), .Z(n14968) );
  XNOR U16454 ( .A(q[5]), .B(DB[271]), .Z(n16822) );
  XNOR U16455 ( .A(q[4]), .B(DB[270]), .Z(n14966) );
  IV U16456 ( .A(n14980), .Z(n16820) );
  XOR U16457 ( .A(n16823), .B(n16824), .Z(n14980) );
  XNOR U16458 ( .A(n14976), .B(n14978), .Z(n16824) );
  XNOR U16459 ( .A(q[0]), .B(DB[266]), .Z(n14978) );
  XNOR U16460 ( .A(q[3]), .B(DB[269]), .Z(n14976) );
  IV U16461 ( .A(n14975), .Z(n16823) );
  XNOR U16462 ( .A(n14973), .B(n16825), .Z(n14975) );
  XNOR U16463 ( .A(q[2]), .B(DB[268]), .Z(n16825) );
  XNOR U16464 ( .A(q[1]), .B(DB[267]), .Z(n14973) );
  XOR U16465 ( .A(n16826), .B(n14938), .Z(n14901) );
  XOR U16466 ( .A(n16827), .B(n14926), .Z(n14938) );
  XNOR U16467 ( .A(q[6]), .B(DB[279]), .Z(n14926) );
  IV U16468 ( .A(n14925), .Z(n16827) );
  XNOR U16469 ( .A(n14923), .B(n16828), .Z(n14925) );
  XNOR U16470 ( .A(q[5]), .B(DB[278]), .Z(n16828) );
  XNOR U16471 ( .A(q[4]), .B(DB[277]), .Z(n14923) );
  IV U16472 ( .A(n14937), .Z(n16826) );
  XOR U16473 ( .A(n16829), .B(n16830), .Z(n14937) );
  XNOR U16474 ( .A(n14933), .B(n14935), .Z(n16830) );
  XNOR U16475 ( .A(q[0]), .B(DB[273]), .Z(n14935) );
  XNOR U16476 ( .A(q[3]), .B(DB[276]), .Z(n14933) );
  IV U16477 ( .A(n14932), .Z(n16829) );
  XNOR U16478 ( .A(n14930), .B(n16831), .Z(n14932) );
  XNOR U16479 ( .A(q[2]), .B(DB[275]), .Z(n16831) );
  XNOR U16480 ( .A(q[1]), .B(DB[274]), .Z(n14930) );
  XOR U16481 ( .A(n16832), .B(n14895), .Z(n14858) );
  XOR U16482 ( .A(n16833), .B(n14883), .Z(n14895) );
  XNOR U16483 ( .A(q[6]), .B(DB[286]), .Z(n14883) );
  IV U16484 ( .A(n14882), .Z(n16833) );
  XNOR U16485 ( .A(n14880), .B(n16834), .Z(n14882) );
  XNOR U16486 ( .A(q[5]), .B(DB[285]), .Z(n16834) );
  XNOR U16487 ( .A(q[4]), .B(DB[284]), .Z(n14880) );
  IV U16488 ( .A(n14894), .Z(n16832) );
  XOR U16489 ( .A(n16835), .B(n16836), .Z(n14894) );
  XNOR U16490 ( .A(n14890), .B(n14892), .Z(n16836) );
  XNOR U16491 ( .A(q[0]), .B(DB[280]), .Z(n14892) );
  XNOR U16492 ( .A(q[3]), .B(DB[283]), .Z(n14890) );
  IV U16493 ( .A(n14889), .Z(n16835) );
  XNOR U16494 ( .A(n14887), .B(n16837), .Z(n14889) );
  XNOR U16495 ( .A(q[2]), .B(DB[282]), .Z(n16837) );
  XNOR U16496 ( .A(q[1]), .B(DB[281]), .Z(n14887) );
  XOR U16497 ( .A(n16838), .B(n14852), .Z(n14815) );
  XOR U16498 ( .A(n16839), .B(n14840), .Z(n14852) );
  XNOR U16499 ( .A(q[6]), .B(DB[293]), .Z(n14840) );
  IV U16500 ( .A(n14839), .Z(n16839) );
  XNOR U16501 ( .A(n14837), .B(n16840), .Z(n14839) );
  XNOR U16502 ( .A(q[5]), .B(DB[292]), .Z(n16840) );
  XNOR U16503 ( .A(q[4]), .B(DB[291]), .Z(n14837) );
  IV U16504 ( .A(n14851), .Z(n16838) );
  XOR U16505 ( .A(n16841), .B(n16842), .Z(n14851) );
  XNOR U16506 ( .A(n14847), .B(n14849), .Z(n16842) );
  XNOR U16507 ( .A(q[0]), .B(DB[287]), .Z(n14849) );
  XNOR U16508 ( .A(q[3]), .B(DB[290]), .Z(n14847) );
  IV U16509 ( .A(n14846), .Z(n16841) );
  XNOR U16510 ( .A(n14844), .B(n16843), .Z(n14846) );
  XNOR U16511 ( .A(q[2]), .B(DB[289]), .Z(n16843) );
  XNOR U16512 ( .A(q[1]), .B(DB[288]), .Z(n14844) );
  XOR U16513 ( .A(n16844), .B(n14809), .Z(n14772) );
  XOR U16514 ( .A(n16845), .B(n14797), .Z(n14809) );
  XNOR U16515 ( .A(q[6]), .B(DB[300]), .Z(n14797) );
  IV U16516 ( .A(n14796), .Z(n16845) );
  XNOR U16517 ( .A(n14794), .B(n16846), .Z(n14796) );
  XNOR U16518 ( .A(q[5]), .B(DB[299]), .Z(n16846) );
  XNOR U16519 ( .A(q[4]), .B(DB[298]), .Z(n14794) );
  IV U16520 ( .A(n14808), .Z(n16844) );
  XOR U16521 ( .A(n16847), .B(n16848), .Z(n14808) );
  XNOR U16522 ( .A(n14804), .B(n14806), .Z(n16848) );
  XNOR U16523 ( .A(q[0]), .B(DB[294]), .Z(n14806) );
  XNOR U16524 ( .A(q[3]), .B(DB[297]), .Z(n14804) );
  IV U16525 ( .A(n14803), .Z(n16847) );
  XNOR U16526 ( .A(n14801), .B(n16849), .Z(n14803) );
  XNOR U16527 ( .A(q[2]), .B(DB[296]), .Z(n16849) );
  XNOR U16528 ( .A(q[1]), .B(DB[295]), .Z(n14801) );
  XOR U16529 ( .A(n16850), .B(n14766), .Z(n14729) );
  XOR U16530 ( .A(n16851), .B(n14754), .Z(n14766) );
  XNOR U16531 ( .A(q[6]), .B(DB[307]), .Z(n14754) );
  IV U16532 ( .A(n14753), .Z(n16851) );
  XNOR U16533 ( .A(n14751), .B(n16852), .Z(n14753) );
  XNOR U16534 ( .A(q[5]), .B(DB[306]), .Z(n16852) );
  XNOR U16535 ( .A(q[4]), .B(DB[305]), .Z(n14751) );
  IV U16536 ( .A(n14765), .Z(n16850) );
  XOR U16537 ( .A(n16853), .B(n16854), .Z(n14765) );
  XNOR U16538 ( .A(n14761), .B(n14763), .Z(n16854) );
  XNOR U16539 ( .A(q[0]), .B(DB[301]), .Z(n14763) );
  XNOR U16540 ( .A(q[3]), .B(DB[304]), .Z(n14761) );
  IV U16541 ( .A(n14760), .Z(n16853) );
  XNOR U16542 ( .A(n14758), .B(n16855), .Z(n14760) );
  XNOR U16543 ( .A(q[2]), .B(DB[303]), .Z(n16855) );
  XNOR U16544 ( .A(q[1]), .B(DB[302]), .Z(n14758) );
  XOR U16545 ( .A(n16856), .B(n14723), .Z(n14686) );
  XOR U16546 ( .A(n16857), .B(n14711), .Z(n14723) );
  XNOR U16547 ( .A(q[6]), .B(DB[314]), .Z(n14711) );
  IV U16548 ( .A(n14710), .Z(n16857) );
  XNOR U16549 ( .A(n14708), .B(n16858), .Z(n14710) );
  XNOR U16550 ( .A(q[5]), .B(DB[313]), .Z(n16858) );
  XNOR U16551 ( .A(q[4]), .B(DB[312]), .Z(n14708) );
  IV U16552 ( .A(n14722), .Z(n16856) );
  XOR U16553 ( .A(n16859), .B(n16860), .Z(n14722) );
  XNOR U16554 ( .A(n14718), .B(n14720), .Z(n16860) );
  XNOR U16555 ( .A(q[0]), .B(DB[308]), .Z(n14720) );
  XNOR U16556 ( .A(q[3]), .B(DB[311]), .Z(n14718) );
  IV U16557 ( .A(n14717), .Z(n16859) );
  XNOR U16558 ( .A(n14715), .B(n16861), .Z(n14717) );
  XNOR U16559 ( .A(q[2]), .B(DB[310]), .Z(n16861) );
  XNOR U16560 ( .A(q[1]), .B(DB[309]), .Z(n14715) );
  XOR U16561 ( .A(n16862), .B(n14680), .Z(n14643) );
  XOR U16562 ( .A(n16863), .B(n14668), .Z(n14680) );
  XNOR U16563 ( .A(q[6]), .B(DB[321]), .Z(n14668) );
  IV U16564 ( .A(n14667), .Z(n16863) );
  XNOR U16565 ( .A(n14665), .B(n16864), .Z(n14667) );
  XNOR U16566 ( .A(q[5]), .B(DB[320]), .Z(n16864) );
  XNOR U16567 ( .A(q[4]), .B(DB[319]), .Z(n14665) );
  IV U16568 ( .A(n14679), .Z(n16862) );
  XOR U16569 ( .A(n16865), .B(n16866), .Z(n14679) );
  XNOR U16570 ( .A(n14675), .B(n14677), .Z(n16866) );
  XNOR U16571 ( .A(q[0]), .B(DB[315]), .Z(n14677) );
  XNOR U16572 ( .A(q[3]), .B(DB[318]), .Z(n14675) );
  IV U16573 ( .A(n14674), .Z(n16865) );
  XNOR U16574 ( .A(n14672), .B(n16867), .Z(n14674) );
  XNOR U16575 ( .A(q[2]), .B(DB[317]), .Z(n16867) );
  XNOR U16576 ( .A(q[1]), .B(DB[316]), .Z(n14672) );
  XOR U16577 ( .A(n16868), .B(n14637), .Z(n14600) );
  XOR U16578 ( .A(n16869), .B(n14625), .Z(n14637) );
  XNOR U16579 ( .A(q[6]), .B(DB[328]), .Z(n14625) );
  IV U16580 ( .A(n14624), .Z(n16869) );
  XNOR U16581 ( .A(n14622), .B(n16870), .Z(n14624) );
  XNOR U16582 ( .A(q[5]), .B(DB[327]), .Z(n16870) );
  XNOR U16583 ( .A(q[4]), .B(DB[326]), .Z(n14622) );
  IV U16584 ( .A(n14636), .Z(n16868) );
  XOR U16585 ( .A(n16871), .B(n16872), .Z(n14636) );
  XNOR U16586 ( .A(n14632), .B(n14634), .Z(n16872) );
  XNOR U16587 ( .A(q[0]), .B(DB[322]), .Z(n14634) );
  XNOR U16588 ( .A(q[3]), .B(DB[325]), .Z(n14632) );
  IV U16589 ( .A(n14631), .Z(n16871) );
  XNOR U16590 ( .A(n14629), .B(n16873), .Z(n14631) );
  XNOR U16591 ( .A(q[2]), .B(DB[324]), .Z(n16873) );
  XNOR U16592 ( .A(q[1]), .B(DB[323]), .Z(n14629) );
  XOR U16593 ( .A(n16874), .B(n14594), .Z(n14557) );
  XOR U16594 ( .A(n16875), .B(n14582), .Z(n14594) );
  XNOR U16595 ( .A(q[6]), .B(DB[335]), .Z(n14582) );
  IV U16596 ( .A(n14581), .Z(n16875) );
  XNOR U16597 ( .A(n14579), .B(n16876), .Z(n14581) );
  XNOR U16598 ( .A(q[5]), .B(DB[334]), .Z(n16876) );
  XNOR U16599 ( .A(q[4]), .B(DB[333]), .Z(n14579) );
  IV U16600 ( .A(n14593), .Z(n16874) );
  XOR U16601 ( .A(n16877), .B(n16878), .Z(n14593) );
  XNOR U16602 ( .A(n14589), .B(n14591), .Z(n16878) );
  XNOR U16603 ( .A(q[0]), .B(DB[329]), .Z(n14591) );
  XNOR U16604 ( .A(q[3]), .B(DB[332]), .Z(n14589) );
  IV U16605 ( .A(n14588), .Z(n16877) );
  XNOR U16606 ( .A(n14586), .B(n16879), .Z(n14588) );
  XNOR U16607 ( .A(q[2]), .B(DB[331]), .Z(n16879) );
  XNOR U16608 ( .A(q[1]), .B(DB[330]), .Z(n14586) );
  XOR U16609 ( .A(n16880), .B(n14551), .Z(n14514) );
  XOR U16610 ( .A(n16881), .B(n14539), .Z(n14551) );
  XNOR U16611 ( .A(q[6]), .B(DB[342]), .Z(n14539) );
  IV U16612 ( .A(n14538), .Z(n16881) );
  XNOR U16613 ( .A(n14536), .B(n16882), .Z(n14538) );
  XNOR U16614 ( .A(q[5]), .B(DB[341]), .Z(n16882) );
  XNOR U16615 ( .A(q[4]), .B(DB[340]), .Z(n14536) );
  IV U16616 ( .A(n14550), .Z(n16880) );
  XOR U16617 ( .A(n16883), .B(n16884), .Z(n14550) );
  XNOR U16618 ( .A(n14546), .B(n14548), .Z(n16884) );
  XNOR U16619 ( .A(q[0]), .B(DB[336]), .Z(n14548) );
  XNOR U16620 ( .A(q[3]), .B(DB[339]), .Z(n14546) );
  IV U16621 ( .A(n14545), .Z(n16883) );
  XNOR U16622 ( .A(n14543), .B(n16885), .Z(n14545) );
  XNOR U16623 ( .A(q[2]), .B(DB[338]), .Z(n16885) );
  XNOR U16624 ( .A(q[1]), .B(DB[337]), .Z(n14543) );
  XOR U16625 ( .A(n16886), .B(n14508), .Z(n14471) );
  XOR U16626 ( .A(n16887), .B(n14496), .Z(n14508) );
  XNOR U16627 ( .A(q[6]), .B(DB[349]), .Z(n14496) );
  IV U16628 ( .A(n14495), .Z(n16887) );
  XNOR U16629 ( .A(n14493), .B(n16888), .Z(n14495) );
  XNOR U16630 ( .A(q[5]), .B(DB[348]), .Z(n16888) );
  XNOR U16631 ( .A(q[4]), .B(DB[347]), .Z(n14493) );
  IV U16632 ( .A(n14507), .Z(n16886) );
  XOR U16633 ( .A(n16889), .B(n16890), .Z(n14507) );
  XNOR U16634 ( .A(n14503), .B(n14505), .Z(n16890) );
  XNOR U16635 ( .A(q[0]), .B(DB[343]), .Z(n14505) );
  XNOR U16636 ( .A(q[3]), .B(DB[346]), .Z(n14503) );
  IV U16637 ( .A(n14502), .Z(n16889) );
  XNOR U16638 ( .A(n14500), .B(n16891), .Z(n14502) );
  XNOR U16639 ( .A(q[2]), .B(DB[345]), .Z(n16891) );
  XNOR U16640 ( .A(q[1]), .B(DB[344]), .Z(n14500) );
  XOR U16641 ( .A(n16892), .B(n14465), .Z(n14428) );
  XOR U16642 ( .A(n16893), .B(n14453), .Z(n14465) );
  XNOR U16643 ( .A(q[6]), .B(DB[356]), .Z(n14453) );
  IV U16644 ( .A(n14452), .Z(n16893) );
  XNOR U16645 ( .A(n14450), .B(n16894), .Z(n14452) );
  XNOR U16646 ( .A(q[5]), .B(DB[355]), .Z(n16894) );
  XNOR U16647 ( .A(q[4]), .B(DB[354]), .Z(n14450) );
  IV U16648 ( .A(n14464), .Z(n16892) );
  XOR U16649 ( .A(n16895), .B(n16896), .Z(n14464) );
  XNOR U16650 ( .A(n14460), .B(n14462), .Z(n16896) );
  XNOR U16651 ( .A(q[0]), .B(DB[350]), .Z(n14462) );
  XNOR U16652 ( .A(q[3]), .B(DB[353]), .Z(n14460) );
  IV U16653 ( .A(n14459), .Z(n16895) );
  XNOR U16654 ( .A(n14457), .B(n16897), .Z(n14459) );
  XNOR U16655 ( .A(q[2]), .B(DB[352]), .Z(n16897) );
  XNOR U16656 ( .A(q[1]), .B(DB[351]), .Z(n14457) );
  XOR U16657 ( .A(n16898), .B(n14422), .Z(n14385) );
  XOR U16658 ( .A(n16899), .B(n14410), .Z(n14422) );
  XNOR U16659 ( .A(q[6]), .B(DB[363]), .Z(n14410) );
  IV U16660 ( .A(n14409), .Z(n16899) );
  XNOR U16661 ( .A(n14407), .B(n16900), .Z(n14409) );
  XNOR U16662 ( .A(q[5]), .B(DB[362]), .Z(n16900) );
  XNOR U16663 ( .A(q[4]), .B(DB[361]), .Z(n14407) );
  IV U16664 ( .A(n14421), .Z(n16898) );
  XOR U16665 ( .A(n16901), .B(n16902), .Z(n14421) );
  XNOR U16666 ( .A(n14417), .B(n14419), .Z(n16902) );
  XNOR U16667 ( .A(q[0]), .B(DB[357]), .Z(n14419) );
  XNOR U16668 ( .A(q[3]), .B(DB[360]), .Z(n14417) );
  IV U16669 ( .A(n14416), .Z(n16901) );
  XNOR U16670 ( .A(n14414), .B(n16903), .Z(n14416) );
  XNOR U16671 ( .A(q[2]), .B(DB[359]), .Z(n16903) );
  XNOR U16672 ( .A(q[1]), .B(DB[358]), .Z(n14414) );
  XOR U16673 ( .A(n16904), .B(n14379), .Z(n14342) );
  XOR U16674 ( .A(n16905), .B(n14367), .Z(n14379) );
  XNOR U16675 ( .A(q[6]), .B(DB[370]), .Z(n14367) );
  IV U16676 ( .A(n14366), .Z(n16905) );
  XNOR U16677 ( .A(n14364), .B(n16906), .Z(n14366) );
  XNOR U16678 ( .A(q[5]), .B(DB[369]), .Z(n16906) );
  XNOR U16679 ( .A(q[4]), .B(DB[368]), .Z(n14364) );
  IV U16680 ( .A(n14378), .Z(n16904) );
  XOR U16681 ( .A(n16907), .B(n16908), .Z(n14378) );
  XNOR U16682 ( .A(n14374), .B(n14376), .Z(n16908) );
  XNOR U16683 ( .A(q[0]), .B(DB[364]), .Z(n14376) );
  XNOR U16684 ( .A(q[3]), .B(DB[367]), .Z(n14374) );
  IV U16685 ( .A(n14373), .Z(n16907) );
  XNOR U16686 ( .A(n14371), .B(n16909), .Z(n14373) );
  XNOR U16687 ( .A(q[2]), .B(DB[366]), .Z(n16909) );
  XNOR U16688 ( .A(q[1]), .B(DB[365]), .Z(n14371) );
  XOR U16689 ( .A(n16910), .B(n14336), .Z(n14299) );
  XOR U16690 ( .A(n16911), .B(n14324), .Z(n14336) );
  XNOR U16691 ( .A(q[6]), .B(DB[377]), .Z(n14324) );
  IV U16692 ( .A(n14323), .Z(n16911) );
  XNOR U16693 ( .A(n14321), .B(n16912), .Z(n14323) );
  XNOR U16694 ( .A(q[5]), .B(DB[376]), .Z(n16912) );
  XNOR U16695 ( .A(q[4]), .B(DB[375]), .Z(n14321) );
  IV U16696 ( .A(n14335), .Z(n16910) );
  XOR U16697 ( .A(n16913), .B(n16914), .Z(n14335) );
  XNOR U16698 ( .A(n14331), .B(n14333), .Z(n16914) );
  XNOR U16699 ( .A(q[0]), .B(DB[371]), .Z(n14333) );
  XNOR U16700 ( .A(q[3]), .B(DB[374]), .Z(n14331) );
  IV U16701 ( .A(n14330), .Z(n16913) );
  XNOR U16702 ( .A(n14328), .B(n16915), .Z(n14330) );
  XNOR U16703 ( .A(q[2]), .B(DB[373]), .Z(n16915) );
  XNOR U16704 ( .A(q[1]), .B(DB[372]), .Z(n14328) );
  XOR U16705 ( .A(n16916), .B(n14293), .Z(n14256) );
  XOR U16706 ( .A(n16917), .B(n14281), .Z(n14293) );
  XNOR U16707 ( .A(q[6]), .B(DB[384]), .Z(n14281) );
  IV U16708 ( .A(n14280), .Z(n16917) );
  XNOR U16709 ( .A(n14278), .B(n16918), .Z(n14280) );
  XNOR U16710 ( .A(q[5]), .B(DB[383]), .Z(n16918) );
  XNOR U16711 ( .A(q[4]), .B(DB[382]), .Z(n14278) );
  IV U16712 ( .A(n14292), .Z(n16916) );
  XOR U16713 ( .A(n16919), .B(n16920), .Z(n14292) );
  XNOR U16714 ( .A(n14288), .B(n14290), .Z(n16920) );
  XNOR U16715 ( .A(q[0]), .B(DB[378]), .Z(n14290) );
  XNOR U16716 ( .A(q[3]), .B(DB[381]), .Z(n14288) );
  IV U16717 ( .A(n14287), .Z(n16919) );
  XNOR U16718 ( .A(n14285), .B(n16921), .Z(n14287) );
  XNOR U16719 ( .A(q[2]), .B(DB[380]), .Z(n16921) );
  XNOR U16720 ( .A(q[1]), .B(DB[379]), .Z(n14285) );
  XOR U16721 ( .A(n16922), .B(n14250), .Z(n14213) );
  XOR U16722 ( .A(n16923), .B(n14238), .Z(n14250) );
  XNOR U16723 ( .A(q[6]), .B(DB[391]), .Z(n14238) );
  IV U16724 ( .A(n14237), .Z(n16923) );
  XNOR U16725 ( .A(n14235), .B(n16924), .Z(n14237) );
  XNOR U16726 ( .A(q[5]), .B(DB[390]), .Z(n16924) );
  XNOR U16727 ( .A(q[4]), .B(DB[389]), .Z(n14235) );
  IV U16728 ( .A(n14249), .Z(n16922) );
  XOR U16729 ( .A(n16925), .B(n16926), .Z(n14249) );
  XNOR U16730 ( .A(n14245), .B(n14247), .Z(n16926) );
  XNOR U16731 ( .A(q[0]), .B(DB[385]), .Z(n14247) );
  XNOR U16732 ( .A(q[3]), .B(DB[388]), .Z(n14245) );
  IV U16733 ( .A(n14244), .Z(n16925) );
  XNOR U16734 ( .A(n14242), .B(n16927), .Z(n14244) );
  XNOR U16735 ( .A(q[2]), .B(DB[387]), .Z(n16927) );
  XNOR U16736 ( .A(q[1]), .B(DB[386]), .Z(n14242) );
  XOR U16737 ( .A(n16928), .B(n14207), .Z(n14170) );
  XOR U16738 ( .A(n16929), .B(n14195), .Z(n14207) );
  XNOR U16739 ( .A(q[6]), .B(DB[398]), .Z(n14195) );
  IV U16740 ( .A(n14194), .Z(n16929) );
  XNOR U16741 ( .A(n14192), .B(n16930), .Z(n14194) );
  XNOR U16742 ( .A(q[5]), .B(DB[397]), .Z(n16930) );
  XNOR U16743 ( .A(q[4]), .B(DB[396]), .Z(n14192) );
  IV U16744 ( .A(n14206), .Z(n16928) );
  XOR U16745 ( .A(n16931), .B(n16932), .Z(n14206) );
  XNOR U16746 ( .A(n14202), .B(n14204), .Z(n16932) );
  XNOR U16747 ( .A(q[0]), .B(DB[392]), .Z(n14204) );
  XNOR U16748 ( .A(q[3]), .B(DB[395]), .Z(n14202) );
  IV U16749 ( .A(n14201), .Z(n16931) );
  XNOR U16750 ( .A(n14199), .B(n16933), .Z(n14201) );
  XNOR U16751 ( .A(q[2]), .B(DB[394]), .Z(n16933) );
  XNOR U16752 ( .A(q[1]), .B(DB[393]), .Z(n14199) );
  XOR U16753 ( .A(n16934), .B(n14164), .Z(n14127) );
  XOR U16754 ( .A(n16935), .B(n14152), .Z(n14164) );
  XNOR U16755 ( .A(q[6]), .B(DB[405]), .Z(n14152) );
  IV U16756 ( .A(n14151), .Z(n16935) );
  XNOR U16757 ( .A(n14149), .B(n16936), .Z(n14151) );
  XNOR U16758 ( .A(q[5]), .B(DB[404]), .Z(n16936) );
  XNOR U16759 ( .A(q[4]), .B(DB[403]), .Z(n14149) );
  IV U16760 ( .A(n14163), .Z(n16934) );
  XOR U16761 ( .A(n16937), .B(n16938), .Z(n14163) );
  XNOR U16762 ( .A(n14159), .B(n14161), .Z(n16938) );
  XNOR U16763 ( .A(q[0]), .B(DB[399]), .Z(n14161) );
  XNOR U16764 ( .A(q[3]), .B(DB[402]), .Z(n14159) );
  IV U16765 ( .A(n14158), .Z(n16937) );
  XNOR U16766 ( .A(n14156), .B(n16939), .Z(n14158) );
  XNOR U16767 ( .A(q[2]), .B(DB[401]), .Z(n16939) );
  XNOR U16768 ( .A(q[1]), .B(DB[400]), .Z(n14156) );
  XOR U16769 ( .A(n16940), .B(n14121), .Z(n14084) );
  XOR U16770 ( .A(n16941), .B(n14109), .Z(n14121) );
  XNOR U16771 ( .A(q[6]), .B(DB[412]), .Z(n14109) );
  IV U16772 ( .A(n14108), .Z(n16941) );
  XNOR U16773 ( .A(n14106), .B(n16942), .Z(n14108) );
  XNOR U16774 ( .A(q[5]), .B(DB[411]), .Z(n16942) );
  XNOR U16775 ( .A(q[4]), .B(DB[410]), .Z(n14106) );
  IV U16776 ( .A(n14120), .Z(n16940) );
  XOR U16777 ( .A(n16943), .B(n16944), .Z(n14120) );
  XNOR U16778 ( .A(n14116), .B(n14118), .Z(n16944) );
  XNOR U16779 ( .A(q[0]), .B(DB[406]), .Z(n14118) );
  XNOR U16780 ( .A(q[3]), .B(DB[409]), .Z(n14116) );
  IV U16781 ( .A(n14115), .Z(n16943) );
  XNOR U16782 ( .A(n14113), .B(n16945), .Z(n14115) );
  XNOR U16783 ( .A(q[2]), .B(DB[408]), .Z(n16945) );
  XNOR U16784 ( .A(q[1]), .B(DB[407]), .Z(n14113) );
  XOR U16785 ( .A(n16946), .B(n14078), .Z(n14041) );
  XOR U16786 ( .A(n16947), .B(n14066), .Z(n14078) );
  XNOR U16787 ( .A(q[6]), .B(DB[419]), .Z(n14066) );
  IV U16788 ( .A(n14065), .Z(n16947) );
  XNOR U16789 ( .A(n14063), .B(n16948), .Z(n14065) );
  XNOR U16790 ( .A(q[5]), .B(DB[418]), .Z(n16948) );
  XNOR U16791 ( .A(q[4]), .B(DB[417]), .Z(n14063) );
  IV U16792 ( .A(n14077), .Z(n16946) );
  XOR U16793 ( .A(n16949), .B(n16950), .Z(n14077) );
  XNOR U16794 ( .A(n14073), .B(n14075), .Z(n16950) );
  XNOR U16795 ( .A(q[0]), .B(DB[413]), .Z(n14075) );
  XNOR U16796 ( .A(q[3]), .B(DB[416]), .Z(n14073) );
  IV U16797 ( .A(n14072), .Z(n16949) );
  XNOR U16798 ( .A(n14070), .B(n16951), .Z(n14072) );
  XNOR U16799 ( .A(q[2]), .B(DB[415]), .Z(n16951) );
  XNOR U16800 ( .A(q[1]), .B(DB[414]), .Z(n14070) );
  XOR U16801 ( .A(n16952), .B(n14035), .Z(n13998) );
  XOR U16802 ( .A(n16953), .B(n14023), .Z(n14035) );
  XNOR U16803 ( .A(q[6]), .B(DB[426]), .Z(n14023) );
  IV U16804 ( .A(n14022), .Z(n16953) );
  XNOR U16805 ( .A(n14020), .B(n16954), .Z(n14022) );
  XNOR U16806 ( .A(q[5]), .B(DB[425]), .Z(n16954) );
  XNOR U16807 ( .A(q[4]), .B(DB[424]), .Z(n14020) );
  IV U16808 ( .A(n14034), .Z(n16952) );
  XOR U16809 ( .A(n16955), .B(n16956), .Z(n14034) );
  XNOR U16810 ( .A(n14030), .B(n14032), .Z(n16956) );
  XNOR U16811 ( .A(q[0]), .B(DB[420]), .Z(n14032) );
  XNOR U16812 ( .A(q[3]), .B(DB[423]), .Z(n14030) );
  IV U16813 ( .A(n14029), .Z(n16955) );
  XNOR U16814 ( .A(n14027), .B(n16957), .Z(n14029) );
  XNOR U16815 ( .A(q[2]), .B(DB[422]), .Z(n16957) );
  XNOR U16816 ( .A(q[1]), .B(DB[421]), .Z(n14027) );
  XOR U16817 ( .A(n16958), .B(n13992), .Z(n13955) );
  XOR U16818 ( .A(n16959), .B(n13980), .Z(n13992) );
  XNOR U16819 ( .A(q[6]), .B(DB[433]), .Z(n13980) );
  IV U16820 ( .A(n13979), .Z(n16959) );
  XNOR U16821 ( .A(n13977), .B(n16960), .Z(n13979) );
  XNOR U16822 ( .A(q[5]), .B(DB[432]), .Z(n16960) );
  XNOR U16823 ( .A(q[4]), .B(DB[431]), .Z(n13977) );
  IV U16824 ( .A(n13991), .Z(n16958) );
  XOR U16825 ( .A(n16961), .B(n16962), .Z(n13991) );
  XNOR U16826 ( .A(n13987), .B(n13989), .Z(n16962) );
  XNOR U16827 ( .A(q[0]), .B(DB[427]), .Z(n13989) );
  XNOR U16828 ( .A(q[3]), .B(DB[430]), .Z(n13987) );
  IV U16829 ( .A(n13986), .Z(n16961) );
  XNOR U16830 ( .A(n13984), .B(n16963), .Z(n13986) );
  XNOR U16831 ( .A(q[2]), .B(DB[429]), .Z(n16963) );
  XNOR U16832 ( .A(q[1]), .B(DB[428]), .Z(n13984) );
  XOR U16833 ( .A(n16964), .B(n13949), .Z(n13912) );
  XOR U16834 ( .A(n16965), .B(n13937), .Z(n13949) );
  XNOR U16835 ( .A(q[6]), .B(DB[440]), .Z(n13937) );
  IV U16836 ( .A(n13936), .Z(n16965) );
  XNOR U16837 ( .A(n13934), .B(n16966), .Z(n13936) );
  XNOR U16838 ( .A(q[5]), .B(DB[439]), .Z(n16966) );
  XNOR U16839 ( .A(q[4]), .B(DB[438]), .Z(n13934) );
  IV U16840 ( .A(n13948), .Z(n16964) );
  XOR U16841 ( .A(n16967), .B(n16968), .Z(n13948) );
  XNOR U16842 ( .A(n13944), .B(n13946), .Z(n16968) );
  XNOR U16843 ( .A(q[0]), .B(DB[434]), .Z(n13946) );
  XNOR U16844 ( .A(q[3]), .B(DB[437]), .Z(n13944) );
  IV U16845 ( .A(n13943), .Z(n16967) );
  XNOR U16846 ( .A(n13941), .B(n16969), .Z(n13943) );
  XNOR U16847 ( .A(q[2]), .B(DB[436]), .Z(n16969) );
  XNOR U16848 ( .A(q[1]), .B(DB[435]), .Z(n13941) );
  XOR U16849 ( .A(n16970), .B(n13906), .Z(n13869) );
  XOR U16850 ( .A(n16971), .B(n13894), .Z(n13906) );
  XNOR U16851 ( .A(q[6]), .B(DB[447]), .Z(n13894) );
  IV U16852 ( .A(n13893), .Z(n16971) );
  XNOR U16853 ( .A(n13891), .B(n16972), .Z(n13893) );
  XNOR U16854 ( .A(q[5]), .B(DB[446]), .Z(n16972) );
  XNOR U16855 ( .A(q[4]), .B(DB[445]), .Z(n13891) );
  IV U16856 ( .A(n13905), .Z(n16970) );
  XOR U16857 ( .A(n16973), .B(n16974), .Z(n13905) );
  XNOR U16858 ( .A(n13901), .B(n13903), .Z(n16974) );
  XNOR U16859 ( .A(q[0]), .B(DB[441]), .Z(n13903) );
  XNOR U16860 ( .A(q[3]), .B(DB[444]), .Z(n13901) );
  IV U16861 ( .A(n13900), .Z(n16973) );
  XNOR U16862 ( .A(n13898), .B(n16975), .Z(n13900) );
  XNOR U16863 ( .A(q[2]), .B(DB[443]), .Z(n16975) );
  XNOR U16864 ( .A(q[1]), .B(DB[442]), .Z(n13898) );
  XOR U16865 ( .A(n16976), .B(n13863), .Z(n13826) );
  XOR U16866 ( .A(n16977), .B(n13851), .Z(n13863) );
  XNOR U16867 ( .A(q[6]), .B(DB[454]), .Z(n13851) );
  IV U16868 ( .A(n13850), .Z(n16977) );
  XNOR U16869 ( .A(n13848), .B(n16978), .Z(n13850) );
  XNOR U16870 ( .A(q[5]), .B(DB[453]), .Z(n16978) );
  XNOR U16871 ( .A(q[4]), .B(DB[452]), .Z(n13848) );
  IV U16872 ( .A(n13862), .Z(n16976) );
  XOR U16873 ( .A(n16979), .B(n16980), .Z(n13862) );
  XNOR U16874 ( .A(n13858), .B(n13860), .Z(n16980) );
  XNOR U16875 ( .A(q[0]), .B(DB[448]), .Z(n13860) );
  XNOR U16876 ( .A(q[3]), .B(DB[451]), .Z(n13858) );
  IV U16877 ( .A(n13857), .Z(n16979) );
  XNOR U16878 ( .A(n13855), .B(n16981), .Z(n13857) );
  XNOR U16879 ( .A(q[2]), .B(DB[450]), .Z(n16981) );
  XNOR U16880 ( .A(q[1]), .B(DB[449]), .Z(n13855) );
  XOR U16881 ( .A(n16982), .B(n13820), .Z(n13783) );
  XOR U16882 ( .A(n16983), .B(n13808), .Z(n13820) );
  XNOR U16883 ( .A(q[6]), .B(DB[461]), .Z(n13808) );
  IV U16884 ( .A(n13807), .Z(n16983) );
  XNOR U16885 ( .A(n13805), .B(n16984), .Z(n13807) );
  XNOR U16886 ( .A(q[5]), .B(DB[460]), .Z(n16984) );
  XNOR U16887 ( .A(q[4]), .B(DB[459]), .Z(n13805) );
  IV U16888 ( .A(n13819), .Z(n16982) );
  XOR U16889 ( .A(n16985), .B(n16986), .Z(n13819) );
  XNOR U16890 ( .A(n13815), .B(n13817), .Z(n16986) );
  XNOR U16891 ( .A(q[0]), .B(DB[455]), .Z(n13817) );
  XNOR U16892 ( .A(q[3]), .B(DB[458]), .Z(n13815) );
  IV U16893 ( .A(n13814), .Z(n16985) );
  XNOR U16894 ( .A(n13812), .B(n16987), .Z(n13814) );
  XNOR U16895 ( .A(q[2]), .B(DB[457]), .Z(n16987) );
  XNOR U16896 ( .A(q[1]), .B(DB[456]), .Z(n13812) );
  XOR U16897 ( .A(n16988), .B(n13777), .Z(n13740) );
  XOR U16898 ( .A(n16989), .B(n13765), .Z(n13777) );
  XNOR U16899 ( .A(q[6]), .B(DB[468]), .Z(n13765) );
  IV U16900 ( .A(n13764), .Z(n16989) );
  XNOR U16901 ( .A(n13762), .B(n16990), .Z(n13764) );
  XNOR U16902 ( .A(q[5]), .B(DB[467]), .Z(n16990) );
  XNOR U16903 ( .A(q[4]), .B(DB[466]), .Z(n13762) );
  IV U16904 ( .A(n13776), .Z(n16988) );
  XOR U16905 ( .A(n16991), .B(n16992), .Z(n13776) );
  XNOR U16906 ( .A(n13772), .B(n13774), .Z(n16992) );
  XNOR U16907 ( .A(q[0]), .B(DB[462]), .Z(n13774) );
  XNOR U16908 ( .A(q[3]), .B(DB[465]), .Z(n13772) );
  IV U16909 ( .A(n13771), .Z(n16991) );
  XNOR U16910 ( .A(n13769), .B(n16993), .Z(n13771) );
  XNOR U16911 ( .A(q[2]), .B(DB[464]), .Z(n16993) );
  XNOR U16912 ( .A(q[1]), .B(DB[463]), .Z(n13769) );
  XOR U16913 ( .A(n16994), .B(n13734), .Z(n13697) );
  XOR U16914 ( .A(n16995), .B(n13722), .Z(n13734) );
  XNOR U16915 ( .A(q[6]), .B(DB[475]), .Z(n13722) );
  IV U16916 ( .A(n13721), .Z(n16995) );
  XNOR U16917 ( .A(n13719), .B(n16996), .Z(n13721) );
  XNOR U16918 ( .A(q[5]), .B(DB[474]), .Z(n16996) );
  XNOR U16919 ( .A(q[4]), .B(DB[473]), .Z(n13719) );
  IV U16920 ( .A(n13733), .Z(n16994) );
  XOR U16921 ( .A(n16997), .B(n16998), .Z(n13733) );
  XNOR U16922 ( .A(n13729), .B(n13731), .Z(n16998) );
  XNOR U16923 ( .A(q[0]), .B(DB[469]), .Z(n13731) );
  XNOR U16924 ( .A(q[3]), .B(DB[472]), .Z(n13729) );
  IV U16925 ( .A(n13728), .Z(n16997) );
  XNOR U16926 ( .A(n13726), .B(n16999), .Z(n13728) );
  XNOR U16927 ( .A(q[2]), .B(DB[471]), .Z(n16999) );
  XNOR U16928 ( .A(q[1]), .B(DB[470]), .Z(n13726) );
  XOR U16929 ( .A(n17000), .B(n13691), .Z(n13654) );
  XOR U16930 ( .A(n17001), .B(n13679), .Z(n13691) );
  XNOR U16931 ( .A(q[6]), .B(DB[482]), .Z(n13679) );
  IV U16932 ( .A(n13678), .Z(n17001) );
  XNOR U16933 ( .A(n13676), .B(n17002), .Z(n13678) );
  XNOR U16934 ( .A(q[5]), .B(DB[481]), .Z(n17002) );
  XNOR U16935 ( .A(q[4]), .B(DB[480]), .Z(n13676) );
  IV U16936 ( .A(n13690), .Z(n17000) );
  XOR U16937 ( .A(n17003), .B(n17004), .Z(n13690) );
  XNOR U16938 ( .A(n13686), .B(n13688), .Z(n17004) );
  XNOR U16939 ( .A(q[0]), .B(DB[476]), .Z(n13688) );
  XNOR U16940 ( .A(q[3]), .B(DB[479]), .Z(n13686) );
  IV U16941 ( .A(n13685), .Z(n17003) );
  XNOR U16942 ( .A(n13683), .B(n17005), .Z(n13685) );
  XNOR U16943 ( .A(q[2]), .B(DB[478]), .Z(n17005) );
  XNOR U16944 ( .A(q[1]), .B(DB[477]), .Z(n13683) );
  XOR U16945 ( .A(n17006), .B(n13648), .Z(n13611) );
  XOR U16946 ( .A(n17007), .B(n13636), .Z(n13648) );
  XNOR U16947 ( .A(q[6]), .B(DB[489]), .Z(n13636) );
  IV U16948 ( .A(n13635), .Z(n17007) );
  XNOR U16949 ( .A(n13633), .B(n17008), .Z(n13635) );
  XNOR U16950 ( .A(q[5]), .B(DB[488]), .Z(n17008) );
  XNOR U16951 ( .A(q[4]), .B(DB[487]), .Z(n13633) );
  IV U16952 ( .A(n13647), .Z(n17006) );
  XOR U16953 ( .A(n17009), .B(n17010), .Z(n13647) );
  XNOR U16954 ( .A(n13643), .B(n13645), .Z(n17010) );
  XNOR U16955 ( .A(q[0]), .B(DB[483]), .Z(n13645) );
  XNOR U16956 ( .A(q[3]), .B(DB[486]), .Z(n13643) );
  IV U16957 ( .A(n13642), .Z(n17009) );
  XNOR U16958 ( .A(n13640), .B(n17011), .Z(n13642) );
  XNOR U16959 ( .A(q[2]), .B(DB[485]), .Z(n17011) );
  XNOR U16960 ( .A(q[1]), .B(DB[484]), .Z(n13640) );
  XOR U16961 ( .A(n17012), .B(n13605), .Z(n13568) );
  XOR U16962 ( .A(n17013), .B(n13593), .Z(n13605) );
  XNOR U16963 ( .A(q[6]), .B(DB[496]), .Z(n13593) );
  IV U16964 ( .A(n13592), .Z(n17013) );
  XNOR U16965 ( .A(n13590), .B(n17014), .Z(n13592) );
  XNOR U16966 ( .A(q[5]), .B(DB[495]), .Z(n17014) );
  XNOR U16967 ( .A(q[4]), .B(DB[494]), .Z(n13590) );
  IV U16968 ( .A(n13604), .Z(n17012) );
  XOR U16969 ( .A(n17015), .B(n17016), .Z(n13604) );
  XNOR U16970 ( .A(n13600), .B(n13602), .Z(n17016) );
  XNOR U16971 ( .A(q[0]), .B(DB[490]), .Z(n13602) );
  XNOR U16972 ( .A(q[3]), .B(DB[493]), .Z(n13600) );
  IV U16973 ( .A(n13599), .Z(n17015) );
  XNOR U16974 ( .A(n13597), .B(n17017), .Z(n13599) );
  XNOR U16975 ( .A(q[2]), .B(DB[492]), .Z(n17017) );
  XNOR U16976 ( .A(q[1]), .B(DB[491]), .Z(n13597) );
  XOR U16977 ( .A(n17018), .B(n13562), .Z(n13525) );
  XOR U16978 ( .A(n17019), .B(n13550), .Z(n13562) );
  XNOR U16979 ( .A(q[6]), .B(DB[503]), .Z(n13550) );
  IV U16980 ( .A(n13549), .Z(n17019) );
  XNOR U16981 ( .A(n13547), .B(n17020), .Z(n13549) );
  XNOR U16982 ( .A(q[5]), .B(DB[502]), .Z(n17020) );
  XNOR U16983 ( .A(q[4]), .B(DB[501]), .Z(n13547) );
  IV U16984 ( .A(n13561), .Z(n17018) );
  XOR U16985 ( .A(n17021), .B(n17022), .Z(n13561) );
  XNOR U16986 ( .A(n13557), .B(n13559), .Z(n17022) );
  XNOR U16987 ( .A(q[0]), .B(DB[497]), .Z(n13559) );
  XNOR U16988 ( .A(q[3]), .B(DB[500]), .Z(n13557) );
  IV U16989 ( .A(n13556), .Z(n17021) );
  XNOR U16990 ( .A(n13554), .B(n17023), .Z(n13556) );
  XNOR U16991 ( .A(q[2]), .B(DB[499]), .Z(n17023) );
  XNOR U16992 ( .A(q[1]), .B(DB[498]), .Z(n13554) );
  XOR U16993 ( .A(n17024), .B(n13519), .Z(n13482) );
  XOR U16994 ( .A(n17025), .B(n13507), .Z(n13519) );
  XNOR U16995 ( .A(q[6]), .B(DB[510]), .Z(n13507) );
  IV U16996 ( .A(n13506), .Z(n17025) );
  XNOR U16997 ( .A(n13504), .B(n17026), .Z(n13506) );
  XNOR U16998 ( .A(q[5]), .B(DB[509]), .Z(n17026) );
  XNOR U16999 ( .A(q[4]), .B(DB[508]), .Z(n13504) );
  IV U17000 ( .A(n13518), .Z(n17024) );
  XOR U17001 ( .A(n17027), .B(n17028), .Z(n13518) );
  XNOR U17002 ( .A(n13514), .B(n13516), .Z(n17028) );
  XNOR U17003 ( .A(q[0]), .B(DB[504]), .Z(n13516) );
  XNOR U17004 ( .A(q[3]), .B(DB[507]), .Z(n13514) );
  IV U17005 ( .A(n13513), .Z(n17027) );
  XNOR U17006 ( .A(n13511), .B(n17029), .Z(n13513) );
  XNOR U17007 ( .A(q[2]), .B(DB[506]), .Z(n17029) );
  XNOR U17008 ( .A(q[1]), .B(DB[505]), .Z(n13511) );
  XOR U17009 ( .A(n17030), .B(n13476), .Z(n13439) );
  XOR U17010 ( .A(n17031), .B(n13464), .Z(n13476) );
  XNOR U17011 ( .A(q[6]), .B(DB[517]), .Z(n13464) );
  IV U17012 ( .A(n13463), .Z(n17031) );
  XNOR U17013 ( .A(n13461), .B(n17032), .Z(n13463) );
  XNOR U17014 ( .A(q[5]), .B(DB[516]), .Z(n17032) );
  XNOR U17015 ( .A(q[4]), .B(DB[515]), .Z(n13461) );
  IV U17016 ( .A(n13475), .Z(n17030) );
  XOR U17017 ( .A(n17033), .B(n17034), .Z(n13475) );
  XNOR U17018 ( .A(n13471), .B(n13473), .Z(n17034) );
  XNOR U17019 ( .A(q[0]), .B(DB[511]), .Z(n13473) );
  XNOR U17020 ( .A(q[3]), .B(DB[514]), .Z(n13471) );
  IV U17021 ( .A(n13470), .Z(n17033) );
  XNOR U17022 ( .A(n13468), .B(n17035), .Z(n13470) );
  XNOR U17023 ( .A(q[2]), .B(DB[513]), .Z(n17035) );
  XNOR U17024 ( .A(q[1]), .B(DB[512]), .Z(n13468) );
  XOR U17025 ( .A(n17036), .B(n13433), .Z(n13396) );
  XOR U17026 ( .A(n17037), .B(n13421), .Z(n13433) );
  XNOR U17027 ( .A(q[6]), .B(DB[524]), .Z(n13421) );
  IV U17028 ( .A(n13420), .Z(n17037) );
  XNOR U17029 ( .A(n13418), .B(n17038), .Z(n13420) );
  XNOR U17030 ( .A(q[5]), .B(DB[523]), .Z(n17038) );
  XNOR U17031 ( .A(q[4]), .B(DB[522]), .Z(n13418) );
  IV U17032 ( .A(n13432), .Z(n17036) );
  XOR U17033 ( .A(n17039), .B(n17040), .Z(n13432) );
  XNOR U17034 ( .A(n13428), .B(n13430), .Z(n17040) );
  XNOR U17035 ( .A(q[0]), .B(DB[518]), .Z(n13430) );
  XNOR U17036 ( .A(q[3]), .B(DB[521]), .Z(n13428) );
  IV U17037 ( .A(n13427), .Z(n17039) );
  XNOR U17038 ( .A(n13425), .B(n17041), .Z(n13427) );
  XNOR U17039 ( .A(q[2]), .B(DB[520]), .Z(n17041) );
  XNOR U17040 ( .A(q[1]), .B(DB[519]), .Z(n13425) );
  XOR U17041 ( .A(n17042), .B(n13390), .Z(n13353) );
  XOR U17042 ( .A(n17043), .B(n13378), .Z(n13390) );
  XNOR U17043 ( .A(q[6]), .B(DB[531]), .Z(n13378) );
  IV U17044 ( .A(n13377), .Z(n17043) );
  XNOR U17045 ( .A(n13375), .B(n17044), .Z(n13377) );
  XNOR U17046 ( .A(q[5]), .B(DB[530]), .Z(n17044) );
  XNOR U17047 ( .A(q[4]), .B(DB[529]), .Z(n13375) );
  IV U17048 ( .A(n13389), .Z(n17042) );
  XOR U17049 ( .A(n17045), .B(n17046), .Z(n13389) );
  XNOR U17050 ( .A(n13385), .B(n13387), .Z(n17046) );
  XNOR U17051 ( .A(q[0]), .B(DB[525]), .Z(n13387) );
  XNOR U17052 ( .A(q[3]), .B(DB[528]), .Z(n13385) );
  IV U17053 ( .A(n13384), .Z(n17045) );
  XNOR U17054 ( .A(n13382), .B(n17047), .Z(n13384) );
  XNOR U17055 ( .A(q[2]), .B(DB[527]), .Z(n17047) );
  XNOR U17056 ( .A(q[1]), .B(DB[526]), .Z(n13382) );
  XOR U17057 ( .A(n17048), .B(n13347), .Z(n13310) );
  XOR U17058 ( .A(n17049), .B(n13335), .Z(n13347) );
  XNOR U17059 ( .A(q[6]), .B(DB[538]), .Z(n13335) );
  IV U17060 ( .A(n13334), .Z(n17049) );
  XNOR U17061 ( .A(n13332), .B(n17050), .Z(n13334) );
  XNOR U17062 ( .A(q[5]), .B(DB[537]), .Z(n17050) );
  XNOR U17063 ( .A(q[4]), .B(DB[536]), .Z(n13332) );
  IV U17064 ( .A(n13346), .Z(n17048) );
  XOR U17065 ( .A(n17051), .B(n17052), .Z(n13346) );
  XNOR U17066 ( .A(n13342), .B(n13344), .Z(n17052) );
  XNOR U17067 ( .A(q[0]), .B(DB[532]), .Z(n13344) );
  XNOR U17068 ( .A(q[3]), .B(DB[535]), .Z(n13342) );
  IV U17069 ( .A(n13341), .Z(n17051) );
  XNOR U17070 ( .A(n13339), .B(n17053), .Z(n13341) );
  XNOR U17071 ( .A(q[2]), .B(DB[534]), .Z(n17053) );
  XNOR U17072 ( .A(q[1]), .B(DB[533]), .Z(n13339) );
  XOR U17073 ( .A(n17054), .B(n13304), .Z(n13267) );
  XOR U17074 ( .A(n17055), .B(n13292), .Z(n13304) );
  XNOR U17075 ( .A(q[6]), .B(DB[545]), .Z(n13292) );
  IV U17076 ( .A(n13291), .Z(n17055) );
  XNOR U17077 ( .A(n13289), .B(n17056), .Z(n13291) );
  XNOR U17078 ( .A(q[5]), .B(DB[544]), .Z(n17056) );
  XNOR U17079 ( .A(q[4]), .B(DB[543]), .Z(n13289) );
  IV U17080 ( .A(n13303), .Z(n17054) );
  XOR U17081 ( .A(n17057), .B(n17058), .Z(n13303) );
  XNOR U17082 ( .A(n13299), .B(n13301), .Z(n17058) );
  XNOR U17083 ( .A(q[0]), .B(DB[539]), .Z(n13301) );
  XNOR U17084 ( .A(q[3]), .B(DB[542]), .Z(n13299) );
  IV U17085 ( .A(n13298), .Z(n17057) );
  XNOR U17086 ( .A(n13296), .B(n17059), .Z(n13298) );
  XNOR U17087 ( .A(q[2]), .B(DB[541]), .Z(n17059) );
  XNOR U17088 ( .A(q[1]), .B(DB[540]), .Z(n13296) );
  XOR U17089 ( .A(n17060), .B(n13261), .Z(n13224) );
  XOR U17090 ( .A(n17061), .B(n13249), .Z(n13261) );
  XNOR U17091 ( .A(q[6]), .B(DB[552]), .Z(n13249) );
  IV U17092 ( .A(n13248), .Z(n17061) );
  XNOR U17093 ( .A(n13246), .B(n17062), .Z(n13248) );
  XNOR U17094 ( .A(q[5]), .B(DB[551]), .Z(n17062) );
  XNOR U17095 ( .A(q[4]), .B(DB[550]), .Z(n13246) );
  IV U17096 ( .A(n13260), .Z(n17060) );
  XOR U17097 ( .A(n17063), .B(n17064), .Z(n13260) );
  XNOR U17098 ( .A(n13256), .B(n13258), .Z(n17064) );
  XNOR U17099 ( .A(q[0]), .B(DB[546]), .Z(n13258) );
  XNOR U17100 ( .A(q[3]), .B(DB[549]), .Z(n13256) );
  IV U17101 ( .A(n13255), .Z(n17063) );
  XNOR U17102 ( .A(n13253), .B(n17065), .Z(n13255) );
  XNOR U17103 ( .A(q[2]), .B(DB[548]), .Z(n17065) );
  XNOR U17104 ( .A(q[1]), .B(DB[547]), .Z(n13253) );
  XOR U17105 ( .A(n17066), .B(n13218), .Z(n13181) );
  XOR U17106 ( .A(n17067), .B(n13206), .Z(n13218) );
  XNOR U17107 ( .A(q[6]), .B(DB[559]), .Z(n13206) );
  IV U17108 ( .A(n13205), .Z(n17067) );
  XNOR U17109 ( .A(n13203), .B(n17068), .Z(n13205) );
  XNOR U17110 ( .A(q[5]), .B(DB[558]), .Z(n17068) );
  XNOR U17111 ( .A(q[4]), .B(DB[557]), .Z(n13203) );
  IV U17112 ( .A(n13217), .Z(n17066) );
  XOR U17113 ( .A(n17069), .B(n17070), .Z(n13217) );
  XNOR U17114 ( .A(n13213), .B(n13215), .Z(n17070) );
  XNOR U17115 ( .A(q[0]), .B(DB[553]), .Z(n13215) );
  XNOR U17116 ( .A(q[3]), .B(DB[556]), .Z(n13213) );
  IV U17117 ( .A(n13212), .Z(n17069) );
  XNOR U17118 ( .A(n13210), .B(n17071), .Z(n13212) );
  XNOR U17119 ( .A(q[2]), .B(DB[555]), .Z(n17071) );
  XNOR U17120 ( .A(q[1]), .B(DB[554]), .Z(n13210) );
  XOR U17121 ( .A(n17072), .B(n13175), .Z(n13138) );
  XOR U17122 ( .A(n17073), .B(n13163), .Z(n13175) );
  XNOR U17123 ( .A(q[6]), .B(DB[566]), .Z(n13163) );
  IV U17124 ( .A(n13162), .Z(n17073) );
  XNOR U17125 ( .A(n13160), .B(n17074), .Z(n13162) );
  XNOR U17126 ( .A(q[5]), .B(DB[565]), .Z(n17074) );
  XNOR U17127 ( .A(q[4]), .B(DB[564]), .Z(n13160) );
  IV U17128 ( .A(n13174), .Z(n17072) );
  XOR U17129 ( .A(n17075), .B(n17076), .Z(n13174) );
  XNOR U17130 ( .A(n13170), .B(n13172), .Z(n17076) );
  XNOR U17131 ( .A(q[0]), .B(DB[560]), .Z(n13172) );
  XNOR U17132 ( .A(q[3]), .B(DB[563]), .Z(n13170) );
  IV U17133 ( .A(n13169), .Z(n17075) );
  XNOR U17134 ( .A(n13167), .B(n17077), .Z(n13169) );
  XNOR U17135 ( .A(q[2]), .B(DB[562]), .Z(n17077) );
  XNOR U17136 ( .A(q[1]), .B(DB[561]), .Z(n13167) );
  XOR U17137 ( .A(n17078), .B(n13132), .Z(n13095) );
  XOR U17138 ( .A(n17079), .B(n13120), .Z(n13132) );
  XNOR U17139 ( .A(q[6]), .B(DB[573]), .Z(n13120) );
  IV U17140 ( .A(n13119), .Z(n17079) );
  XNOR U17141 ( .A(n13117), .B(n17080), .Z(n13119) );
  XNOR U17142 ( .A(q[5]), .B(DB[572]), .Z(n17080) );
  XNOR U17143 ( .A(q[4]), .B(DB[571]), .Z(n13117) );
  IV U17144 ( .A(n13131), .Z(n17078) );
  XOR U17145 ( .A(n17081), .B(n17082), .Z(n13131) );
  XNOR U17146 ( .A(n13127), .B(n13129), .Z(n17082) );
  XNOR U17147 ( .A(q[0]), .B(DB[567]), .Z(n13129) );
  XNOR U17148 ( .A(q[3]), .B(DB[570]), .Z(n13127) );
  IV U17149 ( .A(n13126), .Z(n17081) );
  XNOR U17150 ( .A(n13124), .B(n17083), .Z(n13126) );
  XNOR U17151 ( .A(q[2]), .B(DB[569]), .Z(n17083) );
  XNOR U17152 ( .A(q[1]), .B(DB[568]), .Z(n13124) );
  XOR U17153 ( .A(n17084), .B(n13089), .Z(n13052) );
  XOR U17154 ( .A(n17085), .B(n13077), .Z(n13089) );
  XNOR U17155 ( .A(q[6]), .B(DB[580]), .Z(n13077) );
  IV U17156 ( .A(n13076), .Z(n17085) );
  XNOR U17157 ( .A(n13074), .B(n17086), .Z(n13076) );
  XNOR U17158 ( .A(q[5]), .B(DB[579]), .Z(n17086) );
  XNOR U17159 ( .A(q[4]), .B(DB[578]), .Z(n13074) );
  IV U17160 ( .A(n13088), .Z(n17084) );
  XOR U17161 ( .A(n17087), .B(n17088), .Z(n13088) );
  XNOR U17162 ( .A(n13084), .B(n13086), .Z(n17088) );
  XNOR U17163 ( .A(q[0]), .B(DB[574]), .Z(n13086) );
  XNOR U17164 ( .A(q[3]), .B(DB[577]), .Z(n13084) );
  IV U17165 ( .A(n13083), .Z(n17087) );
  XNOR U17166 ( .A(n13081), .B(n17089), .Z(n13083) );
  XNOR U17167 ( .A(q[2]), .B(DB[576]), .Z(n17089) );
  XNOR U17168 ( .A(q[1]), .B(DB[575]), .Z(n13081) );
  XOR U17169 ( .A(n17090), .B(n13046), .Z(n13009) );
  XOR U17170 ( .A(n17091), .B(n13034), .Z(n13046) );
  XNOR U17171 ( .A(q[6]), .B(DB[587]), .Z(n13034) );
  IV U17172 ( .A(n13033), .Z(n17091) );
  XNOR U17173 ( .A(n13031), .B(n17092), .Z(n13033) );
  XNOR U17174 ( .A(q[5]), .B(DB[586]), .Z(n17092) );
  XNOR U17175 ( .A(q[4]), .B(DB[585]), .Z(n13031) );
  IV U17176 ( .A(n13045), .Z(n17090) );
  XOR U17177 ( .A(n17093), .B(n17094), .Z(n13045) );
  XNOR U17178 ( .A(n13041), .B(n13043), .Z(n17094) );
  XNOR U17179 ( .A(q[0]), .B(DB[581]), .Z(n13043) );
  XNOR U17180 ( .A(q[3]), .B(DB[584]), .Z(n13041) );
  IV U17181 ( .A(n13040), .Z(n17093) );
  XNOR U17182 ( .A(n13038), .B(n17095), .Z(n13040) );
  XNOR U17183 ( .A(q[2]), .B(DB[583]), .Z(n17095) );
  XNOR U17184 ( .A(q[1]), .B(DB[582]), .Z(n13038) );
  XOR U17185 ( .A(n17096), .B(n13003), .Z(n12966) );
  XOR U17186 ( .A(n17097), .B(n12991), .Z(n13003) );
  XNOR U17187 ( .A(q[6]), .B(DB[594]), .Z(n12991) );
  IV U17188 ( .A(n12990), .Z(n17097) );
  XNOR U17189 ( .A(n12988), .B(n17098), .Z(n12990) );
  XNOR U17190 ( .A(q[5]), .B(DB[593]), .Z(n17098) );
  XNOR U17191 ( .A(q[4]), .B(DB[592]), .Z(n12988) );
  IV U17192 ( .A(n13002), .Z(n17096) );
  XOR U17193 ( .A(n17099), .B(n17100), .Z(n13002) );
  XNOR U17194 ( .A(n12998), .B(n13000), .Z(n17100) );
  XNOR U17195 ( .A(q[0]), .B(DB[588]), .Z(n13000) );
  XNOR U17196 ( .A(q[3]), .B(DB[591]), .Z(n12998) );
  IV U17197 ( .A(n12997), .Z(n17099) );
  XNOR U17198 ( .A(n12995), .B(n17101), .Z(n12997) );
  XNOR U17199 ( .A(q[2]), .B(DB[590]), .Z(n17101) );
  XNOR U17200 ( .A(q[1]), .B(DB[589]), .Z(n12995) );
  XOR U17201 ( .A(n17102), .B(n12960), .Z(n12923) );
  XOR U17202 ( .A(n17103), .B(n12948), .Z(n12960) );
  XNOR U17203 ( .A(q[6]), .B(DB[601]), .Z(n12948) );
  IV U17204 ( .A(n12947), .Z(n17103) );
  XNOR U17205 ( .A(n12945), .B(n17104), .Z(n12947) );
  XNOR U17206 ( .A(q[5]), .B(DB[600]), .Z(n17104) );
  XNOR U17207 ( .A(q[4]), .B(DB[599]), .Z(n12945) );
  IV U17208 ( .A(n12959), .Z(n17102) );
  XOR U17209 ( .A(n17105), .B(n17106), .Z(n12959) );
  XNOR U17210 ( .A(n12955), .B(n12957), .Z(n17106) );
  XNOR U17211 ( .A(q[0]), .B(DB[595]), .Z(n12957) );
  XNOR U17212 ( .A(q[3]), .B(DB[598]), .Z(n12955) );
  IV U17213 ( .A(n12954), .Z(n17105) );
  XNOR U17214 ( .A(n12952), .B(n17107), .Z(n12954) );
  XNOR U17215 ( .A(q[2]), .B(DB[597]), .Z(n17107) );
  XNOR U17216 ( .A(q[1]), .B(DB[596]), .Z(n12952) );
  XOR U17217 ( .A(n17108), .B(n12917), .Z(n12880) );
  XOR U17218 ( .A(n17109), .B(n12905), .Z(n12917) );
  XNOR U17219 ( .A(q[6]), .B(DB[608]), .Z(n12905) );
  IV U17220 ( .A(n12904), .Z(n17109) );
  XNOR U17221 ( .A(n12902), .B(n17110), .Z(n12904) );
  XNOR U17222 ( .A(q[5]), .B(DB[607]), .Z(n17110) );
  XNOR U17223 ( .A(q[4]), .B(DB[606]), .Z(n12902) );
  IV U17224 ( .A(n12916), .Z(n17108) );
  XOR U17225 ( .A(n17111), .B(n17112), .Z(n12916) );
  XNOR U17226 ( .A(n12912), .B(n12914), .Z(n17112) );
  XNOR U17227 ( .A(q[0]), .B(DB[602]), .Z(n12914) );
  XNOR U17228 ( .A(q[3]), .B(DB[605]), .Z(n12912) );
  IV U17229 ( .A(n12911), .Z(n17111) );
  XNOR U17230 ( .A(n12909), .B(n17113), .Z(n12911) );
  XNOR U17231 ( .A(q[2]), .B(DB[604]), .Z(n17113) );
  XNOR U17232 ( .A(q[1]), .B(DB[603]), .Z(n12909) );
  XOR U17233 ( .A(n17114), .B(n12874), .Z(n12837) );
  XOR U17234 ( .A(n17115), .B(n12862), .Z(n12874) );
  XNOR U17235 ( .A(q[6]), .B(DB[615]), .Z(n12862) );
  IV U17236 ( .A(n12861), .Z(n17115) );
  XNOR U17237 ( .A(n12859), .B(n17116), .Z(n12861) );
  XNOR U17238 ( .A(q[5]), .B(DB[614]), .Z(n17116) );
  XNOR U17239 ( .A(q[4]), .B(DB[613]), .Z(n12859) );
  IV U17240 ( .A(n12873), .Z(n17114) );
  XOR U17241 ( .A(n17117), .B(n17118), .Z(n12873) );
  XNOR U17242 ( .A(n12869), .B(n12871), .Z(n17118) );
  XNOR U17243 ( .A(q[0]), .B(DB[609]), .Z(n12871) );
  XNOR U17244 ( .A(q[3]), .B(DB[612]), .Z(n12869) );
  IV U17245 ( .A(n12868), .Z(n17117) );
  XNOR U17246 ( .A(n12866), .B(n17119), .Z(n12868) );
  XNOR U17247 ( .A(q[2]), .B(DB[611]), .Z(n17119) );
  XNOR U17248 ( .A(q[1]), .B(DB[610]), .Z(n12866) );
  XOR U17249 ( .A(n17120), .B(n12831), .Z(n12794) );
  XOR U17250 ( .A(n17121), .B(n12819), .Z(n12831) );
  XNOR U17251 ( .A(q[6]), .B(DB[622]), .Z(n12819) );
  IV U17252 ( .A(n12818), .Z(n17121) );
  XNOR U17253 ( .A(n12816), .B(n17122), .Z(n12818) );
  XNOR U17254 ( .A(q[5]), .B(DB[621]), .Z(n17122) );
  XNOR U17255 ( .A(q[4]), .B(DB[620]), .Z(n12816) );
  IV U17256 ( .A(n12830), .Z(n17120) );
  XOR U17257 ( .A(n17123), .B(n17124), .Z(n12830) );
  XNOR U17258 ( .A(n12826), .B(n12828), .Z(n17124) );
  XNOR U17259 ( .A(q[0]), .B(DB[616]), .Z(n12828) );
  XNOR U17260 ( .A(q[3]), .B(DB[619]), .Z(n12826) );
  IV U17261 ( .A(n12825), .Z(n17123) );
  XNOR U17262 ( .A(n12823), .B(n17125), .Z(n12825) );
  XNOR U17263 ( .A(q[2]), .B(DB[618]), .Z(n17125) );
  XNOR U17264 ( .A(q[1]), .B(DB[617]), .Z(n12823) );
  XOR U17265 ( .A(n17126), .B(n12788), .Z(n12751) );
  XOR U17266 ( .A(n17127), .B(n12776), .Z(n12788) );
  XNOR U17267 ( .A(q[6]), .B(DB[629]), .Z(n12776) );
  IV U17268 ( .A(n12775), .Z(n17127) );
  XNOR U17269 ( .A(n12773), .B(n17128), .Z(n12775) );
  XNOR U17270 ( .A(q[5]), .B(DB[628]), .Z(n17128) );
  XNOR U17271 ( .A(q[4]), .B(DB[627]), .Z(n12773) );
  IV U17272 ( .A(n12787), .Z(n17126) );
  XOR U17273 ( .A(n17129), .B(n17130), .Z(n12787) );
  XNOR U17274 ( .A(n12783), .B(n12785), .Z(n17130) );
  XNOR U17275 ( .A(q[0]), .B(DB[623]), .Z(n12785) );
  XNOR U17276 ( .A(q[3]), .B(DB[626]), .Z(n12783) );
  IV U17277 ( .A(n12782), .Z(n17129) );
  XNOR U17278 ( .A(n12780), .B(n17131), .Z(n12782) );
  XNOR U17279 ( .A(q[2]), .B(DB[625]), .Z(n17131) );
  XNOR U17280 ( .A(q[1]), .B(DB[624]), .Z(n12780) );
  XOR U17281 ( .A(n17132), .B(n12745), .Z(n12708) );
  XOR U17282 ( .A(n17133), .B(n12733), .Z(n12745) );
  XNOR U17283 ( .A(q[6]), .B(DB[636]), .Z(n12733) );
  IV U17284 ( .A(n12732), .Z(n17133) );
  XNOR U17285 ( .A(n12730), .B(n17134), .Z(n12732) );
  XNOR U17286 ( .A(q[5]), .B(DB[635]), .Z(n17134) );
  XNOR U17287 ( .A(q[4]), .B(DB[634]), .Z(n12730) );
  IV U17288 ( .A(n12744), .Z(n17132) );
  XOR U17289 ( .A(n17135), .B(n17136), .Z(n12744) );
  XNOR U17290 ( .A(n12740), .B(n12742), .Z(n17136) );
  XNOR U17291 ( .A(q[0]), .B(DB[630]), .Z(n12742) );
  XNOR U17292 ( .A(q[3]), .B(DB[633]), .Z(n12740) );
  IV U17293 ( .A(n12739), .Z(n17135) );
  XNOR U17294 ( .A(n12737), .B(n17137), .Z(n12739) );
  XNOR U17295 ( .A(q[2]), .B(DB[632]), .Z(n17137) );
  XNOR U17296 ( .A(q[1]), .B(DB[631]), .Z(n12737) );
  XOR U17297 ( .A(n17138), .B(n12702), .Z(n12665) );
  XOR U17298 ( .A(n17139), .B(n12690), .Z(n12702) );
  XNOR U17299 ( .A(q[6]), .B(DB[643]), .Z(n12690) );
  IV U17300 ( .A(n12689), .Z(n17139) );
  XNOR U17301 ( .A(n12687), .B(n17140), .Z(n12689) );
  XNOR U17302 ( .A(q[5]), .B(DB[642]), .Z(n17140) );
  XNOR U17303 ( .A(q[4]), .B(DB[641]), .Z(n12687) );
  IV U17304 ( .A(n12701), .Z(n17138) );
  XOR U17305 ( .A(n17141), .B(n17142), .Z(n12701) );
  XNOR U17306 ( .A(n12697), .B(n12699), .Z(n17142) );
  XNOR U17307 ( .A(q[0]), .B(DB[637]), .Z(n12699) );
  XNOR U17308 ( .A(q[3]), .B(DB[640]), .Z(n12697) );
  IV U17309 ( .A(n12696), .Z(n17141) );
  XNOR U17310 ( .A(n12694), .B(n17143), .Z(n12696) );
  XNOR U17311 ( .A(q[2]), .B(DB[639]), .Z(n17143) );
  XNOR U17312 ( .A(q[1]), .B(DB[638]), .Z(n12694) );
  XOR U17313 ( .A(n17144), .B(n12659), .Z(n12622) );
  XOR U17314 ( .A(n17145), .B(n12647), .Z(n12659) );
  XNOR U17315 ( .A(q[6]), .B(DB[650]), .Z(n12647) );
  IV U17316 ( .A(n12646), .Z(n17145) );
  XNOR U17317 ( .A(n12644), .B(n17146), .Z(n12646) );
  XNOR U17318 ( .A(q[5]), .B(DB[649]), .Z(n17146) );
  XNOR U17319 ( .A(q[4]), .B(DB[648]), .Z(n12644) );
  IV U17320 ( .A(n12658), .Z(n17144) );
  XOR U17321 ( .A(n17147), .B(n17148), .Z(n12658) );
  XNOR U17322 ( .A(n12654), .B(n12656), .Z(n17148) );
  XNOR U17323 ( .A(q[0]), .B(DB[644]), .Z(n12656) );
  XNOR U17324 ( .A(q[3]), .B(DB[647]), .Z(n12654) );
  IV U17325 ( .A(n12653), .Z(n17147) );
  XNOR U17326 ( .A(n12651), .B(n17149), .Z(n12653) );
  XNOR U17327 ( .A(q[2]), .B(DB[646]), .Z(n17149) );
  XNOR U17328 ( .A(q[1]), .B(DB[645]), .Z(n12651) );
  XOR U17329 ( .A(n17150), .B(n12616), .Z(n12579) );
  XOR U17330 ( .A(n17151), .B(n12604), .Z(n12616) );
  XNOR U17331 ( .A(q[6]), .B(DB[657]), .Z(n12604) );
  IV U17332 ( .A(n12603), .Z(n17151) );
  XNOR U17333 ( .A(n12601), .B(n17152), .Z(n12603) );
  XNOR U17334 ( .A(q[5]), .B(DB[656]), .Z(n17152) );
  XNOR U17335 ( .A(q[4]), .B(DB[655]), .Z(n12601) );
  IV U17336 ( .A(n12615), .Z(n17150) );
  XOR U17337 ( .A(n17153), .B(n17154), .Z(n12615) );
  XNOR U17338 ( .A(n12611), .B(n12613), .Z(n17154) );
  XNOR U17339 ( .A(q[0]), .B(DB[651]), .Z(n12613) );
  XNOR U17340 ( .A(q[3]), .B(DB[654]), .Z(n12611) );
  IV U17341 ( .A(n12610), .Z(n17153) );
  XNOR U17342 ( .A(n12608), .B(n17155), .Z(n12610) );
  XNOR U17343 ( .A(q[2]), .B(DB[653]), .Z(n17155) );
  XNOR U17344 ( .A(q[1]), .B(DB[652]), .Z(n12608) );
  XOR U17345 ( .A(n17156), .B(n12573), .Z(n12536) );
  XOR U17346 ( .A(n17157), .B(n12561), .Z(n12573) );
  XNOR U17347 ( .A(q[6]), .B(DB[664]), .Z(n12561) );
  IV U17348 ( .A(n12560), .Z(n17157) );
  XNOR U17349 ( .A(n12558), .B(n17158), .Z(n12560) );
  XNOR U17350 ( .A(q[5]), .B(DB[663]), .Z(n17158) );
  XNOR U17351 ( .A(q[4]), .B(DB[662]), .Z(n12558) );
  IV U17352 ( .A(n12572), .Z(n17156) );
  XOR U17353 ( .A(n17159), .B(n17160), .Z(n12572) );
  XNOR U17354 ( .A(n12568), .B(n12570), .Z(n17160) );
  XNOR U17355 ( .A(q[0]), .B(DB[658]), .Z(n12570) );
  XNOR U17356 ( .A(q[3]), .B(DB[661]), .Z(n12568) );
  IV U17357 ( .A(n12567), .Z(n17159) );
  XNOR U17358 ( .A(n12565), .B(n17161), .Z(n12567) );
  XNOR U17359 ( .A(q[2]), .B(DB[660]), .Z(n17161) );
  XNOR U17360 ( .A(q[1]), .B(DB[659]), .Z(n12565) );
  XOR U17361 ( .A(n17162), .B(n12530), .Z(n12493) );
  XOR U17362 ( .A(n17163), .B(n12518), .Z(n12530) );
  XNOR U17363 ( .A(q[6]), .B(DB[671]), .Z(n12518) );
  IV U17364 ( .A(n12517), .Z(n17163) );
  XNOR U17365 ( .A(n12515), .B(n17164), .Z(n12517) );
  XNOR U17366 ( .A(q[5]), .B(DB[670]), .Z(n17164) );
  XNOR U17367 ( .A(q[4]), .B(DB[669]), .Z(n12515) );
  IV U17368 ( .A(n12529), .Z(n17162) );
  XOR U17369 ( .A(n17165), .B(n17166), .Z(n12529) );
  XNOR U17370 ( .A(n12525), .B(n12527), .Z(n17166) );
  XNOR U17371 ( .A(q[0]), .B(DB[665]), .Z(n12527) );
  XNOR U17372 ( .A(q[3]), .B(DB[668]), .Z(n12525) );
  IV U17373 ( .A(n12524), .Z(n17165) );
  XNOR U17374 ( .A(n12522), .B(n17167), .Z(n12524) );
  XNOR U17375 ( .A(q[2]), .B(DB[667]), .Z(n17167) );
  XNOR U17376 ( .A(q[1]), .B(DB[666]), .Z(n12522) );
  XOR U17377 ( .A(n17168), .B(n12487), .Z(n12450) );
  XOR U17378 ( .A(n17169), .B(n12475), .Z(n12487) );
  XNOR U17379 ( .A(q[6]), .B(DB[678]), .Z(n12475) );
  IV U17380 ( .A(n12474), .Z(n17169) );
  XNOR U17381 ( .A(n12472), .B(n17170), .Z(n12474) );
  XNOR U17382 ( .A(q[5]), .B(DB[677]), .Z(n17170) );
  XNOR U17383 ( .A(q[4]), .B(DB[676]), .Z(n12472) );
  IV U17384 ( .A(n12486), .Z(n17168) );
  XOR U17385 ( .A(n17171), .B(n17172), .Z(n12486) );
  XNOR U17386 ( .A(n12482), .B(n12484), .Z(n17172) );
  XNOR U17387 ( .A(q[0]), .B(DB[672]), .Z(n12484) );
  XNOR U17388 ( .A(q[3]), .B(DB[675]), .Z(n12482) );
  IV U17389 ( .A(n12481), .Z(n17171) );
  XNOR U17390 ( .A(n12479), .B(n17173), .Z(n12481) );
  XNOR U17391 ( .A(q[2]), .B(DB[674]), .Z(n17173) );
  XNOR U17392 ( .A(q[1]), .B(DB[673]), .Z(n12479) );
  XOR U17393 ( .A(n17174), .B(n12444), .Z(n12407) );
  XOR U17394 ( .A(n17175), .B(n12432), .Z(n12444) );
  XNOR U17395 ( .A(q[6]), .B(DB[685]), .Z(n12432) );
  IV U17396 ( .A(n12431), .Z(n17175) );
  XNOR U17397 ( .A(n12429), .B(n17176), .Z(n12431) );
  XNOR U17398 ( .A(q[5]), .B(DB[684]), .Z(n17176) );
  XNOR U17399 ( .A(q[4]), .B(DB[683]), .Z(n12429) );
  IV U17400 ( .A(n12443), .Z(n17174) );
  XOR U17401 ( .A(n17177), .B(n17178), .Z(n12443) );
  XNOR U17402 ( .A(n12439), .B(n12441), .Z(n17178) );
  XNOR U17403 ( .A(q[0]), .B(DB[679]), .Z(n12441) );
  XNOR U17404 ( .A(q[3]), .B(DB[682]), .Z(n12439) );
  IV U17405 ( .A(n12438), .Z(n17177) );
  XNOR U17406 ( .A(n12436), .B(n17179), .Z(n12438) );
  XNOR U17407 ( .A(q[2]), .B(DB[681]), .Z(n17179) );
  XNOR U17408 ( .A(q[1]), .B(DB[680]), .Z(n12436) );
  XOR U17409 ( .A(n17180), .B(n12401), .Z(n12364) );
  XOR U17410 ( .A(n17181), .B(n12389), .Z(n12401) );
  XNOR U17411 ( .A(q[6]), .B(DB[692]), .Z(n12389) );
  IV U17412 ( .A(n12388), .Z(n17181) );
  XNOR U17413 ( .A(n12386), .B(n17182), .Z(n12388) );
  XNOR U17414 ( .A(q[5]), .B(DB[691]), .Z(n17182) );
  XNOR U17415 ( .A(q[4]), .B(DB[690]), .Z(n12386) );
  IV U17416 ( .A(n12400), .Z(n17180) );
  XOR U17417 ( .A(n17183), .B(n17184), .Z(n12400) );
  XNOR U17418 ( .A(n12396), .B(n12398), .Z(n17184) );
  XNOR U17419 ( .A(q[0]), .B(DB[686]), .Z(n12398) );
  XNOR U17420 ( .A(q[3]), .B(DB[689]), .Z(n12396) );
  IV U17421 ( .A(n12395), .Z(n17183) );
  XNOR U17422 ( .A(n12393), .B(n17185), .Z(n12395) );
  XNOR U17423 ( .A(q[2]), .B(DB[688]), .Z(n17185) );
  XNOR U17424 ( .A(q[1]), .B(DB[687]), .Z(n12393) );
  XOR U17425 ( .A(n17186), .B(n12358), .Z(n12321) );
  XOR U17426 ( .A(n17187), .B(n12346), .Z(n12358) );
  XNOR U17427 ( .A(q[6]), .B(DB[699]), .Z(n12346) );
  IV U17428 ( .A(n12345), .Z(n17187) );
  XNOR U17429 ( .A(n12343), .B(n17188), .Z(n12345) );
  XNOR U17430 ( .A(q[5]), .B(DB[698]), .Z(n17188) );
  XNOR U17431 ( .A(q[4]), .B(DB[697]), .Z(n12343) );
  IV U17432 ( .A(n12357), .Z(n17186) );
  XOR U17433 ( .A(n17189), .B(n17190), .Z(n12357) );
  XNOR U17434 ( .A(n12353), .B(n12355), .Z(n17190) );
  XNOR U17435 ( .A(q[0]), .B(DB[693]), .Z(n12355) );
  XNOR U17436 ( .A(q[3]), .B(DB[696]), .Z(n12353) );
  IV U17437 ( .A(n12352), .Z(n17189) );
  XNOR U17438 ( .A(n12350), .B(n17191), .Z(n12352) );
  XNOR U17439 ( .A(q[2]), .B(DB[695]), .Z(n17191) );
  XNOR U17440 ( .A(q[1]), .B(DB[694]), .Z(n12350) );
  XOR U17441 ( .A(n17192), .B(n12315), .Z(n12278) );
  XOR U17442 ( .A(n17193), .B(n12303), .Z(n12315) );
  XNOR U17443 ( .A(q[6]), .B(DB[706]), .Z(n12303) );
  IV U17444 ( .A(n12302), .Z(n17193) );
  XNOR U17445 ( .A(n12300), .B(n17194), .Z(n12302) );
  XNOR U17446 ( .A(q[5]), .B(DB[705]), .Z(n17194) );
  XNOR U17447 ( .A(q[4]), .B(DB[704]), .Z(n12300) );
  IV U17448 ( .A(n12314), .Z(n17192) );
  XOR U17449 ( .A(n17195), .B(n17196), .Z(n12314) );
  XNOR U17450 ( .A(n12310), .B(n12312), .Z(n17196) );
  XNOR U17451 ( .A(q[0]), .B(DB[700]), .Z(n12312) );
  XNOR U17452 ( .A(q[3]), .B(DB[703]), .Z(n12310) );
  IV U17453 ( .A(n12309), .Z(n17195) );
  XNOR U17454 ( .A(n12307), .B(n17197), .Z(n12309) );
  XNOR U17455 ( .A(q[2]), .B(DB[702]), .Z(n17197) );
  XNOR U17456 ( .A(q[1]), .B(DB[701]), .Z(n12307) );
  XOR U17457 ( .A(n17198), .B(n12272), .Z(n12235) );
  XOR U17458 ( .A(n17199), .B(n12260), .Z(n12272) );
  XNOR U17459 ( .A(q[6]), .B(DB[713]), .Z(n12260) );
  IV U17460 ( .A(n12259), .Z(n17199) );
  XNOR U17461 ( .A(n12257), .B(n17200), .Z(n12259) );
  XNOR U17462 ( .A(q[5]), .B(DB[712]), .Z(n17200) );
  XNOR U17463 ( .A(q[4]), .B(DB[711]), .Z(n12257) );
  IV U17464 ( .A(n12271), .Z(n17198) );
  XOR U17465 ( .A(n17201), .B(n17202), .Z(n12271) );
  XNOR U17466 ( .A(n12267), .B(n12269), .Z(n17202) );
  XNOR U17467 ( .A(q[0]), .B(DB[707]), .Z(n12269) );
  XNOR U17468 ( .A(q[3]), .B(DB[710]), .Z(n12267) );
  IV U17469 ( .A(n12266), .Z(n17201) );
  XNOR U17470 ( .A(n12264), .B(n17203), .Z(n12266) );
  XNOR U17471 ( .A(q[2]), .B(DB[709]), .Z(n17203) );
  XNOR U17472 ( .A(q[1]), .B(DB[708]), .Z(n12264) );
  XOR U17473 ( .A(n17204), .B(n12229), .Z(n12192) );
  XOR U17474 ( .A(n17205), .B(n12217), .Z(n12229) );
  XNOR U17475 ( .A(q[6]), .B(DB[720]), .Z(n12217) );
  IV U17476 ( .A(n12216), .Z(n17205) );
  XNOR U17477 ( .A(n12214), .B(n17206), .Z(n12216) );
  XNOR U17478 ( .A(q[5]), .B(DB[719]), .Z(n17206) );
  XNOR U17479 ( .A(q[4]), .B(DB[718]), .Z(n12214) );
  IV U17480 ( .A(n12228), .Z(n17204) );
  XOR U17481 ( .A(n17207), .B(n17208), .Z(n12228) );
  XNOR U17482 ( .A(n12224), .B(n12226), .Z(n17208) );
  XNOR U17483 ( .A(q[0]), .B(DB[714]), .Z(n12226) );
  XNOR U17484 ( .A(q[3]), .B(DB[717]), .Z(n12224) );
  IV U17485 ( .A(n12223), .Z(n17207) );
  XNOR U17486 ( .A(n12221), .B(n17209), .Z(n12223) );
  XNOR U17487 ( .A(q[2]), .B(DB[716]), .Z(n17209) );
  XNOR U17488 ( .A(q[1]), .B(DB[715]), .Z(n12221) );
  XOR U17489 ( .A(n17210), .B(n12186), .Z(n12149) );
  XOR U17490 ( .A(n17211), .B(n12174), .Z(n12186) );
  XNOR U17491 ( .A(q[6]), .B(DB[727]), .Z(n12174) );
  IV U17492 ( .A(n12173), .Z(n17211) );
  XNOR U17493 ( .A(n12171), .B(n17212), .Z(n12173) );
  XNOR U17494 ( .A(q[5]), .B(DB[726]), .Z(n17212) );
  XNOR U17495 ( .A(q[4]), .B(DB[725]), .Z(n12171) );
  IV U17496 ( .A(n12185), .Z(n17210) );
  XOR U17497 ( .A(n17213), .B(n17214), .Z(n12185) );
  XNOR U17498 ( .A(n12181), .B(n12183), .Z(n17214) );
  XNOR U17499 ( .A(q[0]), .B(DB[721]), .Z(n12183) );
  XNOR U17500 ( .A(q[3]), .B(DB[724]), .Z(n12181) );
  IV U17501 ( .A(n12180), .Z(n17213) );
  XNOR U17502 ( .A(n12178), .B(n17215), .Z(n12180) );
  XNOR U17503 ( .A(q[2]), .B(DB[723]), .Z(n17215) );
  XNOR U17504 ( .A(q[1]), .B(DB[722]), .Z(n12178) );
  XOR U17505 ( .A(n17216), .B(n12143), .Z(n12106) );
  XOR U17506 ( .A(n17217), .B(n12131), .Z(n12143) );
  XNOR U17507 ( .A(q[6]), .B(DB[734]), .Z(n12131) );
  IV U17508 ( .A(n12130), .Z(n17217) );
  XNOR U17509 ( .A(n12128), .B(n17218), .Z(n12130) );
  XNOR U17510 ( .A(q[5]), .B(DB[733]), .Z(n17218) );
  XNOR U17511 ( .A(q[4]), .B(DB[732]), .Z(n12128) );
  IV U17512 ( .A(n12142), .Z(n17216) );
  XOR U17513 ( .A(n17219), .B(n17220), .Z(n12142) );
  XNOR U17514 ( .A(n12138), .B(n12140), .Z(n17220) );
  XNOR U17515 ( .A(q[0]), .B(DB[728]), .Z(n12140) );
  XNOR U17516 ( .A(q[3]), .B(DB[731]), .Z(n12138) );
  IV U17517 ( .A(n12137), .Z(n17219) );
  XNOR U17518 ( .A(n12135), .B(n17221), .Z(n12137) );
  XNOR U17519 ( .A(q[2]), .B(DB[730]), .Z(n17221) );
  XNOR U17520 ( .A(q[1]), .B(DB[729]), .Z(n12135) );
  XOR U17521 ( .A(n17222), .B(n12100), .Z(n12063) );
  XOR U17522 ( .A(n17223), .B(n12088), .Z(n12100) );
  XNOR U17523 ( .A(q[6]), .B(DB[741]), .Z(n12088) );
  IV U17524 ( .A(n12087), .Z(n17223) );
  XNOR U17525 ( .A(n12085), .B(n17224), .Z(n12087) );
  XNOR U17526 ( .A(q[5]), .B(DB[740]), .Z(n17224) );
  XNOR U17527 ( .A(q[4]), .B(DB[739]), .Z(n12085) );
  IV U17528 ( .A(n12099), .Z(n17222) );
  XOR U17529 ( .A(n17225), .B(n17226), .Z(n12099) );
  XNOR U17530 ( .A(n12095), .B(n12097), .Z(n17226) );
  XNOR U17531 ( .A(q[0]), .B(DB[735]), .Z(n12097) );
  XNOR U17532 ( .A(q[3]), .B(DB[738]), .Z(n12095) );
  IV U17533 ( .A(n12094), .Z(n17225) );
  XNOR U17534 ( .A(n12092), .B(n17227), .Z(n12094) );
  XNOR U17535 ( .A(q[2]), .B(DB[737]), .Z(n17227) );
  XNOR U17536 ( .A(q[1]), .B(DB[736]), .Z(n12092) );
  XOR U17537 ( .A(n17228), .B(n12057), .Z(n12020) );
  XOR U17538 ( .A(n17229), .B(n12045), .Z(n12057) );
  XNOR U17539 ( .A(q[6]), .B(DB[748]), .Z(n12045) );
  IV U17540 ( .A(n12044), .Z(n17229) );
  XNOR U17541 ( .A(n12042), .B(n17230), .Z(n12044) );
  XNOR U17542 ( .A(q[5]), .B(DB[747]), .Z(n17230) );
  XNOR U17543 ( .A(q[4]), .B(DB[746]), .Z(n12042) );
  IV U17544 ( .A(n12056), .Z(n17228) );
  XOR U17545 ( .A(n17231), .B(n17232), .Z(n12056) );
  XNOR U17546 ( .A(n12052), .B(n12054), .Z(n17232) );
  XNOR U17547 ( .A(q[0]), .B(DB[742]), .Z(n12054) );
  XNOR U17548 ( .A(q[3]), .B(DB[745]), .Z(n12052) );
  IV U17549 ( .A(n12051), .Z(n17231) );
  XNOR U17550 ( .A(n12049), .B(n17233), .Z(n12051) );
  XNOR U17551 ( .A(q[2]), .B(DB[744]), .Z(n17233) );
  XNOR U17552 ( .A(q[1]), .B(DB[743]), .Z(n12049) );
  XOR U17553 ( .A(n17234), .B(n12014), .Z(n11977) );
  XOR U17554 ( .A(n17235), .B(n12002), .Z(n12014) );
  XNOR U17555 ( .A(q[6]), .B(DB[755]), .Z(n12002) );
  IV U17556 ( .A(n12001), .Z(n17235) );
  XNOR U17557 ( .A(n11999), .B(n17236), .Z(n12001) );
  XNOR U17558 ( .A(q[5]), .B(DB[754]), .Z(n17236) );
  XNOR U17559 ( .A(q[4]), .B(DB[753]), .Z(n11999) );
  IV U17560 ( .A(n12013), .Z(n17234) );
  XOR U17561 ( .A(n17237), .B(n17238), .Z(n12013) );
  XNOR U17562 ( .A(n12009), .B(n12011), .Z(n17238) );
  XNOR U17563 ( .A(q[0]), .B(DB[749]), .Z(n12011) );
  XNOR U17564 ( .A(q[3]), .B(DB[752]), .Z(n12009) );
  IV U17565 ( .A(n12008), .Z(n17237) );
  XNOR U17566 ( .A(n12006), .B(n17239), .Z(n12008) );
  XNOR U17567 ( .A(q[2]), .B(DB[751]), .Z(n17239) );
  XNOR U17568 ( .A(q[1]), .B(DB[750]), .Z(n12006) );
  XOR U17569 ( .A(n17240), .B(n11971), .Z(n11934) );
  XOR U17570 ( .A(n17241), .B(n11959), .Z(n11971) );
  XNOR U17571 ( .A(q[6]), .B(DB[762]), .Z(n11959) );
  IV U17572 ( .A(n11958), .Z(n17241) );
  XNOR U17573 ( .A(n11956), .B(n17242), .Z(n11958) );
  XNOR U17574 ( .A(q[5]), .B(DB[761]), .Z(n17242) );
  XNOR U17575 ( .A(q[4]), .B(DB[760]), .Z(n11956) );
  IV U17576 ( .A(n11970), .Z(n17240) );
  XOR U17577 ( .A(n17243), .B(n17244), .Z(n11970) );
  XNOR U17578 ( .A(n11966), .B(n11968), .Z(n17244) );
  XNOR U17579 ( .A(q[0]), .B(DB[756]), .Z(n11968) );
  XNOR U17580 ( .A(q[3]), .B(DB[759]), .Z(n11966) );
  IV U17581 ( .A(n11965), .Z(n17243) );
  XNOR U17582 ( .A(n11963), .B(n17245), .Z(n11965) );
  XNOR U17583 ( .A(q[2]), .B(DB[758]), .Z(n17245) );
  XNOR U17584 ( .A(q[1]), .B(DB[757]), .Z(n11963) );
  XOR U17585 ( .A(n17246), .B(n11928), .Z(n11891) );
  XOR U17586 ( .A(n17247), .B(n11916), .Z(n11928) );
  XNOR U17587 ( .A(q[6]), .B(DB[769]), .Z(n11916) );
  IV U17588 ( .A(n11915), .Z(n17247) );
  XNOR U17589 ( .A(n11913), .B(n17248), .Z(n11915) );
  XNOR U17590 ( .A(q[5]), .B(DB[768]), .Z(n17248) );
  XNOR U17591 ( .A(q[4]), .B(DB[767]), .Z(n11913) );
  IV U17592 ( .A(n11927), .Z(n17246) );
  XOR U17593 ( .A(n17249), .B(n17250), .Z(n11927) );
  XNOR U17594 ( .A(n11923), .B(n11925), .Z(n17250) );
  XNOR U17595 ( .A(q[0]), .B(DB[763]), .Z(n11925) );
  XNOR U17596 ( .A(q[3]), .B(DB[766]), .Z(n11923) );
  IV U17597 ( .A(n11922), .Z(n17249) );
  XNOR U17598 ( .A(n11920), .B(n17251), .Z(n11922) );
  XNOR U17599 ( .A(q[2]), .B(DB[765]), .Z(n17251) );
  XNOR U17600 ( .A(q[1]), .B(DB[764]), .Z(n11920) );
  XOR U17601 ( .A(n17252), .B(n11885), .Z(n11848) );
  XOR U17602 ( .A(n17253), .B(n11873), .Z(n11885) );
  XNOR U17603 ( .A(q[6]), .B(DB[776]), .Z(n11873) );
  IV U17604 ( .A(n11872), .Z(n17253) );
  XNOR U17605 ( .A(n11870), .B(n17254), .Z(n11872) );
  XNOR U17606 ( .A(q[5]), .B(DB[775]), .Z(n17254) );
  XNOR U17607 ( .A(q[4]), .B(DB[774]), .Z(n11870) );
  IV U17608 ( .A(n11884), .Z(n17252) );
  XOR U17609 ( .A(n17255), .B(n17256), .Z(n11884) );
  XNOR U17610 ( .A(n11880), .B(n11882), .Z(n17256) );
  XNOR U17611 ( .A(q[0]), .B(DB[770]), .Z(n11882) );
  XNOR U17612 ( .A(q[3]), .B(DB[773]), .Z(n11880) );
  IV U17613 ( .A(n11879), .Z(n17255) );
  XNOR U17614 ( .A(n11877), .B(n17257), .Z(n11879) );
  XNOR U17615 ( .A(q[2]), .B(DB[772]), .Z(n17257) );
  XNOR U17616 ( .A(q[1]), .B(DB[771]), .Z(n11877) );
  XOR U17617 ( .A(n17258), .B(n11842), .Z(n11805) );
  XOR U17618 ( .A(n17259), .B(n11830), .Z(n11842) );
  XNOR U17619 ( .A(q[6]), .B(DB[783]), .Z(n11830) );
  IV U17620 ( .A(n11829), .Z(n17259) );
  XNOR U17621 ( .A(n11827), .B(n17260), .Z(n11829) );
  XNOR U17622 ( .A(q[5]), .B(DB[782]), .Z(n17260) );
  XNOR U17623 ( .A(q[4]), .B(DB[781]), .Z(n11827) );
  IV U17624 ( .A(n11841), .Z(n17258) );
  XOR U17625 ( .A(n17261), .B(n17262), .Z(n11841) );
  XNOR U17626 ( .A(n11837), .B(n11839), .Z(n17262) );
  XNOR U17627 ( .A(q[0]), .B(DB[777]), .Z(n11839) );
  XNOR U17628 ( .A(q[3]), .B(DB[780]), .Z(n11837) );
  IV U17629 ( .A(n11836), .Z(n17261) );
  XNOR U17630 ( .A(n11834), .B(n17263), .Z(n11836) );
  XNOR U17631 ( .A(q[2]), .B(DB[779]), .Z(n17263) );
  XNOR U17632 ( .A(q[1]), .B(DB[778]), .Z(n11834) );
  XOR U17633 ( .A(n17264), .B(n11799), .Z(n11762) );
  XOR U17634 ( .A(n17265), .B(n11787), .Z(n11799) );
  XNOR U17635 ( .A(q[6]), .B(DB[790]), .Z(n11787) );
  IV U17636 ( .A(n11786), .Z(n17265) );
  XNOR U17637 ( .A(n11784), .B(n17266), .Z(n11786) );
  XNOR U17638 ( .A(q[5]), .B(DB[789]), .Z(n17266) );
  XNOR U17639 ( .A(q[4]), .B(DB[788]), .Z(n11784) );
  IV U17640 ( .A(n11798), .Z(n17264) );
  XOR U17641 ( .A(n17267), .B(n17268), .Z(n11798) );
  XNOR U17642 ( .A(n11794), .B(n11796), .Z(n17268) );
  XNOR U17643 ( .A(q[0]), .B(DB[784]), .Z(n11796) );
  XNOR U17644 ( .A(q[3]), .B(DB[787]), .Z(n11794) );
  IV U17645 ( .A(n11793), .Z(n17267) );
  XNOR U17646 ( .A(n11791), .B(n17269), .Z(n11793) );
  XNOR U17647 ( .A(q[2]), .B(DB[786]), .Z(n17269) );
  XNOR U17648 ( .A(q[1]), .B(DB[785]), .Z(n11791) );
  XOR U17649 ( .A(n17270), .B(n11756), .Z(n11719) );
  XOR U17650 ( .A(n17271), .B(n11744), .Z(n11756) );
  XNOR U17651 ( .A(q[6]), .B(DB[797]), .Z(n11744) );
  IV U17652 ( .A(n11743), .Z(n17271) );
  XNOR U17653 ( .A(n11741), .B(n17272), .Z(n11743) );
  XNOR U17654 ( .A(q[5]), .B(DB[796]), .Z(n17272) );
  XNOR U17655 ( .A(q[4]), .B(DB[795]), .Z(n11741) );
  IV U17656 ( .A(n11755), .Z(n17270) );
  XOR U17657 ( .A(n17273), .B(n17274), .Z(n11755) );
  XNOR U17658 ( .A(n11751), .B(n11753), .Z(n17274) );
  XNOR U17659 ( .A(q[0]), .B(DB[791]), .Z(n11753) );
  XNOR U17660 ( .A(q[3]), .B(DB[794]), .Z(n11751) );
  IV U17661 ( .A(n11750), .Z(n17273) );
  XNOR U17662 ( .A(n11748), .B(n17275), .Z(n11750) );
  XNOR U17663 ( .A(q[2]), .B(DB[793]), .Z(n17275) );
  XNOR U17664 ( .A(q[1]), .B(DB[792]), .Z(n11748) );
  XOR U17665 ( .A(n17276), .B(n11713), .Z(n11676) );
  XOR U17666 ( .A(n17277), .B(n11701), .Z(n11713) );
  XNOR U17667 ( .A(q[6]), .B(DB[804]), .Z(n11701) );
  IV U17668 ( .A(n11700), .Z(n17277) );
  XNOR U17669 ( .A(n11698), .B(n17278), .Z(n11700) );
  XNOR U17670 ( .A(q[5]), .B(DB[803]), .Z(n17278) );
  XNOR U17671 ( .A(q[4]), .B(DB[802]), .Z(n11698) );
  IV U17672 ( .A(n11712), .Z(n17276) );
  XOR U17673 ( .A(n17279), .B(n17280), .Z(n11712) );
  XNOR U17674 ( .A(n11708), .B(n11710), .Z(n17280) );
  XNOR U17675 ( .A(q[0]), .B(DB[798]), .Z(n11710) );
  XNOR U17676 ( .A(q[3]), .B(DB[801]), .Z(n11708) );
  IV U17677 ( .A(n11707), .Z(n17279) );
  XNOR U17678 ( .A(n11705), .B(n17281), .Z(n11707) );
  XNOR U17679 ( .A(q[2]), .B(DB[800]), .Z(n17281) );
  XNOR U17680 ( .A(q[1]), .B(DB[799]), .Z(n11705) );
  XOR U17681 ( .A(n17282), .B(n11670), .Z(n11633) );
  XOR U17682 ( .A(n17283), .B(n11658), .Z(n11670) );
  XNOR U17683 ( .A(q[6]), .B(DB[811]), .Z(n11658) );
  IV U17684 ( .A(n11657), .Z(n17283) );
  XNOR U17685 ( .A(n11655), .B(n17284), .Z(n11657) );
  XNOR U17686 ( .A(q[5]), .B(DB[810]), .Z(n17284) );
  XNOR U17687 ( .A(q[4]), .B(DB[809]), .Z(n11655) );
  IV U17688 ( .A(n11669), .Z(n17282) );
  XOR U17689 ( .A(n17285), .B(n17286), .Z(n11669) );
  XNOR U17690 ( .A(n11665), .B(n11667), .Z(n17286) );
  XNOR U17691 ( .A(q[0]), .B(DB[805]), .Z(n11667) );
  XNOR U17692 ( .A(q[3]), .B(DB[808]), .Z(n11665) );
  IV U17693 ( .A(n11664), .Z(n17285) );
  XNOR U17694 ( .A(n11662), .B(n17287), .Z(n11664) );
  XNOR U17695 ( .A(q[2]), .B(DB[807]), .Z(n17287) );
  XNOR U17696 ( .A(q[1]), .B(DB[806]), .Z(n11662) );
  XOR U17697 ( .A(n17288), .B(n11627), .Z(n11590) );
  XOR U17698 ( .A(n17289), .B(n11615), .Z(n11627) );
  XNOR U17699 ( .A(q[6]), .B(DB[818]), .Z(n11615) );
  IV U17700 ( .A(n11614), .Z(n17289) );
  XNOR U17701 ( .A(n11612), .B(n17290), .Z(n11614) );
  XNOR U17702 ( .A(q[5]), .B(DB[817]), .Z(n17290) );
  XNOR U17703 ( .A(q[4]), .B(DB[816]), .Z(n11612) );
  IV U17704 ( .A(n11626), .Z(n17288) );
  XOR U17705 ( .A(n17291), .B(n17292), .Z(n11626) );
  XNOR U17706 ( .A(n11622), .B(n11624), .Z(n17292) );
  XNOR U17707 ( .A(q[0]), .B(DB[812]), .Z(n11624) );
  XNOR U17708 ( .A(q[3]), .B(DB[815]), .Z(n11622) );
  IV U17709 ( .A(n11621), .Z(n17291) );
  XNOR U17710 ( .A(n11619), .B(n17293), .Z(n11621) );
  XNOR U17711 ( .A(q[2]), .B(DB[814]), .Z(n17293) );
  XNOR U17712 ( .A(q[1]), .B(DB[813]), .Z(n11619) );
  XOR U17713 ( .A(n17294), .B(n11584), .Z(n11547) );
  XOR U17714 ( .A(n17295), .B(n11572), .Z(n11584) );
  XNOR U17715 ( .A(q[6]), .B(DB[825]), .Z(n11572) );
  IV U17716 ( .A(n11571), .Z(n17295) );
  XNOR U17717 ( .A(n11569), .B(n17296), .Z(n11571) );
  XNOR U17718 ( .A(q[5]), .B(DB[824]), .Z(n17296) );
  XNOR U17719 ( .A(q[4]), .B(DB[823]), .Z(n11569) );
  IV U17720 ( .A(n11583), .Z(n17294) );
  XOR U17721 ( .A(n17297), .B(n17298), .Z(n11583) );
  XNOR U17722 ( .A(n11579), .B(n11581), .Z(n17298) );
  XNOR U17723 ( .A(q[0]), .B(DB[819]), .Z(n11581) );
  XNOR U17724 ( .A(q[3]), .B(DB[822]), .Z(n11579) );
  IV U17725 ( .A(n11578), .Z(n17297) );
  XNOR U17726 ( .A(n11576), .B(n17299), .Z(n11578) );
  XNOR U17727 ( .A(q[2]), .B(DB[821]), .Z(n17299) );
  XNOR U17728 ( .A(q[1]), .B(DB[820]), .Z(n11576) );
  XOR U17729 ( .A(n17300), .B(n11541), .Z(n11504) );
  XOR U17730 ( .A(n17301), .B(n11529), .Z(n11541) );
  XNOR U17731 ( .A(q[6]), .B(DB[832]), .Z(n11529) );
  IV U17732 ( .A(n11528), .Z(n17301) );
  XNOR U17733 ( .A(n11526), .B(n17302), .Z(n11528) );
  XNOR U17734 ( .A(q[5]), .B(DB[831]), .Z(n17302) );
  XNOR U17735 ( .A(q[4]), .B(DB[830]), .Z(n11526) );
  IV U17736 ( .A(n11540), .Z(n17300) );
  XOR U17737 ( .A(n17303), .B(n17304), .Z(n11540) );
  XNOR U17738 ( .A(n11536), .B(n11538), .Z(n17304) );
  XNOR U17739 ( .A(q[0]), .B(DB[826]), .Z(n11538) );
  XNOR U17740 ( .A(q[3]), .B(DB[829]), .Z(n11536) );
  IV U17741 ( .A(n11535), .Z(n17303) );
  XNOR U17742 ( .A(n11533), .B(n17305), .Z(n11535) );
  XNOR U17743 ( .A(q[2]), .B(DB[828]), .Z(n17305) );
  XNOR U17744 ( .A(q[1]), .B(DB[827]), .Z(n11533) );
  XOR U17745 ( .A(n17306), .B(n11498), .Z(n11461) );
  XOR U17746 ( .A(n17307), .B(n11486), .Z(n11498) );
  XNOR U17747 ( .A(q[6]), .B(DB[839]), .Z(n11486) );
  IV U17748 ( .A(n11485), .Z(n17307) );
  XNOR U17749 ( .A(n11483), .B(n17308), .Z(n11485) );
  XNOR U17750 ( .A(q[5]), .B(DB[838]), .Z(n17308) );
  XNOR U17751 ( .A(q[4]), .B(DB[837]), .Z(n11483) );
  IV U17752 ( .A(n11497), .Z(n17306) );
  XOR U17753 ( .A(n17309), .B(n17310), .Z(n11497) );
  XNOR U17754 ( .A(n11493), .B(n11495), .Z(n17310) );
  XNOR U17755 ( .A(q[0]), .B(DB[833]), .Z(n11495) );
  XNOR U17756 ( .A(q[3]), .B(DB[836]), .Z(n11493) );
  IV U17757 ( .A(n11492), .Z(n17309) );
  XNOR U17758 ( .A(n11490), .B(n17311), .Z(n11492) );
  XNOR U17759 ( .A(q[2]), .B(DB[835]), .Z(n17311) );
  XNOR U17760 ( .A(q[1]), .B(DB[834]), .Z(n11490) );
  XOR U17761 ( .A(n17312), .B(n11455), .Z(n11418) );
  XOR U17762 ( .A(n17313), .B(n11443), .Z(n11455) );
  XNOR U17763 ( .A(q[6]), .B(DB[846]), .Z(n11443) );
  IV U17764 ( .A(n11442), .Z(n17313) );
  XNOR U17765 ( .A(n11440), .B(n17314), .Z(n11442) );
  XNOR U17766 ( .A(q[5]), .B(DB[845]), .Z(n17314) );
  XNOR U17767 ( .A(q[4]), .B(DB[844]), .Z(n11440) );
  IV U17768 ( .A(n11454), .Z(n17312) );
  XOR U17769 ( .A(n17315), .B(n17316), .Z(n11454) );
  XNOR U17770 ( .A(n11450), .B(n11452), .Z(n17316) );
  XNOR U17771 ( .A(q[0]), .B(DB[840]), .Z(n11452) );
  XNOR U17772 ( .A(q[3]), .B(DB[843]), .Z(n11450) );
  IV U17773 ( .A(n11449), .Z(n17315) );
  XNOR U17774 ( .A(n11447), .B(n17317), .Z(n11449) );
  XNOR U17775 ( .A(q[2]), .B(DB[842]), .Z(n17317) );
  XNOR U17776 ( .A(q[1]), .B(DB[841]), .Z(n11447) );
  XOR U17777 ( .A(n17318), .B(n11412), .Z(n11375) );
  XOR U17778 ( .A(n17319), .B(n11400), .Z(n11412) );
  XNOR U17779 ( .A(q[6]), .B(DB[853]), .Z(n11400) );
  IV U17780 ( .A(n11399), .Z(n17319) );
  XNOR U17781 ( .A(n11397), .B(n17320), .Z(n11399) );
  XNOR U17782 ( .A(q[5]), .B(DB[852]), .Z(n17320) );
  XNOR U17783 ( .A(q[4]), .B(DB[851]), .Z(n11397) );
  IV U17784 ( .A(n11411), .Z(n17318) );
  XOR U17785 ( .A(n17321), .B(n17322), .Z(n11411) );
  XNOR U17786 ( .A(n11407), .B(n11409), .Z(n17322) );
  XNOR U17787 ( .A(q[0]), .B(DB[847]), .Z(n11409) );
  XNOR U17788 ( .A(q[3]), .B(DB[850]), .Z(n11407) );
  IV U17789 ( .A(n11406), .Z(n17321) );
  XNOR U17790 ( .A(n11404), .B(n17323), .Z(n11406) );
  XNOR U17791 ( .A(q[2]), .B(DB[849]), .Z(n17323) );
  XNOR U17792 ( .A(q[1]), .B(DB[848]), .Z(n11404) );
  XOR U17793 ( .A(n17324), .B(n11369), .Z(n11332) );
  XOR U17794 ( .A(n17325), .B(n11357), .Z(n11369) );
  XNOR U17795 ( .A(q[6]), .B(DB[860]), .Z(n11357) );
  IV U17796 ( .A(n11356), .Z(n17325) );
  XNOR U17797 ( .A(n11354), .B(n17326), .Z(n11356) );
  XNOR U17798 ( .A(q[5]), .B(DB[859]), .Z(n17326) );
  XNOR U17799 ( .A(q[4]), .B(DB[858]), .Z(n11354) );
  IV U17800 ( .A(n11368), .Z(n17324) );
  XOR U17801 ( .A(n17327), .B(n17328), .Z(n11368) );
  XNOR U17802 ( .A(n11364), .B(n11366), .Z(n17328) );
  XNOR U17803 ( .A(q[0]), .B(DB[854]), .Z(n11366) );
  XNOR U17804 ( .A(q[3]), .B(DB[857]), .Z(n11364) );
  IV U17805 ( .A(n11363), .Z(n17327) );
  XNOR U17806 ( .A(n11361), .B(n17329), .Z(n11363) );
  XNOR U17807 ( .A(q[2]), .B(DB[856]), .Z(n17329) );
  XNOR U17808 ( .A(q[1]), .B(DB[855]), .Z(n11361) );
  XOR U17809 ( .A(n17330), .B(n11326), .Z(n11289) );
  XOR U17810 ( .A(n17331), .B(n11314), .Z(n11326) );
  XNOR U17811 ( .A(q[6]), .B(DB[867]), .Z(n11314) );
  IV U17812 ( .A(n11313), .Z(n17331) );
  XNOR U17813 ( .A(n11311), .B(n17332), .Z(n11313) );
  XNOR U17814 ( .A(q[5]), .B(DB[866]), .Z(n17332) );
  XNOR U17815 ( .A(q[4]), .B(DB[865]), .Z(n11311) );
  IV U17816 ( .A(n11325), .Z(n17330) );
  XOR U17817 ( .A(n17333), .B(n17334), .Z(n11325) );
  XNOR U17818 ( .A(n11321), .B(n11323), .Z(n17334) );
  XNOR U17819 ( .A(q[0]), .B(DB[861]), .Z(n11323) );
  XNOR U17820 ( .A(q[3]), .B(DB[864]), .Z(n11321) );
  IV U17821 ( .A(n11320), .Z(n17333) );
  XNOR U17822 ( .A(n11318), .B(n17335), .Z(n11320) );
  XNOR U17823 ( .A(q[2]), .B(DB[863]), .Z(n17335) );
  XNOR U17824 ( .A(q[1]), .B(DB[862]), .Z(n11318) );
  XOR U17825 ( .A(n17336), .B(n11283), .Z(n11246) );
  XOR U17826 ( .A(n17337), .B(n11271), .Z(n11283) );
  XNOR U17827 ( .A(q[6]), .B(DB[874]), .Z(n11271) );
  IV U17828 ( .A(n11270), .Z(n17337) );
  XNOR U17829 ( .A(n11268), .B(n17338), .Z(n11270) );
  XNOR U17830 ( .A(q[5]), .B(DB[873]), .Z(n17338) );
  XNOR U17831 ( .A(q[4]), .B(DB[872]), .Z(n11268) );
  IV U17832 ( .A(n11282), .Z(n17336) );
  XOR U17833 ( .A(n17339), .B(n17340), .Z(n11282) );
  XNOR U17834 ( .A(n11278), .B(n11280), .Z(n17340) );
  XNOR U17835 ( .A(q[0]), .B(DB[868]), .Z(n11280) );
  XNOR U17836 ( .A(q[3]), .B(DB[871]), .Z(n11278) );
  IV U17837 ( .A(n11277), .Z(n17339) );
  XNOR U17838 ( .A(n11275), .B(n17341), .Z(n11277) );
  XNOR U17839 ( .A(q[2]), .B(DB[870]), .Z(n17341) );
  XNOR U17840 ( .A(q[1]), .B(DB[869]), .Z(n11275) );
  XOR U17841 ( .A(n17342), .B(n11240), .Z(n11203) );
  XOR U17842 ( .A(n17343), .B(n11228), .Z(n11240) );
  XNOR U17843 ( .A(q[6]), .B(DB[881]), .Z(n11228) );
  IV U17844 ( .A(n11227), .Z(n17343) );
  XNOR U17845 ( .A(n11225), .B(n17344), .Z(n11227) );
  XNOR U17846 ( .A(q[5]), .B(DB[880]), .Z(n17344) );
  XNOR U17847 ( .A(q[4]), .B(DB[879]), .Z(n11225) );
  IV U17848 ( .A(n11239), .Z(n17342) );
  XOR U17849 ( .A(n17345), .B(n17346), .Z(n11239) );
  XNOR U17850 ( .A(n11235), .B(n11237), .Z(n17346) );
  XNOR U17851 ( .A(q[0]), .B(DB[875]), .Z(n11237) );
  XNOR U17852 ( .A(q[3]), .B(DB[878]), .Z(n11235) );
  IV U17853 ( .A(n11234), .Z(n17345) );
  XNOR U17854 ( .A(n11232), .B(n17347), .Z(n11234) );
  XNOR U17855 ( .A(q[2]), .B(DB[877]), .Z(n17347) );
  XNOR U17856 ( .A(q[1]), .B(DB[876]), .Z(n11232) );
  XOR U17857 ( .A(n17348), .B(n11197), .Z(n11160) );
  XOR U17858 ( .A(n17349), .B(n11185), .Z(n11197) );
  XNOR U17859 ( .A(q[6]), .B(DB[888]), .Z(n11185) );
  IV U17860 ( .A(n11184), .Z(n17349) );
  XNOR U17861 ( .A(n11182), .B(n17350), .Z(n11184) );
  XNOR U17862 ( .A(q[5]), .B(DB[887]), .Z(n17350) );
  XNOR U17863 ( .A(q[4]), .B(DB[886]), .Z(n11182) );
  IV U17864 ( .A(n11196), .Z(n17348) );
  XOR U17865 ( .A(n17351), .B(n17352), .Z(n11196) );
  XNOR U17866 ( .A(n11192), .B(n11194), .Z(n17352) );
  XNOR U17867 ( .A(q[0]), .B(DB[882]), .Z(n11194) );
  XNOR U17868 ( .A(q[3]), .B(DB[885]), .Z(n11192) );
  IV U17869 ( .A(n11191), .Z(n17351) );
  XNOR U17870 ( .A(n11189), .B(n17353), .Z(n11191) );
  XNOR U17871 ( .A(q[2]), .B(DB[884]), .Z(n17353) );
  XNOR U17872 ( .A(q[1]), .B(DB[883]), .Z(n11189) );
  XOR U17873 ( .A(n17354), .B(n11154), .Z(n11117) );
  XOR U17874 ( .A(n17355), .B(n11142), .Z(n11154) );
  XNOR U17875 ( .A(q[6]), .B(DB[895]), .Z(n11142) );
  IV U17876 ( .A(n11141), .Z(n17355) );
  XNOR U17877 ( .A(n11139), .B(n17356), .Z(n11141) );
  XNOR U17878 ( .A(q[5]), .B(DB[894]), .Z(n17356) );
  XNOR U17879 ( .A(q[4]), .B(DB[893]), .Z(n11139) );
  IV U17880 ( .A(n11153), .Z(n17354) );
  XOR U17881 ( .A(n17357), .B(n17358), .Z(n11153) );
  XNOR U17882 ( .A(n11149), .B(n11151), .Z(n17358) );
  XNOR U17883 ( .A(q[0]), .B(DB[889]), .Z(n11151) );
  XNOR U17884 ( .A(q[3]), .B(DB[892]), .Z(n11149) );
  IV U17885 ( .A(n11148), .Z(n17357) );
  XNOR U17886 ( .A(n11146), .B(n17359), .Z(n11148) );
  XNOR U17887 ( .A(q[2]), .B(DB[891]), .Z(n17359) );
  XNOR U17888 ( .A(q[1]), .B(DB[890]), .Z(n11146) );
  XOR U17889 ( .A(n17360), .B(n11111), .Z(n11074) );
  XOR U17890 ( .A(n17361), .B(n11099), .Z(n11111) );
  XNOR U17891 ( .A(q[6]), .B(DB[902]), .Z(n11099) );
  IV U17892 ( .A(n11098), .Z(n17361) );
  XNOR U17893 ( .A(n11096), .B(n17362), .Z(n11098) );
  XNOR U17894 ( .A(q[5]), .B(DB[901]), .Z(n17362) );
  XNOR U17895 ( .A(q[4]), .B(DB[900]), .Z(n11096) );
  IV U17896 ( .A(n11110), .Z(n17360) );
  XOR U17897 ( .A(n17363), .B(n17364), .Z(n11110) );
  XNOR U17898 ( .A(n11106), .B(n11108), .Z(n17364) );
  XNOR U17899 ( .A(q[0]), .B(DB[896]), .Z(n11108) );
  XNOR U17900 ( .A(q[3]), .B(DB[899]), .Z(n11106) );
  IV U17901 ( .A(n11105), .Z(n17363) );
  XNOR U17902 ( .A(n11103), .B(n17365), .Z(n11105) );
  XNOR U17903 ( .A(q[2]), .B(DB[898]), .Z(n17365) );
  XNOR U17904 ( .A(q[1]), .B(DB[897]), .Z(n11103) );
  XOR U17905 ( .A(n17366), .B(n11068), .Z(n11031) );
  XOR U17906 ( .A(n17367), .B(n11056), .Z(n11068) );
  XNOR U17907 ( .A(q[6]), .B(DB[909]), .Z(n11056) );
  IV U17908 ( .A(n11055), .Z(n17367) );
  XNOR U17909 ( .A(n11053), .B(n17368), .Z(n11055) );
  XNOR U17910 ( .A(q[5]), .B(DB[908]), .Z(n17368) );
  XNOR U17911 ( .A(q[4]), .B(DB[907]), .Z(n11053) );
  IV U17912 ( .A(n11067), .Z(n17366) );
  XOR U17913 ( .A(n17369), .B(n17370), .Z(n11067) );
  XNOR U17914 ( .A(n11063), .B(n11065), .Z(n17370) );
  XNOR U17915 ( .A(q[0]), .B(DB[903]), .Z(n11065) );
  XNOR U17916 ( .A(q[3]), .B(DB[906]), .Z(n11063) );
  IV U17917 ( .A(n11062), .Z(n17369) );
  XNOR U17918 ( .A(n11060), .B(n17371), .Z(n11062) );
  XNOR U17919 ( .A(q[2]), .B(DB[905]), .Z(n17371) );
  XNOR U17920 ( .A(q[1]), .B(DB[904]), .Z(n11060) );
  XOR U17921 ( .A(n17372), .B(n11025), .Z(n10988) );
  XOR U17922 ( .A(n17373), .B(n11013), .Z(n11025) );
  XNOR U17923 ( .A(q[6]), .B(DB[916]), .Z(n11013) );
  IV U17924 ( .A(n11012), .Z(n17373) );
  XNOR U17925 ( .A(n11010), .B(n17374), .Z(n11012) );
  XNOR U17926 ( .A(q[5]), .B(DB[915]), .Z(n17374) );
  XNOR U17927 ( .A(q[4]), .B(DB[914]), .Z(n11010) );
  IV U17928 ( .A(n11024), .Z(n17372) );
  XOR U17929 ( .A(n17375), .B(n17376), .Z(n11024) );
  XNOR U17930 ( .A(n11020), .B(n11022), .Z(n17376) );
  XNOR U17931 ( .A(q[0]), .B(DB[910]), .Z(n11022) );
  XNOR U17932 ( .A(q[3]), .B(DB[913]), .Z(n11020) );
  IV U17933 ( .A(n11019), .Z(n17375) );
  XNOR U17934 ( .A(n11017), .B(n17377), .Z(n11019) );
  XNOR U17935 ( .A(q[2]), .B(DB[912]), .Z(n17377) );
  XNOR U17936 ( .A(q[1]), .B(DB[911]), .Z(n11017) );
  XOR U17937 ( .A(n17378), .B(n10982), .Z(n10945) );
  XOR U17938 ( .A(n17379), .B(n10970), .Z(n10982) );
  XNOR U17939 ( .A(q[6]), .B(DB[923]), .Z(n10970) );
  IV U17940 ( .A(n10969), .Z(n17379) );
  XNOR U17941 ( .A(n10967), .B(n17380), .Z(n10969) );
  XNOR U17942 ( .A(q[5]), .B(DB[922]), .Z(n17380) );
  XNOR U17943 ( .A(q[4]), .B(DB[921]), .Z(n10967) );
  IV U17944 ( .A(n10981), .Z(n17378) );
  XOR U17945 ( .A(n17381), .B(n17382), .Z(n10981) );
  XNOR U17946 ( .A(n10977), .B(n10979), .Z(n17382) );
  XNOR U17947 ( .A(q[0]), .B(DB[917]), .Z(n10979) );
  XNOR U17948 ( .A(q[3]), .B(DB[920]), .Z(n10977) );
  IV U17949 ( .A(n10976), .Z(n17381) );
  XNOR U17950 ( .A(n10974), .B(n17383), .Z(n10976) );
  XNOR U17951 ( .A(q[2]), .B(DB[919]), .Z(n17383) );
  XNOR U17952 ( .A(q[1]), .B(DB[918]), .Z(n10974) );
  XOR U17953 ( .A(n17384), .B(n10939), .Z(n10902) );
  XOR U17954 ( .A(n17385), .B(n10927), .Z(n10939) );
  XNOR U17955 ( .A(q[6]), .B(DB[930]), .Z(n10927) );
  IV U17956 ( .A(n10926), .Z(n17385) );
  XNOR U17957 ( .A(n10924), .B(n17386), .Z(n10926) );
  XNOR U17958 ( .A(q[5]), .B(DB[929]), .Z(n17386) );
  XNOR U17959 ( .A(q[4]), .B(DB[928]), .Z(n10924) );
  IV U17960 ( .A(n10938), .Z(n17384) );
  XOR U17961 ( .A(n17387), .B(n17388), .Z(n10938) );
  XNOR U17962 ( .A(n10934), .B(n10936), .Z(n17388) );
  XNOR U17963 ( .A(q[0]), .B(DB[924]), .Z(n10936) );
  XNOR U17964 ( .A(q[3]), .B(DB[927]), .Z(n10934) );
  IV U17965 ( .A(n10933), .Z(n17387) );
  XNOR U17966 ( .A(n10931), .B(n17389), .Z(n10933) );
  XNOR U17967 ( .A(q[2]), .B(DB[926]), .Z(n17389) );
  XNOR U17968 ( .A(q[1]), .B(DB[925]), .Z(n10931) );
  XOR U17969 ( .A(n17390), .B(n10896), .Z(n10859) );
  XOR U17970 ( .A(n17391), .B(n10884), .Z(n10896) );
  XNOR U17971 ( .A(q[6]), .B(DB[937]), .Z(n10884) );
  IV U17972 ( .A(n10883), .Z(n17391) );
  XNOR U17973 ( .A(n10881), .B(n17392), .Z(n10883) );
  XNOR U17974 ( .A(q[5]), .B(DB[936]), .Z(n17392) );
  XNOR U17975 ( .A(q[4]), .B(DB[935]), .Z(n10881) );
  IV U17976 ( .A(n10895), .Z(n17390) );
  XOR U17977 ( .A(n17393), .B(n17394), .Z(n10895) );
  XNOR U17978 ( .A(n10891), .B(n10893), .Z(n17394) );
  XNOR U17979 ( .A(q[0]), .B(DB[931]), .Z(n10893) );
  XNOR U17980 ( .A(q[3]), .B(DB[934]), .Z(n10891) );
  IV U17981 ( .A(n10890), .Z(n17393) );
  XNOR U17982 ( .A(n10888), .B(n17395), .Z(n10890) );
  XNOR U17983 ( .A(q[2]), .B(DB[933]), .Z(n17395) );
  XNOR U17984 ( .A(q[1]), .B(DB[932]), .Z(n10888) );
  XOR U17985 ( .A(n17396), .B(n10853), .Z(n10816) );
  XOR U17986 ( .A(n17397), .B(n10841), .Z(n10853) );
  XNOR U17987 ( .A(q[6]), .B(DB[944]), .Z(n10841) );
  IV U17988 ( .A(n10840), .Z(n17397) );
  XNOR U17989 ( .A(n10838), .B(n17398), .Z(n10840) );
  XNOR U17990 ( .A(q[5]), .B(DB[943]), .Z(n17398) );
  XNOR U17991 ( .A(q[4]), .B(DB[942]), .Z(n10838) );
  IV U17992 ( .A(n10852), .Z(n17396) );
  XOR U17993 ( .A(n17399), .B(n17400), .Z(n10852) );
  XNOR U17994 ( .A(n10848), .B(n10850), .Z(n17400) );
  XNOR U17995 ( .A(q[0]), .B(DB[938]), .Z(n10850) );
  XNOR U17996 ( .A(q[3]), .B(DB[941]), .Z(n10848) );
  IV U17997 ( .A(n10847), .Z(n17399) );
  XNOR U17998 ( .A(n10845), .B(n17401), .Z(n10847) );
  XNOR U17999 ( .A(q[2]), .B(DB[940]), .Z(n17401) );
  XNOR U18000 ( .A(q[1]), .B(DB[939]), .Z(n10845) );
  XOR U18001 ( .A(n17402), .B(n10810), .Z(n10773) );
  XOR U18002 ( .A(n17403), .B(n10798), .Z(n10810) );
  XNOR U18003 ( .A(q[6]), .B(DB[951]), .Z(n10798) );
  IV U18004 ( .A(n10797), .Z(n17403) );
  XNOR U18005 ( .A(n10795), .B(n17404), .Z(n10797) );
  XNOR U18006 ( .A(q[5]), .B(DB[950]), .Z(n17404) );
  XNOR U18007 ( .A(q[4]), .B(DB[949]), .Z(n10795) );
  IV U18008 ( .A(n10809), .Z(n17402) );
  XOR U18009 ( .A(n17405), .B(n17406), .Z(n10809) );
  XNOR U18010 ( .A(n10805), .B(n10807), .Z(n17406) );
  XNOR U18011 ( .A(q[0]), .B(DB[945]), .Z(n10807) );
  XNOR U18012 ( .A(q[3]), .B(DB[948]), .Z(n10805) );
  IV U18013 ( .A(n10804), .Z(n17405) );
  XNOR U18014 ( .A(n10802), .B(n17407), .Z(n10804) );
  XNOR U18015 ( .A(q[2]), .B(DB[947]), .Z(n17407) );
  XNOR U18016 ( .A(q[1]), .B(DB[946]), .Z(n10802) );
  XOR U18017 ( .A(n17408), .B(n10767), .Z(n10730) );
  XOR U18018 ( .A(n17409), .B(n10755), .Z(n10767) );
  XNOR U18019 ( .A(q[6]), .B(DB[958]), .Z(n10755) );
  IV U18020 ( .A(n10754), .Z(n17409) );
  XNOR U18021 ( .A(n10752), .B(n17410), .Z(n10754) );
  XNOR U18022 ( .A(q[5]), .B(DB[957]), .Z(n17410) );
  XNOR U18023 ( .A(q[4]), .B(DB[956]), .Z(n10752) );
  IV U18024 ( .A(n10766), .Z(n17408) );
  XOR U18025 ( .A(n17411), .B(n17412), .Z(n10766) );
  XNOR U18026 ( .A(n10762), .B(n10764), .Z(n17412) );
  XNOR U18027 ( .A(q[0]), .B(DB[952]), .Z(n10764) );
  XNOR U18028 ( .A(q[3]), .B(DB[955]), .Z(n10762) );
  IV U18029 ( .A(n10761), .Z(n17411) );
  XNOR U18030 ( .A(n10759), .B(n17413), .Z(n10761) );
  XNOR U18031 ( .A(q[2]), .B(DB[954]), .Z(n17413) );
  XNOR U18032 ( .A(q[1]), .B(DB[953]), .Z(n10759) );
  XOR U18033 ( .A(n17414), .B(n10724), .Z(n10687) );
  XOR U18034 ( .A(n17415), .B(n10712), .Z(n10724) );
  XNOR U18035 ( .A(q[6]), .B(DB[965]), .Z(n10712) );
  IV U18036 ( .A(n10711), .Z(n17415) );
  XNOR U18037 ( .A(n10709), .B(n17416), .Z(n10711) );
  XNOR U18038 ( .A(q[5]), .B(DB[964]), .Z(n17416) );
  XNOR U18039 ( .A(q[4]), .B(DB[963]), .Z(n10709) );
  IV U18040 ( .A(n10723), .Z(n17414) );
  XOR U18041 ( .A(n17417), .B(n17418), .Z(n10723) );
  XNOR U18042 ( .A(n10719), .B(n10721), .Z(n17418) );
  XNOR U18043 ( .A(q[0]), .B(DB[959]), .Z(n10721) );
  XNOR U18044 ( .A(q[3]), .B(DB[962]), .Z(n10719) );
  IV U18045 ( .A(n10718), .Z(n17417) );
  XNOR U18046 ( .A(n10716), .B(n17419), .Z(n10718) );
  XNOR U18047 ( .A(q[2]), .B(DB[961]), .Z(n17419) );
  XNOR U18048 ( .A(q[1]), .B(DB[960]), .Z(n10716) );
  XOR U18049 ( .A(n17420), .B(n10681), .Z(n10644) );
  XOR U18050 ( .A(n17421), .B(n10669), .Z(n10681) );
  XNOR U18051 ( .A(q[6]), .B(DB[972]), .Z(n10669) );
  IV U18052 ( .A(n10668), .Z(n17421) );
  XNOR U18053 ( .A(n10666), .B(n17422), .Z(n10668) );
  XNOR U18054 ( .A(q[5]), .B(DB[971]), .Z(n17422) );
  XNOR U18055 ( .A(q[4]), .B(DB[970]), .Z(n10666) );
  IV U18056 ( .A(n10680), .Z(n17420) );
  XOR U18057 ( .A(n17423), .B(n17424), .Z(n10680) );
  XNOR U18058 ( .A(n10676), .B(n10678), .Z(n17424) );
  XNOR U18059 ( .A(q[0]), .B(DB[966]), .Z(n10678) );
  XNOR U18060 ( .A(q[3]), .B(DB[969]), .Z(n10676) );
  IV U18061 ( .A(n10675), .Z(n17423) );
  XNOR U18062 ( .A(n10673), .B(n17425), .Z(n10675) );
  XNOR U18063 ( .A(q[2]), .B(DB[968]), .Z(n17425) );
  XNOR U18064 ( .A(q[1]), .B(DB[967]), .Z(n10673) );
  XOR U18065 ( .A(n17426), .B(n10638), .Z(n10601) );
  XOR U18066 ( .A(n17427), .B(n10626), .Z(n10638) );
  XNOR U18067 ( .A(q[6]), .B(DB[979]), .Z(n10626) );
  IV U18068 ( .A(n10625), .Z(n17427) );
  XNOR U18069 ( .A(n10623), .B(n17428), .Z(n10625) );
  XNOR U18070 ( .A(q[5]), .B(DB[978]), .Z(n17428) );
  XNOR U18071 ( .A(q[4]), .B(DB[977]), .Z(n10623) );
  IV U18072 ( .A(n10637), .Z(n17426) );
  XOR U18073 ( .A(n17429), .B(n17430), .Z(n10637) );
  XNOR U18074 ( .A(n10633), .B(n10635), .Z(n17430) );
  XNOR U18075 ( .A(q[0]), .B(DB[973]), .Z(n10635) );
  XNOR U18076 ( .A(q[3]), .B(DB[976]), .Z(n10633) );
  IV U18077 ( .A(n10632), .Z(n17429) );
  XNOR U18078 ( .A(n10630), .B(n17431), .Z(n10632) );
  XNOR U18079 ( .A(q[2]), .B(DB[975]), .Z(n17431) );
  XNOR U18080 ( .A(q[1]), .B(DB[974]), .Z(n10630) );
  XOR U18081 ( .A(n17432), .B(n10595), .Z(n10558) );
  XOR U18082 ( .A(n17433), .B(n10583), .Z(n10595) );
  XNOR U18083 ( .A(q[6]), .B(DB[986]), .Z(n10583) );
  IV U18084 ( .A(n10582), .Z(n17433) );
  XNOR U18085 ( .A(n10580), .B(n17434), .Z(n10582) );
  XNOR U18086 ( .A(q[5]), .B(DB[985]), .Z(n17434) );
  XNOR U18087 ( .A(q[4]), .B(DB[984]), .Z(n10580) );
  IV U18088 ( .A(n10594), .Z(n17432) );
  XOR U18089 ( .A(n17435), .B(n17436), .Z(n10594) );
  XNOR U18090 ( .A(n10590), .B(n10592), .Z(n17436) );
  XNOR U18091 ( .A(q[0]), .B(DB[980]), .Z(n10592) );
  XNOR U18092 ( .A(q[3]), .B(DB[983]), .Z(n10590) );
  IV U18093 ( .A(n10589), .Z(n17435) );
  XNOR U18094 ( .A(n10587), .B(n17437), .Z(n10589) );
  XNOR U18095 ( .A(q[2]), .B(DB[982]), .Z(n17437) );
  XNOR U18096 ( .A(q[1]), .B(DB[981]), .Z(n10587) );
  XOR U18097 ( .A(n17438), .B(n10552), .Z(n10515) );
  XOR U18098 ( .A(n17439), .B(n10540), .Z(n10552) );
  XNOR U18099 ( .A(q[6]), .B(DB[993]), .Z(n10540) );
  IV U18100 ( .A(n10539), .Z(n17439) );
  XNOR U18101 ( .A(n10537), .B(n17440), .Z(n10539) );
  XNOR U18102 ( .A(q[5]), .B(DB[992]), .Z(n17440) );
  XNOR U18103 ( .A(q[4]), .B(DB[991]), .Z(n10537) );
  IV U18104 ( .A(n10551), .Z(n17438) );
  XOR U18105 ( .A(n17441), .B(n17442), .Z(n10551) );
  XNOR U18106 ( .A(n10547), .B(n10549), .Z(n17442) );
  XNOR U18107 ( .A(q[0]), .B(DB[987]), .Z(n10549) );
  XNOR U18108 ( .A(q[3]), .B(DB[990]), .Z(n10547) );
  IV U18109 ( .A(n10546), .Z(n17441) );
  XNOR U18110 ( .A(n10544), .B(n17443), .Z(n10546) );
  XNOR U18111 ( .A(q[2]), .B(DB[989]), .Z(n17443) );
  XNOR U18112 ( .A(q[1]), .B(DB[988]), .Z(n10544) );
  XOR U18113 ( .A(n17444), .B(n10509), .Z(n10472) );
  XOR U18114 ( .A(n17445), .B(n10497), .Z(n10509) );
  XNOR U18115 ( .A(q[6]), .B(DB[1000]), .Z(n10497) );
  IV U18116 ( .A(n10496), .Z(n17445) );
  XNOR U18117 ( .A(n10494), .B(n17446), .Z(n10496) );
  XNOR U18118 ( .A(q[5]), .B(DB[999]), .Z(n17446) );
  XNOR U18119 ( .A(q[4]), .B(DB[998]), .Z(n10494) );
  IV U18120 ( .A(n10508), .Z(n17444) );
  XOR U18121 ( .A(n17447), .B(n17448), .Z(n10508) );
  XNOR U18122 ( .A(n10504), .B(n10506), .Z(n17448) );
  XNOR U18123 ( .A(q[0]), .B(DB[994]), .Z(n10506) );
  XNOR U18124 ( .A(q[3]), .B(DB[997]), .Z(n10504) );
  IV U18125 ( .A(n10503), .Z(n17447) );
  XNOR U18126 ( .A(n10501), .B(n17449), .Z(n10503) );
  XNOR U18127 ( .A(q[2]), .B(DB[996]), .Z(n17449) );
  XNOR U18128 ( .A(q[1]), .B(DB[995]), .Z(n10501) );
  XOR U18129 ( .A(n17450), .B(n10466), .Z(n10429) );
  XOR U18130 ( .A(n17451), .B(n10454), .Z(n10466) );
  XNOR U18131 ( .A(q[6]), .B(DB[1007]), .Z(n10454) );
  IV U18132 ( .A(n10453), .Z(n17451) );
  XNOR U18133 ( .A(n10451), .B(n17452), .Z(n10453) );
  XNOR U18134 ( .A(q[5]), .B(DB[1006]), .Z(n17452) );
  XNOR U18135 ( .A(q[4]), .B(DB[1005]), .Z(n10451) );
  IV U18136 ( .A(n10465), .Z(n17450) );
  XOR U18137 ( .A(n17453), .B(n17454), .Z(n10465) );
  XNOR U18138 ( .A(n10461), .B(n10463), .Z(n17454) );
  XNOR U18139 ( .A(q[0]), .B(DB[1001]), .Z(n10463) );
  XNOR U18140 ( .A(q[3]), .B(DB[1004]), .Z(n10461) );
  IV U18141 ( .A(n10460), .Z(n17453) );
  XNOR U18142 ( .A(n10458), .B(n17455), .Z(n10460) );
  XNOR U18143 ( .A(q[2]), .B(DB[1003]), .Z(n17455) );
  XNOR U18144 ( .A(q[1]), .B(DB[1002]), .Z(n10458) );
  XOR U18145 ( .A(n17456), .B(n10423), .Z(n10386) );
  XOR U18146 ( .A(n17457), .B(n10411), .Z(n10423) );
  XNOR U18147 ( .A(q[6]), .B(DB[1014]), .Z(n10411) );
  IV U18148 ( .A(n10410), .Z(n17457) );
  XNOR U18149 ( .A(n10408), .B(n17458), .Z(n10410) );
  XNOR U18150 ( .A(q[5]), .B(DB[1013]), .Z(n17458) );
  XNOR U18151 ( .A(q[4]), .B(DB[1012]), .Z(n10408) );
  IV U18152 ( .A(n10422), .Z(n17456) );
  XOR U18153 ( .A(n17459), .B(n17460), .Z(n10422) );
  XNOR U18154 ( .A(n10418), .B(n10420), .Z(n17460) );
  XNOR U18155 ( .A(q[0]), .B(DB[1008]), .Z(n10420) );
  XNOR U18156 ( .A(q[3]), .B(DB[1011]), .Z(n10418) );
  IV U18157 ( .A(n10417), .Z(n17459) );
  XNOR U18158 ( .A(n10415), .B(n17461), .Z(n10417) );
  XNOR U18159 ( .A(q[2]), .B(DB[1010]), .Z(n17461) );
  XNOR U18160 ( .A(q[1]), .B(DB[1009]), .Z(n10415) );
  XOR U18161 ( .A(n17462), .B(n10380), .Z(n10343) );
  XOR U18162 ( .A(n17463), .B(n10368), .Z(n10380) );
  XNOR U18163 ( .A(q[6]), .B(DB[1021]), .Z(n10368) );
  IV U18164 ( .A(n10367), .Z(n17463) );
  XNOR U18165 ( .A(n10365), .B(n17464), .Z(n10367) );
  XNOR U18166 ( .A(q[5]), .B(DB[1020]), .Z(n17464) );
  XNOR U18167 ( .A(q[4]), .B(DB[1019]), .Z(n10365) );
  IV U18168 ( .A(n10379), .Z(n17462) );
  XOR U18169 ( .A(n17465), .B(n17466), .Z(n10379) );
  XNOR U18170 ( .A(n10375), .B(n10377), .Z(n17466) );
  XNOR U18171 ( .A(q[0]), .B(DB[1015]), .Z(n10377) );
  XNOR U18172 ( .A(q[3]), .B(DB[1018]), .Z(n10375) );
  IV U18173 ( .A(n10374), .Z(n17465) );
  XNOR U18174 ( .A(n10372), .B(n17467), .Z(n10374) );
  XNOR U18175 ( .A(q[2]), .B(DB[1017]), .Z(n17467) );
  XNOR U18176 ( .A(q[1]), .B(DB[1016]), .Z(n10372) );
  XOR U18177 ( .A(n17468), .B(n10337), .Z(n10300) );
  XOR U18178 ( .A(n17469), .B(n10325), .Z(n10337) );
  XNOR U18179 ( .A(q[6]), .B(DB[1028]), .Z(n10325) );
  IV U18180 ( .A(n10324), .Z(n17469) );
  XNOR U18181 ( .A(n10322), .B(n17470), .Z(n10324) );
  XNOR U18182 ( .A(q[5]), .B(DB[1027]), .Z(n17470) );
  XNOR U18183 ( .A(q[4]), .B(DB[1026]), .Z(n10322) );
  IV U18184 ( .A(n10336), .Z(n17468) );
  XOR U18185 ( .A(n17471), .B(n17472), .Z(n10336) );
  XNOR U18186 ( .A(n10332), .B(n10334), .Z(n17472) );
  XNOR U18187 ( .A(q[0]), .B(DB[1022]), .Z(n10334) );
  XNOR U18188 ( .A(q[3]), .B(DB[1025]), .Z(n10332) );
  IV U18189 ( .A(n10331), .Z(n17471) );
  XNOR U18190 ( .A(n10329), .B(n17473), .Z(n10331) );
  XNOR U18191 ( .A(q[2]), .B(DB[1024]), .Z(n17473) );
  XNOR U18192 ( .A(q[1]), .B(DB[1023]), .Z(n10329) );
  XOR U18193 ( .A(n17474), .B(n10294), .Z(n10257) );
  XOR U18194 ( .A(n17475), .B(n10282), .Z(n10294) );
  XNOR U18195 ( .A(q[6]), .B(DB[1035]), .Z(n10282) );
  IV U18196 ( .A(n10281), .Z(n17475) );
  XNOR U18197 ( .A(n10279), .B(n17476), .Z(n10281) );
  XNOR U18198 ( .A(q[5]), .B(DB[1034]), .Z(n17476) );
  XNOR U18199 ( .A(q[4]), .B(DB[1033]), .Z(n10279) );
  IV U18200 ( .A(n10293), .Z(n17474) );
  XOR U18201 ( .A(n17477), .B(n17478), .Z(n10293) );
  XNOR U18202 ( .A(n10289), .B(n10291), .Z(n17478) );
  XNOR U18203 ( .A(q[0]), .B(DB[1029]), .Z(n10291) );
  XNOR U18204 ( .A(q[3]), .B(DB[1032]), .Z(n10289) );
  IV U18205 ( .A(n10288), .Z(n17477) );
  XNOR U18206 ( .A(n10286), .B(n17479), .Z(n10288) );
  XNOR U18207 ( .A(q[2]), .B(DB[1031]), .Z(n17479) );
  XNOR U18208 ( .A(q[1]), .B(DB[1030]), .Z(n10286) );
  XOR U18209 ( .A(n17480), .B(n10251), .Z(n10214) );
  XOR U18210 ( .A(n17481), .B(n10239), .Z(n10251) );
  XNOR U18211 ( .A(q[6]), .B(DB[1042]), .Z(n10239) );
  IV U18212 ( .A(n10238), .Z(n17481) );
  XNOR U18213 ( .A(n10236), .B(n17482), .Z(n10238) );
  XNOR U18214 ( .A(q[5]), .B(DB[1041]), .Z(n17482) );
  XNOR U18215 ( .A(q[4]), .B(DB[1040]), .Z(n10236) );
  IV U18216 ( .A(n10250), .Z(n17480) );
  XOR U18217 ( .A(n17483), .B(n17484), .Z(n10250) );
  XNOR U18218 ( .A(n10246), .B(n10248), .Z(n17484) );
  XNOR U18219 ( .A(q[0]), .B(DB[1036]), .Z(n10248) );
  XNOR U18220 ( .A(q[3]), .B(DB[1039]), .Z(n10246) );
  IV U18221 ( .A(n10245), .Z(n17483) );
  XNOR U18222 ( .A(n10243), .B(n17485), .Z(n10245) );
  XNOR U18223 ( .A(q[2]), .B(DB[1038]), .Z(n17485) );
  XNOR U18224 ( .A(q[1]), .B(DB[1037]), .Z(n10243) );
  XOR U18225 ( .A(n17486), .B(n10208), .Z(n10171) );
  XOR U18226 ( .A(n17487), .B(n10196), .Z(n10208) );
  XNOR U18227 ( .A(q[6]), .B(DB[1049]), .Z(n10196) );
  IV U18228 ( .A(n10195), .Z(n17487) );
  XNOR U18229 ( .A(n10193), .B(n17488), .Z(n10195) );
  XNOR U18230 ( .A(q[5]), .B(DB[1048]), .Z(n17488) );
  XNOR U18231 ( .A(q[4]), .B(DB[1047]), .Z(n10193) );
  IV U18232 ( .A(n10207), .Z(n17486) );
  XOR U18233 ( .A(n17489), .B(n17490), .Z(n10207) );
  XNOR U18234 ( .A(n10203), .B(n10205), .Z(n17490) );
  XNOR U18235 ( .A(q[0]), .B(DB[1043]), .Z(n10205) );
  XNOR U18236 ( .A(q[3]), .B(DB[1046]), .Z(n10203) );
  IV U18237 ( .A(n10202), .Z(n17489) );
  XNOR U18238 ( .A(n10200), .B(n17491), .Z(n10202) );
  XNOR U18239 ( .A(q[2]), .B(DB[1045]), .Z(n17491) );
  XNOR U18240 ( .A(q[1]), .B(DB[1044]), .Z(n10200) );
  XOR U18241 ( .A(n17492), .B(n10165), .Z(n10128) );
  XOR U18242 ( .A(n17493), .B(n10153), .Z(n10165) );
  XNOR U18243 ( .A(q[6]), .B(DB[1056]), .Z(n10153) );
  IV U18244 ( .A(n10152), .Z(n17493) );
  XNOR U18245 ( .A(n10150), .B(n17494), .Z(n10152) );
  XNOR U18246 ( .A(q[5]), .B(DB[1055]), .Z(n17494) );
  XNOR U18247 ( .A(q[4]), .B(DB[1054]), .Z(n10150) );
  IV U18248 ( .A(n10164), .Z(n17492) );
  XOR U18249 ( .A(n17495), .B(n17496), .Z(n10164) );
  XNOR U18250 ( .A(n10160), .B(n10162), .Z(n17496) );
  XNOR U18251 ( .A(q[0]), .B(DB[1050]), .Z(n10162) );
  XNOR U18252 ( .A(q[3]), .B(DB[1053]), .Z(n10160) );
  IV U18253 ( .A(n10159), .Z(n17495) );
  XNOR U18254 ( .A(n10157), .B(n17497), .Z(n10159) );
  XNOR U18255 ( .A(q[2]), .B(DB[1052]), .Z(n17497) );
  XNOR U18256 ( .A(q[1]), .B(DB[1051]), .Z(n10157) );
  XOR U18257 ( .A(n17498), .B(n10122), .Z(n10085) );
  XOR U18258 ( .A(n17499), .B(n10110), .Z(n10122) );
  XNOR U18259 ( .A(q[6]), .B(DB[1063]), .Z(n10110) );
  IV U18260 ( .A(n10109), .Z(n17499) );
  XNOR U18261 ( .A(n10107), .B(n17500), .Z(n10109) );
  XNOR U18262 ( .A(q[5]), .B(DB[1062]), .Z(n17500) );
  XNOR U18263 ( .A(q[4]), .B(DB[1061]), .Z(n10107) );
  IV U18264 ( .A(n10121), .Z(n17498) );
  XOR U18265 ( .A(n17501), .B(n17502), .Z(n10121) );
  XNOR U18266 ( .A(n10117), .B(n10119), .Z(n17502) );
  XNOR U18267 ( .A(q[0]), .B(DB[1057]), .Z(n10119) );
  XNOR U18268 ( .A(q[3]), .B(DB[1060]), .Z(n10117) );
  IV U18269 ( .A(n10116), .Z(n17501) );
  XNOR U18270 ( .A(n10114), .B(n17503), .Z(n10116) );
  XNOR U18271 ( .A(q[2]), .B(DB[1059]), .Z(n17503) );
  XNOR U18272 ( .A(q[1]), .B(DB[1058]), .Z(n10114) );
  XOR U18273 ( .A(n17504), .B(n10079), .Z(n10042) );
  XOR U18274 ( .A(n17505), .B(n10067), .Z(n10079) );
  XNOR U18275 ( .A(q[6]), .B(DB[1070]), .Z(n10067) );
  IV U18276 ( .A(n10066), .Z(n17505) );
  XNOR U18277 ( .A(n10064), .B(n17506), .Z(n10066) );
  XNOR U18278 ( .A(q[5]), .B(DB[1069]), .Z(n17506) );
  XNOR U18279 ( .A(q[4]), .B(DB[1068]), .Z(n10064) );
  IV U18280 ( .A(n10078), .Z(n17504) );
  XOR U18281 ( .A(n17507), .B(n17508), .Z(n10078) );
  XNOR U18282 ( .A(n10074), .B(n10076), .Z(n17508) );
  XNOR U18283 ( .A(q[0]), .B(DB[1064]), .Z(n10076) );
  XNOR U18284 ( .A(q[3]), .B(DB[1067]), .Z(n10074) );
  IV U18285 ( .A(n10073), .Z(n17507) );
  XNOR U18286 ( .A(n10071), .B(n17509), .Z(n10073) );
  XNOR U18287 ( .A(q[2]), .B(DB[1066]), .Z(n17509) );
  XNOR U18288 ( .A(q[1]), .B(DB[1065]), .Z(n10071) );
  XOR U18289 ( .A(n17510), .B(n10036), .Z(n9999) );
  XOR U18290 ( .A(n17511), .B(n10024), .Z(n10036) );
  XNOR U18291 ( .A(q[6]), .B(DB[1077]), .Z(n10024) );
  IV U18292 ( .A(n10023), .Z(n17511) );
  XNOR U18293 ( .A(n10021), .B(n17512), .Z(n10023) );
  XNOR U18294 ( .A(q[5]), .B(DB[1076]), .Z(n17512) );
  XNOR U18295 ( .A(q[4]), .B(DB[1075]), .Z(n10021) );
  IV U18296 ( .A(n10035), .Z(n17510) );
  XOR U18297 ( .A(n17513), .B(n17514), .Z(n10035) );
  XNOR U18298 ( .A(n10031), .B(n10033), .Z(n17514) );
  XNOR U18299 ( .A(q[0]), .B(DB[1071]), .Z(n10033) );
  XNOR U18300 ( .A(q[3]), .B(DB[1074]), .Z(n10031) );
  IV U18301 ( .A(n10030), .Z(n17513) );
  XNOR U18302 ( .A(n10028), .B(n17515), .Z(n10030) );
  XNOR U18303 ( .A(q[2]), .B(DB[1073]), .Z(n17515) );
  XNOR U18304 ( .A(q[1]), .B(DB[1072]), .Z(n10028) );
  XOR U18305 ( .A(n17516), .B(n9993), .Z(n9956) );
  XOR U18306 ( .A(n17517), .B(n9981), .Z(n9993) );
  XNOR U18307 ( .A(q[6]), .B(DB[1084]), .Z(n9981) );
  IV U18308 ( .A(n9980), .Z(n17517) );
  XNOR U18309 ( .A(n9978), .B(n17518), .Z(n9980) );
  XNOR U18310 ( .A(q[5]), .B(DB[1083]), .Z(n17518) );
  XNOR U18311 ( .A(q[4]), .B(DB[1082]), .Z(n9978) );
  IV U18312 ( .A(n9992), .Z(n17516) );
  XOR U18313 ( .A(n17519), .B(n17520), .Z(n9992) );
  XNOR U18314 ( .A(n9988), .B(n9990), .Z(n17520) );
  XNOR U18315 ( .A(q[0]), .B(DB[1078]), .Z(n9990) );
  XNOR U18316 ( .A(q[3]), .B(DB[1081]), .Z(n9988) );
  IV U18317 ( .A(n9987), .Z(n17519) );
  XNOR U18318 ( .A(n9985), .B(n17521), .Z(n9987) );
  XNOR U18319 ( .A(q[2]), .B(DB[1080]), .Z(n17521) );
  XNOR U18320 ( .A(q[1]), .B(DB[1079]), .Z(n9985) );
  XOR U18321 ( .A(n17522), .B(n9950), .Z(n9913) );
  XOR U18322 ( .A(n17523), .B(n9938), .Z(n9950) );
  XNOR U18323 ( .A(q[6]), .B(DB[1091]), .Z(n9938) );
  IV U18324 ( .A(n9937), .Z(n17523) );
  XNOR U18325 ( .A(n9935), .B(n17524), .Z(n9937) );
  XNOR U18326 ( .A(q[5]), .B(DB[1090]), .Z(n17524) );
  XNOR U18327 ( .A(q[4]), .B(DB[1089]), .Z(n9935) );
  IV U18328 ( .A(n9949), .Z(n17522) );
  XOR U18329 ( .A(n17525), .B(n17526), .Z(n9949) );
  XNOR U18330 ( .A(n9945), .B(n9947), .Z(n17526) );
  XNOR U18331 ( .A(q[0]), .B(DB[1085]), .Z(n9947) );
  XNOR U18332 ( .A(q[3]), .B(DB[1088]), .Z(n9945) );
  IV U18333 ( .A(n9944), .Z(n17525) );
  XNOR U18334 ( .A(n9942), .B(n17527), .Z(n9944) );
  XNOR U18335 ( .A(q[2]), .B(DB[1087]), .Z(n17527) );
  XNOR U18336 ( .A(q[1]), .B(DB[1086]), .Z(n9942) );
  XOR U18337 ( .A(n17528), .B(n9907), .Z(n9870) );
  XOR U18338 ( .A(n17529), .B(n9895), .Z(n9907) );
  XNOR U18339 ( .A(q[6]), .B(DB[1098]), .Z(n9895) );
  IV U18340 ( .A(n9894), .Z(n17529) );
  XNOR U18341 ( .A(n9892), .B(n17530), .Z(n9894) );
  XNOR U18342 ( .A(q[5]), .B(DB[1097]), .Z(n17530) );
  XNOR U18343 ( .A(q[4]), .B(DB[1096]), .Z(n9892) );
  IV U18344 ( .A(n9906), .Z(n17528) );
  XOR U18345 ( .A(n17531), .B(n17532), .Z(n9906) );
  XNOR U18346 ( .A(n9902), .B(n9904), .Z(n17532) );
  XNOR U18347 ( .A(q[0]), .B(DB[1092]), .Z(n9904) );
  XNOR U18348 ( .A(q[3]), .B(DB[1095]), .Z(n9902) );
  IV U18349 ( .A(n9901), .Z(n17531) );
  XNOR U18350 ( .A(n9899), .B(n17533), .Z(n9901) );
  XNOR U18351 ( .A(q[2]), .B(DB[1094]), .Z(n17533) );
  XNOR U18352 ( .A(q[1]), .B(DB[1093]), .Z(n9899) );
  XOR U18353 ( .A(n17534), .B(n9864), .Z(n9827) );
  XOR U18354 ( .A(n17535), .B(n9852), .Z(n9864) );
  XNOR U18355 ( .A(q[6]), .B(DB[1105]), .Z(n9852) );
  IV U18356 ( .A(n9851), .Z(n17535) );
  XNOR U18357 ( .A(n9849), .B(n17536), .Z(n9851) );
  XNOR U18358 ( .A(q[5]), .B(DB[1104]), .Z(n17536) );
  XNOR U18359 ( .A(q[4]), .B(DB[1103]), .Z(n9849) );
  IV U18360 ( .A(n9863), .Z(n17534) );
  XOR U18361 ( .A(n17537), .B(n17538), .Z(n9863) );
  XNOR U18362 ( .A(n9859), .B(n9861), .Z(n17538) );
  XNOR U18363 ( .A(q[0]), .B(DB[1099]), .Z(n9861) );
  XNOR U18364 ( .A(q[3]), .B(DB[1102]), .Z(n9859) );
  IV U18365 ( .A(n9858), .Z(n17537) );
  XNOR U18366 ( .A(n9856), .B(n17539), .Z(n9858) );
  XNOR U18367 ( .A(q[2]), .B(DB[1101]), .Z(n17539) );
  XNOR U18368 ( .A(q[1]), .B(DB[1100]), .Z(n9856) );
  XOR U18369 ( .A(n17540), .B(n9821), .Z(n9784) );
  XOR U18370 ( .A(n17541), .B(n9809), .Z(n9821) );
  XNOR U18371 ( .A(q[6]), .B(DB[1112]), .Z(n9809) );
  IV U18372 ( .A(n9808), .Z(n17541) );
  XNOR U18373 ( .A(n9806), .B(n17542), .Z(n9808) );
  XNOR U18374 ( .A(q[5]), .B(DB[1111]), .Z(n17542) );
  XNOR U18375 ( .A(q[4]), .B(DB[1110]), .Z(n9806) );
  IV U18376 ( .A(n9820), .Z(n17540) );
  XOR U18377 ( .A(n17543), .B(n17544), .Z(n9820) );
  XNOR U18378 ( .A(n9816), .B(n9818), .Z(n17544) );
  XNOR U18379 ( .A(q[0]), .B(DB[1106]), .Z(n9818) );
  XNOR U18380 ( .A(q[3]), .B(DB[1109]), .Z(n9816) );
  IV U18381 ( .A(n9815), .Z(n17543) );
  XNOR U18382 ( .A(n9813), .B(n17545), .Z(n9815) );
  XNOR U18383 ( .A(q[2]), .B(DB[1108]), .Z(n17545) );
  XNOR U18384 ( .A(q[1]), .B(DB[1107]), .Z(n9813) );
  XOR U18385 ( .A(n17546), .B(n9778), .Z(n9741) );
  XOR U18386 ( .A(n17547), .B(n9766), .Z(n9778) );
  XNOR U18387 ( .A(q[6]), .B(DB[1119]), .Z(n9766) );
  IV U18388 ( .A(n9765), .Z(n17547) );
  XNOR U18389 ( .A(n9763), .B(n17548), .Z(n9765) );
  XNOR U18390 ( .A(q[5]), .B(DB[1118]), .Z(n17548) );
  XNOR U18391 ( .A(q[4]), .B(DB[1117]), .Z(n9763) );
  IV U18392 ( .A(n9777), .Z(n17546) );
  XOR U18393 ( .A(n17549), .B(n17550), .Z(n9777) );
  XNOR U18394 ( .A(n9773), .B(n9775), .Z(n17550) );
  XNOR U18395 ( .A(q[0]), .B(DB[1113]), .Z(n9775) );
  XNOR U18396 ( .A(q[3]), .B(DB[1116]), .Z(n9773) );
  IV U18397 ( .A(n9772), .Z(n17549) );
  XNOR U18398 ( .A(n9770), .B(n17551), .Z(n9772) );
  XNOR U18399 ( .A(q[2]), .B(DB[1115]), .Z(n17551) );
  XNOR U18400 ( .A(q[1]), .B(DB[1114]), .Z(n9770) );
  XOR U18401 ( .A(n17552), .B(n9735), .Z(n9698) );
  XOR U18402 ( .A(n17553), .B(n9723), .Z(n9735) );
  XNOR U18403 ( .A(q[6]), .B(DB[1126]), .Z(n9723) );
  IV U18404 ( .A(n9722), .Z(n17553) );
  XNOR U18405 ( .A(n9720), .B(n17554), .Z(n9722) );
  XNOR U18406 ( .A(q[5]), .B(DB[1125]), .Z(n17554) );
  XNOR U18407 ( .A(q[4]), .B(DB[1124]), .Z(n9720) );
  IV U18408 ( .A(n9734), .Z(n17552) );
  XOR U18409 ( .A(n17555), .B(n17556), .Z(n9734) );
  XNOR U18410 ( .A(n9730), .B(n9732), .Z(n17556) );
  XNOR U18411 ( .A(q[0]), .B(DB[1120]), .Z(n9732) );
  XNOR U18412 ( .A(q[3]), .B(DB[1123]), .Z(n9730) );
  IV U18413 ( .A(n9729), .Z(n17555) );
  XNOR U18414 ( .A(n9727), .B(n17557), .Z(n9729) );
  XNOR U18415 ( .A(q[2]), .B(DB[1122]), .Z(n17557) );
  XNOR U18416 ( .A(q[1]), .B(DB[1121]), .Z(n9727) );
  XOR U18417 ( .A(n17558), .B(n9692), .Z(n9655) );
  XOR U18418 ( .A(n17559), .B(n9680), .Z(n9692) );
  XNOR U18419 ( .A(q[6]), .B(DB[1133]), .Z(n9680) );
  IV U18420 ( .A(n9679), .Z(n17559) );
  XNOR U18421 ( .A(n9677), .B(n17560), .Z(n9679) );
  XNOR U18422 ( .A(q[5]), .B(DB[1132]), .Z(n17560) );
  XNOR U18423 ( .A(q[4]), .B(DB[1131]), .Z(n9677) );
  IV U18424 ( .A(n9691), .Z(n17558) );
  XOR U18425 ( .A(n17561), .B(n17562), .Z(n9691) );
  XNOR U18426 ( .A(n9687), .B(n9689), .Z(n17562) );
  XNOR U18427 ( .A(q[0]), .B(DB[1127]), .Z(n9689) );
  XNOR U18428 ( .A(q[3]), .B(DB[1130]), .Z(n9687) );
  IV U18429 ( .A(n9686), .Z(n17561) );
  XNOR U18430 ( .A(n9684), .B(n17563), .Z(n9686) );
  XNOR U18431 ( .A(q[2]), .B(DB[1129]), .Z(n17563) );
  XNOR U18432 ( .A(q[1]), .B(DB[1128]), .Z(n9684) );
  XOR U18433 ( .A(n17564), .B(n9649), .Z(n9612) );
  XOR U18434 ( .A(n17565), .B(n9637), .Z(n9649) );
  XNOR U18435 ( .A(q[6]), .B(DB[1140]), .Z(n9637) );
  IV U18436 ( .A(n9636), .Z(n17565) );
  XNOR U18437 ( .A(n9634), .B(n17566), .Z(n9636) );
  XNOR U18438 ( .A(q[5]), .B(DB[1139]), .Z(n17566) );
  XNOR U18439 ( .A(q[4]), .B(DB[1138]), .Z(n9634) );
  IV U18440 ( .A(n9648), .Z(n17564) );
  XOR U18441 ( .A(n17567), .B(n17568), .Z(n9648) );
  XNOR U18442 ( .A(n9644), .B(n9646), .Z(n17568) );
  XNOR U18443 ( .A(q[0]), .B(DB[1134]), .Z(n9646) );
  XNOR U18444 ( .A(q[3]), .B(DB[1137]), .Z(n9644) );
  IV U18445 ( .A(n9643), .Z(n17567) );
  XNOR U18446 ( .A(n9641), .B(n17569), .Z(n9643) );
  XNOR U18447 ( .A(q[2]), .B(DB[1136]), .Z(n17569) );
  XNOR U18448 ( .A(q[1]), .B(DB[1135]), .Z(n9641) );
  XOR U18449 ( .A(n17570), .B(n9606), .Z(n9569) );
  XOR U18450 ( .A(n17571), .B(n9594), .Z(n9606) );
  XNOR U18451 ( .A(q[6]), .B(DB[1147]), .Z(n9594) );
  IV U18452 ( .A(n9593), .Z(n17571) );
  XNOR U18453 ( .A(n9591), .B(n17572), .Z(n9593) );
  XNOR U18454 ( .A(q[5]), .B(DB[1146]), .Z(n17572) );
  XNOR U18455 ( .A(q[4]), .B(DB[1145]), .Z(n9591) );
  IV U18456 ( .A(n9605), .Z(n17570) );
  XOR U18457 ( .A(n17573), .B(n17574), .Z(n9605) );
  XNOR U18458 ( .A(n9601), .B(n9603), .Z(n17574) );
  XNOR U18459 ( .A(q[0]), .B(DB[1141]), .Z(n9603) );
  XNOR U18460 ( .A(q[3]), .B(DB[1144]), .Z(n9601) );
  IV U18461 ( .A(n9600), .Z(n17573) );
  XNOR U18462 ( .A(n9598), .B(n17575), .Z(n9600) );
  XNOR U18463 ( .A(q[2]), .B(DB[1143]), .Z(n17575) );
  XNOR U18464 ( .A(q[1]), .B(DB[1142]), .Z(n9598) );
  XOR U18465 ( .A(n17576), .B(n9563), .Z(n9526) );
  XOR U18466 ( .A(n17577), .B(n9551), .Z(n9563) );
  XNOR U18467 ( .A(q[6]), .B(DB[1154]), .Z(n9551) );
  IV U18468 ( .A(n9550), .Z(n17577) );
  XNOR U18469 ( .A(n9548), .B(n17578), .Z(n9550) );
  XNOR U18470 ( .A(q[5]), .B(DB[1153]), .Z(n17578) );
  XNOR U18471 ( .A(q[4]), .B(DB[1152]), .Z(n9548) );
  IV U18472 ( .A(n9562), .Z(n17576) );
  XOR U18473 ( .A(n17579), .B(n17580), .Z(n9562) );
  XNOR U18474 ( .A(n9558), .B(n9560), .Z(n17580) );
  XNOR U18475 ( .A(q[0]), .B(DB[1148]), .Z(n9560) );
  XNOR U18476 ( .A(q[3]), .B(DB[1151]), .Z(n9558) );
  IV U18477 ( .A(n9557), .Z(n17579) );
  XNOR U18478 ( .A(n9555), .B(n17581), .Z(n9557) );
  XNOR U18479 ( .A(q[2]), .B(DB[1150]), .Z(n17581) );
  XNOR U18480 ( .A(q[1]), .B(DB[1149]), .Z(n9555) );
  XOR U18481 ( .A(n17582), .B(n9520), .Z(n9483) );
  XOR U18482 ( .A(n17583), .B(n9508), .Z(n9520) );
  XNOR U18483 ( .A(q[6]), .B(DB[1161]), .Z(n9508) );
  IV U18484 ( .A(n9507), .Z(n17583) );
  XNOR U18485 ( .A(n9505), .B(n17584), .Z(n9507) );
  XNOR U18486 ( .A(q[5]), .B(DB[1160]), .Z(n17584) );
  XNOR U18487 ( .A(q[4]), .B(DB[1159]), .Z(n9505) );
  IV U18488 ( .A(n9519), .Z(n17582) );
  XOR U18489 ( .A(n17585), .B(n17586), .Z(n9519) );
  XNOR U18490 ( .A(n9515), .B(n9517), .Z(n17586) );
  XNOR U18491 ( .A(q[0]), .B(DB[1155]), .Z(n9517) );
  XNOR U18492 ( .A(q[3]), .B(DB[1158]), .Z(n9515) );
  IV U18493 ( .A(n9514), .Z(n17585) );
  XNOR U18494 ( .A(n9512), .B(n17587), .Z(n9514) );
  XNOR U18495 ( .A(q[2]), .B(DB[1157]), .Z(n17587) );
  XNOR U18496 ( .A(q[1]), .B(DB[1156]), .Z(n9512) );
  XOR U18497 ( .A(n17588), .B(n9477), .Z(n9440) );
  XOR U18498 ( .A(n17589), .B(n9465), .Z(n9477) );
  XNOR U18499 ( .A(q[6]), .B(DB[1168]), .Z(n9465) );
  IV U18500 ( .A(n9464), .Z(n17589) );
  XNOR U18501 ( .A(n9462), .B(n17590), .Z(n9464) );
  XNOR U18502 ( .A(q[5]), .B(DB[1167]), .Z(n17590) );
  XNOR U18503 ( .A(q[4]), .B(DB[1166]), .Z(n9462) );
  IV U18504 ( .A(n9476), .Z(n17588) );
  XOR U18505 ( .A(n17591), .B(n17592), .Z(n9476) );
  XNOR U18506 ( .A(n9472), .B(n9474), .Z(n17592) );
  XNOR U18507 ( .A(q[0]), .B(DB[1162]), .Z(n9474) );
  XNOR U18508 ( .A(q[3]), .B(DB[1165]), .Z(n9472) );
  IV U18509 ( .A(n9471), .Z(n17591) );
  XNOR U18510 ( .A(n9469), .B(n17593), .Z(n9471) );
  XNOR U18511 ( .A(q[2]), .B(DB[1164]), .Z(n17593) );
  XNOR U18512 ( .A(q[1]), .B(DB[1163]), .Z(n9469) );
  XOR U18513 ( .A(n17594), .B(n9434), .Z(n9397) );
  XOR U18514 ( .A(n17595), .B(n9422), .Z(n9434) );
  XNOR U18515 ( .A(q[6]), .B(DB[1175]), .Z(n9422) );
  IV U18516 ( .A(n9421), .Z(n17595) );
  XNOR U18517 ( .A(n9419), .B(n17596), .Z(n9421) );
  XNOR U18518 ( .A(q[5]), .B(DB[1174]), .Z(n17596) );
  XNOR U18519 ( .A(q[4]), .B(DB[1173]), .Z(n9419) );
  IV U18520 ( .A(n9433), .Z(n17594) );
  XOR U18521 ( .A(n17597), .B(n17598), .Z(n9433) );
  XNOR U18522 ( .A(n9429), .B(n9431), .Z(n17598) );
  XNOR U18523 ( .A(q[0]), .B(DB[1169]), .Z(n9431) );
  XNOR U18524 ( .A(q[3]), .B(DB[1172]), .Z(n9429) );
  IV U18525 ( .A(n9428), .Z(n17597) );
  XNOR U18526 ( .A(n9426), .B(n17599), .Z(n9428) );
  XNOR U18527 ( .A(q[2]), .B(DB[1171]), .Z(n17599) );
  XNOR U18528 ( .A(q[1]), .B(DB[1170]), .Z(n9426) );
  XOR U18529 ( .A(n17600), .B(n9391), .Z(n9354) );
  XOR U18530 ( .A(n17601), .B(n9379), .Z(n9391) );
  XNOR U18531 ( .A(q[6]), .B(DB[1182]), .Z(n9379) );
  IV U18532 ( .A(n9378), .Z(n17601) );
  XNOR U18533 ( .A(n9376), .B(n17602), .Z(n9378) );
  XNOR U18534 ( .A(q[5]), .B(DB[1181]), .Z(n17602) );
  XNOR U18535 ( .A(q[4]), .B(DB[1180]), .Z(n9376) );
  IV U18536 ( .A(n9390), .Z(n17600) );
  XOR U18537 ( .A(n17603), .B(n17604), .Z(n9390) );
  XNOR U18538 ( .A(n9386), .B(n9388), .Z(n17604) );
  XNOR U18539 ( .A(q[0]), .B(DB[1176]), .Z(n9388) );
  XNOR U18540 ( .A(q[3]), .B(DB[1179]), .Z(n9386) );
  IV U18541 ( .A(n9385), .Z(n17603) );
  XNOR U18542 ( .A(n9383), .B(n17605), .Z(n9385) );
  XNOR U18543 ( .A(q[2]), .B(DB[1178]), .Z(n17605) );
  XNOR U18544 ( .A(q[1]), .B(DB[1177]), .Z(n9383) );
  XOR U18545 ( .A(n17606), .B(n9348), .Z(n9311) );
  XOR U18546 ( .A(n17607), .B(n9336), .Z(n9348) );
  XNOR U18547 ( .A(q[6]), .B(DB[1189]), .Z(n9336) );
  IV U18548 ( .A(n9335), .Z(n17607) );
  XNOR U18549 ( .A(n9333), .B(n17608), .Z(n9335) );
  XNOR U18550 ( .A(q[5]), .B(DB[1188]), .Z(n17608) );
  XNOR U18551 ( .A(q[4]), .B(DB[1187]), .Z(n9333) );
  IV U18552 ( .A(n9347), .Z(n17606) );
  XOR U18553 ( .A(n17609), .B(n17610), .Z(n9347) );
  XNOR U18554 ( .A(n9343), .B(n9345), .Z(n17610) );
  XNOR U18555 ( .A(q[0]), .B(DB[1183]), .Z(n9345) );
  XNOR U18556 ( .A(q[3]), .B(DB[1186]), .Z(n9343) );
  IV U18557 ( .A(n9342), .Z(n17609) );
  XNOR U18558 ( .A(n9340), .B(n17611), .Z(n9342) );
  XNOR U18559 ( .A(q[2]), .B(DB[1185]), .Z(n17611) );
  XNOR U18560 ( .A(q[1]), .B(DB[1184]), .Z(n9340) );
  XOR U18561 ( .A(n17612), .B(n9305), .Z(n9268) );
  XOR U18562 ( .A(n17613), .B(n9293), .Z(n9305) );
  XNOR U18563 ( .A(q[6]), .B(DB[1196]), .Z(n9293) );
  IV U18564 ( .A(n9292), .Z(n17613) );
  XNOR U18565 ( .A(n9290), .B(n17614), .Z(n9292) );
  XNOR U18566 ( .A(q[5]), .B(DB[1195]), .Z(n17614) );
  XNOR U18567 ( .A(q[4]), .B(DB[1194]), .Z(n9290) );
  IV U18568 ( .A(n9304), .Z(n17612) );
  XOR U18569 ( .A(n17615), .B(n17616), .Z(n9304) );
  XNOR U18570 ( .A(n9300), .B(n9302), .Z(n17616) );
  XNOR U18571 ( .A(q[0]), .B(DB[1190]), .Z(n9302) );
  XNOR U18572 ( .A(q[3]), .B(DB[1193]), .Z(n9300) );
  IV U18573 ( .A(n9299), .Z(n17615) );
  XNOR U18574 ( .A(n9297), .B(n17617), .Z(n9299) );
  XNOR U18575 ( .A(q[2]), .B(DB[1192]), .Z(n17617) );
  XNOR U18576 ( .A(q[1]), .B(DB[1191]), .Z(n9297) );
  XOR U18577 ( .A(n17618), .B(n9262), .Z(n9225) );
  XOR U18578 ( .A(n17619), .B(n9250), .Z(n9262) );
  XNOR U18579 ( .A(q[6]), .B(DB[1203]), .Z(n9250) );
  IV U18580 ( .A(n9249), .Z(n17619) );
  XNOR U18581 ( .A(n9247), .B(n17620), .Z(n9249) );
  XNOR U18582 ( .A(q[5]), .B(DB[1202]), .Z(n17620) );
  XNOR U18583 ( .A(q[4]), .B(DB[1201]), .Z(n9247) );
  IV U18584 ( .A(n9261), .Z(n17618) );
  XOR U18585 ( .A(n17621), .B(n17622), .Z(n9261) );
  XNOR U18586 ( .A(n9257), .B(n9259), .Z(n17622) );
  XNOR U18587 ( .A(q[0]), .B(DB[1197]), .Z(n9259) );
  XNOR U18588 ( .A(q[3]), .B(DB[1200]), .Z(n9257) );
  IV U18589 ( .A(n9256), .Z(n17621) );
  XNOR U18590 ( .A(n9254), .B(n17623), .Z(n9256) );
  XNOR U18591 ( .A(q[2]), .B(DB[1199]), .Z(n17623) );
  XNOR U18592 ( .A(q[1]), .B(DB[1198]), .Z(n9254) );
  XOR U18593 ( .A(n17624), .B(n9219), .Z(n9182) );
  XOR U18594 ( .A(n17625), .B(n9207), .Z(n9219) );
  XNOR U18595 ( .A(q[6]), .B(DB[1210]), .Z(n9207) );
  IV U18596 ( .A(n9206), .Z(n17625) );
  XNOR U18597 ( .A(n9204), .B(n17626), .Z(n9206) );
  XNOR U18598 ( .A(q[5]), .B(DB[1209]), .Z(n17626) );
  XNOR U18599 ( .A(q[4]), .B(DB[1208]), .Z(n9204) );
  IV U18600 ( .A(n9218), .Z(n17624) );
  XOR U18601 ( .A(n17627), .B(n17628), .Z(n9218) );
  XNOR U18602 ( .A(n9214), .B(n9216), .Z(n17628) );
  XNOR U18603 ( .A(q[0]), .B(DB[1204]), .Z(n9216) );
  XNOR U18604 ( .A(q[3]), .B(DB[1207]), .Z(n9214) );
  IV U18605 ( .A(n9213), .Z(n17627) );
  XNOR U18606 ( .A(n9211), .B(n17629), .Z(n9213) );
  XNOR U18607 ( .A(q[2]), .B(DB[1206]), .Z(n17629) );
  XNOR U18608 ( .A(q[1]), .B(DB[1205]), .Z(n9211) );
  XOR U18609 ( .A(n17630), .B(n9176), .Z(n9139) );
  XOR U18610 ( .A(n17631), .B(n9164), .Z(n9176) );
  XNOR U18611 ( .A(q[6]), .B(DB[1217]), .Z(n9164) );
  IV U18612 ( .A(n9163), .Z(n17631) );
  XNOR U18613 ( .A(n9161), .B(n17632), .Z(n9163) );
  XNOR U18614 ( .A(q[5]), .B(DB[1216]), .Z(n17632) );
  XNOR U18615 ( .A(q[4]), .B(DB[1215]), .Z(n9161) );
  IV U18616 ( .A(n9175), .Z(n17630) );
  XOR U18617 ( .A(n17633), .B(n17634), .Z(n9175) );
  XNOR U18618 ( .A(n9171), .B(n9173), .Z(n17634) );
  XNOR U18619 ( .A(q[0]), .B(DB[1211]), .Z(n9173) );
  XNOR U18620 ( .A(q[3]), .B(DB[1214]), .Z(n9171) );
  IV U18621 ( .A(n9170), .Z(n17633) );
  XNOR U18622 ( .A(n9168), .B(n17635), .Z(n9170) );
  XNOR U18623 ( .A(q[2]), .B(DB[1213]), .Z(n17635) );
  XNOR U18624 ( .A(q[1]), .B(DB[1212]), .Z(n9168) );
  XOR U18625 ( .A(n17636), .B(n9133), .Z(n9096) );
  XOR U18626 ( .A(n17637), .B(n9121), .Z(n9133) );
  XNOR U18627 ( .A(q[6]), .B(DB[1224]), .Z(n9121) );
  IV U18628 ( .A(n9120), .Z(n17637) );
  XNOR U18629 ( .A(n9118), .B(n17638), .Z(n9120) );
  XNOR U18630 ( .A(q[5]), .B(DB[1223]), .Z(n17638) );
  XNOR U18631 ( .A(q[4]), .B(DB[1222]), .Z(n9118) );
  IV U18632 ( .A(n9132), .Z(n17636) );
  XOR U18633 ( .A(n17639), .B(n17640), .Z(n9132) );
  XNOR U18634 ( .A(n9128), .B(n9130), .Z(n17640) );
  XNOR U18635 ( .A(q[0]), .B(DB[1218]), .Z(n9130) );
  XNOR U18636 ( .A(q[3]), .B(DB[1221]), .Z(n9128) );
  IV U18637 ( .A(n9127), .Z(n17639) );
  XNOR U18638 ( .A(n9125), .B(n17641), .Z(n9127) );
  XNOR U18639 ( .A(q[2]), .B(DB[1220]), .Z(n17641) );
  XNOR U18640 ( .A(q[1]), .B(DB[1219]), .Z(n9125) );
  XOR U18641 ( .A(n17642), .B(n9090), .Z(n9053) );
  XOR U18642 ( .A(n17643), .B(n9078), .Z(n9090) );
  XNOR U18643 ( .A(q[6]), .B(DB[1231]), .Z(n9078) );
  IV U18644 ( .A(n9077), .Z(n17643) );
  XNOR U18645 ( .A(n9075), .B(n17644), .Z(n9077) );
  XNOR U18646 ( .A(q[5]), .B(DB[1230]), .Z(n17644) );
  XNOR U18647 ( .A(q[4]), .B(DB[1229]), .Z(n9075) );
  IV U18648 ( .A(n9089), .Z(n17642) );
  XOR U18649 ( .A(n17645), .B(n17646), .Z(n9089) );
  XNOR U18650 ( .A(n9085), .B(n9087), .Z(n17646) );
  XNOR U18651 ( .A(q[0]), .B(DB[1225]), .Z(n9087) );
  XNOR U18652 ( .A(q[3]), .B(DB[1228]), .Z(n9085) );
  IV U18653 ( .A(n9084), .Z(n17645) );
  XNOR U18654 ( .A(n9082), .B(n17647), .Z(n9084) );
  XNOR U18655 ( .A(q[2]), .B(DB[1227]), .Z(n17647) );
  XNOR U18656 ( .A(q[1]), .B(DB[1226]), .Z(n9082) );
  XOR U18657 ( .A(n17648), .B(n9047), .Z(n9010) );
  XOR U18658 ( .A(n17649), .B(n9035), .Z(n9047) );
  XNOR U18659 ( .A(q[6]), .B(DB[1238]), .Z(n9035) );
  IV U18660 ( .A(n9034), .Z(n17649) );
  XNOR U18661 ( .A(n9032), .B(n17650), .Z(n9034) );
  XNOR U18662 ( .A(q[5]), .B(DB[1237]), .Z(n17650) );
  XNOR U18663 ( .A(q[4]), .B(DB[1236]), .Z(n9032) );
  IV U18664 ( .A(n9046), .Z(n17648) );
  XOR U18665 ( .A(n17651), .B(n17652), .Z(n9046) );
  XNOR U18666 ( .A(n9042), .B(n9044), .Z(n17652) );
  XNOR U18667 ( .A(q[0]), .B(DB[1232]), .Z(n9044) );
  XNOR U18668 ( .A(q[3]), .B(DB[1235]), .Z(n9042) );
  IV U18669 ( .A(n9041), .Z(n17651) );
  XNOR U18670 ( .A(n9039), .B(n17653), .Z(n9041) );
  XNOR U18671 ( .A(q[2]), .B(DB[1234]), .Z(n17653) );
  XNOR U18672 ( .A(q[1]), .B(DB[1233]), .Z(n9039) );
  XOR U18673 ( .A(n17654), .B(n9004), .Z(n8967) );
  XOR U18674 ( .A(n17655), .B(n8992), .Z(n9004) );
  XNOR U18675 ( .A(q[6]), .B(DB[1245]), .Z(n8992) );
  IV U18676 ( .A(n8991), .Z(n17655) );
  XNOR U18677 ( .A(n8989), .B(n17656), .Z(n8991) );
  XNOR U18678 ( .A(q[5]), .B(DB[1244]), .Z(n17656) );
  XNOR U18679 ( .A(q[4]), .B(DB[1243]), .Z(n8989) );
  IV U18680 ( .A(n9003), .Z(n17654) );
  XOR U18681 ( .A(n17657), .B(n17658), .Z(n9003) );
  XNOR U18682 ( .A(n8999), .B(n9001), .Z(n17658) );
  XNOR U18683 ( .A(q[0]), .B(DB[1239]), .Z(n9001) );
  XNOR U18684 ( .A(q[3]), .B(DB[1242]), .Z(n8999) );
  IV U18685 ( .A(n8998), .Z(n17657) );
  XNOR U18686 ( .A(n8996), .B(n17659), .Z(n8998) );
  XNOR U18687 ( .A(q[2]), .B(DB[1241]), .Z(n17659) );
  XNOR U18688 ( .A(q[1]), .B(DB[1240]), .Z(n8996) );
  XOR U18689 ( .A(n17660), .B(n8961), .Z(n8924) );
  XOR U18690 ( .A(n17661), .B(n8949), .Z(n8961) );
  XNOR U18691 ( .A(q[6]), .B(DB[1252]), .Z(n8949) );
  IV U18692 ( .A(n8948), .Z(n17661) );
  XNOR U18693 ( .A(n8946), .B(n17662), .Z(n8948) );
  XNOR U18694 ( .A(q[5]), .B(DB[1251]), .Z(n17662) );
  XNOR U18695 ( .A(q[4]), .B(DB[1250]), .Z(n8946) );
  IV U18696 ( .A(n8960), .Z(n17660) );
  XOR U18697 ( .A(n17663), .B(n17664), .Z(n8960) );
  XNOR U18698 ( .A(n8956), .B(n8958), .Z(n17664) );
  XNOR U18699 ( .A(q[0]), .B(DB[1246]), .Z(n8958) );
  XNOR U18700 ( .A(q[3]), .B(DB[1249]), .Z(n8956) );
  IV U18701 ( .A(n8955), .Z(n17663) );
  XNOR U18702 ( .A(n8953), .B(n17665), .Z(n8955) );
  XNOR U18703 ( .A(q[2]), .B(DB[1248]), .Z(n17665) );
  XNOR U18704 ( .A(q[1]), .B(DB[1247]), .Z(n8953) );
  XOR U18705 ( .A(n17666), .B(n8918), .Z(n8881) );
  XOR U18706 ( .A(n17667), .B(n8906), .Z(n8918) );
  XNOR U18707 ( .A(q[6]), .B(DB[1259]), .Z(n8906) );
  IV U18708 ( .A(n8905), .Z(n17667) );
  XNOR U18709 ( .A(n8903), .B(n17668), .Z(n8905) );
  XNOR U18710 ( .A(q[5]), .B(DB[1258]), .Z(n17668) );
  XNOR U18711 ( .A(q[4]), .B(DB[1257]), .Z(n8903) );
  IV U18712 ( .A(n8917), .Z(n17666) );
  XOR U18713 ( .A(n17669), .B(n17670), .Z(n8917) );
  XNOR U18714 ( .A(n8913), .B(n8915), .Z(n17670) );
  XNOR U18715 ( .A(q[0]), .B(DB[1253]), .Z(n8915) );
  XNOR U18716 ( .A(q[3]), .B(DB[1256]), .Z(n8913) );
  IV U18717 ( .A(n8912), .Z(n17669) );
  XNOR U18718 ( .A(n8910), .B(n17671), .Z(n8912) );
  XNOR U18719 ( .A(q[2]), .B(DB[1255]), .Z(n17671) );
  XNOR U18720 ( .A(q[1]), .B(DB[1254]), .Z(n8910) );
  XOR U18721 ( .A(n17672), .B(n8875), .Z(n8838) );
  XOR U18722 ( .A(n17673), .B(n8863), .Z(n8875) );
  XNOR U18723 ( .A(q[6]), .B(DB[1266]), .Z(n8863) );
  IV U18724 ( .A(n8862), .Z(n17673) );
  XNOR U18725 ( .A(n8860), .B(n17674), .Z(n8862) );
  XNOR U18726 ( .A(q[5]), .B(DB[1265]), .Z(n17674) );
  XNOR U18727 ( .A(q[4]), .B(DB[1264]), .Z(n8860) );
  IV U18728 ( .A(n8874), .Z(n17672) );
  XOR U18729 ( .A(n17675), .B(n17676), .Z(n8874) );
  XNOR U18730 ( .A(n8870), .B(n8872), .Z(n17676) );
  XNOR U18731 ( .A(q[0]), .B(DB[1260]), .Z(n8872) );
  XNOR U18732 ( .A(q[3]), .B(DB[1263]), .Z(n8870) );
  IV U18733 ( .A(n8869), .Z(n17675) );
  XNOR U18734 ( .A(n8867), .B(n17677), .Z(n8869) );
  XNOR U18735 ( .A(q[2]), .B(DB[1262]), .Z(n17677) );
  XNOR U18736 ( .A(q[1]), .B(DB[1261]), .Z(n8867) );
  XOR U18737 ( .A(n17678), .B(n8832), .Z(n8795) );
  XOR U18738 ( .A(n17679), .B(n8820), .Z(n8832) );
  XNOR U18739 ( .A(q[6]), .B(DB[1273]), .Z(n8820) );
  IV U18740 ( .A(n8819), .Z(n17679) );
  XNOR U18741 ( .A(n8817), .B(n17680), .Z(n8819) );
  XNOR U18742 ( .A(q[5]), .B(DB[1272]), .Z(n17680) );
  XNOR U18743 ( .A(q[4]), .B(DB[1271]), .Z(n8817) );
  IV U18744 ( .A(n8831), .Z(n17678) );
  XOR U18745 ( .A(n17681), .B(n17682), .Z(n8831) );
  XNOR U18746 ( .A(n8827), .B(n8829), .Z(n17682) );
  XNOR U18747 ( .A(q[0]), .B(DB[1267]), .Z(n8829) );
  XNOR U18748 ( .A(q[3]), .B(DB[1270]), .Z(n8827) );
  IV U18749 ( .A(n8826), .Z(n17681) );
  XNOR U18750 ( .A(n8824), .B(n17683), .Z(n8826) );
  XNOR U18751 ( .A(q[2]), .B(DB[1269]), .Z(n17683) );
  XNOR U18752 ( .A(q[1]), .B(DB[1268]), .Z(n8824) );
  XOR U18753 ( .A(n17684), .B(n8789), .Z(n8752) );
  XOR U18754 ( .A(n17685), .B(n8777), .Z(n8789) );
  XNOR U18755 ( .A(q[6]), .B(DB[1280]), .Z(n8777) );
  IV U18756 ( .A(n8776), .Z(n17685) );
  XNOR U18757 ( .A(n8774), .B(n17686), .Z(n8776) );
  XNOR U18758 ( .A(q[5]), .B(DB[1279]), .Z(n17686) );
  XNOR U18759 ( .A(q[4]), .B(DB[1278]), .Z(n8774) );
  IV U18760 ( .A(n8788), .Z(n17684) );
  XOR U18761 ( .A(n17687), .B(n17688), .Z(n8788) );
  XNOR U18762 ( .A(n8784), .B(n8786), .Z(n17688) );
  XNOR U18763 ( .A(q[0]), .B(DB[1274]), .Z(n8786) );
  XNOR U18764 ( .A(q[3]), .B(DB[1277]), .Z(n8784) );
  IV U18765 ( .A(n8783), .Z(n17687) );
  XNOR U18766 ( .A(n8781), .B(n17689), .Z(n8783) );
  XNOR U18767 ( .A(q[2]), .B(DB[1276]), .Z(n17689) );
  XNOR U18768 ( .A(q[1]), .B(DB[1275]), .Z(n8781) );
  XOR U18769 ( .A(n17690), .B(n8746), .Z(n8709) );
  XOR U18770 ( .A(n17691), .B(n8734), .Z(n8746) );
  XNOR U18771 ( .A(q[6]), .B(DB[1287]), .Z(n8734) );
  IV U18772 ( .A(n8733), .Z(n17691) );
  XNOR U18773 ( .A(n8731), .B(n17692), .Z(n8733) );
  XNOR U18774 ( .A(q[5]), .B(DB[1286]), .Z(n17692) );
  XNOR U18775 ( .A(q[4]), .B(DB[1285]), .Z(n8731) );
  IV U18776 ( .A(n8745), .Z(n17690) );
  XOR U18777 ( .A(n17693), .B(n17694), .Z(n8745) );
  XNOR U18778 ( .A(n8741), .B(n8743), .Z(n17694) );
  XNOR U18779 ( .A(q[0]), .B(DB[1281]), .Z(n8743) );
  XNOR U18780 ( .A(q[3]), .B(DB[1284]), .Z(n8741) );
  IV U18781 ( .A(n8740), .Z(n17693) );
  XNOR U18782 ( .A(n8738), .B(n17695), .Z(n8740) );
  XNOR U18783 ( .A(q[2]), .B(DB[1283]), .Z(n17695) );
  XNOR U18784 ( .A(q[1]), .B(DB[1282]), .Z(n8738) );
  XOR U18785 ( .A(n17696), .B(n8703), .Z(n8666) );
  XOR U18786 ( .A(n17697), .B(n8691), .Z(n8703) );
  XNOR U18787 ( .A(q[6]), .B(DB[1294]), .Z(n8691) );
  IV U18788 ( .A(n8690), .Z(n17697) );
  XNOR U18789 ( .A(n8688), .B(n17698), .Z(n8690) );
  XNOR U18790 ( .A(q[5]), .B(DB[1293]), .Z(n17698) );
  XNOR U18791 ( .A(q[4]), .B(DB[1292]), .Z(n8688) );
  IV U18792 ( .A(n8702), .Z(n17696) );
  XOR U18793 ( .A(n17699), .B(n17700), .Z(n8702) );
  XNOR U18794 ( .A(n8698), .B(n8700), .Z(n17700) );
  XNOR U18795 ( .A(q[0]), .B(DB[1288]), .Z(n8700) );
  XNOR U18796 ( .A(q[3]), .B(DB[1291]), .Z(n8698) );
  IV U18797 ( .A(n8697), .Z(n17699) );
  XNOR U18798 ( .A(n8695), .B(n17701), .Z(n8697) );
  XNOR U18799 ( .A(q[2]), .B(DB[1290]), .Z(n17701) );
  XNOR U18800 ( .A(q[1]), .B(DB[1289]), .Z(n8695) );
  XOR U18801 ( .A(n17702), .B(n8660), .Z(n8623) );
  XOR U18802 ( .A(n17703), .B(n8648), .Z(n8660) );
  XNOR U18803 ( .A(q[6]), .B(DB[1301]), .Z(n8648) );
  IV U18804 ( .A(n8647), .Z(n17703) );
  XNOR U18805 ( .A(n8645), .B(n17704), .Z(n8647) );
  XNOR U18806 ( .A(q[5]), .B(DB[1300]), .Z(n17704) );
  XNOR U18807 ( .A(q[4]), .B(DB[1299]), .Z(n8645) );
  IV U18808 ( .A(n8659), .Z(n17702) );
  XOR U18809 ( .A(n17705), .B(n17706), .Z(n8659) );
  XNOR U18810 ( .A(n8655), .B(n8657), .Z(n17706) );
  XNOR U18811 ( .A(q[0]), .B(DB[1295]), .Z(n8657) );
  XNOR U18812 ( .A(q[3]), .B(DB[1298]), .Z(n8655) );
  IV U18813 ( .A(n8654), .Z(n17705) );
  XNOR U18814 ( .A(n8652), .B(n17707), .Z(n8654) );
  XNOR U18815 ( .A(q[2]), .B(DB[1297]), .Z(n17707) );
  XNOR U18816 ( .A(q[1]), .B(DB[1296]), .Z(n8652) );
  XOR U18817 ( .A(n17708), .B(n8617), .Z(n8580) );
  XOR U18818 ( .A(n17709), .B(n8605), .Z(n8617) );
  XNOR U18819 ( .A(q[6]), .B(DB[1308]), .Z(n8605) );
  IV U18820 ( .A(n8604), .Z(n17709) );
  XNOR U18821 ( .A(n8602), .B(n17710), .Z(n8604) );
  XNOR U18822 ( .A(q[5]), .B(DB[1307]), .Z(n17710) );
  XNOR U18823 ( .A(q[4]), .B(DB[1306]), .Z(n8602) );
  IV U18824 ( .A(n8616), .Z(n17708) );
  XOR U18825 ( .A(n17711), .B(n17712), .Z(n8616) );
  XNOR U18826 ( .A(n8612), .B(n8614), .Z(n17712) );
  XNOR U18827 ( .A(q[0]), .B(DB[1302]), .Z(n8614) );
  XNOR U18828 ( .A(q[3]), .B(DB[1305]), .Z(n8612) );
  IV U18829 ( .A(n8611), .Z(n17711) );
  XNOR U18830 ( .A(n8609), .B(n17713), .Z(n8611) );
  XNOR U18831 ( .A(q[2]), .B(DB[1304]), .Z(n17713) );
  XNOR U18832 ( .A(q[1]), .B(DB[1303]), .Z(n8609) );
  XOR U18833 ( .A(n17714), .B(n8574), .Z(n8537) );
  XOR U18834 ( .A(n17715), .B(n8562), .Z(n8574) );
  XNOR U18835 ( .A(q[6]), .B(DB[1315]), .Z(n8562) );
  IV U18836 ( .A(n8561), .Z(n17715) );
  XNOR U18837 ( .A(n8559), .B(n17716), .Z(n8561) );
  XNOR U18838 ( .A(q[5]), .B(DB[1314]), .Z(n17716) );
  XNOR U18839 ( .A(q[4]), .B(DB[1313]), .Z(n8559) );
  IV U18840 ( .A(n8573), .Z(n17714) );
  XOR U18841 ( .A(n17717), .B(n17718), .Z(n8573) );
  XNOR U18842 ( .A(n8569), .B(n8571), .Z(n17718) );
  XNOR U18843 ( .A(q[0]), .B(DB[1309]), .Z(n8571) );
  XNOR U18844 ( .A(q[3]), .B(DB[1312]), .Z(n8569) );
  IV U18845 ( .A(n8568), .Z(n17717) );
  XNOR U18846 ( .A(n8566), .B(n17719), .Z(n8568) );
  XNOR U18847 ( .A(q[2]), .B(DB[1311]), .Z(n17719) );
  XNOR U18848 ( .A(q[1]), .B(DB[1310]), .Z(n8566) );
  XOR U18849 ( .A(n17720), .B(n8531), .Z(n8494) );
  XOR U18850 ( .A(n17721), .B(n8519), .Z(n8531) );
  XNOR U18851 ( .A(q[6]), .B(DB[1322]), .Z(n8519) );
  IV U18852 ( .A(n8518), .Z(n17721) );
  XNOR U18853 ( .A(n8516), .B(n17722), .Z(n8518) );
  XNOR U18854 ( .A(q[5]), .B(DB[1321]), .Z(n17722) );
  XNOR U18855 ( .A(q[4]), .B(DB[1320]), .Z(n8516) );
  IV U18856 ( .A(n8530), .Z(n17720) );
  XOR U18857 ( .A(n17723), .B(n17724), .Z(n8530) );
  XNOR U18858 ( .A(n8526), .B(n8528), .Z(n17724) );
  XNOR U18859 ( .A(q[0]), .B(DB[1316]), .Z(n8528) );
  XNOR U18860 ( .A(q[3]), .B(DB[1319]), .Z(n8526) );
  IV U18861 ( .A(n8525), .Z(n17723) );
  XNOR U18862 ( .A(n8523), .B(n17725), .Z(n8525) );
  XNOR U18863 ( .A(q[2]), .B(DB[1318]), .Z(n17725) );
  XNOR U18864 ( .A(q[1]), .B(DB[1317]), .Z(n8523) );
  XOR U18865 ( .A(n17726), .B(n8488), .Z(n8451) );
  XOR U18866 ( .A(n17727), .B(n8476), .Z(n8488) );
  XNOR U18867 ( .A(q[6]), .B(DB[1329]), .Z(n8476) );
  IV U18868 ( .A(n8475), .Z(n17727) );
  XNOR U18869 ( .A(n8473), .B(n17728), .Z(n8475) );
  XNOR U18870 ( .A(q[5]), .B(DB[1328]), .Z(n17728) );
  XNOR U18871 ( .A(q[4]), .B(DB[1327]), .Z(n8473) );
  IV U18872 ( .A(n8487), .Z(n17726) );
  XOR U18873 ( .A(n17729), .B(n17730), .Z(n8487) );
  XNOR U18874 ( .A(n8483), .B(n8485), .Z(n17730) );
  XNOR U18875 ( .A(q[0]), .B(DB[1323]), .Z(n8485) );
  XNOR U18876 ( .A(q[3]), .B(DB[1326]), .Z(n8483) );
  IV U18877 ( .A(n8482), .Z(n17729) );
  XNOR U18878 ( .A(n8480), .B(n17731), .Z(n8482) );
  XNOR U18879 ( .A(q[2]), .B(DB[1325]), .Z(n17731) );
  XNOR U18880 ( .A(q[1]), .B(DB[1324]), .Z(n8480) );
  XOR U18881 ( .A(n17732), .B(n8445), .Z(n8408) );
  XOR U18882 ( .A(n17733), .B(n8433), .Z(n8445) );
  XNOR U18883 ( .A(q[6]), .B(DB[1336]), .Z(n8433) );
  IV U18884 ( .A(n8432), .Z(n17733) );
  XNOR U18885 ( .A(n8430), .B(n17734), .Z(n8432) );
  XNOR U18886 ( .A(q[5]), .B(DB[1335]), .Z(n17734) );
  XNOR U18887 ( .A(q[4]), .B(DB[1334]), .Z(n8430) );
  IV U18888 ( .A(n8444), .Z(n17732) );
  XOR U18889 ( .A(n17735), .B(n17736), .Z(n8444) );
  XNOR U18890 ( .A(n8440), .B(n8442), .Z(n17736) );
  XNOR U18891 ( .A(q[0]), .B(DB[1330]), .Z(n8442) );
  XNOR U18892 ( .A(q[3]), .B(DB[1333]), .Z(n8440) );
  IV U18893 ( .A(n8439), .Z(n17735) );
  XNOR U18894 ( .A(n8437), .B(n17737), .Z(n8439) );
  XNOR U18895 ( .A(q[2]), .B(DB[1332]), .Z(n17737) );
  XNOR U18896 ( .A(q[1]), .B(DB[1331]), .Z(n8437) );
  XOR U18897 ( .A(n17738), .B(n8402), .Z(n8365) );
  XOR U18898 ( .A(n17739), .B(n8390), .Z(n8402) );
  XNOR U18899 ( .A(q[6]), .B(DB[1343]), .Z(n8390) );
  IV U18900 ( .A(n8389), .Z(n17739) );
  XNOR U18901 ( .A(n8387), .B(n17740), .Z(n8389) );
  XNOR U18902 ( .A(q[5]), .B(DB[1342]), .Z(n17740) );
  XNOR U18903 ( .A(q[4]), .B(DB[1341]), .Z(n8387) );
  IV U18904 ( .A(n8401), .Z(n17738) );
  XOR U18905 ( .A(n17741), .B(n17742), .Z(n8401) );
  XNOR U18906 ( .A(n8397), .B(n8399), .Z(n17742) );
  XNOR U18907 ( .A(q[0]), .B(DB[1337]), .Z(n8399) );
  XNOR U18908 ( .A(q[3]), .B(DB[1340]), .Z(n8397) );
  IV U18909 ( .A(n8396), .Z(n17741) );
  XNOR U18910 ( .A(n8394), .B(n17743), .Z(n8396) );
  XNOR U18911 ( .A(q[2]), .B(DB[1339]), .Z(n17743) );
  XNOR U18912 ( .A(q[1]), .B(DB[1338]), .Z(n8394) );
  XOR U18913 ( .A(n17744), .B(n8359), .Z(n8322) );
  XOR U18914 ( .A(n17745), .B(n8347), .Z(n8359) );
  XNOR U18915 ( .A(q[6]), .B(DB[1350]), .Z(n8347) );
  IV U18916 ( .A(n8346), .Z(n17745) );
  XNOR U18917 ( .A(n8344), .B(n17746), .Z(n8346) );
  XNOR U18918 ( .A(q[5]), .B(DB[1349]), .Z(n17746) );
  XNOR U18919 ( .A(q[4]), .B(DB[1348]), .Z(n8344) );
  IV U18920 ( .A(n8358), .Z(n17744) );
  XOR U18921 ( .A(n17747), .B(n17748), .Z(n8358) );
  XNOR U18922 ( .A(n8354), .B(n8356), .Z(n17748) );
  XNOR U18923 ( .A(q[0]), .B(DB[1344]), .Z(n8356) );
  XNOR U18924 ( .A(q[3]), .B(DB[1347]), .Z(n8354) );
  IV U18925 ( .A(n8353), .Z(n17747) );
  XNOR U18926 ( .A(n8351), .B(n17749), .Z(n8353) );
  XNOR U18927 ( .A(q[2]), .B(DB[1346]), .Z(n17749) );
  XNOR U18928 ( .A(q[1]), .B(DB[1345]), .Z(n8351) );
  XOR U18929 ( .A(n17750), .B(n8316), .Z(n8279) );
  XOR U18930 ( .A(n17751), .B(n8304), .Z(n8316) );
  XNOR U18931 ( .A(q[6]), .B(DB[1357]), .Z(n8304) );
  IV U18932 ( .A(n8303), .Z(n17751) );
  XNOR U18933 ( .A(n8301), .B(n17752), .Z(n8303) );
  XNOR U18934 ( .A(q[5]), .B(DB[1356]), .Z(n17752) );
  XNOR U18935 ( .A(q[4]), .B(DB[1355]), .Z(n8301) );
  IV U18936 ( .A(n8315), .Z(n17750) );
  XOR U18937 ( .A(n17753), .B(n17754), .Z(n8315) );
  XNOR U18938 ( .A(n8311), .B(n8313), .Z(n17754) );
  XNOR U18939 ( .A(q[0]), .B(DB[1351]), .Z(n8313) );
  XNOR U18940 ( .A(q[3]), .B(DB[1354]), .Z(n8311) );
  IV U18941 ( .A(n8310), .Z(n17753) );
  XNOR U18942 ( .A(n8308), .B(n17755), .Z(n8310) );
  XNOR U18943 ( .A(q[2]), .B(DB[1353]), .Z(n17755) );
  XNOR U18944 ( .A(q[1]), .B(DB[1352]), .Z(n8308) );
  XOR U18945 ( .A(n17756), .B(n8273), .Z(n8236) );
  XOR U18946 ( .A(n17757), .B(n8261), .Z(n8273) );
  XNOR U18947 ( .A(q[6]), .B(DB[1364]), .Z(n8261) );
  IV U18948 ( .A(n8260), .Z(n17757) );
  XNOR U18949 ( .A(n8258), .B(n17758), .Z(n8260) );
  XNOR U18950 ( .A(q[5]), .B(DB[1363]), .Z(n17758) );
  XNOR U18951 ( .A(q[4]), .B(DB[1362]), .Z(n8258) );
  IV U18952 ( .A(n8272), .Z(n17756) );
  XOR U18953 ( .A(n17759), .B(n17760), .Z(n8272) );
  XNOR U18954 ( .A(n8268), .B(n8270), .Z(n17760) );
  XNOR U18955 ( .A(q[0]), .B(DB[1358]), .Z(n8270) );
  XNOR U18956 ( .A(q[3]), .B(DB[1361]), .Z(n8268) );
  IV U18957 ( .A(n8267), .Z(n17759) );
  XNOR U18958 ( .A(n8265), .B(n17761), .Z(n8267) );
  XNOR U18959 ( .A(q[2]), .B(DB[1360]), .Z(n17761) );
  XNOR U18960 ( .A(q[1]), .B(DB[1359]), .Z(n8265) );
  XOR U18961 ( .A(n17762), .B(n8230), .Z(n8193) );
  XOR U18962 ( .A(n17763), .B(n8218), .Z(n8230) );
  XNOR U18963 ( .A(q[6]), .B(DB[1371]), .Z(n8218) );
  IV U18964 ( .A(n8217), .Z(n17763) );
  XNOR U18965 ( .A(n8215), .B(n17764), .Z(n8217) );
  XNOR U18966 ( .A(q[5]), .B(DB[1370]), .Z(n17764) );
  XNOR U18967 ( .A(q[4]), .B(DB[1369]), .Z(n8215) );
  IV U18968 ( .A(n8229), .Z(n17762) );
  XOR U18969 ( .A(n17765), .B(n17766), .Z(n8229) );
  XNOR U18970 ( .A(n8225), .B(n8227), .Z(n17766) );
  XNOR U18971 ( .A(q[0]), .B(DB[1365]), .Z(n8227) );
  XNOR U18972 ( .A(q[3]), .B(DB[1368]), .Z(n8225) );
  IV U18973 ( .A(n8224), .Z(n17765) );
  XNOR U18974 ( .A(n8222), .B(n17767), .Z(n8224) );
  XNOR U18975 ( .A(q[2]), .B(DB[1367]), .Z(n17767) );
  XNOR U18976 ( .A(q[1]), .B(DB[1366]), .Z(n8222) );
  XOR U18977 ( .A(n17768), .B(n8187), .Z(n8150) );
  XOR U18978 ( .A(n17769), .B(n8175), .Z(n8187) );
  XNOR U18979 ( .A(q[6]), .B(DB[1378]), .Z(n8175) );
  IV U18980 ( .A(n8174), .Z(n17769) );
  XNOR U18981 ( .A(n8172), .B(n17770), .Z(n8174) );
  XNOR U18982 ( .A(q[5]), .B(DB[1377]), .Z(n17770) );
  XNOR U18983 ( .A(q[4]), .B(DB[1376]), .Z(n8172) );
  IV U18984 ( .A(n8186), .Z(n17768) );
  XOR U18985 ( .A(n17771), .B(n17772), .Z(n8186) );
  XNOR U18986 ( .A(n8182), .B(n8184), .Z(n17772) );
  XNOR U18987 ( .A(q[0]), .B(DB[1372]), .Z(n8184) );
  XNOR U18988 ( .A(q[3]), .B(DB[1375]), .Z(n8182) );
  IV U18989 ( .A(n8181), .Z(n17771) );
  XNOR U18990 ( .A(n8179), .B(n17773), .Z(n8181) );
  XNOR U18991 ( .A(q[2]), .B(DB[1374]), .Z(n17773) );
  XNOR U18992 ( .A(q[1]), .B(DB[1373]), .Z(n8179) );
  XOR U18993 ( .A(n17774), .B(n8144), .Z(n8107) );
  XOR U18994 ( .A(n17775), .B(n8132), .Z(n8144) );
  XNOR U18995 ( .A(q[6]), .B(DB[1385]), .Z(n8132) );
  IV U18996 ( .A(n8131), .Z(n17775) );
  XNOR U18997 ( .A(n8129), .B(n17776), .Z(n8131) );
  XNOR U18998 ( .A(q[5]), .B(DB[1384]), .Z(n17776) );
  XNOR U18999 ( .A(q[4]), .B(DB[1383]), .Z(n8129) );
  IV U19000 ( .A(n8143), .Z(n17774) );
  XOR U19001 ( .A(n17777), .B(n17778), .Z(n8143) );
  XNOR U19002 ( .A(n8139), .B(n8141), .Z(n17778) );
  XNOR U19003 ( .A(q[0]), .B(DB[1379]), .Z(n8141) );
  XNOR U19004 ( .A(q[3]), .B(DB[1382]), .Z(n8139) );
  IV U19005 ( .A(n8138), .Z(n17777) );
  XNOR U19006 ( .A(n8136), .B(n17779), .Z(n8138) );
  XNOR U19007 ( .A(q[2]), .B(DB[1381]), .Z(n17779) );
  XNOR U19008 ( .A(q[1]), .B(DB[1380]), .Z(n8136) );
  XOR U19009 ( .A(n17780), .B(n8101), .Z(n8064) );
  XOR U19010 ( .A(n17781), .B(n8089), .Z(n8101) );
  XNOR U19011 ( .A(q[6]), .B(DB[1392]), .Z(n8089) );
  IV U19012 ( .A(n8088), .Z(n17781) );
  XNOR U19013 ( .A(n8086), .B(n17782), .Z(n8088) );
  XNOR U19014 ( .A(q[5]), .B(DB[1391]), .Z(n17782) );
  XNOR U19015 ( .A(q[4]), .B(DB[1390]), .Z(n8086) );
  IV U19016 ( .A(n8100), .Z(n17780) );
  XOR U19017 ( .A(n17783), .B(n17784), .Z(n8100) );
  XNOR U19018 ( .A(n8096), .B(n8098), .Z(n17784) );
  XNOR U19019 ( .A(q[0]), .B(DB[1386]), .Z(n8098) );
  XNOR U19020 ( .A(q[3]), .B(DB[1389]), .Z(n8096) );
  IV U19021 ( .A(n8095), .Z(n17783) );
  XNOR U19022 ( .A(n8093), .B(n17785), .Z(n8095) );
  XNOR U19023 ( .A(q[2]), .B(DB[1388]), .Z(n17785) );
  XNOR U19024 ( .A(q[1]), .B(DB[1387]), .Z(n8093) );
  XOR U19025 ( .A(n17786), .B(n8058), .Z(n8021) );
  XOR U19026 ( .A(n17787), .B(n8046), .Z(n8058) );
  XNOR U19027 ( .A(q[6]), .B(DB[1399]), .Z(n8046) );
  IV U19028 ( .A(n8045), .Z(n17787) );
  XNOR U19029 ( .A(n8043), .B(n17788), .Z(n8045) );
  XNOR U19030 ( .A(q[5]), .B(DB[1398]), .Z(n17788) );
  XNOR U19031 ( .A(q[4]), .B(DB[1397]), .Z(n8043) );
  IV U19032 ( .A(n8057), .Z(n17786) );
  XOR U19033 ( .A(n17789), .B(n17790), .Z(n8057) );
  XNOR U19034 ( .A(n8053), .B(n8055), .Z(n17790) );
  XNOR U19035 ( .A(q[0]), .B(DB[1393]), .Z(n8055) );
  XNOR U19036 ( .A(q[3]), .B(DB[1396]), .Z(n8053) );
  IV U19037 ( .A(n8052), .Z(n17789) );
  XNOR U19038 ( .A(n8050), .B(n17791), .Z(n8052) );
  XNOR U19039 ( .A(q[2]), .B(DB[1395]), .Z(n17791) );
  XNOR U19040 ( .A(q[1]), .B(DB[1394]), .Z(n8050) );
  XOR U19041 ( .A(n17792), .B(n8015), .Z(n7978) );
  XOR U19042 ( .A(n17793), .B(n8003), .Z(n8015) );
  XNOR U19043 ( .A(q[6]), .B(DB[1406]), .Z(n8003) );
  IV U19044 ( .A(n8002), .Z(n17793) );
  XNOR U19045 ( .A(n8000), .B(n17794), .Z(n8002) );
  XNOR U19046 ( .A(q[5]), .B(DB[1405]), .Z(n17794) );
  XNOR U19047 ( .A(q[4]), .B(DB[1404]), .Z(n8000) );
  IV U19048 ( .A(n8014), .Z(n17792) );
  XOR U19049 ( .A(n17795), .B(n17796), .Z(n8014) );
  XNOR U19050 ( .A(n8010), .B(n8012), .Z(n17796) );
  XNOR U19051 ( .A(q[0]), .B(DB[1400]), .Z(n8012) );
  XNOR U19052 ( .A(q[3]), .B(DB[1403]), .Z(n8010) );
  IV U19053 ( .A(n8009), .Z(n17795) );
  XNOR U19054 ( .A(n8007), .B(n17797), .Z(n8009) );
  XNOR U19055 ( .A(q[2]), .B(DB[1402]), .Z(n17797) );
  XNOR U19056 ( .A(q[1]), .B(DB[1401]), .Z(n8007) );
  XOR U19057 ( .A(n17798), .B(n7972), .Z(n7935) );
  XOR U19058 ( .A(n17799), .B(n7960), .Z(n7972) );
  XNOR U19059 ( .A(q[6]), .B(DB[1413]), .Z(n7960) );
  IV U19060 ( .A(n7959), .Z(n17799) );
  XNOR U19061 ( .A(n7957), .B(n17800), .Z(n7959) );
  XNOR U19062 ( .A(q[5]), .B(DB[1412]), .Z(n17800) );
  XNOR U19063 ( .A(q[4]), .B(DB[1411]), .Z(n7957) );
  IV U19064 ( .A(n7971), .Z(n17798) );
  XOR U19065 ( .A(n17801), .B(n17802), .Z(n7971) );
  XNOR U19066 ( .A(n7967), .B(n7969), .Z(n17802) );
  XNOR U19067 ( .A(q[0]), .B(DB[1407]), .Z(n7969) );
  XNOR U19068 ( .A(q[3]), .B(DB[1410]), .Z(n7967) );
  IV U19069 ( .A(n7966), .Z(n17801) );
  XNOR U19070 ( .A(n7964), .B(n17803), .Z(n7966) );
  XNOR U19071 ( .A(q[2]), .B(DB[1409]), .Z(n17803) );
  XNOR U19072 ( .A(q[1]), .B(DB[1408]), .Z(n7964) );
  XOR U19073 ( .A(n17804), .B(n7929), .Z(n7892) );
  XOR U19074 ( .A(n17805), .B(n7917), .Z(n7929) );
  XNOR U19075 ( .A(q[6]), .B(DB[1420]), .Z(n7917) );
  IV U19076 ( .A(n7916), .Z(n17805) );
  XNOR U19077 ( .A(n7914), .B(n17806), .Z(n7916) );
  XNOR U19078 ( .A(q[5]), .B(DB[1419]), .Z(n17806) );
  XNOR U19079 ( .A(q[4]), .B(DB[1418]), .Z(n7914) );
  IV U19080 ( .A(n7928), .Z(n17804) );
  XOR U19081 ( .A(n17807), .B(n17808), .Z(n7928) );
  XNOR U19082 ( .A(n7924), .B(n7926), .Z(n17808) );
  XNOR U19083 ( .A(q[0]), .B(DB[1414]), .Z(n7926) );
  XNOR U19084 ( .A(q[3]), .B(DB[1417]), .Z(n7924) );
  IV U19085 ( .A(n7923), .Z(n17807) );
  XNOR U19086 ( .A(n7921), .B(n17809), .Z(n7923) );
  XNOR U19087 ( .A(q[2]), .B(DB[1416]), .Z(n17809) );
  XNOR U19088 ( .A(q[1]), .B(DB[1415]), .Z(n7921) );
  XOR U19089 ( .A(n17810), .B(n7886), .Z(n7849) );
  XOR U19090 ( .A(n17811), .B(n7874), .Z(n7886) );
  XNOR U19091 ( .A(q[6]), .B(DB[1427]), .Z(n7874) );
  IV U19092 ( .A(n7873), .Z(n17811) );
  XNOR U19093 ( .A(n7871), .B(n17812), .Z(n7873) );
  XNOR U19094 ( .A(q[5]), .B(DB[1426]), .Z(n17812) );
  XNOR U19095 ( .A(q[4]), .B(DB[1425]), .Z(n7871) );
  IV U19096 ( .A(n7885), .Z(n17810) );
  XOR U19097 ( .A(n17813), .B(n17814), .Z(n7885) );
  XNOR U19098 ( .A(n7881), .B(n7883), .Z(n17814) );
  XNOR U19099 ( .A(q[0]), .B(DB[1421]), .Z(n7883) );
  XNOR U19100 ( .A(q[3]), .B(DB[1424]), .Z(n7881) );
  IV U19101 ( .A(n7880), .Z(n17813) );
  XNOR U19102 ( .A(n7878), .B(n17815), .Z(n7880) );
  XNOR U19103 ( .A(q[2]), .B(DB[1423]), .Z(n17815) );
  XNOR U19104 ( .A(q[1]), .B(DB[1422]), .Z(n7878) );
  XOR U19105 ( .A(n17816), .B(n7843), .Z(n7806) );
  XOR U19106 ( .A(n17817), .B(n7831), .Z(n7843) );
  XNOR U19107 ( .A(q[6]), .B(DB[1434]), .Z(n7831) );
  IV U19108 ( .A(n7830), .Z(n17817) );
  XNOR U19109 ( .A(n7828), .B(n17818), .Z(n7830) );
  XNOR U19110 ( .A(q[5]), .B(DB[1433]), .Z(n17818) );
  XNOR U19111 ( .A(q[4]), .B(DB[1432]), .Z(n7828) );
  IV U19112 ( .A(n7842), .Z(n17816) );
  XOR U19113 ( .A(n17819), .B(n17820), .Z(n7842) );
  XNOR U19114 ( .A(n7838), .B(n7840), .Z(n17820) );
  XNOR U19115 ( .A(q[0]), .B(DB[1428]), .Z(n7840) );
  XNOR U19116 ( .A(q[3]), .B(DB[1431]), .Z(n7838) );
  IV U19117 ( .A(n7837), .Z(n17819) );
  XNOR U19118 ( .A(n7835), .B(n17821), .Z(n7837) );
  XNOR U19119 ( .A(q[2]), .B(DB[1430]), .Z(n17821) );
  XNOR U19120 ( .A(q[1]), .B(DB[1429]), .Z(n7835) );
  XOR U19121 ( .A(n17822), .B(n7800), .Z(n7763) );
  XOR U19122 ( .A(n17823), .B(n7788), .Z(n7800) );
  XNOR U19123 ( .A(q[6]), .B(DB[1441]), .Z(n7788) );
  IV U19124 ( .A(n7787), .Z(n17823) );
  XNOR U19125 ( .A(n7785), .B(n17824), .Z(n7787) );
  XNOR U19126 ( .A(q[5]), .B(DB[1440]), .Z(n17824) );
  XNOR U19127 ( .A(q[4]), .B(DB[1439]), .Z(n7785) );
  IV U19128 ( .A(n7799), .Z(n17822) );
  XOR U19129 ( .A(n17825), .B(n17826), .Z(n7799) );
  XNOR U19130 ( .A(n7795), .B(n7797), .Z(n17826) );
  XNOR U19131 ( .A(q[0]), .B(DB[1435]), .Z(n7797) );
  XNOR U19132 ( .A(q[3]), .B(DB[1438]), .Z(n7795) );
  IV U19133 ( .A(n7794), .Z(n17825) );
  XNOR U19134 ( .A(n7792), .B(n17827), .Z(n7794) );
  XNOR U19135 ( .A(q[2]), .B(DB[1437]), .Z(n17827) );
  XNOR U19136 ( .A(q[1]), .B(DB[1436]), .Z(n7792) );
  XOR U19137 ( .A(n17828), .B(n7757), .Z(n7720) );
  XOR U19138 ( .A(n17829), .B(n7745), .Z(n7757) );
  XNOR U19139 ( .A(q[6]), .B(DB[1448]), .Z(n7745) );
  IV U19140 ( .A(n7744), .Z(n17829) );
  XNOR U19141 ( .A(n7742), .B(n17830), .Z(n7744) );
  XNOR U19142 ( .A(q[5]), .B(DB[1447]), .Z(n17830) );
  XNOR U19143 ( .A(q[4]), .B(DB[1446]), .Z(n7742) );
  IV U19144 ( .A(n7756), .Z(n17828) );
  XOR U19145 ( .A(n17831), .B(n17832), .Z(n7756) );
  XNOR U19146 ( .A(n7752), .B(n7754), .Z(n17832) );
  XNOR U19147 ( .A(q[0]), .B(DB[1442]), .Z(n7754) );
  XNOR U19148 ( .A(q[3]), .B(DB[1445]), .Z(n7752) );
  IV U19149 ( .A(n7751), .Z(n17831) );
  XNOR U19150 ( .A(n7749), .B(n17833), .Z(n7751) );
  XNOR U19151 ( .A(q[2]), .B(DB[1444]), .Z(n17833) );
  XNOR U19152 ( .A(q[1]), .B(DB[1443]), .Z(n7749) );
  XOR U19153 ( .A(n17834), .B(n7714), .Z(n7677) );
  XOR U19154 ( .A(n17835), .B(n7702), .Z(n7714) );
  XNOR U19155 ( .A(q[6]), .B(DB[1455]), .Z(n7702) );
  IV U19156 ( .A(n7701), .Z(n17835) );
  XNOR U19157 ( .A(n7699), .B(n17836), .Z(n7701) );
  XNOR U19158 ( .A(q[5]), .B(DB[1454]), .Z(n17836) );
  XNOR U19159 ( .A(q[4]), .B(DB[1453]), .Z(n7699) );
  IV U19160 ( .A(n7713), .Z(n17834) );
  XOR U19161 ( .A(n17837), .B(n17838), .Z(n7713) );
  XNOR U19162 ( .A(n7709), .B(n7711), .Z(n17838) );
  XNOR U19163 ( .A(q[0]), .B(DB[1449]), .Z(n7711) );
  XNOR U19164 ( .A(q[3]), .B(DB[1452]), .Z(n7709) );
  IV U19165 ( .A(n7708), .Z(n17837) );
  XNOR U19166 ( .A(n7706), .B(n17839), .Z(n7708) );
  XNOR U19167 ( .A(q[2]), .B(DB[1451]), .Z(n17839) );
  XNOR U19168 ( .A(q[1]), .B(DB[1450]), .Z(n7706) );
  XOR U19169 ( .A(n17840), .B(n7671), .Z(n7634) );
  XOR U19170 ( .A(n17841), .B(n7659), .Z(n7671) );
  XNOR U19171 ( .A(q[6]), .B(DB[1462]), .Z(n7659) );
  IV U19172 ( .A(n7658), .Z(n17841) );
  XNOR U19173 ( .A(n7656), .B(n17842), .Z(n7658) );
  XNOR U19174 ( .A(q[5]), .B(DB[1461]), .Z(n17842) );
  XNOR U19175 ( .A(q[4]), .B(DB[1460]), .Z(n7656) );
  IV U19176 ( .A(n7670), .Z(n17840) );
  XOR U19177 ( .A(n17843), .B(n17844), .Z(n7670) );
  XNOR U19178 ( .A(n7666), .B(n7668), .Z(n17844) );
  XNOR U19179 ( .A(q[0]), .B(DB[1456]), .Z(n7668) );
  XNOR U19180 ( .A(q[3]), .B(DB[1459]), .Z(n7666) );
  IV U19181 ( .A(n7665), .Z(n17843) );
  XNOR U19182 ( .A(n7663), .B(n17845), .Z(n7665) );
  XNOR U19183 ( .A(q[2]), .B(DB[1458]), .Z(n17845) );
  XNOR U19184 ( .A(q[1]), .B(DB[1457]), .Z(n7663) );
  XOR U19185 ( .A(n17846), .B(n7628), .Z(n7591) );
  XOR U19186 ( .A(n17847), .B(n7616), .Z(n7628) );
  XNOR U19187 ( .A(q[6]), .B(DB[1469]), .Z(n7616) );
  IV U19188 ( .A(n7615), .Z(n17847) );
  XNOR U19189 ( .A(n7613), .B(n17848), .Z(n7615) );
  XNOR U19190 ( .A(q[5]), .B(DB[1468]), .Z(n17848) );
  XNOR U19191 ( .A(q[4]), .B(DB[1467]), .Z(n7613) );
  IV U19192 ( .A(n7627), .Z(n17846) );
  XOR U19193 ( .A(n17849), .B(n17850), .Z(n7627) );
  XNOR U19194 ( .A(n7623), .B(n7625), .Z(n17850) );
  XNOR U19195 ( .A(q[0]), .B(DB[1463]), .Z(n7625) );
  XNOR U19196 ( .A(q[3]), .B(DB[1466]), .Z(n7623) );
  IV U19197 ( .A(n7622), .Z(n17849) );
  XNOR U19198 ( .A(n7620), .B(n17851), .Z(n7622) );
  XNOR U19199 ( .A(q[2]), .B(DB[1465]), .Z(n17851) );
  XNOR U19200 ( .A(q[1]), .B(DB[1464]), .Z(n7620) );
  XOR U19201 ( .A(n17852), .B(n7585), .Z(n7548) );
  XOR U19202 ( .A(n17853), .B(n7573), .Z(n7585) );
  XNOR U19203 ( .A(q[6]), .B(DB[1476]), .Z(n7573) );
  IV U19204 ( .A(n7572), .Z(n17853) );
  XNOR U19205 ( .A(n7570), .B(n17854), .Z(n7572) );
  XNOR U19206 ( .A(q[5]), .B(DB[1475]), .Z(n17854) );
  XNOR U19207 ( .A(q[4]), .B(DB[1474]), .Z(n7570) );
  IV U19208 ( .A(n7584), .Z(n17852) );
  XOR U19209 ( .A(n17855), .B(n17856), .Z(n7584) );
  XNOR U19210 ( .A(n7580), .B(n7582), .Z(n17856) );
  XNOR U19211 ( .A(q[0]), .B(DB[1470]), .Z(n7582) );
  XNOR U19212 ( .A(q[3]), .B(DB[1473]), .Z(n7580) );
  IV U19213 ( .A(n7579), .Z(n17855) );
  XNOR U19214 ( .A(n7577), .B(n17857), .Z(n7579) );
  XNOR U19215 ( .A(q[2]), .B(DB[1472]), .Z(n17857) );
  XNOR U19216 ( .A(q[1]), .B(DB[1471]), .Z(n7577) );
  XOR U19217 ( .A(n17858), .B(n7542), .Z(n7505) );
  XOR U19218 ( .A(n17859), .B(n7530), .Z(n7542) );
  XNOR U19219 ( .A(q[6]), .B(DB[1483]), .Z(n7530) );
  IV U19220 ( .A(n7529), .Z(n17859) );
  XNOR U19221 ( .A(n7527), .B(n17860), .Z(n7529) );
  XNOR U19222 ( .A(q[5]), .B(DB[1482]), .Z(n17860) );
  XNOR U19223 ( .A(q[4]), .B(DB[1481]), .Z(n7527) );
  IV U19224 ( .A(n7541), .Z(n17858) );
  XOR U19225 ( .A(n17861), .B(n17862), .Z(n7541) );
  XNOR U19226 ( .A(n7537), .B(n7539), .Z(n17862) );
  XNOR U19227 ( .A(q[0]), .B(DB[1477]), .Z(n7539) );
  XNOR U19228 ( .A(q[3]), .B(DB[1480]), .Z(n7537) );
  IV U19229 ( .A(n7536), .Z(n17861) );
  XNOR U19230 ( .A(n7534), .B(n17863), .Z(n7536) );
  XNOR U19231 ( .A(q[2]), .B(DB[1479]), .Z(n17863) );
  XNOR U19232 ( .A(q[1]), .B(DB[1478]), .Z(n7534) );
  XOR U19233 ( .A(n17864), .B(n7499), .Z(n7462) );
  XOR U19234 ( .A(n17865), .B(n7487), .Z(n7499) );
  XNOR U19235 ( .A(q[6]), .B(DB[1490]), .Z(n7487) );
  IV U19236 ( .A(n7486), .Z(n17865) );
  XNOR U19237 ( .A(n7484), .B(n17866), .Z(n7486) );
  XNOR U19238 ( .A(q[5]), .B(DB[1489]), .Z(n17866) );
  XNOR U19239 ( .A(q[4]), .B(DB[1488]), .Z(n7484) );
  IV U19240 ( .A(n7498), .Z(n17864) );
  XOR U19241 ( .A(n17867), .B(n17868), .Z(n7498) );
  XNOR U19242 ( .A(n7494), .B(n7496), .Z(n17868) );
  XNOR U19243 ( .A(q[0]), .B(DB[1484]), .Z(n7496) );
  XNOR U19244 ( .A(q[3]), .B(DB[1487]), .Z(n7494) );
  IV U19245 ( .A(n7493), .Z(n17867) );
  XNOR U19246 ( .A(n7491), .B(n17869), .Z(n7493) );
  XNOR U19247 ( .A(q[2]), .B(DB[1486]), .Z(n17869) );
  XNOR U19248 ( .A(q[1]), .B(DB[1485]), .Z(n7491) );
  XOR U19249 ( .A(n17870), .B(n7456), .Z(n7419) );
  XOR U19250 ( .A(n17871), .B(n7444), .Z(n7456) );
  XNOR U19251 ( .A(q[6]), .B(DB[1497]), .Z(n7444) );
  IV U19252 ( .A(n7443), .Z(n17871) );
  XNOR U19253 ( .A(n7441), .B(n17872), .Z(n7443) );
  XNOR U19254 ( .A(q[5]), .B(DB[1496]), .Z(n17872) );
  XNOR U19255 ( .A(q[4]), .B(DB[1495]), .Z(n7441) );
  IV U19256 ( .A(n7455), .Z(n17870) );
  XOR U19257 ( .A(n17873), .B(n17874), .Z(n7455) );
  XNOR U19258 ( .A(n7451), .B(n7453), .Z(n17874) );
  XNOR U19259 ( .A(q[0]), .B(DB[1491]), .Z(n7453) );
  XNOR U19260 ( .A(q[3]), .B(DB[1494]), .Z(n7451) );
  IV U19261 ( .A(n7450), .Z(n17873) );
  XNOR U19262 ( .A(n7448), .B(n17875), .Z(n7450) );
  XNOR U19263 ( .A(q[2]), .B(DB[1493]), .Z(n17875) );
  XNOR U19264 ( .A(q[1]), .B(DB[1492]), .Z(n7448) );
  XOR U19265 ( .A(n17876), .B(n7413), .Z(n7376) );
  XOR U19266 ( .A(n17877), .B(n7401), .Z(n7413) );
  XNOR U19267 ( .A(q[6]), .B(DB[1504]), .Z(n7401) );
  IV U19268 ( .A(n7400), .Z(n17877) );
  XNOR U19269 ( .A(n7398), .B(n17878), .Z(n7400) );
  XNOR U19270 ( .A(q[5]), .B(DB[1503]), .Z(n17878) );
  XNOR U19271 ( .A(q[4]), .B(DB[1502]), .Z(n7398) );
  IV U19272 ( .A(n7412), .Z(n17876) );
  XOR U19273 ( .A(n17879), .B(n17880), .Z(n7412) );
  XNOR U19274 ( .A(n7408), .B(n7410), .Z(n17880) );
  XNOR U19275 ( .A(q[0]), .B(DB[1498]), .Z(n7410) );
  XNOR U19276 ( .A(q[3]), .B(DB[1501]), .Z(n7408) );
  IV U19277 ( .A(n7407), .Z(n17879) );
  XNOR U19278 ( .A(n7405), .B(n17881), .Z(n7407) );
  XNOR U19279 ( .A(q[2]), .B(DB[1500]), .Z(n17881) );
  XNOR U19280 ( .A(q[1]), .B(DB[1499]), .Z(n7405) );
  XOR U19281 ( .A(n17882), .B(n7370), .Z(n7333) );
  XOR U19282 ( .A(n17883), .B(n7358), .Z(n7370) );
  XNOR U19283 ( .A(q[6]), .B(DB[1511]), .Z(n7358) );
  IV U19284 ( .A(n7357), .Z(n17883) );
  XNOR U19285 ( .A(n7355), .B(n17884), .Z(n7357) );
  XNOR U19286 ( .A(q[5]), .B(DB[1510]), .Z(n17884) );
  XNOR U19287 ( .A(q[4]), .B(DB[1509]), .Z(n7355) );
  IV U19288 ( .A(n7369), .Z(n17882) );
  XOR U19289 ( .A(n17885), .B(n17886), .Z(n7369) );
  XNOR U19290 ( .A(n7365), .B(n7367), .Z(n17886) );
  XNOR U19291 ( .A(q[0]), .B(DB[1505]), .Z(n7367) );
  XNOR U19292 ( .A(q[3]), .B(DB[1508]), .Z(n7365) );
  IV U19293 ( .A(n7364), .Z(n17885) );
  XNOR U19294 ( .A(n7362), .B(n17887), .Z(n7364) );
  XNOR U19295 ( .A(q[2]), .B(DB[1507]), .Z(n17887) );
  XNOR U19296 ( .A(q[1]), .B(DB[1506]), .Z(n7362) );
  XOR U19297 ( .A(n17888), .B(n7327), .Z(n7290) );
  XOR U19298 ( .A(n17889), .B(n7315), .Z(n7327) );
  XNOR U19299 ( .A(q[6]), .B(DB[1518]), .Z(n7315) );
  IV U19300 ( .A(n7314), .Z(n17889) );
  XNOR U19301 ( .A(n7312), .B(n17890), .Z(n7314) );
  XNOR U19302 ( .A(q[5]), .B(DB[1517]), .Z(n17890) );
  XNOR U19303 ( .A(q[4]), .B(DB[1516]), .Z(n7312) );
  IV U19304 ( .A(n7326), .Z(n17888) );
  XOR U19305 ( .A(n17891), .B(n17892), .Z(n7326) );
  XNOR U19306 ( .A(n7322), .B(n7324), .Z(n17892) );
  XNOR U19307 ( .A(q[0]), .B(DB[1512]), .Z(n7324) );
  XNOR U19308 ( .A(q[3]), .B(DB[1515]), .Z(n7322) );
  IV U19309 ( .A(n7321), .Z(n17891) );
  XNOR U19310 ( .A(n7319), .B(n17893), .Z(n7321) );
  XNOR U19311 ( .A(q[2]), .B(DB[1514]), .Z(n17893) );
  XNOR U19312 ( .A(q[1]), .B(DB[1513]), .Z(n7319) );
  XOR U19313 ( .A(n17894), .B(n7284), .Z(n7247) );
  XOR U19314 ( .A(n17895), .B(n7272), .Z(n7284) );
  XNOR U19315 ( .A(q[6]), .B(DB[1525]), .Z(n7272) );
  IV U19316 ( .A(n7271), .Z(n17895) );
  XNOR U19317 ( .A(n7269), .B(n17896), .Z(n7271) );
  XNOR U19318 ( .A(q[5]), .B(DB[1524]), .Z(n17896) );
  XNOR U19319 ( .A(q[4]), .B(DB[1523]), .Z(n7269) );
  IV U19320 ( .A(n7283), .Z(n17894) );
  XOR U19321 ( .A(n17897), .B(n17898), .Z(n7283) );
  XNOR U19322 ( .A(n7279), .B(n7281), .Z(n17898) );
  XNOR U19323 ( .A(q[0]), .B(DB[1519]), .Z(n7281) );
  XNOR U19324 ( .A(q[3]), .B(DB[1522]), .Z(n7279) );
  IV U19325 ( .A(n7278), .Z(n17897) );
  XNOR U19326 ( .A(n7276), .B(n17899), .Z(n7278) );
  XNOR U19327 ( .A(q[2]), .B(DB[1521]), .Z(n17899) );
  XNOR U19328 ( .A(q[1]), .B(DB[1520]), .Z(n7276) );
  XOR U19329 ( .A(n17900), .B(n7241), .Z(n7204) );
  XOR U19330 ( .A(n17901), .B(n7229), .Z(n7241) );
  XNOR U19331 ( .A(q[6]), .B(DB[1532]), .Z(n7229) );
  IV U19332 ( .A(n7228), .Z(n17901) );
  XNOR U19333 ( .A(n7226), .B(n17902), .Z(n7228) );
  XNOR U19334 ( .A(q[5]), .B(DB[1531]), .Z(n17902) );
  XNOR U19335 ( .A(q[4]), .B(DB[1530]), .Z(n7226) );
  IV U19336 ( .A(n7240), .Z(n17900) );
  XOR U19337 ( .A(n17903), .B(n17904), .Z(n7240) );
  XNOR U19338 ( .A(n7236), .B(n7238), .Z(n17904) );
  XNOR U19339 ( .A(q[0]), .B(DB[1526]), .Z(n7238) );
  XNOR U19340 ( .A(q[3]), .B(DB[1529]), .Z(n7236) );
  IV U19341 ( .A(n7235), .Z(n17903) );
  XNOR U19342 ( .A(n7233), .B(n17905), .Z(n7235) );
  XNOR U19343 ( .A(q[2]), .B(DB[1528]), .Z(n17905) );
  XNOR U19344 ( .A(q[1]), .B(DB[1527]), .Z(n7233) );
  XOR U19345 ( .A(n17906), .B(n7198), .Z(n7161) );
  XOR U19346 ( .A(n17907), .B(n7186), .Z(n7198) );
  XNOR U19347 ( .A(q[6]), .B(DB[1539]), .Z(n7186) );
  IV U19348 ( .A(n7185), .Z(n17907) );
  XNOR U19349 ( .A(n7183), .B(n17908), .Z(n7185) );
  XNOR U19350 ( .A(q[5]), .B(DB[1538]), .Z(n17908) );
  XNOR U19351 ( .A(q[4]), .B(DB[1537]), .Z(n7183) );
  IV U19352 ( .A(n7197), .Z(n17906) );
  XOR U19353 ( .A(n17909), .B(n17910), .Z(n7197) );
  XNOR U19354 ( .A(n7193), .B(n7195), .Z(n17910) );
  XNOR U19355 ( .A(q[0]), .B(DB[1533]), .Z(n7195) );
  XNOR U19356 ( .A(q[3]), .B(DB[1536]), .Z(n7193) );
  IV U19357 ( .A(n7192), .Z(n17909) );
  XNOR U19358 ( .A(n7190), .B(n17911), .Z(n7192) );
  XNOR U19359 ( .A(q[2]), .B(DB[1535]), .Z(n17911) );
  XNOR U19360 ( .A(q[1]), .B(DB[1534]), .Z(n7190) );
  XOR U19361 ( .A(n17912), .B(n7155), .Z(n7118) );
  XOR U19362 ( .A(n17913), .B(n7143), .Z(n7155) );
  XNOR U19363 ( .A(q[6]), .B(DB[1546]), .Z(n7143) );
  IV U19364 ( .A(n7142), .Z(n17913) );
  XNOR U19365 ( .A(n7140), .B(n17914), .Z(n7142) );
  XNOR U19366 ( .A(q[5]), .B(DB[1545]), .Z(n17914) );
  XNOR U19367 ( .A(q[4]), .B(DB[1544]), .Z(n7140) );
  IV U19368 ( .A(n7154), .Z(n17912) );
  XOR U19369 ( .A(n17915), .B(n17916), .Z(n7154) );
  XNOR U19370 ( .A(n7150), .B(n7152), .Z(n17916) );
  XNOR U19371 ( .A(q[0]), .B(DB[1540]), .Z(n7152) );
  XNOR U19372 ( .A(q[3]), .B(DB[1543]), .Z(n7150) );
  IV U19373 ( .A(n7149), .Z(n17915) );
  XNOR U19374 ( .A(n7147), .B(n17917), .Z(n7149) );
  XNOR U19375 ( .A(q[2]), .B(DB[1542]), .Z(n17917) );
  XNOR U19376 ( .A(q[1]), .B(DB[1541]), .Z(n7147) );
  XOR U19377 ( .A(n17918), .B(n7112), .Z(n7075) );
  XOR U19378 ( .A(n17919), .B(n7100), .Z(n7112) );
  XNOR U19379 ( .A(q[6]), .B(DB[1553]), .Z(n7100) );
  IV U19380 ( .A(n7099), .Z(n17919) );
  XNOR U19381 ( .A(n7097), .B(n17920), .Z(n7099) );
  XNOR U19382 ( .A(q[5]), .B(DB[1552]), .Z(n17920) );
  XNOR U19383 ( .A(q[4]), .B(DB[1551]), .Z(n7097) );
  IV U19384 ( .A(n7111), .Z(n17918) );
  XOR U19385 ( .A(n17921), .B(n17922), .Z(n7111) );
  XNOR U19386 ( .A(n7107), .B(n7109), .Z(n17922) );
  XNOR U19387 ( .A(q[0]), .B(DB[1547]), .Z(n7109) );
  XNOR U19388 ( .A(q[3]), .B(DB[1550]), .Z(n7107) );
  IV U19389 ( .A(n7106), .Z(n17921) );
  XNOR U19390 ( .A(n7104), .B(n17923), .Z(n7106) );
  XNOR U19391 ( .A(q[2]), .B(DB[1549]), .Z(n17923) );
  XNOR U19392 ( .A(q[1]), .B(DB[1548]), .Z(n7104) );
  XOR U19393 ( .A(n17924), .B(n7069), .Z(n7032) );
  XOR U19394 ( .A(n17925), .B(n7057), .Z(n7069) );
  XNOR U19395 ( .A(q[6]), .B(DB[1560]), .Z(n7057) );
  IV U19396 ( .A(n7056), .Z(n17925) );
  XNOR U19397 ( .A(n7054), .B(n17926), .Z(n7056) );
  XNOR U19398 ( .A(q[5]), .B(DB[1559]), .Z(n17926) );
  XNOR U19399 ( .A(q[4]), .B(DB[1558]), .Z(n7054) );
  IV U19400 ( .A(n7068), .Z(n17924) );
  XOR U19401 ( .A(n17927), .B(n17928), .Z(n7068) );
  XNOR U19402 ( .A(n7064), .B(n7066), .Z(n17928) );
  XNOR U19403 ( .A(q[0]), .B(DB[1554]), .Z(n7066) );
  XNOR U19404 ( .A(q[3]), .B(DB[1557]), .Z(n7064) );
  IV U19405 ( .A(n7063), .Z(n17927) );
  XNOR U19406 ( .A(n7061), .B(n17929), .Z(n7063) );
  XNOR U19407 ( .A(q[2]), .B(DB[1556]), .Z(n17929) );
  XNOR U19408 ( .A(q[1]), .B(DB[1555]), .Z(n7061) );
  XOR U19409 ( .A(n17930), .B(n7026), .Z(n6989) );
  XOR U19410 ( .A(n17931), .B(n7014), .Z(n7026) );
  XNOR U19411 ( .A(q[6]), .B(DB[1567]), .Z(n7014) );
  IV U19412 ( .A(n7013), .Z(n17931) );
  XNOR U19413 ( .A(n7011), .B(n17932), .Z(n7013) );
  XNOR U19414 ( .A(q[5]), .B(DB[1566]), .Z(n17932) );
  XNOR U19415 ( .A(q[4]), .B(DB[1565]), .Z(n7011) );
  IV U19416 ( .A(n7025), .Z(n17930) );
  XOR U19417 ( .A(n17933), .B(n17934), .Z(n7025) );
  XNOR U19418 ( .A(n7021), .B(n7023), .Z(n17934) );
  XNOR U19419 ( .A(q[0]), .B(DB[1561]), .Z(n7023) );
  XNOR U19420 ( .A(q[3]), .B(DB[1564]), .Z(n7021) );
  IV U19421 ( .A(n7020), .Z(n17933) );
  XNOR U19422 ( .A(n7018), .B(n17935), .Z(n7020) );
  XNOR U19423 ( .A(q[2]), .B(DB[1563]), .Z(n17935) );
  XNOR U19424 ( .A(q[1]), .B(DB[1562]), .Z(n7018) );
  XOR U19425 ( .A(n17936), .B(n6983), .Z(n6946) );
  XOR U19426 ( .A(n17937), .B(n6971), .Z(n6983) );
  XNOR U19427 ( .A(q[6]), .B(DB[1574]), .Z(n6971) );
  IV U19428 ( .A(n6970), .Z(n17937) );
  XNOR U19429 ( .A(n6968), .B(n17938), .Z(n6970) );
  XNOR U19430 ( .A(q[5]), .B(DB[1573]), .Z(n17938) );
  XNOR U19431 ( .A(q[4]), .B(DB[1572]), .Z(n6968) );
  IV U19432 ( .A(n6982), .Z(n17936) );
  XOR U19433 ( .A(n17939), .B(n17940), .Z(n6982) );
  XNOR U19434 ( .A(n6978), .B(n6980), .Z(n17940) );
  XNOR U19435 ( .A(q[0]), .B(DB[1568]), .Z(n6980) );
  XNOR U19436 ( .A(q[3]), .B(DB[1571]), .Z(n6978) );
  IV U19437 ( .A(n6977), .Z(n17939) );
  XNOR U19438 ( .A(n6975), .B(n17941), .Z(n6977) );
  XNOR U19439 ( .A(q[2]), .B(DB[1570]), .Z(n17941) );
  XNOR U19440 ( .A(q[1]), .B(DB[1569]), .Z(n6975) );
  XOR U19441 ( .A(n17942), .B(n6940), .Z(n6903) );
  XOR U19442 ( .A(n17943), .B(n6928), .Z(n6940) );
  XNOR U19443 ( .A(q[6]), .B(DB[1581]), .Z(n6928) );
  IV U19444 ( .A(n6927), .Z(n17943) );
  XNOR U19445 ( .A(n6925), .B(n17944), .Z(n6927) );
  XNOR U19446 ( .A(q[5]), .B(DB[1580]), .Z(n17944) );
  XNOR U19447 ( .A(q[4]), .B(DB[1579]), .Z(n6925) );
  IV U19448 ( .A(n6939), .Z(n17942) );
  XOR U19449 ( .A(n17945), .B(n17946), .Z(n6939) );
  XNOR U19450 ( .A(n6935), .B(n6937), .Z(n17946) );
  XNOR U19451 ( .A(q[0]), .B(DB[1575]), .Z(n6937) );
  XNOR U19452 ( .A(q[3]), .B(DB[1578]), .Z(n6935) );
  IV U19453 ( .A(n6934), .Z(n17945) );
  XNOR U19454 ( .A(n6932), .B(n17947), .Z(n6934) );
  XNOR U19455 ( .A(q[2]), .B(DB[1577]), .Z(n17947) );
  XNOR U19456 ( .A(q[1]), .B(DB[1576]), .Z(n6932) );
  XOR U19457 ( .A(n17948), .B(n6897), .Z(n6860) );
  XOR U19458 ( .A(n17949), .B(n6885), .Z(n6897) );
  XNOR U19459 ( .A(q[6]), .B(DB[1588]), .Z(n6885) );
  IV U19460 ( .A(n6884), .Z(n17949) );
  XNOR U19461 ( .A(n6882), .B(n17950), .Z(n6884) );
  XNOR U19462 ( .A(q[5]), .B(DB[1587]), .Z(n17950) );
  XNOR U19463 ( .A(q[4]), .B(DB[1586]), .Z(n6882) );
  IV U19464 ( .A(n6896), .Z(n17948) );
  XOR U19465 ( .A(n17951), .B(n17952), .Z(n6896) );
  XNOR U19466 ( .A(n6892), .B(n6894), .Z(n17952) );
  XNOR U19467 ( .A(q[0]), .B(DB[1582]), .Z(n6894) );
  XNOR U19468 ( .A(q[3]), .B(DB[1585]), .Z(n6892) );
  IV U19469 ( .A(n6891), .Z(n17951) );
  XNOR U19470 ( .A(n6889), .B(n17953), .Z(n6891) );
  XNOR U19471 ( .A(q[2]), .B(DB[1584]), .Z(n17953) );
  XNOR U19472 ( .A(q[1]), .B(DB[1583]), .Z(n6889) );
  XOR U19473 ( .A(n17954), .B(n6854), .Z(n6817) );
  XOR U19474 ( .A(n17955), .B(n6842), .Z(n6854) );
  XNOR U19475 ( .A(q[6]), .B(DB[1595]), .Z(n6842) );
  IV U19476 ( .A(n6841), .Z(n17955) );
  XNOR U19477 ( .A(n6839), .B(n17956), .Z(n6841) );
  XNOR U19478 ( .A(q[5]), .B(DB[1594]), .Z(n17956) );
  XNOR U19479 ( .A(q[4]), .B(DB[1593]), .Z(n6839) );
  IV U19480 ( .A(n6853), .Z(n17954) );
  XOR U19481 ( .A(n17957), .B(n17958), .Z(n6853) );
  XNOR U19482 ( .A(n6849), .B(n6851), .Z(n17958) );
  XNOR U19483 ( .A(q[0]), .B(DB[1589]), .Z(n6851) );
  XNOR U19484 ( .A(q[3]), .B(DB[1592]), .Z(n6849) );
  IV U19485 ( .A(n6848), .Z(n17957) );
  XNOR U19486 ( .A(n6846), .B(n17959), .Z(n6848) );
  XNOR U19487 ( .A(q[2]), .B(DB[1591]), .Z(n17959) );
  XNOR U19488 ( .A(q[1]), .B(DB[1590]), .Z(n6846) );
  XOR U19489 ( .A(n17960), .B(n6811), .Z(n6774) );
  XOR U19490 ( .A(n17961), .B(n6799), .Z(n6811) );
  XNOR U19491 ( .A(q[6]), .B(DB[1602]), .Z(n6799) );
  IV U19492 ( .A(n6798), .Z(n17961) );
  XNOR U19493 ( .A(n6796), .B(n17962), .Z(n6798) );
  XNOR U19494 ( .A(q[5]), .B(DB[1601]), .Z(n17962) );
  XNOR U19495 ( .A(q[4]), .B(DB[1600]), .Z(n6796) );
  IV U19496 ( .A(n6810), .Z(n17960) );
  XOR U19497 ( .A(n17963), .B(n17964), .Z(n6810) );
  XNOR U19498 ( .A(n6806), .B(n6808), .Z(n17964) );
  XNOR U19499 ( .A(q[0]), .B(DB[1596]), .Z(n6808) );
  XNOR U19500 ( .A(q[3]), .B(DB[1599]), .Z(n6806) );
  IV U19501 ( .A(n6805), .Z(n17963) );
  XNOR U19502 ( .A(n6803), .B(n17965), .Z(n6805) );
  XNOR U19503 ( .A(q[2]), .B(DB[1598]), .Z(n17965) );
  XNOR U19504 ( .A(q[1]), .B(DB[1597]), .Z(n6803) );
  XOR U19505 ( .A(n17966), .B(n6768), .Z(n6731) );
  XOR U19506 ( .A(n17967), .B(n6756), .Z(n6768) );
  XNOR U19507 ( .A(q[6]), .B(DB[1609]), .Z(n6756) );
  IV U19508 ( .A(n6755), .Z(n17967) );
  XNOR U19509 ( .A(n6753), .B(n17968), .Z(n6755) );
  XNOR U19510 ( .A(q[5]), .B(DB[1608]), .Z(n17968) );
  XNOR U19511 ( .A(q[4]), .B(DB[1607]), .Z(n6753) );
  IV U19512 ( .A(n6767), .Z(n17966) );
  XOR U19513 ( .A(n17969), .B(n17970), .Z(n6767) );
  XNOR U19514 ( .A(n6763), .B(n6765), .Z(n17970) );
  XNOR U19515 ( .A(q[0]), .B(DB[1603]), .Z(n6765) );
  XNOR U19516 ( .A(q[3]), .B(DB[1606]), .Z(n6763) );
  IV U19517 ( .A(n6762), .Z(n17969) );
  XNOR U19518 ( .A(n6760), .B(n17971), .Z(n6762) );
  XNOR U19519 ( .A(q[2]), .B(DB[1605]), .Z(n17971) );
  XNOR U19520 ( .A(q[1]), .B(DB[1604]), .Z(n6760) );
  XOR U19521 ( .A(n17972), .B(n6725), .Z(n6688) );
  XOR U19522 ( .A(n17973), .B(n6713), .Z(n6725) );
  XNOR U19523 ( .A(q[6]), .B(DB[1616]), .Z(n6713) );
  IV U19524 ( .A(n6712), .Z(n17973) );
  XNOR U19525 ( .A(n6710), .B(n17974), .Z(n6712) );
  XNOR U19526 ( .A(q[5]), .B(DB[1615]), .Z(n17974) );
  XNOR U19527 ( .A(q[4]), .B(DB[1614]), .Z(n6710) );
  IV U19528 ( .A(n6724), .Z(n17972) );
  XOR U19529 ( .A(n17975), .B(n17976), .Z(n6724) );
  XNOR U19530 ( .A(n6720), .B(n6722), .Z(n17976) );
  XNOR U19531 ( .A(q[0]), .B(DB[1610]), .Z(n6722) );
  XNOR U19532 ( .A(q[3]), .B(DB[1613]), .Z(n6720) );
  IV U19533 ( .A(n6719), .Z(n17975) );
  XNOR U19534 ( .A(n6717), .B(n17977), .Z(n6719) );
  XNOR U19535 ( .A(q[2]), .B(DB[1612]), .Z(n17977) );
  XNOR U19536 ( .A(q[1]), .B(DB[1611]), .Z(n6717) );
  XOR U19537 ( .A(n17978), .B(n6682), .Z(n6645) );
  XOR U19538 ( .A(n17979), .B(n6670), .Z(n6682) );
  XNOR U19539 ( .A(q[6]), .B(DB[1623]), .Z(n6670) );
  IV U19540 ( .A(n6669), .Z(n17979) );
  XNOR U19541 ( .A(n6667), .B(n17980), .Z(n6669) );
  XNOR U19542 ( .A(q[5]), .B(DB[1622]), .Z(n17980) );
  XNOR U19543 ( .A(q[4]), .B(DB[1621]), .Z(n6667) );
  IV U19544 ( .A(n6681), .Z(n17978) );
  XOR U19545 ( .A(n17981), .B(n17982), .Z(n6681) );
  XNOR U19546 ( .A(n6677), .B(n6679), .Z(n17982) );
  XNOR U19547 ( .A(q[0]), .B(DB[1617]), .Z(n6679) );
  XNOR U19548 ( .A(q[3]), .B(DB[1620]), .Z(n6677) );
  IV U19549 ( .A(n6676), .Z(n17981) );
  XNOR U19550 ( .A(n6674), .B(n17983), .Z(n6676) );
  XNOR U19551 ( .A(q[2]), .B(DB[1619]), .Z(n17983) );
  XNOR U19552 ( .A(q[1]), .B(DB[1618]), .Z(n6674) );
  XOR U19553 ( .A(n17984), .B(n6639), .Z(n6602) );
  XOR U19554 ( .A(n17985), .B(n6627), .Z(n6639) );
  XNOR U19555 ( .A(q[6]), .B(DB[1630]), .Z(n6627) );
  IV U19556 ( .A(n6626), .Z(n17985) );
  XNOR U19557 ( .A(n6624), .B(n17986), .Z(n6626) );
  XNOR U19558 ( .A(q[5]), .B(DB[1629]), .Z(n17986) );
  XNOR U19559 ( .A(q[4]), .B(DB[1628]), .Z(n6624) );
  IV U19560 ( .A(n6638), .Z(n17984) );
  XOR U19561 ( .A(n17987), .B(n17988), .Z(n6638) );
  XNOR U19562 ( .A(n6634), .B(n6636), .Z(n17988) );
  XNOR U19563 ( .A(q[0]), .B(DB[1624]), .Z(n6636) );
  XNOR U19564 ( .A(q[3]), .B(DB[1627]), .Z(n6634) );
  IV U19565 ( .A(n6633), .Z(n17987) );
  XNOR U19566 ( .A(n6631), .B(n17989), .Z(n6633) );
  XNOR U19567 ( .A(q[2]), .B(DB[1626]), .Z(n17989) );
  XNOR U19568 ( .A(q[1]), .B(DB[1625]), .Z(n6631) );
  XOR U19569 ( .A(n17990), .B(n6596), .Z(n6559) );
  XOR U19570 ( .A(n17991), .B(n6584), .Z(n6596) );
  XNOR U19571 ( .A(q[6]), .B(DB[1637]), .Z(n6584) );
  IV U19572 ( .A(n6583), .Z(n17991) );
  XNOR U19573 ( .A(n6581), .B(n17992), .Z(n6583) );
  XNOR U19574 ( .A(q[5]), .B(DB[1636]), .Z(n17992) );
  XNOR U19575 ( .A(q[4]), .B(DB[1635]), .Z(n6581) );
  IV U19576 ( .A(n6595), .Z(n17990) );
  XOR U19577 ( .A(n17993), .B(n17994), .Z(n6595) );
  XNOR U19578 ( .A(n6591), .B(n6593), .Z(n17994) );
  XNOR U19579 ( .A(q[0]), .B(DB[1631]), .Z(n6593) );
  XNOR U19580 ( .A(q[3]), .B(DB[1634]), .Z(n6591) );
  IV U19581 ( .A(n6590), .Z(n17993) );
  XNOR U19582 ( .A(n6588), .B(n17995), .Z(n6590) );
  XNOR U19583 ( .A(q[2]), .B(DB[1633]), .Z(n17995) );
  XNOR U19584 ( .A(q[1]), .B(DB[1632]), .Z(n6588) );
  XOR U19585 ( .A(n17996), .B(n6553), .Z(n6516) );
  XOR U19586 ( .A(n17997), .B(n6541), .Z(n6553) );
  XNOR U19587 ( .A(q[6]), .B(DB[1644]), .Z(n6541) );
  IV U19588 ( .A(n6540), .Z(n17997) );
  XNOR U19589 ( .A(n6538), .B(n17998), .Z(n6540) );
  XNOR U19590 ( .A(q[5]), .B(DB[1643]), .Z(n17998) );
  XNOR U19591 ( .A(q[4]), .B(DB[1642]), .Z(n6538) );
  IV U19592 ( .A(n6552), .Z(n17996) );
  XOR U19593 ( .A(n17999), .B(n18000), .Z(n6552) );
  XNOR U19594 ( .A(n6548), .B(n6550), .Z(n18000) );
  XNOR U19595 ( .A(q[0]), .B(DB[1638]), .Z(n6550) );
  XNOR U19596 ( .A(q[3]), .B(DB[1641]), .Z(n6548) );
  IV U19597 ( .A(n6547), .Z(n17999) );
  XNOR U19598 ( .A(n6545), .B(n18001), .Z(n6547) );
  XNOR U19599 ( .A(q[2]), .B(DB[1640]), .Z(n18001) );
  XNOR U19600 ( .A(q[1]), .B(DB[1639]), .Z(n6545) );
  XOR U19601 ( .A(n18002), .B(n6510), .Z(n6473) );
  XOR U19602 ( .A(n18003), .B(n6498), .Z(n6510) );
  XNOR U19603 ( .A(q[6]), .B(DB[1651]), .Z(n6498) );
  IV U19604 ( .A(n6497), .Z(n18003) );
  XNOR U19605 ( .A(n6495), .B(n18004), .Z(n6497) );
  XNOR U19606 ( .A(q[5]), .B(DB[1650]), .Z(n18004) );
  XNOR U19607 ( .A(q[4]), .B(DB[1649]), .Z(n6495) );
  IV U19608 ( .A(n6509), .Z(n18002) );
  XOR U19609 ( .A(n18005), .B(n18006), .Z(n6509) );
  XNOR U19610 ( .A(n6505), .B(n6507), .Z(n18006) );
  XNOR U19611 ( .A(q[0]), .B(DB[1645]), .Z(n6507) );
  XNOR U19612 ( .A(q[3]), .B(DB[1648]), .Z(n6505) );
  IV U19613 ( .A(n6504), .Z(n18005) );
  XNOR U19614 ( .A(n6502), .B(n18007), .Z(n6504) );
  XNOR U19615 ( .A(q[2]), .B(DB[1647]), .Z(n18007) );
  XNOR U19616 ( .A(q[1]), .B(DB[1646]), .Z(n6502) );
  XOR U19617 ( .A(n18008), .B(n6467), .Z(n6430) );
  XOR U19618 ( .A(n18009), .B(n6455), .Z(n6467) );
  XNOR U19619 ( .A(q[6]), .B(DB[1658]), .Z(n6455) );
  IV U19620 ( .A(n6454), .Z(n18009) );
  XNOR U19621 ( .A(n6452), .B(n18010), .Z(n6454) );
  XNOR U19622 ( .A(q[5]), .B(DB[1657]), .Z(n18010) );
  XNOR U19623 ( .A(q[4]), .B(DB[1656]), .Z(n6452) );
  IV U19624 ( .A(n6466), .Z(n18008) );
  XOR U19625 ( .A(n18011), .B(n18012), .Z(n6466) );
  XNOR U19626 ( .A(n6462), .B(n6464), .Z(n18012) );
  XNOR U19627 ( .A(q[0]), .B(DB[1652]), .Z(n6464) );
  XNOR U19628 ( .A(q[3]), .B(DB[1655]), .Z(n6462) );
  IV U19629 ( .A(n6461), .Z(n18011) );
  XNOR U19630 ( .A(n6459), .B(n18013), .Z(n6461) );
  XNOR U19631 ( .A(q[2]), .B(DB[1654]), .Z(n18013) );
  XNOR U19632 ( .A(q[1]), .B(DB[1653]), .Z(n6459) );
  XOR U19633 ( .A(n18014), .B(n6424), .Z(n6387) );
  XOR U19634 ( .A(n18015), .B(n6412), .Z(n6424) );
  XNOR U19635 ( .A(q[6]), .B(DB[1665]), .Z(n6412) );
  IV U19636 ( .A(n6411), .Z(n18015) );
  XNOR U19637 ( .A(n6409), .B(n18016), .Z(n6411) );
  XNOR U19638 ( .A(q[5]), .B(DB[1664]), .Z(n18016) );
  XNOR U19639 ( .A(q[4]), .B(DB[1663]), .Z(n6409) );
  IV U19640 ( .A(n6423), .Z(n18014) );
  XOR U19641 ( .A(n18017), .B(n18018), .Z(n6423) );
  XNOR U19642 ( .A(n6419), .B(n6421), .Z(n18018) );
  XNOR U19643 ( .A(q[0]), .B(DB[1659]), .Z(n6421) );
  XNOR U19644 ( .A(q[3]), .B(DB[1662]), .Z(n6419) );
  IV U19645 ( .A(n6418), .Z(n18017) );
  XNOR U19646 ( .A(n6416), .B(n18019), .Z(n6418) );
  XNOR U19647 ( .A(q[2]), .B(DB[1661]), .Z(n18019) );
  XNOR U19648 ( .A(q[1]), .B(DB[1660]), .Z(n6416) );
  XOR U19649 ( .A(n18020), .B(n6381), .Z(n6344) );
  XOR U19650 ( .A(n18021), .B(n6369), .Z(n6381) );
  XNOR U19651 ( .A(q[6]), .B(DB[1672]), .Z(n6369) );
  IV U19652 ( .A(n6368), .Z(n18021) );
  XNOR U19653 ( .A(n6366), .B(n18022), .Z(n6368) );
  XNOR U19654 ( .A(q[5]), .B(DB[1671]), .Z(n18022) );
  XNOR U19655 ( .A(q[4]), .B(DB[1670]), .Z(n6366) );
  IV U19656 ( .A(n6380), .Z(n18020) );
  XOR U19657 ( .A(n18023), .B(n18024), .Z(n6380) );
  XNOR U19658 ( .A(n6376), .B(n6378), .Z(n18024) );
  XNOR U19659 ( .A(q[0]), .B(DB[1666]), .Z(n6378) );
  XNOR U19660 ( .A(q[3]), .B(DB[1669]), .Z(n6376) );
  IV U19661 ( .A(n6375), .Z(n18023) );
  XNOR U19662 ( .A(n6373), .B(n18025), .Z(n6375) );
  XNOR U19663 ( .A(q[2]), .B(DB[1668]), .Z(n18025) );
  XNOR U19664 ( .A(q[1]), .B(DB[1667]), .Z(n6373) );
  XOR U19665 ( .A(n18026), .B(n6338), .Z(n6301) );
  XOR U19666 ( .A(n18027), .B(n6326), .Z(n6338) );
  XNOR U19667 ( .A(q[6]), .B(DB[1679]), .Z(n6326) );
  IV U19668 ( .A(n6325), .Z(n18027) );
  XNOR U19669 ( .A(n6323), .B(n18028), .Z(n6325) );
  XNOR U19670 ( .A(q[5]), .B(DB[1678]), .Z(n18028) );
  XNOR U19671 ( .A(q[4]), .B(DB[1677]), .Z(n6323) );
  IV U19672 ( .A(n6337), .Z(n18026) );
  XOR U19673 ( .A(n18029), .B(n18030), .Z(n6337) );
  XNOR U19674 ( .A(n6333), .B(n6335), .Z(n18030) );
  XNOR U19675 ( .A(q[0]), .B(DB[1673]), .Z(n6335) );
  XNOR U19676 ( .A(q[3]), .B(DB[1676]), .Z(n6333) );
  IV U19677 ( .A(n6332), .Z(n18029) );
  XNOR U19678 ( .A(n6330), .B(n18031), .Z(n6332) );
  XNOR U19679 ( .A(q[2]), .B(DB[1675]), .Z(n18031) );
  XNOR U19680 ( .A(q[1]), .B(DB[1674]), .Z(n6330) );
  XOR U19681 ( .A(n18032), .B(n6295), .Z(n6258) );
  XOR U19682 ( .A(n18033), .B(n6283), .Z(n6295) );
  XNOR U19683 ( .A(q[6]), .B(DB[1686]), .Z(n6283) );
  IV U19684 ( .A(n6282), .Z(n18033) );
  XNOR U19685 ( .A(n6280), .B(n18034), .Z(n6282) );
  XNOR U19686 ( .A(q[5]), .B(DB[1685]), .Z(n18034) );
  XNOR U19687 ( .A(q[4]), .B(DB[1684]), .Z(n6280) );
  IV U19688 ( .A(n6294), .Z(n18032) );
  XOR U19689 ( .A(n18035), .B(n18036), .Z(n6294) );
  XNOR U19690 ( .A(n6290), .B(n6292), .Z(n18036) );
  XNOR U19691 ( .A(q[0]), .B(DB[1680]), .Z(n6292) );
  XNOR U19692 ( .A(q[3]), .B(DB[1683]), .Z(n6290) );
  IV U19693 ( .A(n6289), .Z(n18035) );
  XNOR U19694 ( .A(n6287), .B(n18037), .Z(n6289) );
  XNOR U19695 ( .A(q[2]), .B(DB[1682]), .Z(n18037) );
  XNOR U19696 ( .A(q[1]), .B(DB[1681]), .Z(n6287) );
  XOR U19697 ( .A(n18038), .B(n6252), .Z(n6215) );
  XOR U19698 ( .A(n18039), .B(n6240), .Z(n6252) );
  XNOR U19699 ( .A(q[6]), .B(DB[1693]), .Z(n6240) );
  IV U19700 ( .A(n6239), .Z(n18039) );
  XNOR U19701 ( .A(n6237), .B(n18040), .Z(n6239) );
  XNOR U19702 ( .A(q[5]), .B(DB[1692]), .Z(n18040) );
  XNOR U19703 ( .A(q[4]), .B(DB[1691]), .Z(n6237) );
  IV U19704 ( .A(n6251), .Z(n18038) );
  XOR U19705 ( .A(n18041), .B(n18042), .Z(n6251) );
  XNOR U19706 ( .A(n6247), .B(n6249), .Z(n18042) );
  XNOR U19707 ( .A(q[0]), .B(DB[1687]), .Z(n6249) );
  XNOR U19708 ( .A(q[3]), .B(DB[1690]), .Z(n6247) );
  IV U19709 ( .A(n6246), .Z(n18041) );
  XNOR U19710 ( .A(n6244), .B(n18043), .Z(n6246) );
  XNOR U19711 ( .A(q[2]), .B(DB[1689]), .Z(n18043) );
  XNOR U19712 ( .A(q[1]), .B(DB[1688]), .Z(n6244) );
  XOR U19713 ( .A(n18044), .B(n6209), .Z(n6172) );
  XOR U19714 ( .A(n18045), .B(n6197), .Z(n6209) );
  XNOR U19715 ( .A(q[6]), .B(DB[1700]), .Z(n6197) );
  IV U19716 ( .A(n6196), .Z(n18045) );
  XNOR U19717 ( .A(n6194), .B(n18046), .Z(n6196) );
  XNOR U19718 ( .A(q[5]), .B(DB[1699]), .Z(n18046) );
  XNOR U19719 ( .A(q[4]), .B(DB[1698]), .Z(n6194) );
  IV U19720 ( .A(n6208), .Z(n18044) );
  XOR U19721 ( .A(n18047), .B(n18048), .Z(n6208) );
  XNOR U19722 ( .A(n6204), .B(n6206), .Z(n18048) );
  XNOR U19723 ( .A(q[0]), .B(DB[1694]), .Z(n6206) );
  XNOR U19724 ( .A(q[3]), .B(DB[1697]), .Z(n6204) );
  IV U19725 ( .A(n6203), .Z(n18047) );
  XNOR U19726 ( .A(n6201), .B(n18049), .Z(n6203) );
  XNOR U19727 ( .A(q[2]), .B(DB[1696]), .Z(n18049) );
  XNOR U19728 ( .A(q[1]), .B(DB[1695]), .Z(n6201) );
  XOR U19729 ( .A(n18050), .B(n6166), .Z(n6129) );
  XOR U19730 ( .A(n18051), .B(n6154), .Z(n6166) );
  XNOR U19731 ( .A(q[6]), .B(DB[1707]), .Z(n6154) );
  IV U19732 ( .A(n6153), .Z(n18051) );
  XNOR U19733 ( .A(n6151), .B(n18052), .Z(n6153) );
  XNOR U19734 ( .A(q[5]), .B(DB[1706]), .Z(n18052) );
  XNOR U19735 ( .A(q[4]), .B(DB[1705]), .Z(n6151) );
  IV U19736 ( .A(n6165), .Z(n18050) );
  XOR U19737 ( .A(n18053), .B(n18054), .Z(n6165) );
  XNOR U19738 ( .A(n6161), .B(n6163), .Z(n18054) );
  XNOR U19739 ( .A(q[0]), .B(DB[1701]), .Z(n6163) );
  XNOR U19740 ( .A(q[3]), .B(DB[1704]), .Z(n6161) );
  IV U19741 ( .A(n6160), .Z(n18053) );
  XNOR U19742 ( .A(n6158), .B(n18055), .Z(n6160) );
  XNOR U19743 ( .A(q[2]), .B(DB[1703]), .Z(n18055) );
  XNOR U19744 ( .A(q[1]), .B(DB[1702]), .Z(n6158) );
  XOR U19745 ( .A(n18056), .B(n6123), .Z(n6086) );
  XOR U19746 ( .A(n18057), .B(n6111), .Z(n6123) );
  XNOR U19747 ( .A(q[6]), .B(DB[1714]), .Z(n6111) );
  IV U19748 ( .A(n6110), .Z(n18057) );
  XNOR U19749 ( .A(n6108), .B(n18058), .Z(n6110) );
  XNOR U19750 ( .A(q[5]), .B(DB[1713]), .Z(n18058) );
  XNOR U19751 ( .A(q[4]), .B(DB[1712]), .Z(n6108) );
  IV U19752 ( .A(n6122), .Z(n18056) );
  XOR U19753 ( .A(n18059), .B(n18060), .Z(n6122) );
  XNOR U19754 ( .A(n6118), .B(n6120), .Z(n18060) );
  XNOR U19755 ( .A(q[0]), .B(DB[1708]), .Z(n6120) );
  XNOR U19756 ( .A(q[3]), .B(DB[1711]), .Z(n6118) );
  IV U19757 ( .A(n6117), .Z(n18059) );
  XNOR U19758 ( .A(n6115), .B(n18061), .Z(n6117) );
  XNOR U19759 ( .A(q[2]), .B(DB[1710]), .Z(n18061) );
  XNOR U19760 ( .A(q[1]), .B(DB[1709]), .Z(n6115) );
  XOR U19761 ( .A(n18062), .B(n6080), .Z(n6043) );
  XOR U19762 ( .A(n18063), .B(n6068), .Z(n6080) );
  XNOR U19763 ( .A(q[6]), .B(DB[1721]), .Z(n6068) );
  IV U19764 ( .A(n6067), .Z(n18063) );
  XNOR U19765 ( .A(n6065), .B(n18064), .Z(n6067) );
  XNOR U19766 ( .A(q[5]), .B(DB[1720]), .Z(n18064) );
  XNOR U19767 ( .A(q[4]), .B(DB[1719]), .Z(n6065) );
  IV U19768 ( .A(n6079), .Z(n18062) );
  XOR U19769 ( .A(n18065), .B(n18066), .Z(n6079) );
  XNOR U19770 ( .A(n6075), .B(n6077), .Z(n18066) );
  XNOR U19771 ( .A(q[0]), .B(DB[1715]), .Z(n6077) );
  XNOR U19772 ( .A(q[3]), .B(DB[1718]), .Z(n6075) );
  IV U19773 ( .A(n6074), .Z(n18065) );
  XNOR U19774 ( .A(n6072), .B(n18067), .Z(n6074) );
  XNOR U19775 ( .A(q[2]), .B(DB[1717]), .Z(n18067) );
  XNOR U19776 ( .A(q[1]), .B(DB[1716]), .Z(n6072) );
  XOR U19777 ( .A(n18068), .B(n6037), .Z(n6000) );
  XOR U19778 ( .A(n18069), .B(n6025), .Z(n6037) );
  XNOR U19779 ( .A(q[6]), .B(DB[1728]), .Z(n6025) );
  IV U19780 ( .A(n6024), .Z(n18069) );
  XNOR U19781 ( .A(n6022), .B(n18070), .Z(n6024) );
  XNOR U19782 ( .A(q[5]), .B(DB[1727]), .Z(n18070) );
  XNOR U19783 ( .A(q[4]), .B(DB[1726]), .Z(n6022) );
  IV U19784 ( .A(n6036), .Z(n18068) );
  XOR U19785 ( .A(n18071), .B(n18072), .Z(n6036) );
  XNOR U19786 ( .A(n6032), .B(n6034), .Z(n18072) );
  XNOR U19787 ( .A(q[0]), .B(DB[1722]), .Z(n6034) );
  XNOR U19788 ( .A(q[3]), .B(DB[1725]), .Z(n6032) );
  IV U19789 ( .A(n6031), .Z(n18071) );
  XNOR U19790 ( .A(n6029), .B(n18073), .Z(n6031) );
  XNOR U19791 ( .A(q[2]), .B(DB[1724]), .Z(n18073) );
  XNOR U19792 ( .A(q[1]), .B(DB[1723]), .Z(n6029) );
  XOR U19793 ( .A(n18074), .B(n5994), .Z(n5957) );
  XOR U19794 ( .A(n18075), .B(n5982), .Z(n5994) );
  XNOR U19795 ( .A(q[6]), .B(DB[1735]), .Z(n5982) );
  IV U19796 ( .A(n5981), .Z(n18075) );
  XNOR U19797 ( .A(n5979), .B(n18076), .Z(n5981) );
  XNOR U19798 ( .A(q[5]), .B(DB[1734]), .Z(n18076) );
  XNOR U19799 ( .A(q[4]), .B(DB[1733]), .Z(n5979) );
  IV U19800 ( .A(n5993), .Z(n18074) );
  XOR U19801 ( .A(n18077), .B(n18078), .Z(n5993) );
  XNOR U19802 ( .A(n5989), .B(n5991), .Z(n18078) );
  XNOR U19803 ( .A(q[0]), .B(DB[1729]), .Z(n5991) );
  XNOR U19804 ( .A(q[3]), .B(DB[1732]), .Z(n5989) );
  IV U19805 ( .A(n5988), .Z(n18077) );
  XNOR U19806 ( .A(n5986), .B(n18079), .Z(n5988) );
  XNOR U19807 ( .A(q[2]), .B(DB[1731]), .Z(n18079) );
  XNOR U19808 ( .A(q[1]), .B(DB[1730]), .Z(n5986) );
  XOR U19809 ( .A(n18080), .B(n5951), .Z(n5914) );
  XOR U19810 ( .A(n18081), .B(n5939), .Z(n5951) );
  XNOR U19811 ( .A(q[6]), .B(DB[1742]), .Z(n5939) );
  IV U19812 ( .A(n5938), .Z(n18081) );
  XNOR U19813 ( .A(n5936), .B(n18082), .Z(n5938) );
  XNOR U19814 ( .A(q[5]), .B(DB[1741]), .Z(n18082) );
  XNOR U19815 ( .A(q[4]), .B(DB[1740]), .Z(n5936) );
  IV U19816 ( .A(n5950), .Z(n18080) );
  XOR U19817 ( .A(n18083), .B(n18084), .Z(n5950) );
  XNOR U19818 ( .A(n5946), .B(n5948), .Z(n18084) );
  XNOR U19819 ( .A(q[0]), .B(DB[1736]), .Z(n5948) );
  XNOR U19820 ( .A(q[3]), .B(DB[1739]), .Z(n5946) );
  IV U19821 ( .A(n5945), .Z(n18083) );
  XNOR U19822 ( .A(n5943), .B(n18085), .Z(n5945) );
  XNOR U19823 ( .A(q[2]), .B(DB[1738]), .Z(n18085) );
  XNOR U19824 ( .A(q[1]), .B(DB[1737]), .Z(n5943) );
  XOR U19825 ( .A(n18086), .B(n5908), .Z(n5871) );
  XOR U19826 ( .A(n18087), .B(n5896), .Z(n5908) );
  XNOR U19827 ( .A(q[6]), .B(DB[1749]), .Z(n5896) );
  IV U19828 ( .A(n5895), .Z(n18087) );
  XNOR U19829 ( .A(n5893), .B(n18088), .Z(n5895) );
  XNOR U19830 ( .A(q[5]), .B(DB[1748]), .Z(n18088) );
  XNOR U19831 ( .A(q[4]), .B(DB[1747]), .Z(n5893) );
  IV U19832 ( .A(n5907), .Z(n18086) );
  XOR U19833 ( .A(n18089), .B(n18090), .Z(n5907) );
  XNOR U19834 ( .A(n5903), .B(n5905), .Z(n18090) );
  XNOR U19835 ( .A(q[0]), .B(DB[1743]), .Z(n5905) );
  XNOR U19836 ( .A(q[3]), .B(DB[1746]), .Z(n5903) );
  IV U19837 ( .A(n5902), .Z(n18089) );
  XNOR U19838 ( .A(n5900), .B(n18091), .Z(n5902) );
  XNOR U19839 ( .A(q[2]), .B(DB[1745]), .Z(n18091) );
  XNOR U19840 ( .A(q[1]), .B(DB[1744]), .Z(n5900) );
  XOR U19841 ( .A(n18092), .B(n5865), .Z(n5828) );
  XOR U19842 ( .A(n18093), .B(n5853), .Z(n5865) );
  XNOR U19843 ( .A(q[6]), .B(DB[1756]), .Z(n5853) );
  IV U19844 ( .A(n5852), .Z(n18093) );
  XNOR U19845 ( .A(n5850), .B(n18094), .Z(n5852) );
  XNOR U19846 ( .A(q[5]), .B(DB[1755]), .Z(n18094) );
  XNOR U19847 ( .A(q[4]), .B(DB[1754]), .Z(n5850) );
  IV U19848 ( .A(n5864), .Z(n18092) );
  XOR U19849 ( .A(n18095), .B(n18096), .Z(n5864) );
  XNOR U19850 ( .A(n5860), .B(n5862), .Z(n18096) );
  XNOR U19851 ( .A(q[0]), .B(DB[1750]), .Z(n5862) );
  XNOR U19852 ( .A(q[3]), .B(DB[1753]), .Z(n5860) );
  IV U19853 ( .A(n5859), .Z(n18095) );
  XNOR U19854 ( .A(n5857), .B(n18097), .Z(n5859) );
  XNOR U19855 ( .A(q[2]), .B(DB[1752]), .Z(n18097) );
  XNOR U19856 ( .A(q[1]), .B(DB[1751]), .Z(n5857) );
  XOR U19857 ( .A(n18098), .B(n5822), .Z(n5785) );
  XOR U19858 ( .A(n18099), .B(n5810), .Z(n5822) );
  XNOR U19859 ( .A(q[6]), .B(DB[1763]), .Z(n5810) );
  IV U19860 ( .A(n5809), .Z(n18099) );
  XNOR U19861 ( .A(n5807), .B(n18100), .Z(n5809) );
  XNOR U19862 ( .A(q[5]), .B(DB[1762]), .Z(n18100) );
  XNOR U19863 ( .A(q[4]), .B(DB[1761]), .Z(n5807) );
  IV U19864 ( .A(n5821), .Z(n18098) );
  XOR U19865 ( .A(n18101), .B(n18102), .Z(n5821) );
  XNOR U19866 ( .A(n5817), .B(n5819), .Z(n18102) );
  XNOR U19867 ( .A(q[0]), .B(DB[1757]), .Z(n5819) );
  XNOR U19868 ( .A(q[3]), .B(DB[1760]), .Z(n5817) );
  IV U19869 ( .A(n5816), .Z(n18101) );
  XNOR U19870 ( .A(n5814), .B(n18103), .Z(n5816) );
  XNOR U19871 ( .A(q[2]), .B(DB[1759]), .Z(n18103) );
  XNOR U19872 ( .A(q[1]), .B(DB[1758]), .Z(n5814) );
  XOR U19873 ( .A(n18104), .B(n5779), .Z(n5742) );
  XOR U19874 ( .A(n18105), .B(n5767), .Z(n5779) );
  XNOR U19875 ( .A(q[6]), .B(DB[1770]), .Z(n5767) );
  IV U19876 ( .A(n5766), .Z(n18105) );
  XNOR U19877 ( .A(n5764), .B(n18106), .Z(n5766) );
  XNOR U19878 ( .A(q[5]), .B(DB[1769]), .Z(n18106) );
  XNOR U19879 ( .A(q[4]), .B(DB[1768]), .Z(n5764) );
  IV U19880 ( .A(n5778), .Z(n18104) );
  XOR U19881 ( .A(n18107), .B(n18108), .Z(n5778) );
  XNOR U19882 ( .A(n5774), .B(n5776), .Z(n18108) );
  XNOR U19883 ( .A(q[0]), .B(DB[1764]), .Z(n5776) );
  XNOR U19884 ( .A(q[3]), .B(DB[1767]), .Z(n5774) );
  IV U19885 ( .A(n5773), .Z(n18107) );
  XNOR U19886 ( .A(n5771), .B(n18109), .Z(n5773) );
  XNOR U19887 ( .A(q[2]), .B(DB[1766]), .Z(n18109) );
  XNOR U19888 ( .A(q[1]), .B(DB[1765]), .Z(n5771) );
  XOR U19889 ( .A(n18110), .B(n5736), .Z(n5699) );
  XOR U19890 ( .A(n18111), .B(n5724), .Z(n5736) );
  XNOR U19891 ( .A(q[6]), .B(DB[1777]), .Z(n5724) );
  IV U19892 ( .A(n5723), .Z(n18111) );
  XNOR U19893 ( .A(n5721), .B(n18112), .Z(n5723) );
  XNOR U19894 ( .A(q[5]), .B(DB[1776]), .Z(n18112) );
  XNOR U19895 ( .A(q[4]), .B(DB[1775]), .Z(n5721) );
  IV U19896 ( .A(n5735), .Z(n18110) );
  XOR U19897 ( .A(n18113), .B(n18114), .Z(n5735) );
  XNOR U19898 ( .A(n5731), .B(n5733), .Z(n18114) );
  XNOR U19899 ( .A(q[0]), .B(DB[1771]), .Z(n5733) );
  XNOR U19900 ( .A(q[3]), .B(DB[1774]), .Z(n5731) );
  IV U19901 ( .A(n5730), .Z(n18113) );
  XNOR U19902 ( .A(n5728), .B(n18115), .Z(n5730) );
  XNOR U19903 ( .A(q[2]), .B(DB[1773]), .Z(n18115) );
  XNOR U19904 ( .A(q[1]), .B(DB[1772]), .Z(n5728) );
  XOR U19905 ( .A(n18116), .B(n5693), .Z(n5655) );
  XOR U19906 ( .A(n18117), .B(n5681), .Z(n5693) );
  XNOR U19907 ( .A(q[6]), .B(DB[1784]), .Z(n5681) );
  IV U19908 ( .A(n5680), .Z(n18117) );
  XNOR U19909 ( .A(n5678), .B(n18118), .Z(n5680) );
  XNOR U19910 ( .A(q[5]), .B(DB[1783]), .Z(n18118) );
  XNOR U19911 ( .A(q[4]), .B(DB[1782]), .Z(n5678) );
  IV U19912 ( .A(n5692), .Z(n18116) );
  XOR U19913 ( .A(n18119), .B(n18120), .Z(n5692) );
  XNOR U19914 ( .A(n5688), .B(n5690), .Z(n18120) );
  XNOR U19915 ( .A(q[0]), .B(DB[1778]), .Z(n5690) );
  XNOR U19916 ( .A(q[3]), .B(DB[1781]), .Z(n5688) );
  IV U19917 ( .A(n5687), .Z(n18119) );
  XNOR U19918 ( .A(n5685), .B(n18121), .Z(n5687) );
  XNOR U19919 ( .A(q[2]), .B(DB[1780]), .Z(n18121) );
  XNOR U19920 ( .A(q[1]), .B(DB[1779]), .Z(n5685) );
endmodule

