`define DIR_ROT 0
`define DIR_VEC 1

`define MOD_CIR 1
`define MOD_LIN 0
`define MOD_HYP -1