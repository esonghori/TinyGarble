
module matrixMultSeq ( clk, rst, x, y, o );
  input [287:0] x;
  input [287:0] y;
  output [287:0] o;
  input clk, rst;
  wire   n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906;
  wire   [31:0] sum;
  wire   [1:0] i;
  wire   [1:0] k;
  wire   [1:0] j;

  DFF \i_reg[0]  ( .D(n1011), .CLK(clk), .RST(rst), .Q(i[0]) );
  DFF \sum_reg[0]  ( .D(n1010), .CLK(clk), .RST(rst), .Q(sum[0]) );
  DFF \sum_reg[1]  ( .D(n1009), .CLK(clk), .RST(rst), .Q(sum[1]) );
  DFF \sum_reg[2]  ( .D(n1008), .CLK(clk), .RST(rst), .Q(sum[2]) );
  DFF \sum_reg[3]  ( .D(n1007), .CLK(clk), .RST(rst), .Q(sum[3]) );
  DFF \sum_reg[4]  ( .D(n1006), .CLK(clk), .RST(rst), .Q(sum[4]) );
  DFF \sum_reg[5]  ( .D(n1005), .CLK(clk), .RST(rst), .Q(sum[5]) );
  DFF \sum_reg[6]  ( .D(n1004), .CLK(clk), .RST(rst), .Q(sum[6]) );
  DFF \sum_reg[7]  ( .D(n1003), .CLK(clk), .RST(rst), .Q(sum[7]) );
  DFF \sum_reg[8]  ( .D(n1002), .CLK(clk), .RST(rst), .Q(sum[8]) );
  DFF \sum_reg[9]  ( .D(n1001), .CLK(clk), .RST(rst), .Q(sum[9]) );
  DFF \sum_reg[10]  ( .D(n1000), .CLK(clk), .RST(rst), .Q(sum[10]) );
  DFF \sum_reg[11]  ( .D(n999), .CLK(clk), .RST(rst), .Q(sum[11]) );
  DFF \sum_reg[12]  ( .D(n998), .CLK(clk), .RST(rst), .Q(sum[12]) );
  DFF \sum_reg[13]  ( .D(n997), .CLK(clk), .RST(rst), .Q(sum[13]) );
  DFF \sum_reg[14]  ( .D(n996), .CLK(clk), .RST(rst), .Q(sum[14]) );
  DFF \sum_reg[15]  ( .D(n995), .CLK(clk), .RST(rst), .Q(sum[15]) );
  DFF \sum_reg[16]  ( .D(n994), .CLK(clk), .RST(rst), .Q(sum[16]) );
  DFF \sum_reg[17]  ( .D(n993), .CLK(clk), .RST(rst), .Q(sum[17]) );
  DFF \sum_reg[18]  ( .D(n992), .CLK(clk), .RST(rst), .Q(sum[18]) );
  DFF \sum_reg[19]  ( .D(n991), .CLK(clk), .RST(rst), .Q(sum[19]) );
  DFF \sum_reg[20]  ( .D(n990), .CLK(clk), .RST(rst), .Q(sum[20]) );
  DFF \sum_reg[21]  ( .D(n989), .CLK(clk), .RST(rst), .Q(sum[21]) );
  DFF \sum_reg[22]  ( .D(n988), .CLK(clk), .RST(rst), .Q(sum[22]) );
  DFF \sum_reg[23]  ( .D(n987), .CLK(clk), .RST(rst), .Q(sum[23]) );
  DFF \sum_reg[24]  ( .D(n986), .CLK(clk), .RST(rst), .Q(sum[24]) );
  DFF \sum_reg[25]  ( .D(n985), .CLK(clk), .RST(rst), .Q(sum[25]) );
  DFF \sum_reg[26]  ( .D(n984), .CLK(clk), .RST(rst), .Q(sum[26]) );
  DFF \sum_reg[27]  ( .D(n983), .CLK(clk), .RST(rst), .Q(sum[27]) );
  DFF \sum_reg[28]  ( .D(n982), .CLK(clk), .RST(rst), .Q(sum[28]) );
  DFF \sum_reg[29]  ( .D(n981), .CLK(clk), .RST(rst), .Q(sum[29]) );
  DFF \sum_reg[30]  ( .D(n980), .CLK(clk), .RST(rst), .Q(sum[30]) );
  DFF \sum_reg[31]  ( .D(n979), .CLK(clk), .RST(rst), .Q(sum[31]) );
  DFF \k_reg[1]  ( .D(n978), .CLK(clk), .RST(rst), .Q(k[1]) );
  DFF \k_reg[0]  ( .D(n977), .CLK(clk), .RST(rst), .Q(k[0]) );
  DFF \j_reg[1]  ( .D(n976), .CLK(clk), .RST(rst), .Q(j[1]) );
  DFF \j_reg[0]  ( .D(n975), .CLK(clk), .RST(rst), .Q(j[0]) );
  DFF \i_reg[1]  ( .D(n974), .CLK(clk), .RST(rst), .Q(i[1]) );
  DFF \oij_reg[0][2][0]  ( .D(n973), .CLK(clk), .RST(rst), .Q(o[64]) );
  DFF \oij_reg[0][2][1]  ( .D(n972), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oij_reg[0][2][2]  ( .D(n971), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oij_reg[0][2][3]  ( .D(n970), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oij_reg[0][2][4]  ( .D(n969), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oij_reg[0][2][5]  ( .D(n968), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oij_reg[0][2][6]  ( .D(n967), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oij_reg[0][2][7]  ( .D(n966), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oij_reg[0][2][8]  ( .D(n965), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oij_reg[0][2][9]  ( .D(n964), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oij_reg[0][2][10]  ( .D(n963), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oij_reg[0][2][11]  ( .D(n962), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oij_reg[0][2][12]  ( .D(n961), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oij_reg[0][2][13]  ( .D(n960), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oij_reg[0][2][14]  ( .D(n959), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oij_reg[0][2][15]  ( .D(n958), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oij_reg[0][2][16]  ( .D(n957), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oij_reg[0][2][17]  ( .D(n956), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oij_reg[0][2][18]  ( .D(n955), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oij_reg[0][2][19]  ( .D(n954), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oij_reg[0][2][20]  ( .D(n953), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oij_reg[0][2][21]  ( .D(n952), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oij_reg[0][2][22]  ( .D(n951), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oij_reg[0][2][23]  ( .D(n950), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oij_reg[0][2][24]  ( .D(n949), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oij_reg[0][2][25]  ( .D(n948), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oij_reg[0][2][26]  ( .D(n947), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oij_reg[0][2][27]  ( .D(n946), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oij_reg[0][2][28]  ( .D(n945), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oij_reg[0][2][29]  ( .D(n944), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oij_reg[0][2][30]  ( .D(n943), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oij_reg[0][2][31]  ( .D(n942), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oij_reg[1][2][0]  ( .D(n941), .CLK(clk), .RST(rst), .Q(o[160]) );
  DFF \oij_reg[1][2][1]  ( .D(n940), .CLK(clk), .RST(rst), .Q(o[161]) );
  DFF \oij_reg[1][2][2]  ( .D(n939), .CLK(clk), .RST(rst), .Q(o[162]) );
  DFF \oij_reg[1][2][3]  ( .D(n938), .CLK(clk), .RST(rst), .Q(o[163]) );
  DFF \oij_reg[1][2][4]  ( .D(n937), .CLK(clk), .RST(rst), .Q(o[164]) );
  DFF \oij_reg[1][2][5]  ( .D(n936), .CLK(clk), .RST(rst), .Q(o[165]) );
  DFF \oij_reg[1][2][6]  ( .D(n935), .CLK(clk), .RST(rst), .Q(o[166]) );
  DFF \oij_reg[1][2][7]  ( .D(n934), .CLK(clk), .RST(rst), .Q(o[167]) );
  DFF \oij_reg[1][2][8]  ( .D(n933), .CLK(clk), .RST(rst), .Q(o[168]) );
  DFF \oij_reg[1][2][9]  ( .D(n932), .CLK(clk), .RST(rst), .Q(o[169]) );
  DFF \oij_reg[1][2][10]  ( .D(n931), .CLK(clk), .RST(rst), .Q(o[170]) );
  DFF \oij_reg[1][2][11]  ( .D(n930), .CLK(clk), .RST(rst), .Q(o[171]) );
  DFF \oij_reg[1][2][12]  ( .D(n929), .CLK(clk), .RST(rst), .Q(o[172]) );
  DFF \oij_reg[1][2][13]  ( .D(n928), .CLK(clk), .RST(rst), .Q(o[173]) );
  DFF \oij_reg[1][2][14]  ( .D(n927), .CLK(clk), .RST(rst), .Q(o[174]) );
  DFF \oij_reg[1][2][15]  ( .D(n926), .CLK(clk), .RST(rst), .Q(o[175]) );
  DFF \oij_reg[1][2][16]  ( .D(n925), .CLK(clk), .RST(rst), .Q(o[176]) );
  DFF \oij_reg[1][2][17]  ( .D(n924), .CLK(clk), .RST(rst), .Q(o[177]) );
  DFF \oij_reg[1][2][18]  ( .D(n923), .CLK(clk), .RST(rst), .Q(o[178]) );
  DFF \oij_reg[1][2][19]  ( .D(n922), .CLK(clk), .RST(rst), .Q(o[179]) );
  DFF \oij_reg[1][2][20]  ( .D(n921), .CLK(clk), .RST(rst), .Q(o[180]) );
  DFF \oij_reg[1][2][21]  ( .D(n920), .CLK(clk), .RST(rst), .Q(o[181]) );
  DFF \oij_reg[1][2][22]  ( .D(n919), .CLK(clk), .RST(rst), .Q(o[182]) );
  DFF \oij_reg[1][2][23]  ( .D(n918), .CLK(clk), .RST(rst), .Q(o[183]) );
  DFF \oij_reg[1][2][24]  ( .D(n917), .CLK(clk), .RST(rst), .Q(o[184]) );
  DFF \oij_reg[1][2][25]  ( .D(n916), .CLK(clk), .RST(rst), .Q(o[185]) );
  DFF \oij_reg[1][2][26]  ( .D(n915), .CLK(clk), .RST(rst), .Q(o[186]) );
  DFF \oij_reg[1][2][27]  ( .D(n914), .CLK(clk), .RST(rst), .Q(o[187]) );
  DFF \oij_reg[1][2][28]  ( .D(n913), .CLK(clk), .RST(rst), .Q(o[188]) );
  DFF \oij_reg[1][2][29]  ( .D(n912), .CLK(clk), .RST(rst), .Q(o[189]) );
  DFF \oij_reg[1][2][30]  ( .D(n911), .CLK(clk), .RST(rst), .Q(o[190]) );
  DFF \oij_reg[1][2][31]  ( .D(n910), .CLK(clk), .RST(rst), .Q(o[191]) );
  DFF \oij_reg[2][2][0]  ( .D(n909), .CLK(clk), .RST(rst), .Q(o[256]) );
  DFF \oij_reg[2][2][1]  ( .D(n908), .CLK(clk), .RST(rst), .Q(o[257]) );
  DFF \oij_reg[2][2][2]  ( .D(n907), .CLK(clk), .RST(rst), .Q(o[258]) );
  DFF \oij_reg[2][2][3]  ( .D(n906), .CLK(clk), .RST(rst), .Q(o[259]) );
  DFF \oij_reg[2][2][4]  ( .D(n905), .CLK(clk), .RST(rst), .Q(o[260]) );
  DFF \oij_reg[2][2][5]  ( .D(n904), .CLK(clk), .RST(rst), .Q(o[261]) );
  DFF \oij_reg[2][2][6]  ( .D(n903), .CLK(clk), .RST(rst), .Q(o[262]) );
  DFF \oij_reg[2][2][7]  ( .D(n902), .CLK(clk), .RST(rst), .Q(o[263]) );
  DFF \oij_reg[2][2][8]  ( .D(n901), .CLK(clk), .RST(rst), .Q(o[264]) );
  DFF \oij_reg[2][2][9]  ( .D(n900), .CLK(clk), .RST(rst), .Q(o[265]) );
  DFF \oij_reg[2][2][10]  ( .D(n899), .CLK(clk), .RST(rst), .Q(o[266]) );
  DFF \oij_reg[2][2][11]  ( .D(n898), .CLK(clk), .RST(rst), .Q(o[267]) );
  DFF \oij_reg[2][2][12]  ( .D(n897), .CLK(clk), .RST(rst), .Q(o[268]) );
  DFF \oij_reg[2][2][13]  ( .D(n896), .CLK(clk), .RST(rst), .Q(o[269]) );
  DFF \oij_reg[2][2][14]  ( .D(n895), .CLK(clk), .RST(rst), .Q(o[270]) );
  DFF \oij_reg[2][2][15]  ( .D(n894), .CLK(clk), .RST(rst), .Q(o[271]) );
  DFF \oij_reg[2][2][16]  ( .D(n893), .CLK(clk), .RST(rst), .Q(o[272]) );
  DFF \oij_reg[2][2][17]  ( .D(n892), .CLK(clk), .RST(rst), .Q(o[273]) );
  DFF \oij_reg[2][2][18]  ( .D(n891), .CLK(clk), .RST(rst), .Q(o[274]) );
  DFF \oij_reg[2][2][19]  ( .D(n890), .CLK(clk), .RST(rst), .Q(o[275]) );
  DFF \oij_reg[2][2][20]  ( .D(n889), .CLK(clk), .RST(rst), .Q(o[276]) );
  DFF \oij_reg[2][2][21]  ( .D(n888), .CLK(clk), .RST(rst), .Q(o[277]) );
  DFF \oij_reg[2][2][22]  ( .D(n887), .CLK(clk), .RST(rst), .Q(o[278]) );
  DFF \oij_reg[2][2][23]  ( .D(n886), .CLK(clk), .RST(rst), .Q(o[279]) );
  DFF \oij_reg[2][2][24]  ( .D(n885), .CLK(clk), .RST(rst), .Q(o[280]) );
  DFF \oij_reg[2][2][25]  ( .D(n884), .CLK(clk), .RST(rst), .Q(o[281]) );
  DFF \oij_reg[2][2][26]  ( .D(n883), .CLK(clk), .RST(rst), .Q(o[282]) );
  DFF \oij_reg[2][2][27]  ( .D(n882), .CLK(clk), .RST(rst), .Q(o[283]) );
  DFF \oij_reg[2][2][28]  ( .D(n881), .CLK(clk), .RST(rst), .Q(o[284]) );
  DFF \oij_reg[2][2][29]  ( .D(n880), .CLK(clk), .RST(rst), .Q(o[285]) );
  DFF \oij_reg[2][2][30]  ( .D(n879), .CLK(clk), .RST(rst), .Q(o[286]) );
  DFF \oij_reg[2][2][31]  ( .D(n878), .CLK(clk), .RST(rst), .Q(o[287]) );
  DFF \oij_reg[0][0][0]  ( .D(n877), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oij_reg[0][0][1]  ( .D(n876), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oij_reg[0][0][2]  ( .D(n875), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oij_reg[0][0][3]  ( .D(n874), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oij_reg[0][0][4]  ( .D(n873), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oij_reg[0][0][5]  ( .D(n872), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oij_reg[0][0][6]  ( .D(n871), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oij_reg[0][0][7]  ( .D(n870), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oij_reg[0][0][8]  ( .D(n869), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oij_reg[0][0][9]  ( .D(n868), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oij_reg[0][0][10]  ( .D(n867), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oij_reg[0][0][11]  ( .D(n866), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oij_reg[0][0][12]  ( .D(n865), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oij_reg[0][0][13]  ( .D(n864), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oij_reg[0][0][14]  ( .D(n863), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oij_reg[0][0][15]  ( .D(n862), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oij_reg[0][0][16]  ( .D(n861), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oij_reg[0][0][17]  ( .D(n860), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oij_reg[0][0][18]  ( .D(n859), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oij_reg[0][0][19]  ( .D(n858), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oij_reg[0][0][20]  ( .D(n857), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oij_reg[0][0][21]  ( .D(n856), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oij_reg[0][0][22]  ( .D(n855), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oij_reg[0][0][23]  ( .D(n854), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oij_reg[0][0][24]  ( .D(n853), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oij_reg[0][0][25]  ( .D(n852), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oij_reg[0][0][26]  ( .D(n851), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oij_reg[0][0][27]  ( .D(n850), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oij_reg[0][0][28]  ( .D(n849), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oij_reg[0][0][29]  ( .D(n848), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oij_reg[0][0][30]  ( .D(n847), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oij_reg[0][0][31]  ( .D(n846), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oij_reg[1][0][0]  ( .D(n845), .CLK(clk), .RST(rst), .Q(o[96]) );
  DFF \oij_reg[1][0][1]  ( .D(n844), .CLK(clk), .RST(rst), .Q(o[97]) );
  DFF \oij_reg[1][0][2]  ( .D(n843), .CLK(clk), .RST(rst), .Q(o[98]) );
  DFF \oij_reg[1][0][3]  ( .D(n842), .CLK(clk), .RST(rst), .Q(o[99]) );
  DFF \oij_reg[1][0][4]  ( .D(n841), .CLK(clk), .RST(rst), .Q(o[100]) );
  DFF \oij_reg[1][0][5]  ( .D(n840), .CLK(clk), .RST(rst), .Q(o[101]) );
  DFF \oij_reg[1][0][6]  ( .D(n839), .CLK(clk), .RST(rst), .Q(o[102]) );
  DFF \oij_reg[1][0][7]  ( .D(n838), .CLK(clk), .RST(rst), .Q(o[103]) );
  DFF \oij_reg[1][0][8]  ( .D(n837), .CLK(clk), .RST(rst), .Q(o[104]) );
  DFF \oij_reg[1][0][9]  ( .D(n836), .CLK(clk), .RST(rst), .Q(o[105]) );
  DFF \oij_reg[1][0][10]  ( .D(n835), .CLK(clk), .RST(rst), .Q(o[106]) );
  DFF \oij_reg[1][0][11]  ( .D(n834), .CLK(clk), .RST(rst), .Q(o[107]) );
  DFF \oij_reg[1][0][12]  ( .D(n833), .CLK(clk), .RST(rst), .Q(o[108]) );
  DFF \oij_reg[1][0][13]  ( .D(n832), .CLK(clk), .RST(rst), .Q(o[109]) );
  DFF \oij_reg[1][0][14]  ( .D(n831), .CLK(clk), .RST(rst), .Q(o[110]) );
  DFF \oij_reg[1][0][15]  ( .D(n830), .CLK(clk), .RST(rst), .Q(o[111]) );
  DFF \oij_reg[1][0][16]  ( .D(n829), .CLK(clk), .RST(rst), .Q(o[112]) );
  DFF \oij_reg[1][0][17]  ( .D(n828), .CLK(clk), .RST(rst), .Q(o[113]) );
  DFF \oij_reg[1][0][18]  ( .D(n827), .CLK(clk), .RST(rst), .Q(o[114]) );
  DFF \oij_reg[1][0][19]  ( .D(n826), .CLK(clk), .RST(rst), .Q(o[115]) );
  DFF \oij_reg[1][0][20]  ( .D(n825), .CLK(clk), .RST(rst), .Q(o[116]) );
  DFF \oij_reg[1][0][21]  ( .D(n824), .CLK(clk), .RST(rst), .Q(o[117]) );
  DFF \oij_reg[1][0][22]  ( .D(n823), .CLK(clk), .RST(rst), .Q(o[118]) );
  DFF \oij_reg[1][0][23]  ( .D(n822), .CLK(clk), .RST(rst), .Q(o[119]) );
  DFF \oij_reg[1][0][24]  ( .D(n821), .CLK(clk), .RST(rst), .Q(o[120]) );
  DFF \oij_reg[1][0][25]  ( .D(n820), .CLK(clk), .RST(rst), .Q(o[121]) );
  DFF \oij_reg[1][0][26]  ( .D(n819), .CLK(clk), .RST(rst), .Q(o[122]) );
  DFF \oij_reg[1][0][27]  ( .D(n818), .CLK(clk), .RST(rst), .Q(o[123]) );
  DFF \oij_reg[1][0][28]  ( .D(n817), .CLK(clk), .RST(rst), .Q(o[124]) );
  DFF \oij_reg[1][0][29]  ( .D(n816), .CLK(clk), .RST(rst), .Q(o[125]) );
  DFF \oij_reg[1][0][30]  ( .D(n815), .CLK(clk), .RST(rst), .Q(o[126]) );
  DFF \oij_reg[1][0][31]  ( .D(n814), .CLK(clk), .RST(rst), .Q(o[127]) );
  DFF \oij_reg[2][0][0]  ( .D(n813), .CLK(clk), .RST(rst), .Q(o[192]) );
  DFF \oij_reg[2][0][1]  ( .D(n812), .CLK(clk), .RST(rst), .Q(o[193]) );
  DFF \oij_reg[2][0][2]  ( .D(n811), .CLK(clk), .RST(rst), .Q(o[194]) );
  DFF \oij_reg[2][0][3]  ( .D(n810), .CLK(clk), .RST(rst), .Q(o[195]) );
  DFF \oij_reg[2][0][4]  ( .D(n809), .CLK(clk), .RST(rst), .Q(o[196]) );
  DFF \oij_reg[2][0][5]  ( .D(n808), .CLK(clk), .RST(rst), .Q(o[197]) );
  DFF \oij_reg[2][0][6]  ( .D(n807), .CLK(clk), .RST(rst), .Q(o[198]) );
  DFF \oij_reg[2][0][7]  ( .D(n806), .CLK(clk), .RST(rst), .Q(o[199]) );
  DFF \oij_reg[2][0][8]  ( .D(n805), .CLK(clk), .RST(rst), .Q(o[200]) );
  DFF \oij_reg[2][0][9]  ( .D(n804), .CLK(clk), .RST(rst), .Q(o[201]) );
  DFF \oij_reg[2][0][10]  ( .D(n803), .CLK(clk), .RST(rst), .Q(o[202]) );
  DFF \oij_reg[2][0][11]  ( .D(n802), .CLK(clk), .RST(rst), .Q(o[203]) );
  DFF \oij_reg[2][0][12]  ( .D(n801), .CLK(clk), .RST(rst), .Q(o[204]) );
  DFF \oij_reg[2][0][13]  ( .D(n800), .CLK(clk), .RST(rst), .Q(o[205]) );
  DFF \oij_reg[2][0][14]  ( .D(n799), .CLK(clk), .RST(rst), .Q(o[206]) );
  DFF \oij_reg[2][0][15]  ( .D(n798), .CLK(clk), .RST(rst), .Q(o[207]) );
  DFF \oij_reg[2][0][16]  ( .D(n797), .CLK(clk), .RST(rst), .Q(o[208]) );
  DFF \oij_reg[2][0][17]  ( .D(n796), .CLK(clk), .RST(rst), .Q(o[209]) );
  DFF \oij_reg[2][0][18]  ( .D(n795), .CLK(clk), .RST(rst), .Q(o[210]) );
  DFF \oij_reg[2][0][19]  ( .D(n794), .CLK(clk), .RST(rst), .Q(o[211]) );
  DFF \oij_reg[2][0][20]  ( .D(n793), .CLK(clk), .RST(rst), .Q(o[212]) );
  DFF \oij_reg[2][0][21]  ( .D(n792), .CLK(clk), .RST(rst), .Q(o[213]) );
  DFF \oij_reg[2][0][22]  ( .D(n791), .CLK(clk), .RST(rst), .Q(o[214]) );
  DFF \oij_reg[2][0][23]  ( .D(n790), .CLK(clk), .RST(rst), .Q(o[215]) );
  DFF \oij_reg[2][0][24]  ( .D(n789), .CLK(clk), .RST(rst), .Q(o[216]) );
  DFF \oij_reg[2][0][25]  ( .D(n788), .CLK(clk), .RST(rst), .Q(o[217]) );
  DFF \oij_reg[2][0][26]  ( .D(n787), .CLK(clk), .RST(rst), .Q(o[218]) );
  DFF \oij_reg[2][0][27]  ( .D(n786), .CLK(clk), .RST(rst), .Q(o[219]) );
  DFF \oij_reg[2][0][28]  ( .D(n785), .CLK(clk), .RST(rst), .Q(o[220]) );
  DFF \oij_reg[2][0][29]  ( .D(n784), .CLK(clk), .RST(rst), .Q(o[221]) );
  DFF \oij_reg[2][0][30]  ( .D(n783), .CLK(clk), .RST(rst), .Q(o[222]) );
  DFF \oij_reg[2][0][31]  ( .D(n782), .CLK(clk), .RST(rst), .Q(o[223]) );
  DFF \oij_reg[0][1][0]  ( .D(n781), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oij_reg[0][1][1]  ( .D(n780), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oij_reg[0][1][2]  ( .D(n779), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oij_reg[0][1][3]  ( .D(n778), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oij_reg[0][1][4]  ( .D(n777), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oij_reg[0][1][5]  ( .D(n776), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oij_reg[0][1][6]  ( .D(n775), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oij_reg[0][1][7]  ( .D(n774), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oij_reg[0][1][8]  ( .D(n773), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oij_reg[0][1][9]  ( .D(n772), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oij_reg[0][1][10]  ( .D(n771), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oij_reg[0][1][11]  ( .D(n770), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oij_reg[0][1][12]  ( .D(n769), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oij_reg[0][1][13]  ( .D(n768), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oij_reg[0][1][14]  ( .D(n767), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oij_reg[0][1][15]  ( .D(n766), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oij_reg[0][1][16]  ( .D(n765), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oij_reg[0][1][17]  ( .D(n764), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oij_reg[0][1][18]  ( .D(n763), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oij_reg[0][1][19]  ( .D(n762), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oij_reg[0][1][20]  ( .D(n761), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oij_reg[0][1][21]  ( .D(n760), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oij_reg[0][1][22]  ( .D(n759), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oij_reg[0][1][23]  ( .D(n758), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oij_reg[0][1][24]  ( .D(n757), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oij_reg[0][1][25]  ( .D(n756), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oij_reg[0][1][26]  ( .D(n755), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oij_reg[0][1][27]  ( .D(n754), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oij_reg[0][1][28]  ( .D(n753), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oij_reg[0][1][29]  ( .D(n752), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oij_reg[0][1][30]  ( .D(n751), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oij_reg[0][1][31]  ( .D(n750), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oij_reg[1][1][0]  ( .D(n749), .CLK(clk), .RST(rst), .Q(o[128]) );
  DFF \oij_reg[1][1][1]  ( .D(n748), .CLK(clk), .RST(rst), .Q(o[129]) );
  DFF \oij_reg[1][1][2]  ( .D(n747), .CLK(clk), .RST(rst), .Q(o[130]) );
  DFF \oij_reg[1][1][3]  ( .D(n746), .CLK(clk), .RST(rst), .Q(o[131]) );
  DFF \oij_reg[1][1][4]  ( .D(n745), .CLK(clk), .RST(rst), .Q(o[132]) );
  DFF \oij_reg[1][1][5]  ( .D(n744), .CLK(clk), .RST(rst), .Q(o[133]) );
  DFF \oij_reg[1][1][6]  ( .D(n743), .CLK(clk), .RST(rst), .Q(o[134]) );
  DFF \oij_reg[1][1][7]  ( .D(n742), .CLK(clk), .RST(rst), .Q(o[135]) );
  DFF \oij_reg[1][1][8]  ( .D(n741), .CLK(clk), .RST(rst), .Q(o[136]) );
  DFF \oij_reg[1][1][9]  ( .D(n740), .CLK(clk), .RST(rst), .Q(o[137]) );
  DFF \oij_reg[1][1][10]  ( .D(n739), .CLK(clk), .RST(rst), .Q(o[138]) );
  DFF \oij_reg[1][1][11]  ( .D(n738), .CLK(clk), .RST(rst), .Q(o[139]) );
  DFF \oij_reg[1][1][12]  ( .D(n737), .CLK(clk), .RST(rst), .Q(o[140]) );
  DFF \oij_reg[1][1][13]  ( .D(n736), .CLK(clk), .RST(rst), .Q(o[141]) );
  DFF \oij_reg[1][1][14]  ( .D(n735), .CLK(clk), .RST(rst), .Q(o[142]) );
  DFF \oij_reg[1][1][15]  ( .D(n734), .CLK(clk), .RST(rst), .Q(o[143]) );
  DFF \oij_reg[1][1][16]  ( .D(n733), .CLK(clk), .RST(rst), .Q(o[144]) );
  DFF \oij_reg[1][1][17]  ( .D(n732), .CLK(clk), .RST(rst), .Q(o[145]) );
  DFF \oij_reg[1][1][18]  ( .D(n731), .CLK(clk), .RST(rst), .Q(o[146]) );
  DFF \oij_reg[1][1][19]  ( .D(n730), .CLK(clk), .RST(rst), .Q(o[147]) );
  DFF \oij_reg[1][1][20]  ( .D(n729), .CLK(clk), .RST(rst), .Q(o[148]) );
  DFF \oij_reg[1][1][21]  ( .D(n728), .CLK(clk), .RST(rst), .Q(o[149]) );
  DFF \oij_reg[1][1][22]  ( .D(n727), .CLK(clk), .RST(rst), .Q(o[150]) );
  DFF \oij_reg[1][1][23]  ( .D(n726), .CLK(clk), .RST(rst), .Q(o[151]) );
  DFF \oij_reg[1][1][24]  ( .D(n725), .CLK(clk), .RST(rst), .Q(o[152]) );
  DFF \oij_reg[1][1][25]  ( .D(n724), .CLK(clk), .RST(rst), .Q(o[153]) );
  DFF \oij_reg[1][1][26]  ( .D(n723), .CLK(clk), .RST(rst), .Q(o[154]) );
  DFF \oij_reg[1][1][27]  ( .D(n722), .CLK(clk), .RST(rst), .Q(o[155]) );
  DFF \oij_reg[1][1][28]  ( .D(n721), .CLK(clk), .RST(rst), .Q(o[156]) );
  DFF \oij_reg[1][1][29]  ( .D(n720), .CLK(clk), .RST(rst), .Q(o[157]) );
  DFF \oij_reg[1][1][30]  ( .D(n719), .CLK(clk), .RST(rst), .Q(o[158]) );
  DFF \oij_reg[1][1][31]  ( .D(n718), .CLK(clk), .RST(rst), .Q(o[159]) );
  DFF \oij_reg[2][1][0]  ( .D(n717), .CLK(clk), .RST(rst), .Q(o[224]) );
  DFF \oij_reg[2][1][1]  ( .D(n716), .CLK(clk), .RST(rst), .Q(o[225]) );
  DFF \oij_reg[2][1][2]  ( .D(n715), .CLK(clk), .RST(rst), .Q(o[226]) );
  DFF \oij_reg[2][1][3]  ( .D(n714), .CLK(clk), .RST(rst), .Q(o[227]) );
  DFF \oij_reg[2][1][4]  ( .D(n713), .CLK(clk), .RST(rst), .Q(o[228]) );
  DFF \oij_reg[2][1][5]  ( .D(n712), .CLK(clk), .RST(rst), .Q(o[229]) );
  DFF \oij_reg[2][1][6]  ( .D(n711), .CLK(clk), .RST(rst), .Q(o[230]) );
  DFF \oij_reg[2][1][7]  ( .D(n710), .CLK(clk), .RST(rst), .Q(o[231]) );
  DFF \oij_reg[2][1][8]  ( .D(n709), .CLK(clk), .RST(rst), .Q(o[232]) );
  DFF \oij_reg[2][1][9]  ( .D(n708), .CLK(clk), .RST(rst), .Q(o[233]) );
  DFF \oij_reg[2][1][10]  ( .D(n707), .CLK(clk), .RST(rst), .Q(o[234]) );
  DFF \oij_reg[2][1][11]  ( .D(n706), .CLK(clk), .RST(rst), .Q(o[235]) );
  DFF \oij_reg[2][1][12]  ( .D(n705), .CLK(clk), .RST(rst), .Q(o[236]) );
  DFF \oij_reg[2][1][13]  ( .D(n704), .CLK(clk), .RST(rst), .Q(o[237]) );
  DFF \oij_reg[2][1][14]  ( .D(n703), .CLK(clk), .RST(rst), .Q(o[238]) );
  DFF \oij_reg[2][1][15]  ( .D(n702), .CLK(clk), .RST(rst), .Q(o[239]) );
  DFF \oij_reg[2][1][16]  ( .D(n701), .CLK(clk), .RST(rst), .Q(o[240]) );
  DFF \oij_reg[2][1][17]  ( .D(n700), .CLK(clk), .RST(rst), .Q(o[241]) );
  DFF \oij_reg[2][1][18]  ( .D(n699), .CLK(clk), .RST(rst), .Q(o[242]) );
  DFF \oij_reg[2][1][19]  ( .D(n698), .CLK(clk), .RST(rst), .Q(o[243]) );
  DFF \oij_reg[2][1][20]  ( .D(n697), .CLK(clk), .RST(rst), .Q(o[244]) );
  DFF \oij_reg[2][1][21]  ( .D(n696), .CLK(clk), .RST(rst), .Q(o[245]) );
  DFF \oij_reg[2][1][22]  ( .D(n695), .CLK(clk), .RST(rst), .Q(o[246]) );
  DFF \oij_reg[2][1][23]  ( .D(n694), .CLK(clk), .RST(rst), .Q(o[247]) );
  DFF \oij_reg[2][1][24]  ( .D(n693), .CLK(clk), .RST(rst), .Q(o[248]) );
  DFF \oij_reg[2][1][25]  ( .D(n692), .CLK(clk), .RST(rst), .Q(o[249]) );
  DFF \oij_reg[2][1][26]  ( .D(n691), .CLK(clk), .RST(rst), .Q(o[250]) );
  DFF \oij_reg[2][1][27]  ( .D(n690), .CLK(clk), .RST(rst), .Q(o[251]) );
  DFF \oij_reg[2][1][28]  ( .D(n689), .CLK(clk), .RST(rst), .Q(o[252]) );
  DFF \oij_reg[2][1][29]  ( .D(n688), .CLK(clk), .RST(rst), .Q(o[253]) );
  DFF \oij_reg[2][1][30]  ( .D(n687), .CLK(clk), .RST(rst), .Q(o[254]) );
  DFF \oij_reg[2][1][31]  ( .D(n686), .CLK(clk), .RST(rst), .Q(o[255]) );
  IV U3241 ( .A(n3838), .Z(n3235) );
  IV U3242 ( .A(n3841), .Z(n3236) );
  IV U3243 ( .A(n9904), .Z(n3237) );
  IV U3244 ( .A(i[1]), .Z(n3872) );
  IV U3245 ( .A(j[0]), .Z(n3917) );
  IV U3246 ( .A(i[0]), .Z(n3875) );
  NOR U3247 ( .A(n3875), .B(n3872), .Z(n9904) );
  IV U3248 ( .A(k[1]), .Z(n3906) );
  NOR U3249 ( .A(n9904), .B(n3906), .Z(n3852) );
  IV U3250 ( .A(n3852), .Z(n3238) );
  NOR U3251 ( .A(k[0]), .B(n3238), .Z(n3846) );
  IV U3252 ( .A(n3846), .Z(n3845) );
  NOR U3253 ( .A(j[1]), .B(n3845), .Z(n3239) );
  IV U3254 ( .A(n3239), .Z(n3240) );
  NOR U3255 ( .A(n3917), .B(n3240), .Z(n3241) );
  IV U3256 ( .A(n3241), .Z(n3375) );
  NOR U3257 ( .A(n3872), .B(n3375), .Z(n3305) );
  IV U3258 ( .A(n3305), .Z(n3304) );
  NOR U3259 ( .A(sum[31]), .B(n3304), .Z(n3243) );
  NOR U3260 ( .A(n3305), .B(o[255]), .Z(n3242) );
  NOR U3261 ( .A(n3243), .B(n3242), .Z(n686) );
  NOR U3262 ( .A(sum[30]), .B(n3304), .Z(n3245) );
  NOR U3263 ( .A(n3305), .B(o[254]), .Z(n3244) );
  NOR U3264 ( .A(n3245), .B(n3244), .Z(n687) );
  NOR U3265 ( .A(sum[29]), .B(n3304), .Z(n3247) );
  NOR U3266 ( .A(n3305), .B(o[253]), .Z(n3246) );
  NOR U3267 ( .A(n3247), .B(n3246), .Z(n688) );
  NOR U3268 ( .A(sum[28]), .B(n3304), .Z(n3249) );
  NOR U3269 ( .A(n3305), .B(o[252]), .Z(n3248) );
  NOR U3270 ( .A(n3249), .B(n3248), .Z(n689) );
  NOR U3271 ( .A(sum[27]), .B(n3304), .Z(n3251) );
  NOR U3272 ( .A(n3305), .B(o[251]), .Z(n3250) );
  NOR U3273 ( .A(n3251), .B(n3250), .Z(n690) );
  NOR U3274 ( .A(sum[26]), .B(n3304), .Z(n3253) );
  NOR U3275 ( .A(n3305), .B(o[250]), .Z(n3252) );
  NOR U3276 ( .A(n3253), .B(n3252), .Z(n691) );
  NOR U3277 ( .A(sum[25]), .B(n3304), .Z(n3255) );
  NOR U3278 ( .A(n3305), .B(o[249]), .Z(n3254) );
  NOR U3279 ( .A(n3255), .B(n3254), .Z(n692) );
  NOR U3280 ( .A(sum[24]), .B(n3304), .Z(n3257) );
  NOR U3281 ( .A(n3305), .B(o[248]), .Z(n3256) );
  NOR U3282 ( .A(n3257), .B(n3256), .Z(n693) );
  NOR U3283 ( .A(sum[23]), .B(n3304), .Z(n3259) );
  NOR U3284 ( .A(n3305), .B(o[247]), .Z(n3258) );
  NOR U3285 ( .A(n3259), .B(n3258), .Z(n694) );
  NOR U3286 ( .A(sum[22]), .B(n3304), .Z(n3261) );
  NOR U3287 ( .A(n3305), .B(o[246]), .Z(n3260) );
  NOR U3288 ( .A(n3261), .B(n3260), .Z(n695) );
  NOR U3289 ( .A(sum[21]), .B(n3304), .Z(n3263) );
  NOR U3290 ( .A(n3305), .B(o[245]), .Z(n3262) );
  NOR U3291 ( .A(n3263), .B(n3262), .Z(n696) );
  NOR U3292 ( .A(sum[20]), .B(n3304), .Z(n3265) );
  NOR U3293 ( .A(n3305), .B(o[244]), .Z(n3264) );
  NOR U3294 ( .A(n3265), .B(n3264), .Z(n697) );
  NOR U3295 ( .A(sum[19]), .B(n3304), .Z(n3267) );
  NOR U3296 ( .A(n3305), .B(o[243]), .Z(n3266) );
  NOR U3297 ( .A(n3267), .B(n3266), .Z(n698) );
  NOR U3298 ( .A(sum[18]), .B(n3304), .Z(n3269) );
  NOR U3299 ( .A(n3305), .B(o[242]), .Z(n3268) );
  NOR U3300 ( .A(n3269), .B(n3268), .Z(n699) );
  NOR U3301 ( .A(sum[17]), .B(n3304), .Z(n3271) );
  NOR U3302 ( .A(n3305), .B(o[241]), .Z(n3270) );
  NOR U3303 ( .A(n3271), .B(n3270), .Z(n700) );
  NOR U3304 ( .A(sum[16]), .B(n3304), .Z(n3273) );
  NOR U3305 ( .A(n3305), .B(o[240]), .Z(n3272) );
  NOR U3306 ( .A(n3273), .B(n3272), .Z(n701) );
  NOR U3307 ( .A(sum[15]), .B(n3304), .Z(n3275) );
  NOR U3308 ( .A(n3305), .B(o[239]), .Z(n3274) );
  NOR U3309 ( .A(n3275), .B(n3274), .Z(n702) );
  NOR U3310 ( .A(sum[14]), .B(n3304), .Z(n3277) );
  NOR U3311 ( .A(n3305), .B(o[238]), .Z(n3276) );
  NOR U3312 ( .A(n3277), .B(n3276), .Z(n703) );
  NOR U3313 ( .A(sum[13]), .B(n3304), .Z(n3279) );
  NOR U3314 ( .A(n3305), .B(o[237]), .Z(n3278) );
  NOR U3315 ( .A(n3279), .B(n3278), .Z(n704) );
  NOR U3316 ( .A(sum[12]), .B(n3304), .Z(n3281) );
  NOR U3317 ( .A(n3305), .B(o[236]), .Z(n3280) );
  NOR U3318 ( .A(n3281), .B(n3280), .Z(n705) );
  NOR U3319 ( .A(sum[11]), .B(n3304), .Z(n3283) );
  NOR U3320 ( .A(n3305), .B(o[235]), .Z(n3282) );
  NOR U3321 ( .A(n3283), .B(n3282), .Z(n706) );
  NOR U3322 ( .A(sum[10]), .B(n3304), .Z(n3285) );
  NOR U3323 ( .A(n3305), .B(o[234]), .Z(n3284) );
  NOR U3324 ( .A(n3285), .B(n3284), .Z(n707) );
  NOR U3325 ( .A(sum[9]), .B(n3304), .Z(n3287) );
  NOR U3326 ( .A(n3305), .B(o[233]), .Z(n3286) );
  NOR U3327 ( .A(n3287), .B(n3286), .Z(n708) );
  NOR U3328 ( .A(sum[8]), .B(n3304), .Z(n3289) );
  NOR U3329 ( .A(n3305), .B(o[232]), .Z(n3288) );
  NOR U3330 ( .A(n3289), .B(n3288), .Z(n709) );
  NOR U3331 ( .A(sum[7]), .B(n3304), .Z(n3291) );
  NOR U3332 ( .A(n3305), .B(o[231]), .Z(n3290) );
  NOR U3333 ( .A(n3291), .B(n3290), .Z(n710) );
  NOR U3334 ( .A(sum[6]), .B(n3304), .Z(n3293) );
  NOR U3335 ( .A(n3305), .B(o[230]), .Z(n3292) );
  NOR U3336 ( .A(n3293), .B(n3292), .Z(n711) );
  NOR U3337 ( .A(sum[5]), .B(n3304), .Z(n3295) );
  NOR U3338 ( .A(n3305), .B(o[229]), .Z(n3294) );
  NOR U3339 ( .A(n3295), .B(n3294), .Z(n712) );
  NOR U3340 ( .A(sum[4]), .B(n3304), .Z(n3297) );
  NOR U3341 ( .A(n3305), .B(o[228]), .Z(n3296) );
  NOR U3342 ( .A(n3297), .B(n3296), .Z(n713) );
  NOR U3343 ( .A(sum[3]), .B(n3304), .Z(n3299) );
  NOR U3344 ( .A(n3305), .B(o[227]), .Z(n3298) );
  NOR U3345 ( .A(n3299), .B(n3298), .Z(n714) );
  NOR U3346 ( .A(sum[2]), .B(n3304), .Z(n3301) );
  NOR U3347 ( .A(n3305), .B(o[226]), .Z(n3300) );
  NOR U3348 ( .A(n3301), .B(n3300), .Z(n715) );
  NOR U3349 ( .A(sum[1]), .B(n3304), .Z(n3303) );
  NOR U3350 ( .A(n3305), .B(o[225]), .Z(n3302) );
  NOR U3351 ( .A(n3303), .B(n3302), .Z(n716) );
  NOR U3352 ( .A(sum[0]), .B(n3304), .Z(n3307) );
  NOR U3353 ( .A(n3305), .B(o[224]), .Z(n3306) );
  NOR U3354 ( .A(n3307), .B(n3306), .Z(n717) );
  NOR U3355 ( .A(n3875), .B(n3375), .Z(n3371) );
  IV U3356 ( .A(n3371), .Z(n3370) );
  NOR U3357 ( .A(sum[31]), .B(n3370), .Z(n3309) );
  NOR U3358 ( .A(n3371), .B(o[159]), .Z(n3308) );
  NOR U3359 ( .A(n3309), .B(n3308), .Z(n718) );
  NOR U3360 ( .A(sum[30]), .B(n3370), .Z(n3311) );
  NOR U3361 ( .A(n3371), .B(o[158]), .Z(n3310) );
  NOR U3362 ( .A(n3311), .B(n3310), .Z(n719) );
  NOR U3363 ( .A(sum[29]), .B(n3370), .Z(n3313) );
  NOR U3364 ( .A(n3371), .B(o[157]), .Z(n3312) );
  NOR U3365 ( .A(n3313), .B(n3312), .Z(n720) );
  NOR U3366 ( .A(sum[28]), .B(n3370), .Z(n3315) );
  NOR U3367 ( .A(n3371), .B(o[156]), .Z(n3314) );
  NOR U3368 ( .A(n3315), .B(n3314), .Z(n721) );
  NOR U3369 ( .A(sum[27]), .B(n3370), .Z(n3317) );
  NOR U3370 ( .A(n3371), .B(o[155]), .Z(n3316) );
  NOR U3371 ( .A(n3317), .B(n3316), .Z(n722) );
  NOR U3372 ( .A(sum[26]), .B(n3370), .Z(n3319) );
  NOR U3373 ( .A(n3371), .B(o[154]), .Z(n3318) );
  NOR U3374 ( .A(n3319), .B(n3318), .Z(n723) );
  NOR U3375 ( .A(sum[25]), .B(n3370), .Z(n3321) );
  NOR U3376 ( .A(n3371), .B(o[153]), .Z(n3320) );
  NOR U3377 ( .A(n3321), .B(n3320), .Z(n724) );
  NOR U3378 ( .A(sum[24]), .B(n3370), .Z(n3323) );
  NOR U3379 ( .A(n3371), .B(o[152]), .Z(n3322) );
  NOR U3380 ( .A(n3323), .B(n3322), .Z(n725) );
  NOR U3381 ( .A(sum[23]), .B(n3370), .Z(n3325) );
  NOR U3382 ( .A(n3371), .B(o[151]), .Z(n3324) );
  NOR U3383 ( .A(n3325), .B(n3324), .Z(n726) );
  NOR U3384 ( .A(sum[22]), .B(n3370), .Z(n3327) );
  NOR U3385 ( .A(n3371), .B(o[150]), .Z(n3326) );
  NOR U3386 ( .A(n3327), .B(n3326), .Z(n727) );
  NOR U3387 ( .A(sum[21]), .B(n3370), .Z(n3329) );
  NOR U3388 ( .A(n3371), .B(o[149]), .Z(n3328) );
  NOR U3389 ( .A(n3329), .B(n3328), .Z(n728) );
  NOR U3390 ( .A(sum[20]), .B(n3370), .Z(n3331) );
  NOR U3391 ( .A(n3371), .B(o[148]), .Z(n3330) );
  NOR U3392 ( .A(n3331), .B(n3330), .Z(n729) );
  NOR U3393 ( .A(sum[19]), .B(n3370), .Z(n3333) );
  NOR U3394 ( .A(n3371), .B(o[147]), .Z(n3332) );
  NOR U3395 ( .A(n3333), .B(n3332), .Z(n730) );
  NOR U3396 ( .A(sum[18]), .B(n3370), .Z(n3335) );
  NOR U3397 ( .A(n3371), .B(o[146]), .Z(n3334) );
  NOR U3398 ( .A(n3335), .B(n3334), .Z(n731) );
  NOR U3399 ( .A(sum[17]), .B(n3370), .Z(n3337) );
  NOR U3400 ( .A(n3371), .B(o[145]), .Z(n3336) );
  NOR U3401 ( .A(n3337), .B(n3336), .Z(n732) );
  NOR U3402 ( .A(sum[16]), .B(n3370), .Z(n3339) );
  NOR U3403 ( .A(n3371), .B(o[144]), .Z(n3338) );
  NOR U3404 ( .A(n3339), .B(n3338), .Z(n733) );
  NOR U3405 ( .A(sum[15]), .B(n3370), .Z(n3341) );
  NOR U3406 ( .A(n3371), .B(o[143]), .Z(n3340) );
  NOR U3407 ( .A(n3341), .B(n3340), .Z(n734) );
  NOR U3408 ( .A(sum[14]), .B(n3370), .Z(n3343) );
  NOR U3409 ( .A(n3371), .B(o[142]), .Z(n3342) );
  NOR U3410 ( .A(n3343), .B(n3342), .Z(n735) );
  NOR U3411 ( .A(sum[13]), .B(n3370), .Z(n3345) );
  NOR U3412 ( .A(n3371), .B(o[141]), .Z(n3344) );
  NOR U3413 ( .A(n3345), .B(n3344), .Z(n736) );
  NOR U3414 ( .A(sum[12]), .B(n3370), .Z(n3347) );
  NOR U3415 ( .A(n3371), .B(o[140]), .Z(n3346) );
  NOR U3416 ( .A(n3347), .B(n3346), .Z(n737) );
  NOR U3417 ( .A(sum[11]), .B(n3370), .Z(n3349) );
  NOR U3418 ( .A(n3371), .B(o[139]), .Z(n3348) );
  NOR U3419 ( .A(n3349), .B(n3348), .Z(n738) );
  NOR U3420 ( .A(sum[10]), .B(n3370), .Z(n3351) );
  NOR U3421 ( .A(n3371), .B(o[138]), .Z(n3350) );
  NOR U3422 ( .A(n3351), .B(n3350), .Z(n739) );
  NOR U3423 ( .A(sum[9]), .B(n3370), .Z(n3353) );
  NOR U3424 ( .A(n3371), .B(o[137]), .Z(n3352) );
  NOR U3425 ( .A(n3353), .B(n3352), .Z(n740) );
  NOR U3426 ( .A(sum[8]), .B(n3370), .Z(n3355) );
  NOR U3427 ( .A(n3371), .B(o[136]), .Z(n3354) );
  NOR U3428 ( .A(n3355), .B(n3354), .Z(n741) );
  NOR U3429 ( .A(sum[7]), .B(n3370), .Z(n3357) );
  NOR U3430 ( .A(n3371), .B(o[135]), .Z(n3356) );
  NOR U3431 ( .A(n3357), .B(n3356), .Z(n742) );
  NOR U3432 ( .A(sum[6]), .B(n3370), .Z(n3359) );
  NOR U3433 ( .A(n3371), .B(o[134]), .Z(n3358) );
  NOR U3434 ( .A(n3359), .B(n3358), .Z(n743) );
  NOR U3435 ( .A(sum[5]), .B(n3370), .Z(n3361) );
  NOR U3436 ( .A(n3371), .B(o[133]), .Z(n3360) );
  NOR U3437 ( .A(n3361), .B(n3360), .Z(n744) );
  NOR U3438 ( .A(sum[4]), .B(n3370), .Z(n3363) );
  NOR U3439 ( .A(n3371), .B(o[132]), .Z(n3362) );
  NOR U3440 ( .A(n3363), .B(n3362), .Z(n745) );
  NOR U3441 ( .A(sum[3]), .B(n3370), .Z(n3365) );
  NOR U3442 ( .A(n3371), .B(o[131]), .Z(n3364) );
  NOR U3443 ( .A(n3365), .B(n3364), .Z(n746) );
  NOR U3444 ( .A(sum[2]), .B(n3370), .Z(n3367) );
  NOR U3445 ( .A(n3371), .B(o[130]), .Z(n3366) );
  NOR U3446 ( .A(n3367), .B(n3366), .Z(n747) );
  NOR U3447 ( .A(sum[1]), .B(n3370), .Z(n3369) );
  NOR U3448 ( .A(n3371), .B(o[129]), .Z(n3368) );
  NOR U3449 ( .A(n3369), .B(n3368), .Z(n748) );
  NOR U3450 ( .A(sum[0]), .B(n3370), .Z(n3373) );
  NOR U3451 ( .A(n3371), .B(o[128]), .Z(n3372) );
  NOR U3452 ( .A(n3373), .B(n3372), .Z(n749) );
  NOR U3453 ( .A(i[0]), .B(i[1]), .Z(n3374) );
  IV U3454 ( .A(n3374), .Z(n3866) );
  NOR U3455 ( .A(n3866), .B(n3375), .Z(n3439) );
  IV U3456 ( .A(n3439), .Z(n3438) );
  NOR U3457 ( .A(sum[31]), .B(n3438), .Z(n3377) );
  NOR U3458 ( .A(n3439), .B(o[63]), .Z(n3376) );
  NOR U3459 ( .A(n3377), .B(n3376), .Z(n750) );
  NOR U3460 ( .A(sum[30]), .B(n3438), .Z(n3379) );
  NOR U3461 ( .A(n3439), .B(o[62]), .Z(n3378) );
  NOR U3462 ( .A(n3379), .B(n3378), .Z(n751) );
  NOR U3463 ( .A(sum[29]), .B(n3438), .Z(n3381) );
  NOR U3464 ( .A(n3439), .B(o[61]), .Z(n3380) );
  NOR U3465 ( .A(n3381), .B(n3380), .Z(n752) );
  NOR U3466 ( .A(sum[28]), .B(n3438), .Z(n3383) );
  NOR U3467 ( .A(n3439), .B(o[60]), .Z(n3382) );
  NOR U3468 ( .A(n3383), .B(n3382), .Z(n753) );
  NOR U3469 ( .A(sum[27]), .B(n3438), .Z(n3385) );
  NOR U3470 ( .A(n3439), .B(o[59]), .Z(n3384) );
  NOR U3471 ( .A(n3385), .B(n3384), .Z(n754) );
  NOR U3472 ( .A(sum[26]), .B(n3438), .Z(n3387) );
  NOR U3473 ( .A(n3439), .B(o[58]), .Z(n3386) );
  NOR U3474 ( .A(n3387), .B(n3386), .Z(n755) );
  NOR U3475 ( .A(sum[25]), .B(n3438), .Z(n3389) );
  NOR U3476 ( .A(n3439), .B(o[57]), .Z(n3388) );
  NOR U3477 ( .A(n3389), .B(n3388), .Z(n756) );
  NOR U3478 ( .A(sum[24]), .B(n3438), .Z(n3391) );
  NOR U3479 ( .A(n3439), .B(o[56]), .Z(n3390) );
  NOR U3480 ( .A(n3391), .B(n3390), .Z(n757) );
  NOR U3481 ( .A(sum[23]), .B(n3438), .Z(n3393) );
  NOR U3482 ( .A(n3439), .B(o[55]), .Z(n3392) );
  NOR U3483 ( .A(n3393), .B(n3392), .Z(n758) );
  NOR U3484 ( .A(sum[22]), .B(n3438), .Z(n3395) );
  NOR U3485 ( .A(n3439), .B(o[54]), .Z(n3394) );
  NOR U3486 ( .A(n3395), .B(n3394), .Z(n759) );
  NOR U3487 ( .A(sum[21]), .B(n3438), .Z(n3397) );
  NOR U3488 ( .A(n3439), .B(o[53]), .Z(n3396) );
  NOR U3489 ( .A(n3397), .B(n3396), .Z(n760) );
  NOR U3490 ( .A(sum[20]), .B(n3438), .Z(n3399) );
  NOR U3491 ( .A(n3439), .B(o[52]), .Z(n3398) );
  NOR U3492 ( .A(n3399), .B(n3398), .Z(n761) );
  NOR U3493 ( .A(sum[19]), .B(n3438), .Z(n3401) );
  NOR U3494 ( .A(n3439), .B(o[51]), .Z(n3400) );
  NOR U3495 ( .A(n3401), .B(n3400), .Z(n762) );
  NOR U3496 ( .A(sum[18]), .B(n3438), .Z(n3403) );
  NOR U3497 ( .A(n3439), .B(o[50]), .Z(n3402) );
  NOR U3498 ( .A(n3403), .B(n3402), .Z(n763) );
  NOR U3499 ( .A(sum[17]), .B(n3438), .Z(n3405) );
  NOR U3500 ( .A(n3439), .B(o[49]), .Z(n3404) );
  NOR U3501 ( .A(n3405), .B(n3404), .Z(n764) );
  NOR U3502 ( .A(sum[16]), .B(n3438), .Z(n3407) );
  NOR U3503 ( .A(n3439), .B(o[48]), .Z(n3406) );
  NOR U3504 ( .A(n3407), .B(n3406), .Z(n765) );
  NOR U3505 ( .A(sum[15]), .B(n3438), .Z(n3409) );
  NOR U3506 ( .A(n3439), .B(o[47]), .Z(n3408) );
  NOR U3507 ( .A(n3409), .B(n3408), .Z(n766) );
  NOR U3508 ( .A(sum[14]), .B(n3438), .Z(n3411) );
  NOR U3509 ( .A(n3439), .B(o[46]), .Z(n3410) );
  NOR U3510 ( .A(n3411), .B(n3410), .Z(n767) );
  NOR U3511 ( .A(sum[13]), .B(n3438), .Z(n3413) );
  NOR U3512 ( .A(n3439), .B(o[45]), .Z(n3412) );
  NOR U3513 ( .A(n3413), .B(n3412), .Z(n768) );
  NOR U3514 ( .A(sum[12]), .B(n3438), .Z(n3415) );
  NOR U3515 ( .A(n3439), .B(o[44]), .Z(n3414) );
  NOR U3516 ( .A(n3415), .B(n3414), .Z(n769) );
  NOR U3517 ( .A(sum[11]), .B(n3438), .Z(n3417) );
  NOR U3518 ( .A(n3439), .B(o[43]), .Z(n3416) );
  NOR U3519 ( .A(n3417), .B(n3416), .Z(n770) );
  NOR U3520 ( .A(sum[10]), .B(n3438), .Z(n3419) );
  NOR U3521 ( .A(n3439), .B(o[42]), .Z(n3418) );
  NOR U3522 ( .A(n3419), .B(n3418), .Z(n771) );
  NOR U3523 ( .A(sum[9]), .B(n3438), .Z(n3421) );
  NOR U3524 ( .A(n3439), .B(o[41]), .Z(n3420) );
  NOR U3525 ( .A(n3421), .B(n3420), .Z(n772) );
  NOR U3526 ( .A(sum[8]), .B(n3438), .Z(n3423) );
  NOR U3527 ( .A(n3439), .B(o[40]), .Z(n3422) );
  NOR U3528 ( .A(n3423), .B(n3422), .Z(n773) );
  NOR U3529 ( .A(sum[7]), .B(n3438), .Z(n3425) );
  NOR U3530 ( .A(n3439), .B(o[39]), .Z(n3424) );
  NOR U3531 ( .A(n3425), .B(n3424), .Z(n774) );
  NOR U3532 ( .A(sum[6]), .B(n3438), .Z(n3427) );
  NOR U3533 ( .A(n3439), .B(o[38]), .Z(n3426) );
  NOR U3534 ( .A(n3427), .B(n3426), .Z(n775) );
  NOR U3535 ( .A(sum[5]), .B(n3438), .Z(n3429) );
  NOR U3536 ( .A(n3439), .B(o[37]), .Z(n3428) );
  NOR U3537 ( .A(n3429), .B(n3428), .Z(n776) );
  NOR U3538 ( .A(sum[4]), .B(n3438), .Z(n3431) );
  NOR U3539 ( .A(n3439), .B(o[36]), .Z(n3430) );
  NOR U3540 ( .A(n3431), .B(n3430), .Z(n777) );
  NOR U3541 ( .A(sum[3]), .B(n3438), .Z(n3433) );
  NOR U3542 ( .A(n3439), .B(o[35]), .Z(n3432) );
  NOR U3543 ( .A(n3433), .B(n3432), .Z(n778) );
  NOR U3544 ( .A(sum[2]), .B(n3438), .Z(n3435) );
  NOR U3545 ( .A(n3439), .B(o[34]), .Z(n3434) );
  NOR U3546 ( .A(n3435), .B(n3434), .Z(n779) );
  NOR U3547 ( .A(sum[1]), .B(n3438), .Z(n3437) );
  NOR U3548 ( .A(n3439), .B(o[33]), .Z(n3436) );
  NOR U3549 ( .A(n3437), .B(n3436), .Z(n780) );
  NOR U3550 ( .A(sum[0]), .B(n3438), .Z(n3441) );
  NOR U3551 ( .A(n3439), .B(o[32]), .Z(n3440) );
  NOR U3552 ( .A(n3441), .B(n3440), .Z(n781) );
  NOR U3553 ( .A(j[0]), .B(j[1]), .Z(n3442) );
  IV U3554 ( .A(n3442), .Z(n3911) );
  NOR U3555 ( .A(n3911), .B(n3845), .Z(n3443) );
  IV U3556 ( .A(n3443), .Z(n3576) );
  NOR U3557 ( .A(n3872), .B(n3576), .Z(n3507) );
  IV U3558 ( .A(n3507), .Z(n3506) );
  NOR U3559 ( .A(sum[31]), .B(n3506), .Z(n3445) );
  NOR U3560 ( .A(n3507), .B(o[223]), .Z(n3444) );
  NOR U3561 ( .A(n3445), .B(n3444), .Z(n782) );
  NOR U3562 ( .A(sum[30]), .B(n3506), .Z(n3447) );
  NOR U3563 ( .A(n3507), .B(o[222]), .Z(n3446) );
  NOR U3564 ( .A(n3447), .B(n3446), .Z(n783) );
  NOR U3565 ( .A(sum[29]), .B(n3506), .Z(n3449) );
  NOR U3566 ( .A(n3507), .B(o[221]), .Z(n3448) );
  NOR U3567 ( .A(n3449), .B(n3448), .Z(n784) );
  NOR U3568 ( .A(sum[28]), .B(n3506), .Z(n3451) );
  NOR U3569 ( .A(n3507), .B(o[220]), .Z(n3450) );
  NOR U3570 ( .A(n3451), .B(n3450), .Z(n785) );
  NOR U3571 ( .A(sum[27]), .B(n3506), .Z(n3453) );
  NOR U3572 ( .A(n3507), .B(o[219]), .Z(n3452) );
  NOR U3573 ( .A(n3453), .B(n3452), .Z(n786) );
  NOR U3574 ( .A(sum[26]), .B(n3506), .Z(n3455) );
  NOR U3575 ( .A(n3507), .B(o[218]), .Z(n3454) );
  NOR U3576 ( .A(n3455), .B(n3454), .Z(n787) );
  NOR U3577 ( .A(sum[25]), .B(n3506), .Z(n3457) );
  NOR U3578 ( .A(n3507), .B(o[217]), .Z(n3456) );
  NOR U3579 ( .A(n3457), .B(n3456), .Z(n788) );
  NOR U3580 ( .A(sum[24]), .B(n3506), .Z(n3459) );
  NOR U3581 ( .A(n3507), .B(o[216]), .Z(n3458) );
  NOR U3582 ( .A(n3459), .B(n3458), .Z(n789) );
  NOR U3583 ( .A(sum[23]), .B(n3506), .Z(n3461) );
  NOR U3584 ( .A(n3507), .B(o[215]), .Z(n3460) );
  NOR U3585 ( .A(n3461), .B(n3460), .Z(n790) );
  NOR U3586 ( .A(sum[22]), .B(n3506), .Z(n3463) );
  NOR U3587 ( .A(n3507), .B(o[214]), .Z(n3462) );
  NOR U3588 ( .A(n3463), .B(n3462), .Z(n791) );
  NOR U3589 ( .A(sum[21]), .B(n3506), .Z(n3465) );
  NOR U3590 ( .A(n3507), .B(o[213]), .Z(n3464) );
  NOR U3591 ( .A(n3465), .B(n3464), .Z(n792) );
  NOR U3592 ( .A(sum[20]), .B(n3506), .Z(n3467) );
  NOR U3593 ( .A(n3507), .B(o[212]), .Z(n3466) );
  NOR U3594 ( .A(n3467), .B(n3466), .Z(n793) );
  NOR U3595 ( .A(sum[19]), .B(n3506), .Z(n3469) );
  NOR U3596 ( .A(n3507), .B(o[211]), .Z(n3468) );
  NOR U3597 ( .A(n3469), .B(n3468), .Z(n794) );
  NOR U3598 ( .A(sum[18]), .B(n3506), .Z(n3471) );
  NOR U3599 ( .A(n3507), .B(o[210]), .Z(n3470) );
  NOR U3600 ( .A(n3471), .B(n3470), .Z(n795) );
  NOR U3601 ( .A(sum[17]), .B(n3506), .Z(n3473) );
  NOR U3602 ( .A(n3507), .B(o[209]), .Z(n3472) );
  NOR U3603 ( .A(n3473), .B(n3472), .Z(n796) );
  NOR U3604 ( .A(sum[16]), .B(n3506), .Z(n3475) );
  NOR U3605 ( .A(n3507), .B(o[208]), .Z(n3474) );
  NOR U3606 ( .A(n3475), .B(n3474), .Z(n797) );
  NOR U3607 ( .A(sum[15]), .B(n3506), .Z(n3477) );
  NOR U3608 ( .A(n3507), .B(o[207]), .Z(n3476) );
  NOR U3609 ( .A(n3477), .B(n3476), .Z(n798) );
  NOR U3610 ( .A(sum[14]), .B(n3506), .Z(n3479) );
  NOR U3611 ( .A(n3507), .B(o[206]), .Z(n3478) );
  NOR U3612 ( .A(n3479), .B(n3478), .Z(n799) );
  NOR U3613 ( .A(sum[13]), .B(n3506), .Z(n3481) );
  NOR U3614 ( .A(n3507), .B(o[205]), .Z(n3480) );
  NOR U3615 ( .A(n3481), .B(n3480), .Z(n800) );
  NOR U3616 ( .A(sum[12]), .B(n3506), .Z(n3483) );
  NOR U3617 ( .A(n3507), .B(o[204]), .Z(n3482) );
  NOR U3618 ( .A(n3483), .B(n3482), .Z(n801) );
  NOR U3619 ( .A(sum[11]), .B(n3506), .Z(n3485) );
  NOR U3620 ( .A(n3507), .B(o[203]), .Z(n3484) );
  NOR U3621 ( .A(n3485), .B(n3484), .Z(n802) );
  NOR U3622 ( .A(sum[10]), .B(n3506), .Z(n3487) );
  NOR U3623 ( .A(n3507), .B(o[202]), .Z(n3486) );
  NOR U3624 ( .A(n3487), .B(n3486), .Z(n803) );
  NOR U3625 ( .A(sum[9]), .B(n3506), .Z(n3489) );
  NOR U3626 ( .A(n3507), .B(o[201]), .Z(n3488) );
  NOR U3627 ( .A(n3489), .B(n3488), .Z(n804) );
  NOR U3628 ( .A(sum[8]), .B(n3506), .Z(n3491) );
  NOR U3629 ( .A(n3507), .B(o[200]), .Z(n3490) );
  NOR U3630 ( .A(n3491), .B(n3490), .Z(n805) );
  NOR U3631 ( .A(sum[7]), .B(n3506), .Z(n3493) );
  NOR U3632 ( .A(n3507), .B(o[199]), .Z(n3492) );
  NOR U3633 ( .A(n3493), .B(n3492), .Z(n806) );
  NOR U3634 ( .A(sum[6]), .B(n3506), .Z(n3495) );
  NOR U3635 ( .A(n3507), .B(o[198]), .Z(n3494) );
  NOR U3636 ( .A(n3495), .B(n3494), .Z(n807) );
  NOR U3637 ( .A(sum[5]), .B(n3506), .Z(n3497) );
  NOR U3638 ( .A(n3507), .B(o[197]), .Z(n3496) );
  NOR U3639 ( .A(n3497), .B(n3496), .Z(n808) );
  NOR U3640 ( .A(sum[4]), .B(n3506), .Z(n3499) );
  NOR U3641 ( .A(n3507), .B(o[196]), .Z(n3498) );
  NOR U3642 ( .A(n3499), .B(n3498), .Z(n809) );
  NOR U3643 ( .A(sum[3]), .B(n3506), .Z(n3501) );
  NOR U3644 ( .A(n3507), .B(o[195]), .Z(n3500) );
  NOR U3645 ( .A(n3501), .B(n3500), .Z(n810) );
  NOR U3646 ( .A(sum[2]), .B(n3506), .Z(n3503) );
  NOR U3647 ( .A(n3507), .B(o[194]), .Z(n3502) );
  NOR U3648 ( .A(n3503), .B(n3502), .Z(n811) );
  NOR U3649 ( .A(sum[1]), .B(n3506), .Z(n3505) );
  NOR U3650 ( .A(n3507), .B(o[193]), .Z(n3504) );
  NOR U3651 ( .A(n3505), .B(n3504), .Z(n812) );
  NOR U3652 ( .A(sum[0]), .B(n3506), .Z(n3509) );
  NOR U3653 ( .A(n3507), .B(o[192]), .Z(n3508) );
  NOR U3654 ( .A(n3509), .B(n3508), .Z(n813) );
  NOR U3655 ( .A(n3875), .B(n3576), .Z(n3573) );
  IV U3656 ( .A(n3573), .Z(n3572) );
  NOR U3657 ( .A(sum[31]), .B(n3572), .Z(n3511) );
  NOR U3658 ( .A(n3573), .B(o[127]), .Z(n3510) );
  NOR U3659 ( .A(n3511), .B(n3510), .Z(n814) );
  NOR U3660 ( .A(sum[30]), .B(n3572), .Z(n3513) );
  NOR U3661 ( .A(n3573), .B(o[126]), .Z(n3512) );
  NOR U3662 ( .A(n3513), .B(n3512), .Z(n815) );
  NOR U3663 ( .A(sum[29]), .B(n3572), .Z(n3515) );
  NOR U3664 ( .A(n3573), .B(o[125]), .Z(n3514) );
  NOR U3665 ( .A(n3515), .B(n3514), .Z(n816) );
  NOR U3666 ( .A(sum[28]), .B(n3572), .Z(n3517) );
  NOR U3667 ( .A(n3573), .B(o[124]), .Z(n3516) );
  NOR U3668 ( .A(n3517), .B(n3516), .Z(n817) );
  NOR U3669 ( .A(sum[27]), .B(n3572), .Z(n3519) );
  NOR U3670 ( .A(n3573), .B(o[123]), .Z(n3518) );
  NOR U3671 ( .A(n3519), .B(n3518), .Z(n818) );
  NOR U3672 ( .A(sum[26]), .B(n3572), .Z(n3521) );
  NOR U3673 ( .A(n3573), .B(o[122]), .Z(n3520) );
  NOR U3674 ( .A(n3521), .B(n3520), .Z(n819) );
  NOR U3675 ( .A(sum[25]), .B(n3572), .Z(n3523) );
  NOR U3676 ( .A(n3573), .B(o[121]), .Z(n3522) );
  NOR U3677 ( .A(n3523), .B(n3522), .Z(n820) );
  NOR U3678 ( .A(sum[24]), .B(n3572), .Z(n3525) );
  NOR U3679 ( .A(n3573), .B(o[120]), .Z(n3524) );
  NOR U3680 ( .A(n3525), .B(n3524), .Z(n821) );
  NOR U3681 ( .A(sum[23]), .B(n3572), .Z(n3527) );
  NOR U3682 ( .A(n3573), .B(o[119]), .Z(n3526) );
  NOR U3683 ( .A(n3527), .B(n3526), .Z(n822) );
  NOR U3684 ( .A(sum[22]), .B(n3572), .Z(n3529) );
  NOR U3685 ( .A(n3573), .B(o[118]), .Z(n3528) );
  NOR U3686 ( .A(n3529), .B(n3528), .Z(n823) );
  NOR U3687 ( .A(sum[21]), .B(n3572), .Z(n3531) );
  NOR U3688 ( .A(n3573), .B(o[117]), .Z(n3530) );
  NOR U3689 ( .A(n3531), .B(n3530), .Z(n824) );
  NOR U3690 ( .A(sum[20]), .B(n3572), .Z(n3533) );
  NOR U3691 ( .A(n3573), .B(o[116]), .Z(n3532) );
  NOR U3692 ( .A(n3533), .B(n3532), .Z(n825) );
  NOR U3693 ( .A(sum[19]), .B(n3572), .Z(n3535) );
  NOR U3694 ( .A(n3573), .B(o[115]), .Z(n3534) );
  NOR U3695 ( .A(n3535), .B(n3534), .Z(n826) );
  NOR U3696 ( .A(sum[18]), .B(n3572), .Z(n3537) );
  NOR U3697 ( .A(n3573), .B(o[114]), .Z(n3536) );
  NOR U3698 ( .A(n3537), .B(n3536), .Z(n827) );
  NOR U3699 ( .A(sum[17]), .B(n3572), .Z(n3539) );
  NOR U3700 ( .A(n3573), .B(o[113]), .Z(n3538) );
  NOR U3701 ( .A(n3539), .B(n3538), .Z(n828) );
  NOR U3702 ( .A(sum[16]), .B(n3572), .Z(n3541) );
  NOR U3703 ( .A(n3573), .B(o[112]), .Z(n3540) );
  NOR U3704 ( .A(n3541), .B(n3540), .Z(n829) );
  NOR U3705 ( .A(sum[15]), .B(n3572), .Z(n3543) );
  NOR U3706 ( .A(n3573), .B(o[111]), .Z(n3542) );
  NOR U3707 ( .A(n3543), .B(n3542), .Z(n830) );
  NOR U3708 ( .A(sum[14]), .B(n3572), .Z(n3545) );
  NOR U3709 ( .A(n3573), .B(o[110]), .Z(n3544) );
  NOR U3710 ( .A(n3545), .B(n3544), .Z(n831) );
  NOR U3711 ( .A(sum[13]), .B(n3572), .Z(n3547) );
  NOR U3712 ( .A(n3573), .B(o[109]), .Z(n3546) );
  NOR U3713 ( .A(n3547), .B(n3546), .Z(n832) );
  NOR U3714 ( .A(sum[12]), .B(n3572), .Z(n3549) );
  NOR U3715 ( .A(n3573), .B(o[108]), .Z(n3548) );
  NOR U3716 ( .A(n3549), .B(n3548), .Z(n833) );
  NOR U3717 ( .A(sum[11]), .B(n3572), .Z(n3551) );
  NOR U3718 ( .A(n3573), .B(o[107]), .Z(n3550) );
  NOR U3719 ( .A(n3551), .B(n3550), .Z(n834) );
  NOR U3720 ( .A(sum[10]), .B(n3572), .Z(n3553) );
  NOR U3721 ( .A(n3573), .B(o[106]), .Z(n3552) );
  NOR U3722 ( .A(n3553), .B(n3552), .Z(n835) );
  NOR U3723 ( .A(sum[9]), .B(n3572), .Z(n3555) );
  NOR U3724 ( .A(n3573), .B(o[105]), .Z(n3554) );
  NOR U3725 ( .A(n3555), .B(n3554), .Z(n836) );
  NOR U3726 ( .A(sum[8]), .B(n3572), .Z(n3557) );
  NOR U3727 ( .A(n3573), .B(o[104]), .Z(n3556) );
  NOR U3728 ( .A(n3557), .B(n3556), .Z(n837) );
  NOR U3729 ( .A(sum[7]), .B(n3572), .Z(n3559) );
  NOR U3730 ( .A(n3573), .B(o[103]), .Z(n3558) );
  NOR U3731 ( .A(n3559), .B(n3558), .Z(n838) );
  NOR U3732 ( .A(sum[6]), .B(n3572), .Z(n3561) );
  NOR U3733 ( .A(n3573), .B(o[102]), .Z(n3560) );
  NOR U3734 ( .A(n3561), .B(n3560), .Z(n839) );
  NOR U3735 ( .A(sum[5]), .B(n3572), .Z(n3563) );
  NOR U3736 ( .A(n3573), .B(o[101]), .Z(n3562) );
  NOR U3737 ( .A(n3563), .B(n3562), .Z(n840) );
  NOR U3738 ( .A(sum[4]), .B(n3572), .Z(n3565) );
  NOR U3739 ( .A(n3573), .B(o[100]), .Z(n3564) );
  NOR U3740 ( .A(n3565), .B(n3564), .Z(n841) );
  NOR U3741 ( .A(sum[3]), .B(n3572), .Z(n3567) );
  NOR U3742 ( .A(n3573), .B(o[99]), .Z(n3566) );
  NOR U3743 ( .A(n3567), .B(n3566), .Z(n842) );
  NOR U3744 ( .A(sum[2]), .B(n3572), .Z(n3569) );
  NOR U3745 ( .A(n3573), .B(o[98]), .Z(n3568) );
  NOR U3746 ( .A(n3569), .B(n3568), .Z(n843) );
  NOR U3747 ( .A(sum[1]), .B(n3572), .Z(n3571) );
  NOR U3748 ( .A(n3573), .B(o[97]), .Z(n3570) );
  NOR U3749 ( .A(n3571), .B(n3570), .Z(n844) );
  NOR U3750 ( .A(sum[0]), .B(n3572), .Z(n3575) );
  NOR U3751 ( .A(n3573), .B(o[96]), .Z(n3574) );
  NOR U3752 ( .A(n3575), .B(n3574), .Z(n845) );
  NOR U3753 ( .A(n3866), .B(n3576), .Z(n3640) );
  IV U3754 ( .A(n3640), .Z(n3639) );
  NOR U3755 ( .A(sum[31]), .B(n3639), .Z(n3578) );
  NOR U3756 ( .A(n3640), .B(o[31]), .Z(n3577) );
  NOR U3757 ( .A(n3578), .B(n3577), .Z(n846) );
  NOR U3758 ( .A(sum[30]), .B(n3639), .Z(n3580) );
  NOR U3759 ( .A(n3640), .B(o[30]), .Z(n3579) );
  NOR U3760 ( .A(n3580), .B(n3579), .Z(n847) );
  NOR U3761 ( .A(sum[29]), .B(n3639), .Z(n3582) );
  NOR U3762 ( .A(n3640), .B(o[29]), .Z(n3581) );
  NOR U3763 ( .A(n3582), .B(n3581), .Z(n848) );
  NOR U3764 ( .A(sum[28]), .B(n3639), .Z(n3584) );
  NOR U3765 ( .A(n3640), .B(o[28]), .Z(n3583) );
  NOR U3766 ( .A(n3584), .B(n3583), .Z(n849) );
  NOR U3767 ( .A(sum[27]), .B(n3639), .Z(n3586) );
  NOR U3768 ( .A(n3640), .B(o[27]), .Z(n3585) );
  NOR U3769 ( .A(n3586), .B(n3585), .Z(n850) );
  NOR U3770 ( .A(sum[26]), .B(n3639), .Z(n3588) );
  NOR U3771 ( .A(n3640), .B(o[26]), .Z(n3587) );
  NOR U3772 ( .A(n3588), .B(n3587), .Z(n851) );
  NOR U3773 ( .A(sum[25]), .B(n3639), .Z(n3590) );
  NOR U3774 ( .A(n3640), .B(o[25]), .Z(n3589) );
  NOR U3775 ( .A(n3590), .B(n3589), .Z(n852) );
  NOR U3776 ( .A(sum[24]), .B(n3639), .Z(n3592) );
  NOR U3777 ( .A(n3640), .B(o[24]), .Z(n3591) );
  NOR U3778 ( .A(n3592), .B(n3591), .Z(n853) );
  NOR U3779 ( .A(sum[23]), .B(n3639), .Z(n3594) );
  NOR U3780 ( .A(n3640), .B(o[23]), .Z(n3593) );
  NOR U3781 ( .A(n3594), .B(n3593), .Z(n854) );
  NOR U3782 ( .A(sum[22]), .B(n3639), .Z(n3596) );
  NOR U3783 ( .A(n3640), .B(o[22]), .Z(n3595) );
  NOR U3784 ( .A(n3596), .B(n3595), .Z(n855) );
  NOR U3785 ( .A(sum[21]), .B(n3639), .Z(n3598) );
  NOR U3786 ( .A(n3640), .B(o[21]), .Z(n3597) );
  NOR U3787 ( .A(n3598), .B(n3597), .Z(n856) );
  NOR U3788 ( .A(sum[20]), .B(n3639), .Z(n3600) );
  NOR U3789 ( .A(n3640), .B(o[20]), .Z(n3599) );
  NOR U3790 ( .A(n3600), .B(n3599), .Z(n857) );
  NOR U3791 ( .A(sum[19]), .B(n3639), .Z(n3602) );
  NOR U3792 ( .A(n3640), .B(o[19]), .Z(n3601) );
  NOR U3793 ( .A(n3602), .B(n3601), .Z(n858) );
  NOR U3794 ( .A(sum[18]), .B(n3639), .Z(n3604) );
  NOR U3795 ( .A(n3640), .B(o[18]), .Z(n3603) );
  NOR U3796 ( .A(n3604), .B(n3603), .Z(n859) );
  NOR U3797 ( .A(sum[17]), .B(n3639), .Z(n3606) );
  NOR U3798 ( .A(n3640), .B(o[17]), .Z(n3605) );
  NOR U3799 ( .A(n3606), .B(n3605), .Z(n860) );
  NOR U3800 ( .A(sum[16]), .B(n3639), .Z(n3608) );
  NOR U3801 ( .A(n3640), .B(o[16]), .Z(n3607) );
  NOR U3802 ( .A(n3608), .B(n3607), .Z(n861) );
  NOR U3803 ( .A(sum[15]), .B(n3639), .Z(n3610) );
  NOR U3804 ( .A(n3640), .B(o[15]), .Z(n3609) );
  NOR U3805 ( .A(n3610), .B(n3609), .Z(n862) );
  NOR U3806 ( .A(sum[14]), .B(n3639), .Z(n3612) );
  NOR U3807 ( .A(n3640), .B(o[14]), .Z(n3611) );
  NOR U3808 ( .A(n3612), .B(n3611), .Z(n863) );
  NOR U3809 ( .A(sum[13]), .B(n3639), .Z(n3614) );
  NOR U3810 ( .A(n3640), .B(o[13]), .Z(n3613) );
  NOR U3811 ( .A(n3614), .B(n3613), .Z(n864) );
  NOR U3812 ( .A(sum[12]), .B(n3639), .Z(n3616) );
  NOR U3813 ( .A(n3640), .B(o[12]), .Z(n3615) );
  NOR U3814 ( .A(n3616), .B(n3615), .Z(n865) );
  NOR U3815 ( .A(sum[11]), .B(n3639), .Z(n3618) );
  NOR U3816 ( .A(n3640), .B(o[11]), .Z(n3617) );
  NOR U3817 ( .A(n3618), .B(n3617), .Z(n866) );
  NOR U3818 ( .A(sum[10]), .B(n3639), .Z(n3620) );
  NOR U3819 ( .A(n3640), .B(o[10]), .Z(n3619) );
  NOR U3820 ( .A(n3620), .B(n3619), .Z(n867) );
  NOR U3821 ( .A(sum[9]), .B(n3639), .Z(n3622) );
  NOR U3822 ( .A(n3640), .B(o[9]), .Z(n3621) );
  NOR U3823 ( .A(n3622), .B(n3621), .Z(n868) );
  NOR U3824 ( .A(sum[8]), .B(n3639), .Z(n3624) );
  NOR U3825 ( .A(n3640), .B(o[8]), .Z(n3623) );
  NOR U3826 ( .A(n3624), .B(n3623), .Z(n869) );
  NOR U3827 ( .A(sum[7]), .B(n3639), .Z(n3626) );
  NOR U3828 ( .A(n3640), .B(o[7]), .Z(n3625) );
  NOR U3829 ( .A(n3626), .B(n3625), .Z(n870) );
  NOR U3830 ( .A(sum[6]), .B(n3639), .Z(n3628) );
  NOR U3831 ( .A(n3640), .B(o[6]), .Z(n3627) );
  NOR U3832 ( .A(n3628), .B(n3627), .Z(n871) );
  NOR U3833 ( .A(sum[5]), .B(n3639), .Z(n3630) );
  NOR U3834 ( .A(n3640), .B(o[5]), .Z(n3629) );
  NOR U3835 ( .A(n3630), .B(n3629), .Z(n872) );
  NOR U3836 ( .A(sum[4]), .B(n3639), .Z(n3632) );
  NOR U3837 ( .A(n3640), .B(o[4]), .Z(n3631) );
  NOR U3838 ( .A(n3632), .B(n3631), .Z(n873) );
  NOR U3839 ( .A(sum[3]), .B(n3639), .Z(n3634) );
  NOR U3840 ( .A(n3640), .B(o[3]), .Z(n3633) );
  NOR U3841 ( .A(n3634), .B(n3633), .Z(n874) );
  NOR U3842 ( .A(sum[2]), .B(n3639), .Z(n3636) );
  NOR U3843 ( .A(n3640), .B(o[2]), .Z(n3635) );
  NOR U3844 ( .A(n3636), .B(n3635), .Z(n875) );
  NOR U3845 ( .A(sum[1]), .B(n3639), .Z(n3638) );
  NOR U3846 ( .A(n3640), .B(o[1]), .Z(n3637) );
  NOR U3847 ( .A(n3638), .B(n3637), .Z(n876) );
  NOR U3848 ( .A(sum[0]), .B(n3639), .Z(n3642) );
  NOR U3849 ( .A(n3640), .B(o[0]), .Z(n3641) );
  NOR U3850 ( .A(n3642), .B(n3641), .Z(n877) );
  IV U3851 ( .A(j[1]), .Z(n3921) );
  NOR U3852 ( .A(n3921), .B(n3845), .Z(n3643) );
  IV U3853 ( .A(n3643), .Z(n3644) );
  NOR U3854 ( .A(j[0]), .B(n3644), .Z(n9906) );
  IV U3855 ( .A(n9906), .Z(n3775) );
  NOR U3856 ( .A(n3872), .B(n3775), .Z(n3708) );
  IV U3857 ( .A(n3708), .Z(n3707) );
  NOR U3858 ( .A(sum[31]), .B(n3707), .Z(n3646) );
  NOR U3859 ( .A(n3708), .B(o[287]), .Z(n3645) );
  NOR U3860 ( .A(n3646), .B(n3645), .Z(n878) );
  NOR U3861 ( .A(sum[30]), .B(n3707), .Z(n3648) );
  NOR U3862 ( .A(n3708), .B(o[286]), .Z(n3647) );
  NOR U3863 ( .A(n3648), .B(n3647), .Z(n879) );
  NOR U3864 ( .A(sum[29]), .B(n3707), .Z(n3650) );
  NOR U3865 ( .A(n3708), .B(o[285]), .Z(n3649) );
  NOR U3866 ( .A(n3650), .B(n3649), .Z(n880) );
  NOR U3867 ( .A(sum[28]), .B(n3707), .Z(n3652) );
  NOR U3868 ( .A(n3708), .B(o[284]), .Z(n3651) );
  NOR U3869 ( .A(n3652), .B(n3651), .Z(n881) );
  NOR U3870 ( .A(sum[27]), .B(n3707), .Z(n3654) );
  NOR U3871 ( .A(n3708), .B(o[283]), .Z(n3653) );
  NOR U3872 ( .A(n3654), .B(n3653), .Z(n882) );
  NOR U3873 ( .A(sum[26]), .B(n3707), .Z(n3656) );
  NOR U3874 ( .A(n3708), .B(o[282]), .Z(n3655) );
  NOR U3875 ( .A(n3656), .B(n3655), .Z(n883) );
  NOR U3876 ( .A(sum[25]), .B(n3707), .Z(n3658) );
  NOR U3877 ( .A(n3708), .B(o[281]), .Z(n3657) );
  NOR U3878 ( .A(n3658), .B(n3657), .Z(n884) );
  NOR U3879 ( .A(sum[24]), .B(n3707), .Z(n3660) );
  NOR U3880 ( .A(n3708), .B(o[280]), .Z(n3659) );
  NOR U3881 ( .A(n3660), .B(n3659), .Z(n885) );
  NOR U3882 ( .A(sum[23]), .B(n3707), .Z(n3662) );
  NOR U3883 ( .A(n3708), .B(o[279]), .Z(n3661) );
  NOR U3884 ( .A(n3662), .B(n3661), .Z(n886) );
  NOR U3885 ( .A(sum[22]), .B(n3707), .Z(n3664) );
  NOR U3886 ( .A(n3708), .B(o[278]), .Z(n3663) );
  NOR U3887 ( .A(n3664), .B(n3663), .Z(n887) );
  NOR U3888 ( .A(sum[21]), .B(n3707), .Z(n3666) );
  NOR U3889 ( .A(n3708), .B(o[277]), .Z(n3665) );
  NOR U3890 ( .A(n3666), .B(n3665), .Z(n888) );
  NOR U3891 ( .A(sum[20]), .B(n3707), .Z(n3668) );
  NOR U3892 ( .A(n3708), .B(o[276]), .Z(n3667) );
  NOR U3893 ( .A(n3668), .B(n3667), .Z(n889) );
  NOR U3894 ( .A(sum[19]), .B(n3707), .Z(n3670) );
  NOR U3895 ( .A(n3708), .B(o[275]), .Z(n3669) );
  NOR U3896 ( .A(n3670), .B(n3669), .Z(n890) );
  NOR U3897 ( .A(sum[18]), .B(n3707), .Z(n3672) );
  NOR U3898 ( .A(n3708), .B(o[274]), .Z(n3671) );
  NOR U3899 ( .A(n3672), .B(n3671), .Z(n891) );
  NOR U3900 ( .A(sum[17]), .B(n3707), .Z(n3674) );
  NOR U3901 ( .A(n3708), .B(o[273]), .Z(n3673) );
  NOR U3902 ( .A(n3674), .B(n3673), .Z(n892) );
  NOR U3903 ( .A(sum[16]), .B(n3707), .Z(n3676) );
  NOR U3904 ( .A(n3708), .B(o[272]), .Z(n3675) );
  NOR U3905 ( .A(n3676), .B(n3675), .Z(n893) );
  NOR U3906 ( .A(sum[15]), .B(n3707), .Z(n3678) );
  NOR U3907 ( .A(n3708), .B(o[271]), .Z(n3677) );
  NOR U3908 ( .A(n3678), .B(n3677), .Z(n894) );
  NOR U3909 ( .A(sum[14]), .B(n3707), .Z(n3680) );
  NOR U3910 ( .A(n3708), .B(o[270]), .Z(n3679) );
  NOR U3911 ( .A(n3680), .B(n3679), .Z(n895) );
  NOR U3912 ( .A(sum[13]), .B(n3707), .Z(n3682) );
  NOR U3913 ( .A(n3708), .B(o[269]), .Z(n3681) );
  NOR U3914 ( .A(n3682), .B(n3681), .Z(n896) );
  NOR U3915 ( .A(sum[12]), .B(n3707), .Z(n3684) );
  NOR U3916 ( .A(n3708), .B(o[268]), .Z(n3683) );
  NOR U3917 ( .A(n3684), .B(n3683), .Z(n897) );
  NOR U3918 ( .A(sum[11]), .B(n3707), .Z(n3686) );
  NOR U3919 ( .A(n3708), .B(o[267]), .Z(n3685) );
  NOR U3920 ( .A(n3686), .B(n3685), .Z(n898) );
  NOR U3921 ( .A(sum[10]), .B(n3707), .Z(n3688) );
  NOR U3922 ( .A(n3708), .B(o[266]), .Z(n3687) );
  NOR U3923 ( .A(n3688), .B(n3687), .Z(n899) );
  NOR U3924 ( .A(sum[9]), .B(n3707), .Z(n3690) );
  NOR U3925 ( .A(n3708), .B(o[265]), .Z(n3689) );
  NOR U3926 ( .A(n3690), .B(n3689), .Z(n900) );
  NOR U3927 ( .A(sum[8]), .B(n3707), .Z(n3692) );
  NOR U3928 ( .A(n3708), .B(o[264]), .Z(n3691) );
  NOR U3929 ( .A(n3692), .B(n3691), .Z(n901) );
  NOR U3930 ( .A(sum[7]), .B(n3707), .Z(n3694) );
  NOR U3931 ( .A(n3708), .B(o[263]), .Z(n3693) );
  NOR U3932 ( .A(n3694), .B(n3693), .Z(n902) );
  NOR U3933 ( .A(sum[6]), .B(n3707), .Z(n3696) );
  NOR U3934 ( .A(n3708), .B(o[262]), .Z(n3695) );
  NOR U3935 ( .A(n3696), .B(n3695), .Z(n903) );
  NOR U3936 ( .A(sum[5]), .B(n3707), .Z(n3698) );
  NOR U3937 ( .A(n3708), .B(o[261]), .Z(n3697) );
  NOR U3938 ( .A(n3698), .B(n3697), .Z(n904) );
  NOR U3939 ( .A(sum[4]), .B(n3707), .Z(n3700) );
  NOR U3940 ( .A(n3708), .B(o[260]), .Z(n3699) );
  NOR U3941 ( .A(n3700), .B(n3699), .Z(n905) );
  NOR U3942 ( .A(sum[3]), .B(n3707), .Z(n3702) );
  NOR U3943 ( .A(n3708), .B(o[259]), .Z(n3701) );
  NOR U3944 ( .A(n3702), .B(n3701), .Z(n906) );
  NOR U3945 ( .A(sum[2]), .B(n3707), .Z(n3704) );
  NOR U3946 ( .A(n3708), .B(o[258]), .Z(n3703) );
  NOR U3947 ( .A(n3704), .B(n3703), .Z(n907) );
  NOR U3948 ( .A(sum[1]), .B(n3707), .Z(n3706) );
  NOR U3949 ( .A(n3708), .B(o[257]), .Z(n3705) );
  NOR U3950 ( .A(n3706), .B(n3705), .Z(n908) );
  NOR U3951 ( .A(sum[0]), .B(n3707), .Z(n3710) );
  NOR U3952 ( .A(n3708), .B(o[256]), .Z(n3709) );
  NOR U3953 ( .A(n3710), .B(n3709), .Z(n909) );
  NOR U3954 ( .A(n3875), .B(n3775), .Z(n3841) );
  NOR U3955 ( .A(sum[31]), .B(n3236), .Z(n3712) );
  NOR U3956 ( .A(n3841), .B(o[191]), .Z(n3711) );
  NOR U3957 ( .A(n3712), .B(n3711), .Z(n910) );
  NOR U3958 ( .A(sum[30]), .B(n3236), .Z(n3714) );
  NOR U3959 ( .A(n3841), .B(o[190]), .Z(n3713) );
  NOR U3960 ( .A(n3714), .B(n3713), .Z(n911) );
  NOR U3961 ( .A(sum[29]), .B(n3236), .Z(n3716) );
  NOR U3962 ( .A(n3841), .B(o[189]), .Z(n3715) );
  NOR U3963 ( .A(n3716), .B(n3715), .Z(n912) );
  NOR U3964 ( .A(sum[28]), .B(n3236), .Z(n3718) );
  NOR U3965 ( .A(n3841), .B(o[188]), .Z(n3717) );
  NOR U3966 ( .A(n3718), .B(n3717), .Z(n913) );
  NOR U3967 ( .A(sum[27]), .B(n3236), .Z(n3720) );
  NOR U3968 ( .A(n3841), .B(o[187]), .Z(n3719) );
  NOR U3969 ( .A(n3720), .B(n3719), .Z(n914) );
  NOR U3970 ( .A(sum[26]), .B(n3236), .Z(n3722) );
  NOR U3971 ( .A(n3841), .B(o[186]), .Z(n3721) );
  NOR U3972 ( .A(n3722), .B(n3721), .Z(n915) );
  NOR U3973 ( .A(sum[25]), .B(n3236), .Z(n3724) );
  NOR U3974 ( .A(n3841), .B(o[185]), .Z(n3723) );
  NOR U3975 ( .A(n3724), .B(n3723), .Z(n916) );
  NOR U3976 ( .A(sum[24]), .B(n3236), .Z(n3726) );
  NOR U3977 ( .A(n3841), .B(o[184]), .Z(n3725) );
  NOR U3978 ( .A(n3726), .B(n3725), .Z(n917) );
  NOR U3979 ( .A(sum[23]), .B(n3236), .Z(n3728) );
  NOR U3980 ( .A(n3841), .B(o[183]), .Z(n3727) );
  NOR U3981 ( .A(n3728), .B(n3727), .Z(n918) );
  NOR U3982 ( .A(sum[22]), .B(n3236), .Z(n3730) );
  NOR U3983 ( .A(n3841), .B(o[182]), .Z(n3729) );
  NOR U3984 ( .A(n3730), .B(n3729), .Z(n919) );
  NOR U3985 ( .A(sum[21]), .B(n3236), .Z(n3732) );
  NOR U3986 ( .A(n3841), .B(o[181]), .Z(n3731) );
  NOR U3987 ( .A(n3732), .B(n3731), .Z(n920) );
  NOR U3988 ( .A(sum[20]), .B(n3236), .Z(n3734) );
  NOR U3989 ( .A(n3841), .B(o[180]), .Z(n3733) );
  NOR U3990 ( .A(n3734), .B(n3733), .Z(n921) );
  NOR U3991 ( .A(sum[19]), .B(n3236), .Z(n3736) );
  NOR U3992 ( .A(n3841), .B(o[179]), .Z(n3735) );
  NOR U3993 ( .A(n3736), .B(n3735), .Z(n922) );
  NOR U3994 ( .A(sum[18]), .B(n3236), .Z(n3738) );
  NOR U3995 ( .A(n3841), .B(o[178]), .Z(n3737) );
  NOR U3996 ( .A(n3738), .B(n3737), .Z(n923) );
  NOR U3997 ( .A(sum[17]), .B(n3236), .Z(n3740) );
  NOR U3998 ( .A(n3841), .B(o[177]), .Z(n3739) );
  NOR U3999 ( .A(n3740), .B(n3739), .Z(n924) );
  NOR U4000 ( .A(sum[16]), .B(n3236), .Z(n3742) );
  NOR U4001 ( .A(n3841), .B(o[176]), .Z(n3741) );
  NOR U4002 ( .A(n3742), .B(n3741), .Z(n925) );
  NOR U4003 ( .A(sum[15]), .B(n3236), .Z(n3744) );
  NOR U4004 ( .A(n3841), .B(o[175]), .Z(n3743) );
  NOR U4005 ( .A(n3744), .B(n3743), .Z(n926) );
  NOR U4006 ( .A(sum[14]), .B(n3236), .Z(n3746) );
  NOR U4007 ( .A(n3841), .B(o[174]), .Z(n3745) );
  NOR U4008 ( .A(n3746), .B(n3745), .Z(n927) );
  NOR U4009 ( .A(sum[13]), .B(n3236), .Z(n3748) );
  NOR U4010 ( .A(n3841), .B(o[173]), .Z(n3747) );
  NOR U4011 ( .A(n3748), .B(n3747), .Z(n928) );
  NOR U4012 ( .A(sum[12]), .B(n3236), .Z(n3750) );
  NOR U4013 ( .A(n3841), .B(o[172]), .Z(n3749) );
  NOR U4014 ( .A(n3750), .B(n3749), .Z(n929) );
  NOR U4015 ( .A(sum[11]), .B(n3236), .Z(n3752) );
  NOR U4016 ( .A(n3841), .B(o[171]), .Z(n3751) );
  NOR U4017 ( .A(n3752), .B(n3751), .Z(n930) );
  NOR U4018 ( .A(sum[10]), .B(n3236), .Z(n3754) );
  NOR U4019 ( .A(n3841), .B(o[170]), .Z(n3753) );
  NOR U4020 ( .A(n3754), .B(n3753), .Z(n931) );
  NOR U4021 ( .A(sum[9]), .B(n3236), .Z(n3756) );
  NOR U4022 ( .A(n3841), .B(o[169]), .Z(n3755) );
  NOR U4023 ( .A(n3756), .B(n3755), .Z(n932) );
  NOR U4024 ( .A(sum[8]), .B(n3236), .Z(n3758) );
  NOR U4025 ( .A(n3841), .B(o[168]), .Z(n3757) );
  NOR U4026 ( .A(n3758), .B(n3757), .Z(n933) );
  NOR U4027 ( .A(sum[7]), .B(n3236), .Z(n3760) );
  NOR U4028 ( .A(n3841), .B(o[167]), .Z(n3759) );
  NOR U4029 ( .A(n3760), .B(n3759), .Z(n934) );
  NOR U4030 ( .A(sum[6]), .B(n3236), .Z(n3762) );
  NOR U4031 ( .A(n3841), .B(o[166]), .Z(n3761) );
  NOR U4032 ( .A(n3762), .B(n3761), .Z(n935) );
  NOR U4033 ( .A(sum[5]), .B(n3236), .Z(n3764) );
  NOR U4034 ( .A(n3841), .B(o[165]), .Z(n3763) );
  NOR U4035 ( .A(n3764), .B(n3763), .Z(n936) );
  NOR U4036 ( .A(sum[4]), .B(n3236), .Z(n3766) );
  NOR U4037 ( .A(n3841), .B(o[164]), .Z(n3765) );
  NOR U4038 ( .A(n3766), .B(n3765), .Z(n937) );
  NOR U4039 ( .A(sum[3]), .B(n3236), .Z(n3768) );
  NOR U4040 ( .A(n3841), .B(o[163]), .Z(n3767) );
  NOR U4041 ( .A(n3768), .B(n3767), .Z(n938) );
  NOR U4042 ( .A(sum[2]), .B(n3236), .Z(n3770) );
  NOR U4043 ( .A(n3841), .B(o[162]), .Z(n3769) );
  NOR U4044 ( .A(n3770), .B(n3769), .Z(n939) );
  NOR U4045 ( .A(sum[1]), .B(n3236), .Z(n3772) );
  NOR U4046 ( .A(n3841), .B(o[161]), .Z(n3771) );
  NOR U4047 ( .A(n3772), .B(n3771), .Z(n940) );
  NOR U4048 ( .A(sum[0]), .B(n3236), .Z(n3774) );
  NOR U4049 ( .A(n3841), .B(o[160]), .Z(n3773) );
  NOR U4050 ( .A(n3774), .B(n3773), .Z(n941) );
  NOR U4051 ( .A(n3866), .B(n3775), .Z(n3838) );
  NOR U4052 ( .A(sum[31]), .B(n3235), .Z(n3777) );
  NOR U4053 ( .A(n3838), .B(o[95]), .Z(n3776) );
  NOR U4054 ( .A(n3777), .B(n3776), .Z(n942) );
  NOR U4055 ( .A(sum[30]), .B(n3235), .Z(n3779) );
  NOR U4056 ( .A(n3838), .B(o[94]), .Z(n3778) );
  NOR U4057 ( .A(n3779), .B(n3778), .Z(n943) );
  NOR U4058 ( .A(sum[29]), .B(n3235), .Z(n3781) );
  NOR U4059 ( .A(n3838), .B(o[93]), .Z(n3780) );
  NOR U4060 ( .A(n3781), .B(n3780), .Z(n944) );
  NOR U4061 ( .A(sum[28]), .B(n3235), .Z(n3783) );
  NOR U4062 ( .A(n3838), .B(o[92]), .Z(n3782) );
  NOR U4063 ( .A(n3783), .B(n3782), .Z(n945) );
  NOR U4064 ( .A(sum[27]), .B(n3235), .Z(n3785) );
  NOR U4065 ( .A(n3838), .B(o[91]), .Z(n3784) );
  NOR U4066 ( .A(n3785), .B(n3784), .Z(n946) );
  NOR U4067 ( .A(sum[26]), .B(n3235), .Z(n3787) );
  NOR U4068 ( .A(n3838), .B(o[90]), .Z(n3786) );
  NOR U4069 ( .A(n3787), .B(n3786), .Z(n947) );
  NOR U4070 ( .A(sum[25]), .B(n3235), .Z(n3789) );
  NOR U4071 ( .A(n3838), .B(o[89]), .Z(n3788) );
  NOR U4072 ( .A(n3789), .B(n3788), .Z(n948) );
  NOR U4073 ( .A(sum[24]), .B(n3235), .Z(n3791) );
  NOR U4074 ( .A(n3838), .B(o[88]), .Z(n3790) );
  NOR U4075 ( .A(n3791), .B(n3790), .Z(n949) );
  NOR U4076 ( .A(sum[23]), .B(n3235), .Z(n3793) );
  NOR U4077 ( .A(n3838), .B(o[87]), .Z(n3792) );
  NOR U4078 ( .A(n3793), .B(n3792), .Z(n950) );
  NOR U4079 ( .A(sum[22]), .B(n3235), .Z(n3795) );
  NOR U4080 ( .A(n3838), .B(o[86]), .Z(n3794) );
  NOR U4081 ( .A(n3795), .B(n3794), .Z(n951) );
  NOR U4082 ( .A(sum[21]), .B(n3235), .Z(n3797) );
  NOR U4083 ( .A(n3838), .B(o[85]), .Z(n3796) );
  NOR U4084 ( .A(n3797), .B(n3796), .Z(n952) );
  NOR U4085 ( .A(sum[20]), .B(n3235), .Z(n3799) );
  NOR U4086 ( .A(n3838), .B(o[84]), .Z(n3798) );
  NOR U4087 ( .A(n3799), .B(n3798), .Z(n953) );
  NOR U4088 ( .A(sum[19]), .B(n3235), .Z(n3801) );
  NOR U4089 ( .A(n3838), .B(o[83]), .Z(n3800) );
  NOR U4090 ( .A(n3801), .B(n3800), .Z(n954) );
  NOR U4091 ( .A(sum[18]), .B(n3235), .Z(n3803) );
  NOR U4092 ( .A(n3838), .B(o[82]), .Z(n3802) );
  NOR U4093 ( .A(n3803), .B(n3802), .Z(n955) );
  NOR U4094 ( .A(sum[17]), .B(n3235), .Z(n3805) );
  NOR U4095 ( .A(n3838), .B(o[81]), .Z(n3804) );
  NOR U4096 ( .A(n3805), .B(n3804), .Z(n956) );
  NOR U4097 ( .A(sum[16]), .B(n3235), .Z(n3807) );
  NOR U4098 ( .A(n3838), .B(o[80]), .Z(n3806) );
  NOR U4099 ( .A(n3807), .B(n3806), .Z(n957) );
  NOR U4100 ( .A(sum[15]), .B(n3235), .Z(n3809) );
  NOR U4101 ( .A(n3838), .B(o[79]), .Z(n3808) );
  NOR U4102 ( .A(n3809), .B(n3808), .Z(n958) );
  NOR U4103 ( .A(sum[14]), .B(n3235), .Z(n3811) );
  NOR U4104 ( .A(n3838), .B(o[78]), .Z(n3810) );
  NOR U4105 ( .A(n3811), .B(n3810), .Z(n959) );
  NOR U4106 ( .A(sum[13]), .B(n3235), .Z(n3813) );
  NOR U4107 ( .A(n3838), .B(o[77]), .Z(n3812) );
  NOR U4108 ( .A(n3813), .B(n3812), .Z(n960) );
  NOR U4109 ( .A(sum[12]), .B(n3235), .Z(n3815) );
  NOR U4110 ( .A(n3838), .B(o[76]), .Z(n3814) );
  NOR U4111 ( .A(n3815), .B(n3814), .Z(n961) );
  NOR U4112 ( .A(sum[11]), .B(n3235), .Z(n3817) );
  NOR U4113 ( .A(n3838), .B(o[75]), .Z(n3816) );
  NOR U4114 ( .A(n3817), .B(n3816), .Z(n962) );
  NOR U4115 ( .A(sum[10]), .B(n3235), .Z(n3819) );
  NOR U4116 ( .A(n3838), .B(o[74]), .Z(n3818) );
  NOR U4117 ( .A(n3819), .B(n3818), .Z(n963) );
  NOR U4118 ( .A(sum[9]), .B(n3235), .Z(n3821) );
  NOR U4119 ( .A(n3838), .B(o[73]), .Z(n3820) );
  NOR U4120 ( .A(n3821), .B(n3820), .Z(n964) );
  NOR U4121 ( .A(sum[8]), .B(n3235), .Z(n3823) );
  NOR U4122 ( .A(n3838), .B(o[72]), .Z(n3822) );
  NOR U4123 ( .A(n3823), .B(n3822), .Z(n965) );
  NOR U4124 ( .A(sum[7]), .B(n3235), .Z(n3825) );
  NOR U4125 ( .A(n3838), .B(o[71]), .Z(n3824) );
  NOR U4126 ( .A(n3825), .B(n3824), .Z(n966) );
  NOR U4127 ( .A(sum[6]), .B(n3235), .Z(n3827) );
  NOR U4128 ( .A(n3838), .B(o[70]), .Z(n3826) );
  NOR U4129 ( .A(n3827), .B(n3826), .Z(n967) );
  NOR U4130 ( .A(sum[5]), .B(n3235), .Z(n3829) );
  NOR U4131 ( .A(n3838), .B(o[69]), .Z(n3828) );
  NOR U4132 ( .A(n3829), .B(n3828), .Z(n968) );
  NOR U4133 ( .A(sum[4]), .B(n3235), .Z(n3831) );
  NOR U4134 ( .A(n3838), .B(o[68]), .Z(n3830) );
  NOR U4135 ( .A(n3831), .B(n3830), .Z(n969) );
  NOR U4136 ( .A(sum[3]), .B(n3235), .Z(n3833) );
  NOR U4137 ( .A(n3838), .B(o[67]), .Z(n3832) );
  NOR U4138 ( .A(n3833), .B(n3832), .Z(n970) );
  NOR U4139 ( .A(sum[2]), .B(n3235), .Z(n3835) );
  NOR U4140 ( .A(n3838), .B(o[66]), .Z(n3834) );
  NOR U4141 ( .A(n3835), .B(n3834), .Z(n971) );
  NOR U4142 ( .A(sum[1]), .B(n3235), .Z(n3837) );
  NOR U4143 ( .A(n3838), .B(o[65]), .Z(n3836) );
  NOR U4144 ( .A(n3837), .B(n3836), .Z(n972) );
  NOR U4145 ( .A(sum[0]), .B(n3235), .Z(n3840) );
  NOR U4146 ( .A(n3838), .B(o[64]), .Z(n3839) );
  NOR U4147 ( .A(n3840), .B(n3839), .Z(n973) );
  NOR U4148 ( .A(i[1]), .B(n3841), .Z(n3842) );
  IV U4149 ( .A(n3842), .Z(n974) );
  XOR U4150 ( .A(n3846), .B(n3917), .Z(n3844) );
  NOR U4151 ( .A(j[0]), .B(n3921), .Z(n3843) );
  NOR U4152 ( .A(n3844), .B(n3843), .Z(n975) );
  NOR U4153 ( .A(j[0]), .B(n3845), .Z(n3848) );
  XOR U4154 ( .A(n3921), .B(n3846), .Z(n3847) );
  NOR U4155 ( .A(n3848), .B(n3847), .Z(n976) );
  NOR U4156 ( .A(k[0]), .B(k[1]), .Z(n3857) );
  NOR U4157 ( .A(n9904), .B(n3857), .Z(n3850) );
  NOR U4158 ( .A(k[0]), .B(n3237), .Z(n3849) );
  NOR U4159 ( .A(n3850), .B(n3849), .Z(n977) );
  NOR U4160 ( .A(k[1]), .B(n3850), .Z(n3851) );
  NOR U4161 ( .A(n3852), .B(n3851), .Z(n978) );
  NOR U4162 ( .A(sum[31]), .B(n3237), .Z(n9752) );
  IV U4163 ( .A(x[245]), .Z(n3854) );
  IV U4164 ( .A(k[0]), .Z(n3918) );
  NOR U4165 ( .A(n3872), .B(n3918), .Z(n3853) );
  IV U4166 ( .A(n3853), .Z(n6057) );
  NOR U4167 ( .A(n3854), .B(n6057), .Z(n3897) );
  NOR U4168 ( .A(n3875), .B(n3918), .Z(n3855) );
  IV U4169 ( .A(n3855), .Z(n6051) );
  IV U4170 ( .A(x[149]), .Z(n3856) );
  NOR U4171 ( .A(n6051), .B(n3856), .Z(n3894) );
  IV U4172 ( .A(n3857), .Z(n3922) );
  NOR U4173 ( .A(n3922), .B(n3866), .Z(n3858) );
  IV U4174 ( .A(n3858), .Z(n6052) );
  IV U4175 ( .A(x[21]), .Z(n3859) );
  NOR U4176 ( .A(n6052), .B(n3859), .Z(n3891) );
  NOR U4177 ( .A(n3906), .B(n3866), .Z(n3860) );
  IV U4178 ( .A(n3860), .Z(n6059) );
  IV U4179 ( .A(x[85]), .Z(n3861) );
  NOR U4180 ( .A(n6059), .B(n3861), .Z(n3888) );
  NOR U4181 ( .A(n3875), .B(n3906), .Z(n3862) );
  IV U4182 ( .A(n3862), .Z(n6048) );
  IV U4183 ( .A(x[181]), .Z(n3863) );
  NOR U4184 ( .A(n6048), .B(n3863), .Z(n3885) );
  NOR U4185 ( .A(n3872), .B(n3922), .Z(n3864) );
  IV U4186 ( .A(n3864), .Z(n6055) );
  IV U4187 ( .A(x[213]), .Z(n3865) );
  NOR U4188 ( .A(n6055), .B(n3865), .Z(n3870) );
  NOR U4189 ( .A(n3918), .B(n3866), .Z(n3867) );
  IV U4190 ( .A(n3867), .Z(n6067) );
  IV U4191 ( .A(x[53]), .Z(n3868) );
  NOR U4192 ( .A(n6067), .B(n3868), .Z(n3869) );
  NOR U4193 ( .A(n3870), .B(n3869), .Z(n3871) );
  IV U4194 ( .A(n3871), .Z(n3882) );
  NOR U4195 ( .A(n3872), .B(n3906), .Z(n3873) );
  IV U4196 ( .A(n3873), .Z(n6065) );
  IV U4197 ( .A(x[277]), .Z(n3874) );
  NOR U4198 ( .A(n6065), .B(n3874), .Z(n3879) );
  NOR U4199 ( .A(n3875), .B(n3922), .Z(n3876) );
  IV U4200 ( .A(n3876), .Z(n6061) );
  IV U4201 ( .A(x[117]), .Z(n3877) );
  NOR U4202 ( .A(n6061), .B(n3877), .Z(n3878) );
  NOR U4203 ( .A(n3879), .B(n3878), .Z(n3880) );
  IV U4204 ( .A(n3880), .Z(n3881) );
  NOR U4205 ( .A(n3882), .B(n3881), .Z(n3883) );
  IV U4206 ( .A(n3883), .Z(n3884) );
  NOR U4207 ( .A(n3885), .B(n3884), .Z(n3886) );
  IV U4208 ( .A(n3886), .Z(n3887) );
  NOR U4209 ( .A(n3888), .B(n3887), .Z(n3889) );
  IV U4210 ( .A(n3889), .Z(n3890) );
  NOR U4211 ( .A(n3891), .B(n3890), .Z(n3892) );
  IV U4212 ( .A(n3892), .Z(n3893) );
  NOR U4213 ( .A(n3894), .B(n3893), .Z(n3895) );
  IV U4214 ( .A(n3895), .Z(n3896) );
  NOR U4215 ( .A(n3897), .B(n3896), .Z(n7772) );
  IV U4216 ( .A(y[264]), .Z(n3899) );
  NOR U4217 ( .A(n3906), .B(n3921), .Z(n3898) );
  IV U4218 ( .A(n3898), .Z(n6197) );
  NOR U4219 ( .A(n3899), .B(n6197), .Z(n3944) );
  NOR U4220 ( .A(n3918), .B(n3921), .Z(n3900) );
  IV U4221 ( .A(n3900), .Z(n6199) );
  IV U4222 ( .A(y[168]), .Z(n3901) );
  NOR U4223 ( .A(n6199), .B(n3901), .Z(n3941) );
  IV U4224 ( .A(y[40]), .Z(n3903) );
  NOR U4225 ( .A(n3922), .B(n3917), .Z(n3902) );
  IV U4226 ( .A(n3902), .Z(n6207) );
  NOR U4227 ( .A(n3903), .B(n6207), .Z(n3938) );
  NOR U4228 ( .A(n3906), .B(n3911), .Z(n3904) );
  IV U4229 ( .A(n3904), .Z(n6203) );
  IV U4230 ( .A(y[200]), .Z(n3905) );
  NOR U4231 ( .A(n6203), .B(n3905), .Z(n3935) );
  NOR U4232 ( .A(n3906), .B(n3917), .Z(n3907) );
  IV U4233 ( .A(n3907), .Z(n6205) );
  IV U4234 ( .A(y[232]), .Z(n3908) );
  NOR U4235 ( .A(n6205), .B(n3908), .Z(n3932) );
  NOR U4236 ( .A(n3922), .B(n3911), .Z(n3909) );
  IV U4237 ( .A(n3909), .Z(n6200) );
  IV U4238 ( .A(y[8]), .Z(n3910) );
  NOR U4239 ( .A(n6200), .B(n3910), .Z(n3915) );
  NOR U4240 ( .A(n3918), .B(n3911), .Z(n3912) );
  IV U4241 ( .A(n3912), .Z(n6209) );
  IV U4242 ( .A(y[104]), .Z(n3913) );
  NOR U4243 ( .A(n6209), .B(n3913), .Z(n3914) );
  NOR U4244 ( .A(n3915), .B(n3914), .Z(n3916) );
  IV U4245 ( .A(n3916), .Z(n3929) );
  NOR U4246 ( .A(n3918), .B(n3917), .Z(n3919) );
  IV U4247 ( .A(n3919), .Z(n6214) );
  IV U4248 ( .A(y[136]), .Z(n3920) );
  NOR U4249 ( .A(n6214), .B(n3920), .Z(n3926) );
  NOR U4250 ( .A(n3922), .B(n3921), .Z(n3923) );
  IV U4251 ( .A(n3923), .Z(n6216) );
  IV U4252 ( .A(y[72]), .Z(n3924) );
  NOR U4253 ( .A(n6216), .B(n3924), .Z(n3925) );
  NOR U4254 ( .A(n3926), .B(n3925), .Z(n3927) );
  IV U4255 ( .A(n3927), .Z(n3928) );
  NOR U4256 ( .A(n3929), .B(n3928), .Z(n3930) );
  IV U4257 ( .A(n3930), .Z(n3931) );
  NOR U4258 ( .A(n3932), .B(n3931), .Z(n3933) );
  IV U4259 ( .A(n3933), .Z(n3934) );
  NOR U4260 ( .A(n3935), .B(n3934), .Z(n3936) );
  IV U4261 ( .A(n3936), .Z(n3937) );
  NOR U4262 ( .A(n3938), .B(n3937), .Z(n3939) );
  IV U4263 ( .A(n3939), .Z(n3940) );
  NOR U4264 ( .A(n3941), .B(n3940), .Z(n3942) );
  IV U4265 ( .A(n3942), .Z(n3943) );
  NOR U4266 ( .A(n3944), .B(n3943), .Z(n9202) );
  NOR U4267 ( .A(n7772), .B(n9202), .Z(n5920) );
  IV U4268 ( .A(y[280]), .Z(n3945) );
  NOR U4269 ( .A(n3945), .B(n6197), .Z(n3976) );
  IV U4270 ( .A(y[152]), .Z(n3946) );
  NOR U4271 ( .A(n6214), .B(n3946), .Z(n3973) );
  IV U4272 ( .A(y[24]), .Z(n3947) );
  NOR U4273 ( .A(n3947), .B(n6200), .Z(n3970) );
  IV U4274 ( .A(y[216]), .Z(n3948) );
  NOR U4275 ( .A(n6203), .B(n3948), .Z(n3967) );
  IV U4276 ( .A(y[248]), .Z(n3949) );
  NOR U4277 ( .A(n6205), .B(n3949), .Z(n3964) );
  IV U4278 ( .A(y[88]), .Z(n3950) );
  NOR U4279 ( .A(n6216), .B(n3950), .Z(n3953) );
  IV U4280 ( .A(y[56]), .Z(n3951) );
  NOR U4281 ( .A(n6207), .B(n3951), .Z(n3952) );
  NOR U4282 ( .A(n3953), .B(n3952), .Z(n3954) );
  IV U4283 ( .A(n3954), .Z(n3961) );
  IV U4284 ( .A(y[184]), .Z(n3955) );
  NOR U4285 ( .A(n3955), .B(n6199), .Z(n3958) );
  IV U4286 ( .A(y[120]), .Z(n3956) );
  NOR U4287 ( .A(n3956), .B(n6209), .Z(n3957) );
  NOR U4288 ( .A(n3958), .B(n3957), .Z(n3959) );
  IV U4289 ( .A(n3959), .Z(n3960) );
  NOR U4290 ( .A(n3961), .B(n3960), .Z(n3962) );
  IV U4291 ( .A(n3962), .Z(n3963) );
  NOR U4292 ( .A(n3964), .B(n3963), .Z(n3965) );
  IV U4293 ( .A(n3965), .Z(n3966) );
  NOR U4294 ( .A(n3967), .B(n3966), .Z(n3968) );
  IV U4295 ( .A(n3968), .Z(n3969) );
  NOR U4296 ( .A(n3970), .B(n3969), .Z(n3971) );
  IV U4297 ( .A(n3971), .Z(n3972) );
  NOR U4298 ( .A(n3973), .B(n3972), .Z(n3974) );
  IV U4299 ( .A(n3974), .Z(n3975) );
  NOR U4300 ( .A(n3976), .B(n3975), .Z(n7167) );
  IV U4301 ( .A(x[165]), .Z(n3977) );
  NOR U4302 ( .A(n6048), .B(n3977), .Z(n4008) );
  IV U4303 ( .A(x[261]), .Z(n3978) );
  NOR U4304 ( .A(n6065), .B(n3978), .Z(n4005) );
  IV U4305 ( .A(x[5]), .Z(n3979) );
  NOR U4306 ( .A(n3979), .B(n6052), .Z(n4002) );
  IV U4307 ( .A(x[37]), .Z(n3980) );
  NOR U4308 ( .A(n6067), .B(n3980), .Z(n3999) );
  IV U4309 ( .A(x[229]), .Z(n3981) );
  NOR U4310 ( .A(n6057), .B(n3981), .Z(n3996) );
  IV U4311 ( .A(x[69]), .Z(n3982) );
  NOR U4312 ( .A(n6059), .B(n3982), .Z(n3985) );
  IV U4313 ( .A(x[197]), .Z(n3983) );
  NOR U4314 ( .A(n6055), .B(n3983), .Z(n3984) );
  NOR U4315 ( .A(n3985), .B(n3984), .Z(n3986) );
  IV U4316 ( .A(n3986), .Z(n3993) );
  IV U4317 ( .A(x[133]), .Z(n3987) );
  NOR U4318 ( .A(n6051), .B(n3987), .Z(n3990) );
  IV U4319 ( .A(x[101]), .Z(n3988) );
  NOR U4320 ( .A(n6061), .B(n3988), .Z(n3989) );
  NOR U4321 ( .A(n3990), .B(n3989), .Z(n3991) );
  IV U4322 ( .A(n3991), .Z(n3992) );
  NOR U4323 ( .A(n3993), .B(n3992), .Z(n3994) );
  IV U4324 ( .A(n3994), .Z(n3995) );
  NOR U4325 ( .A(n3996), .B(n3995), .Z(n3997) );
  IV U4326 ( .A(n3997), .Z(n3998) );
  NOR U4327 ( .A(n3999), .B(n3998), .Z(n4000) );
  IV U4328 ( .A(n4000), .Z(n4001) );
  NOR U4329 ( .A(n4002), .B(n4001), .Z(n4003) );
  IV U4330 ( .A(n4003), .Z(n4004) );
  NOR U4331 ( .A(n4005), .B(n4004), .Z(n4006) );
  IV U4332 ( .A(n4006), .Z(n4007) );
  NOR U4333 ( .A(n4008), .B(n4007), .Z(n9388) );
  NOR U4334 ( .A(n7167), .B(n9388), .Z(n4009) );
  IV U4335 ( .A(n4009), .Z(n5921) );
  XOR U4336 ( .A(n5920), .B(n5921), .Z(n5924) );
  IV U4337 ( .A(x[184]), .Z(n4010) );
  NOR U4338 ( .A(n6048), .B(n4010), .Z(n4041) );
  IV U4339 ( .A(x[152]), .Z(n4011) );
  NOR U4340 ( .A(n6051), .B(n4011), .Z(n4038) );
  IV U4341 ( .A(x[24]), .Z(n4012) );
  NOR U4342 ( .A(n4012), .B(n6052), .Z(n4035) );
  IV U4343 ( .A(x[56]), .Z(n4013) );
  NOR U4344 ( .A(n6067), .B(n4013), .Z(n4032) );
  IV U4345 ( .A(x[248]), .Z(n4014) );
  NOR U4346 ( .A(n6057), .B(n4014), .Z(n4029) );
  IV U4347 ( .A(x[216]), .Z(n4015) );
  NOR U4348 ( .A(n6055), .B(n4015), .Z(n4018) );
  IV U4349 ( .A(x[120]), .Z(n4016) );
  NOR U4350 ( .A(n6061), .B(n4016), .Z(n4017) );
  NOR U4351 ( .A(n4018), .B(n4017), .Z(n4019) );
  IV U4352 ( .A(n4019), .Z(n4026) );
  IV U4353 ( .A(x[88]), .Z(n4020) );
  NOR U4354 ( .A(n6059), .B(n4020), .Z(n4023) );
  IV U4355 ( .A(x[280]), .Z(n4021) );
  NOR U4356 ( .A(n4021), .B(n6065), .Z(n4022) );
  NOR U4357 ( .A(n4023), .B(n4022), .Z(n4024) );
  IV U4358 ( .A(n4024), .Z(n4025) );
  NOR U4359 ( .A(n4026), .B(n4025), .Z(n4027) );
  IV U4360 ( .A(n4027), .Z(n4028) );
  NOR U4361 ( .A(n4029), .B(n4028), .Z(n4030) );
  IV U4362 ( .A(n4030), .Z(n4031) );
  NOR U4363 ( .A(n4032), .B(n4031), .Z(n4033) );
  IV U4364 ( .A(n4033), .Z(n4034) );
  NOR U4365 ( .A(n4035), .B(n4034), .Z(n4036) );
  IV U4366 ( .A(n4036), .Z(n4037) );
  NOR U4367 ( .A(n4038), .B(n4037), .Z(n4039) );
  IV U4368 ( .A(n4039), .Z(n4040) );
  NOR U4369 ( .A(n4041), .B(n4040), .Z(n7225) );
  IV U4370 ( .A(y[261]), .Z(n4042) );
  NOR U4371 ( .A(n4042), .B(n6197), .Z(n4073) );
  IV U4372 ( .A(y[133]), .Z(n4043) );
  NOR U4373 ( .A(n6214), .B(n4043), .Z(n4070) );
  IV U4374 ( .A(y[5]), .Z(n4044) );
  NOR U4375 ( .A(n4044), .B(n6200), .Z(n4067) );
  IV U4376 ( .A(y[69]), .Z(n4045) );
  NOR U4377 ( .A(n6216), .B(n4045), .Z(n4064) );
  IV U4378 ( .A(y[229]), .Z(n4046) );
  NOR U4379 ( .A(n6205), .B(n4046), .Z(n4061) );
  IV U4380 ( .A(y[197]), .Z(n4047) );
  NOR U4381 ( .A(n6203), .B(n4047), .Z(n4050) );
  IV U4382 ( .A(y[37]), .Z(n4048) );
  NOR U4383 ( .A(n6207), .B(n4048), .Z(n4049) );
  NOR U4384 ( .A(n4050), .B(n4049), .Z(n4051) );
  IV U4385 ( .A(n4051), .Z(n4058) );
  IV U4386 ( .A(y[165]), .Z(n4052) );
  NOR U4387 ( .A(n4052), .B(n6199), .Z(n4055) );
  IV U4388 ( .A(y[101]), .Z(n4053) );
  NOR U4389 ( .A(n4053), .B(n6209), .Z(n4054) );
  NOR U4390 ( .A(n4055), .B(n4054), .Z(n4056) );
  IV U4391 ( .A(n4056), .Z(n4057) );
  NOR U4392 ( .A(n4058), .B(n4057), .Z(n4059) );
  IV U4393 ( .A(n4059), .Z(n4060) );
  NOR U4394 ( .A(n4061), .B(n4060), .Z(n4062) );
  IV U4395 ( .A(n4062), .Z(n4063) );
  NOR U4396 ( .A(n4064), .B(n4063), .Z(n4065) );
  IV U4397 ( .A(n4065), .Z(n4066) );
  NOR U4398 ( .A(n4067), .B(n4066), .Z(n4068) );
  IV U4399 ( .A(n4068), .Z(n4069) );
  NOR U4400 ( .A(n4070), .B(n4069), .Z(n4071) );
  IV U4401 ( .A(n4071), .Z(n4072) );
  NOR U4402 ( .A(n4073), .B(n4072), .Z(n9414) );
  NOR U4403 ( .A(n7225), .B(n9414), .Z(n4074) );
  IV U4404 ( .A(n4074), .Z(n5923) );
  XOR U4405 ( .A(n5924), .B(n5923), .Z(n5933) );
  IV U4406 ( .A(x[267]), .Z(n4075) );
  NOR U4407 ( .A(n4075), .B(n6065), .Z(n4106) );
  IV U4408 ( .A(x[139]), .Z(n4076) );
  NOR U4409 ( .A(n6051), .B(n4076), .Z(n4103) );
  IV U4410 ( .A(x[203]), .Z(n4077) );
  NOR U4411 ( .A(n4077), .B(n6055), .Z(n4100) );
  IV U4412 ( .A(x[75]), .Z(n4078) );
  NOR U4413 ( .A(n6059), .B(n4078), .Z(n4097) );
  IV U4414 ( .A(x[235]), .Z(n4079) );
  NOR U4415 ( .A(n6057), .B(n4079), .Z(n4094) );
  IV U4416 ( .A(x[11]), .Z(n4080) );
  NOR U4417 ( .A(n6052), .B(n4080), .Z(n4083) );
  IV U4418 ( .A(x[107]), .Z(n4081) );
  NOR U4419 ( .A(n6061), .B(n4081), .Z(n4082) );
  NOR U4420 ( .A(n4083), .B(n4082), .Z(n4084) );
  IV U4421 ( .A(n4084), .Z(n4091) );
  IV U4422 ( .A(x[43]), .Z(n4085) );
  NOR U4423 ( .A(n6067), .B(n4085), .Z(n4088) );
  IV U4424 ( .A(x[171]), .Z(n4086) );
  NOR U4425 ( .A(n4086), .B(n6048), .Z(n4087) );
  NOR U4426 ( .A(n4088), .B(n4087), .Z(n4089) );
  IV U4427 ( .A(n4089), .Z(n4090) );
  NOR U4428 ( .A(n4091), .B(n4090), .Z(n4092) );
  IV U4429 ( .A(n4092), .Z(n4093) );
  NOR U4430 ( .A(n4094), .B(n4093), .Z(n4095) );
  IV U4431 ( .A(n4095), .Z(n4096) );
  NOR U4432 ( .A(n4097), .B(n4096), .Z(n4098) );
  IV U4433 ( .A(n4098), .Z(n4099) );
  NOR U4434 ( .A(n4100), .B(n4099), .Z(n4101) );
  IV U4435 ( .A(n4101), .Z(n4102) );
  NOR U4436 ( .A(n4103), .B(n4102), .Z(n4104) );
  IV U4437 ( .A(n4104), .Z(n4105) );
  NOR U4438 ( .A(n4106), .B(n4105), .Z(n9034) );
  IV U4439 ( .A(y[242]), .Z(n4107) );
  NOR U4440 ( .A(n4107), .B(n6205), .Z(n4138) );
  IV U4441 ( .A(y[274]), .Z(n4108) );
  NOR U4442 ( .A(n6197), .B(n4108), .Z(n4135) );
  IV U4443 ( .A(y[82]), .Z(n4109) );
  NOR U4444 ( .A(n6216), .B(n4109), .Z(n4132) );
  IV U4445 ( .A(y[210]), .Z(n4110) );
  NOR U4446 ( .A(n6203), .B(n4110), .Z(n4129) );
  IV U4447 ( .A(y[50]), .Z(n4111) );
  NOR U4448 ( .A(n6207), .B(n4111), .Z(n4126) );
  IV U4449 ( .A(y[18]), .Z(n4112) );
  NOR U4450 ( .A(n6200), .B(n4112), .Z(n4115) );
  IV U4451 ( .A(y[114]), .Z(n4113) );
  NOR U4452 ( .A(n6209), .B(n4113), .Z(n4114) );
  NOR U4453 ( .A(n4115), .B(n4114), .Z(n4116) );
  IV U4454 ( .A(n4116), .Z(n4123) );
  IV U4455 ( .A(y[146]), .Z(n4117) );
  NOR U4456 ( .A(n6214), .B(n4117), .Z(n4120) );
  IV U4457 ( .A(y[178]), .Z(n4118) );
  NOR U4458 ( .A(n6199), .B(n4118), .Z(n4119) );
  NOR U4459 ( .A(n4120), .B(n4119), .Z(n4121) );
  IV U4460 ( .A(n4121), .Z(n4122) );
  NOR U4461 ( .A(n4123), .B(n4122), .Z(n4124) );
  IV U4462 ( .A(n4124), .Z(n4125) );
  NOR U4463 ( .A(n4126), .B(n4125), .Z(n4127) );
  IV U4464 ( .A(n4127), .Z(n4128) );
  NOR U4465 ( .A(n4129), .B(n4128), .Z(n4130) );
  IV U4466 ( .A(n4130), .Z(n4131) );
  NOR U4467 ( .A(n4132), .B(n4131), .Z(n4133) );
  IV U4468 ( .A(n4133), .Z(n4134) );
  NOR U4469 ( .A(n4135), .B(n4134), .Z(n4136) );
  IV U4470 ( .A(n4136), .Z(n4137) );
  NOR U4471 ( .A(n4138), .B(n4137), .Z(n8228) );
  NOR U4472 ( .A(n9034), .B(n8228), .Z(n5931) );
  IV U4473 ( .A(n5931), .Z(n8226) );
  IV U4474 ( .A(y[166]), .Z(n4139) );
  NOR U4475 ( .A(n6199), .B(n4139), .Z(n4170) );
  IV U4476 ( .A(y[134]), .Z(n4140) );
  NOR U4477 ( .A(n6214), .B(n4140), .Z(n4167) );
  IV U4478 ( .A(y[6]), .Z(n4141) );
  NOR U4479 ( .A(n6200), .B(n4141), .Z(n4164) );
  IV U4480 ( .A(y[198]), .Z(n4142) );
  NOR U4481 ( .A(n6203), .B(n4142), .Z(n4161) );
  IV U4482 ( .A(y[230]), .Z(n4143) );
  NOR U4483 ( .A(n6205), .B(n4143), .Z(n4158) );
  IV U4484 ( .A(y[70]), .Z(n4144) );
  NOR U4485 ( .A(n6216), .B(n4144), .Z(n4147) );
  IV U4486 ( .A(y[102]), .Z(n4145) );
  NOR U4487 ( .A(n6209), .B(n4145), .Z(n4146) );
  NOR U4488 ( .A(n4147), .B(n4146), .Z(n4148) );
  IV U4489 ( .A(n4148), .Z(n4155) );
  IV U4490 ( .A(y[38]), .Z(n4149) );
  NOR U4491 ( .A(n6207), .B(n4149), .Z(n4152) );
  IV U4492 ( .A(y[262]), .Z(n4150) );
  NOR U4493 ( .A(n6197), .B(n4150), .Z(n4151) );
  NOR U4494 ( .A(n4152), .B(n4151), .Z(n4153) );
  IV U4495 ( .A(n4153), .Z(n4154) );
  NOR U4496 ( .A(n4155), .B(n4154), .Z(n4156) );
  IV U4497 ( .A(n4156), .Z(n4157) );
  NOR U4498 ( .A(n4158), .B(n4157), .Z(n4159) );
  IV U4499 ( .A(n4159), .Z(n4160) );
  NOR U4500 ( .A(n4161), .B(n4160), .Z(n4162) );
  IV U4501 ( .A(n4162), .Z(n4163) );
  NOR U4502 ( .A(n4164), .B(n4163), .Z(n4165) );
  IV U4503 ( .A(n4165), .Z(n4166) );
  NOR U4504 ( .A(n4167), .B(n4166), .Z(n4168) );
  IV U4505 ( .A(n4168), .Z(n4169) );
  NOR U4506 ( .A(n4170), .B(n4169), .Z(n9429) );
  IV U4507 ( .A(x[247]), .Z(n4171) );
  NOR U4508 ( .A(n6057), .B(n4171), .Z(n4202) );
  IV U4509 ( .A(x[279]), .Z(n4172) );
  NOR U4510 ( .A(n6065), .B(n4172), .Z(n4199) );
  IV U4511 ( .A(x[23]), .Z(n4173) );
  NOR U4512 ( .A(n6052), .B(n4173), .Z(n4196) );
  IV U4513 ( .A(x[215]), .Z(n4174) );
  NOR U4514 ( .A(n6055), .B(n4174), .Z(n4193) );
  IV U4515 ( .A(x[183]), .Z(n4175) );
  NOR U4516 ( .A(n6048), .B(n4175), .Z(n4190) );
  IV U4517 ( .A(x[55]), .Z(n4176) );
  NOR U4518 ( .A(n6067), .B(n4176), .Z(n4179) );
  IV U4519 ( .A(x[119]), .Z(n4177) );
  NOR U4520 ( .A(n6061), .B(n4177), .Z(n4178) );
  NOR U4521 ( .A(n4179), .B(n4178), .Z(n4180) );
  IV U4522 ( .A(n4180), .Z(n4187) );
  IV U4523 ( .A(x[87]), .Z(n4181) );
  NOR U4524 ( .A(n6059), .B(n4181), .Z(n4184) );
  IV U4525 ( .A(x[151]), .Z(n4182) );
  NOR U4526 ( .A(n4182), .B(n6051), .Z(n4183) );
  NOR U4527 ( .A(n4184), .B(n4183), .Z(n4185) );
  IV U4528 ( .A(n4185), .Z(n4186) );
  NOR U4529 ( .A(n4187), .B(n4186), .Z(n4188) );
  IV U4530 ( .A(n4188), .Z(n4189) );
  NOR U4531 ( .A(n4190), .B(n4189), .Z(n4191) );
  IV U4532 ( .A(n4191), .Z(n4192) );
  NOR U4533 ( .A(n4193), .B(n4192), .Z(n4194) );
  IV U4534 ( .A(n4194), .Z(n4195) );
  NOR U4535 ( .A(n4196), .B(n4195), .Z(n4197) );
  IV U4536 ( .A(n4197), .Z(n4198) );
  NOR U4537 ( .A(n4199), .B(n4198), .Z(n4200) );
  IV U4538 ( .A(n4200), .Z(n4201) );
  NOR U4539 ( .A(n4202), .B(n4201), .Z(n7314) );
  NOR U4540 ( .A(n9429), .B(n7314), .Z(n5930) );
  XOR U4541 ( .A(n8226), .B(n5930), .Z(n5932) );
  XOR U4542 ( .A(n5933), .B(n5932), .Z(n4694) );
  IV U4543 ( .A(y[239]), .Z(n4203) );
  NOR U4544 ( .A(n4203), .B(n6205), .Z(n4234) );
  IV U4545 ( .A(y[143]), .Z(n4204) );
  NOR U4546 ( .A(n6214), .B(n4204), .Z(n4231) );
  IV U4547 ( .A(y[79]), .Z(n4205) );
  NOR U4548 ( .A(n6216), .B(n4205), .Z(n4228) );
  IV U4549 ( .A(y[207]), .Z(n4206) );
  NOR U4550 ( .A(n6203), .B(n4206), .Z(n4225) );
  IV U4551 ( .A(y[271]), .Z(n4207) );
  NOR U4552 ( .A(n6197), .B(n4207), .Z(n4222) );
  IV U4553 ( .A(y[15]), .Z(n4208) );
  NOR U4554 ( .A(n6200), .B(n4208), .Z(n4211) );
  IV U4555 ( .A(y[111]), .Z(n4209) );
  NOR U4556 ( .A(n6209), .B(n4209), .Z(n4210) );
  NOR U4557 ( .A(n4211), .B(n4210), .Z(n4212) );
  IV U4558 ( .A(n4212), .Z(n4219) );
  IV U4559 ( .A(y[175]), .Z(n4213) );
  NOR U4560 ( .A(n6199), .B(n4213), .Z(n4216) );
  IV U4561 ( .A(y[47]), .Z(n4214) );
  NOR U4562 ( .A(n6207), .B(n4214), .Z(n4215) );
  NOR U4563 ( .A(n4216), .B(n4215), .Z(n4217) );
  IV U4564 ( .A(n4217), .Z(n4218) );
  NOR U4565 ( .A(n4219), .B(n4218), .Z(n4220) );
  IV U4566 ( .A(n4220), .Z(n4221) );
  NOR U4567 ( .A(n4222), .B(n4221), .Z(n4223) );
  IV U4568 ( .A(n4223), .Z(n4224) );
  NOR U4569 ( .A(n4225), .B(n4224), .Z(n4226) );
  IV U4570 ( .A(n4226), .Z(n4227) );
  NOR U4571 ( .A(n4228), .B(n4227), .Z(n4229) );
  IV U4572 ( .A(n4229), .Z(n4230) );
  NOR U4573 ( .A(n4231), .B(n4230), .Z(n4232) );
  IV U4574 ( .A(n4232), .Z(n4233) );
  NOR U4575 ( .A(n4234), .B(n4233), .Z(n8582) );
  IV U4576 ( .A(x[174]), .Z(n4235) );
  NOR U4577 ( .A(n6048), .B(n4235), .Z(n4266) );
  IV U4578 ( .A(x[270]), .Z(n4236) );
  NOR U4579 ( .A(n6065), .B(n4236), .Z(n4263) );
  IV U4580 ( .A(x[206]), .Z(n4237) );
  NOR U4581 ( .A(n4237), .B(n6055), .Z(n4260) );
  IV U4582 ( .A(x[78]), .Z(n4238) );
  NOR U4583 ( .A(n6059), .B(n4238), .Z(n4257) );
  IV U4584 ( .A(x[238]), .Z(n4239) );
  NOR U4585 ( .A(n6057), .B(n4239), .Z(n4254) );
  IV U4586 ( .A(x[14]), .Z(n4240) );
  NOR U4587 ( .A(n6052), .B(n4240), .Z(n4243) );
  IV U4588 ( .A(x[110]), .Z(n4241) );
  NOR U4589 ( .A(n6061), .B(n4241), .Z(n4242) );
  NOR U4590 ( .A(n4243), .B(n4242), .Z(n4244) );
  IV U4591 ( .A(n4244), .Z(n4251) );
  IV U4592 ( .A(x[142]), .Z(n4245) );
  NOR U4593 ( .A(n4245), .B(n6051), .Z(n4248) );
  IV U4594 ( .A(x[46]), .Z(n4246) );
  NOR U4595 ( .A(n4246), .B(n6067), .Z(n4247) );
  NOR U4596 ( .A(n4248), .B(n4247), .Z(n4249) );
  IV U4597 ( .A(n4249), .Z(n4250) );
  NOR U4598 ( .A(n4251), .B(n4250), .Z(n4252) );
  IV U4599 ( .A(n4252), .Z(n4253) );
  NOR U4600 ( .A(n4254), .B(n4253), .Z(n4255) );
  IV U4601 ( .A(n4255), .Z(n4256) );
  NOR U4602 ( .A(n4257), .B(n4256), .Z(n4258) );
  IV U4603 ( .A(n4258), .Z(n4259) );
  NOR U4604 ( .A(n4260), .B(n4259), .Z(n4261) );
  IV U4605 ( .A(n4261), .Z(n4262) );
  NOR U4606 ( .A(n4263), .B(n4262), .Z(n4264) );
  IV U4607 ( .A(n4264), .Z(n4265) );
  NOR U4608 ( .A(n4266), .B(n4265), .Z(n8729) );
  NOR U4609 ( .A(n8582), .B(n8729), .Z(n6012) );
  IV U4610 ( .A(x[257]), .Z(n4267) );
  NOR U4611 ( .A(n6065), .B(n4267), .Z(n4298) );
  IV U4612 ( .A(x[129]), .Z(n4268) );
  NOR U4613 ( .A(n6051), .B(n4268), .Z(n4295) );
  IV U4614 ( .A(x[33]), .Z(n4269) );
  NOR U4615 ( .A(n4269), .B(n6067), .Z(n4292) );
  IV U4616 ( .A(x[193]), .Z(n4270) );
  NOR U4617 ( .A(n6055), .B(n4270), .Z(n4289) );
  IV U4618 ( .A(x[225]), .Z(n4271) );
  NOR U4619 ( .A(n6057), .B(n4271), .Z(n4286) );
  IV U4620 ( .A(x[1]), .Z(n4272) );
  NOR U4621 ( .A(n6052), .B(n4272), .Z(n4275) );
  IV U4622 ( .A(x[97]), .Z(n4273) );
  NOR U4623 ( .A(n6061), .B(n4273), .Z(n4274) );
  NOR U4624 ( .A(n4275), .B(n4274), .Z(n4276) );
  IV U4625 ( .A(n4276), .Z(n4283) );
  IV U4626 ( .A(x[65]), .Z(n4277) );
  NOR U4627 ( .A(n6059), .B(n4277), .Z(n4280) );
  IV U4628 ( .A(x[161]), .Z(n4278) );
  NOR U4629 ( .A(n4278), .B(n6048), .Z(n4279) );
  NOR U4630 ( .A(n4280), .B(n4279), .Z(n4281) );
  IV U4631 ( .A(n4281), .Z(n4282) );
  NOR U4632 ( .A(n4283), .B(n4282), .Z(n4284) );
  IV U4633 ( .A(n4284), .Z(n4285) );
  NOR U4634 ( .A(n4286), .B(n4285), .Z(n4287) );
  IV U4635 ( .A(n4287), .Z(n4288) );
  NOR U4636 ( .A(n4289), .B(n4288), .Z(n4290) );
  IV U4637 ( .A(n4290), .Z(n4291) );
  NOR U4638 ( .A(n4292), .B(n4291), .Z(n4293) );
  IV U4639 ( .A(n4293), .Z(n4294) );
  NOR U4640 ( .A(n4295), .B(n4294), .Z(n4296) );
  IV U4641 ( .A(n4296), .Z(n4297) );
  NOR U4642 ( .A(n4298), .B(n4297), .Z(n9599) );
  IV U4643 ( .A(y[252]), .Z(n4299) );
  NOR U4644 ( .A(n6205), .B(n4299), .Z(n4330) );
  IV U4645 ( .A(y[284]), .Z(n4300) );
  NOR U4646 ( .A(n6197), .B(n4300), .Z(n4327) );
  IV U4647 ( .A(y[124]), .Z(n4301) );
  NOR U4648 ( .A(n6209), .B(n4301), .Z(n4324) );
  IV U4649 ( .A(y[60]), .Z(n4302) );
  NOR U4650 ( .A(n6207), .B(n4302), .Z(n4321) );
  IV U4651 ( .A(y[188]), .Z(n4303) );
  NOR U4652 ( .A(n6199), .B(n4303), .Z(n4318) );
  IV U4653 ( .A(y[220]), .Z(n4304) );
  NOR U4654 ( .A(n6203), .B(n4304), .Z(n4307) );
  IV U4655 ( .A(y[92]), .Z(n4305) );
  NOR U4656 ( .A(n6216), .B(n4305), .Z(n4306) );
  NOR U4657 ( .A(n4307), .B(n4306), .Z(n4308) );
  IV U4658 ( .A(n4308), .Z(n4315) );
  IV U4659 ( .A(y[156]), .Z(n4309) );
  NOR U4660 ( .A(n6214), .B(n4309), .Z(n4312) );
  IV U4661 ( .A(y[28]), .Z(n4310) );
  NOR U4662 ( .A(n6200), .B(n4310), .Z(n4311) );
  NOR U4663 ( .A(n4312), .B(n4311), .Z(n4313) );
  IV U4664 ( .A(n4313), .Z(n4314) );
  NOR U4665 ( .A(n4315), .B(n4314), .Z(n4316) );
  IV U4666 ( .A(n4316), .Z(n4317) );
  NOR U4667 ( .A(n4318), .B(n4317), .Z(n4319) );
  IV U4668 ( .A(n4319), .Z(n4320) );
  NOR U4669 ( .A(n4321), .B(n4320), .Z(n4322) );
  IV U4670 ( .A(n4322), .Z(n4323) );
  NOR U4671 ( .A(n4324), .B(n4323), .Z(n4325) );
  IV U4672 ( .A(n4325), .Z(n4326) );
  NOR U4673 ( .A(n4327), .B(n4326), .Z(n4328) );
  IV U4674 ( .A(n4328), .Z(n4329) );
  NOR U4675 ( .A(n4330), .B(n4329), .Z(n6368) );
  NOR U4676 ( .A(n9599), .B(n6368), .Z(n4331) );
  IV U4677 ( .A(n4331), .Z(n6013) );
  XOR U4678 ( .A(n6012), .B(n6013), .Z(n6016) );
  IV U4679 ( .A(x[250]), .Z(n4332) );
  NOR U4680 ( .A(n4332), .B(n6057), .Z(n4363) );
  IV U4681 ( .A(x[186]), .Z(n4333) );
  NOR U4682 ( .A(n6048), .B(n4333), .Z(n4360) );
  IV U4683 ( .A(x[122]), .Z(n4334) );
  NOR U4684 ( .A(n4334), .B(n6061), .Z(n4357) );
  IV U4685 ( .A(x[90]), .Z(n4335) );
  NOR U4686 ( .A(n6059), .B(n4335), .Z(n4354) );
  IV U4687 ( .A(x[282]), .Z(n4336) );
  NOR U4688 ( .A(n6065), .B(n4336), .Z(n4351) );
  IV U4689 ( .A(x[218]), .Z(n4337) );
  NOR U4690 ( .A(n6055), .B(n4337), .Z(n4340) );
  IV U4691 ( .A(x[58]), .Z(n4338) );
  NOR U4692 ( .A(n6067), .B(n4338), .Z(n4339) );
  NOR U4693 ( .A(n4340), .B(n4339), .Z(n4341) );
  IV U4694 ( .A(n4341), .Z(n4348) );
  IV U4695 ( .A(x[154]), .Z(n4342) );
  NOR U4696 ( .A(n6051), .B(n4342), .Z(n4345) );
  IV U4697 ( .A(x[26]), .Z(n4343) );
  NOR U4698 ( .A(n6052), .B(n4343), .Z(n4344) );
  NOR U4699 ( .A(n4345), .B(n4344), .Z(n4346) );
  IV U4700 ( .A(n4346), .Z(n4347) );
  NOR U4701 ( .A(n4348), .B(n4347), .Z(n4349) );
  IV U4702 ( .A(n4349), .Z(n4350) );
  NOR U4703 ( .A(n4351), .B(n4350), .Z(n4352) );
  IV U4704 ( .A(n4352), .Z(n4353) );
  NOR U4705 ( .A(n4354), .B(n4353), .Z(n4355) );
  IV U4706 ( .A(n4355), .Z(n4356) );
  NOR U4707 ( .A(n4357), .B(n4356), .Z(n4358) );
  IV U4708 ( .A(n4358), .Z(n4359) );
  NOR U4709 ( .A(n4360), .B(n4359), .Z(n4361) );
  IV U4710 ( .A(n4361), .Z(n4362) );
  NOR U4711 ( .A(n4363), .B(n4362), .Z(n6728) );
  IV U4712 ( .A(y[227]), .Z(n4364) );
  NOR U4713 ( .A(n4364), .B(n6205), .Z(n4395) );
  IV U4714 ( .A(y[259]), .Z(n4365) );
  NOR U4715 ( .A(n6197), .B(n4365), .Z(n4392) );
  IV U4716 ( .A(y[99]), .Z(n4366) );
  NOR U4717 ( .A(n4366), .B(n6209), .Z(n4389) );
  IV U4718 ( .A(y[67]), .Z(n4367) );
  NOR U4719 ( .A(n6216), .B(n4367), .Z(n4386) );
  IV U4720 ( .A(y[163]), .Z(n4368) );
  NOR U4721 ( .A(n6199), .B(n4368), .Z(n4383) );
  IV U4722 ( .A(y[195]), .Z(n4369) );
  NOR U4723 ( .A(n6203), .B(n4369), .Z(n4372) );
  IV U4724 ( .A(y[35]), .Z(n4370) );
  NOR U4725 ( .A(n6207), .B(n4370), .Z(n4371) );
  NOR U4726 ( .A(n4372), .B(n4371), .Z(n4373) );
  IV U4727 ( .A(n4373), .Z(n4380) );
  IV U4728 ( .A(y[131]), .Z(n4374) );
  NOR U4729 ( .A(n6214), .B(n4374), .Z(n4377) );
  IV U4730 ( .A(y[3]), .Z(n4375) );
  NOR U4731 ( .A(n6200), .B(n4375), .Z(n4376) );
  NOR U4732 ( .A(n4377), .B(n4376), .Z(n4378) );
  IV U4733 ( .A(n4378), .Z(n4379) );
  NOR U4734 ( .A(n4380), .B(n4379), .Z(n4381) );
  IV U4735 ( .A(n4381), .Z(n4382) );
  NOR U4736 ( .A(n4383), .B(n4382), .Z(n4384) );
  IV U4737 ( .A(n4384), .Z(n4385) );
  NOR U4738 ( .A(n4386), .B(n4385), .Z(n4387) );
  IV U4739 ( .A(n4387), .Z(n4388) );
  NOR U4740 ( .A(n4389), .B(n4388), .Z(n4390) );
  IV U4741 ( .A(n4390), .Z(n4391) );
  NOR U4742 ( .A(n4392), .B(n4391), .Z(n4393) );
  IV U4743 ( .A(n4393), .Z(n4394) );
  NOR U4744 ( .A(n4395), .B(n4394), .Z(n9490) );
  NOR U4745 ( .A(n6728), .B(n9490), .Z(n4396) );
  IV U4746 ( .A(n4396), .Z(n6015) );
  XOR U4747 ( .A(n6016), .B(n6015), .Z(n6348) );
  IV U4748 ( .A(x[240]), .Z(n4397) );
  NOR U4749 ( .A(n4397), .B(n6057), .Z(n4428) );
  IV U4750 ( .A(x[176]), .Z(n4398) );
  NOR U4751 ( .A(n6048), .B(n4398), .Z(n4425) );
  IV U4752 ( .A(x[16]), .Z(n4399) );
  NOR U4753 ( .A(n6052), .B(n4399), .Z(n4422) );
  IV U4754 ( .A(x[80]), .Z(n4400) );
  NOR U4755 ( .A(n6059), .B(n4400), .Z(n4419) );
  IV U4756 ( .A(x[208]), .Z(n4401) );
  NOR U4757 ( .A(n6055), .B(n4401), .Z(n4416) );
  IV U4758 ( .A(x[48]), .Z(n4402) );
  NOR U4759 ( .A(n6067), .B(n4402), .Z(n4405) );
  IV U4760 ( .A(x[112]), .Z(n4403) );
  NOR U4761 ( .A(n6061), .B(n4403), .Z(n4404) );
  NOR U4762 ( .A(n4405), .B(n4404), .Z(n4406) );
  IV U4763 ( .A(n4406), .Z(n4413) );
  IV U4764 ( .A(x[144]), .Z(n4407) );
  NOR U4765 ( .A(n6051), .B(n4407), .Z(n4410) );
  IV U4766 ( .A(x[272]), .Z(n4408) );
  NOR U4767 ( .A(n6065), .B(n4408), .Z(n4409) );
  NOR U4768 ( .A(n4410), .B(n4409), .Z(n4411) );
  IV U4769 ( .A(n4411), .Z(n4412) );
  NOR U4770 ( .A(n4413), .B(n4412), .Z(n4414) );
  IV U4771 ( .A(n4414), .Z(n4415) );
  NOR U4772 ( .A(n4416), .B(n4415), .Z(n4417) );
  IV U4773 ( .A(n4417), .Z(n4418) );
  NOR U4774 ( .A(n4419), .B(n4418), .Z(n4420) );
  IV U4775 ( .A(n4420), .Z(n4421) );
  NOR U4776 ( .A(n4422), .B(n4421), .Z(n4423) );
  IV U4777 ( .A(n4423), .Z(n4424) );
  NOR U4778 ( .A(n4425), .B(n4424), .Z(n4426) );
  IV U4779 ( .A(n4426), .Z(n4427) );
  NOR U4780 ( .A(n4428), .B(n4427), .Z(n8499) );
  IV U4781 ( .A(y[269]), .Z(n4429) );
  NOR U4782 ( .A(n6197), .B(n4429), .Z(n4460) );
  IV U4783 ( .A(y[173]), .Z(n4430) );
  NOR U4784 ( .A(n6199), .B(n4430), .Z(n4457) );
  IV U4785 ( .A(y[45]), .Z(n4431) );
  NOR U4786 ( .A(n4431), .B(n6207), .Z(n4454) );
  IV U4787 ( .A(y[13]), .Z(n4432) );
  NOR U4788 ( .A(n6200), .B(n4432), .Z(n4451) );
  IV U4789 ( .A(y[237]), .Z(n4433) );
  NOR U4790 ( .A(n6205), .B(n4433), .Z(n4448) );
  IV U4791 ( .A(y[77]), .Z(n4434) );
  NOR U4792 ( .A(n6216), .B(n4434), .Z(n4437) );
  IV U4793 ( .A(y[109]), .Z(n4435) );
  NOR U4794 ( .A(n6209), .B(n4435), .Z(n4436) );
  NOR U4795 ( .A(n4437), .B(n4436), .Z(n4438) );
  IV U4796 ( .A(n4438), .Z(n4445) );
  IV U4797 ( .A(y[205]), .Z(n4439) );
  NOR U4798 ( .A(n6203), .B(n4439), .Z(n4442) );
  IV U4799 ( .A(y[141]), .Z(n4440) );
  NOR U4800 ( .A(n4440), .B(n6214), .Z(n4441) );
  NOR U4801 ( .A(n4442), .B(n4441), .Z(n4443) );
  IV U4802 ( .A(n4443), .Z(n4444) );
  NOR U4803 ( .A(n4445), .B(n4444), .Z(n4446) );
  IV U4804 ( .A(n4446), .Z(n4447) );
  NOR U4805 ( .A(n4448), .B(n4447), .Z(n4449) );
  IV U4806 ( .A(n4449), .Z(n4450) );
  NOR U4807 ( .A(n4451), .B(n4450), .Z(n4452) );
  IV U4808 ( .A(n4452), .Z(n4453) );
  NOR U4809 ( .A(n4454), .B(n4453), .Z(n4455) );
  IV U4810 ( .A(n4455), .Z(n4456) );
  NOR U4811 ( .A(n4457), .B(n4456), .Z(n4458) );
  IV U4812 ( .A(n4458), .Z(n4459) );
  NOR U4813 ( .A(n4460), .B(n4459), .Z(n8862) );
  NOR U4814 ( .A(n8499), .B(n8862), .Z(n6346) );
  IV U4815 ( .A(y[187]), .Z(n4461) );
  NOR U4816 ( .A(n4461), .B(n6199), .Z(n4492) );
  IV U4817 ( .A(y[155]), .Z(n4462) );
  NOR U4818 ( .A(n6214), .B(n4462), .Z(n4489) );
  IV U4819 ( .A(y[27]), .Z(n4463) );
  NOR U4820 ( .A(n6200), .B(n4463), .Z(n4486) );
  IV U4821 ( .A(y[219]), .Z(n4464) );
  NOR U4822 ( .A(n6203), .B(n4464), .Z(n4483) );
  IV U4823 ( .A(y[251]), .Z(n4465) );
  NOR U4824 ( .A(n6205), .B(n4465), .Z(n4480) );
  IV U4825 ( .A(y[91]), .Z(n4466) );
  NOR U4826 ( .A(n6216), .B(n4466), .Z(n4469) );
  IV U4827 ( .A(y[59]), .Z(n4467) );
  NOR U4828 ( .A(n6207), .B(n4467), .Z(n4468) );
  NOR U4829 ( .A(n4469), .B(n4468), .Z(n4470) );
  IV U4830 ( .A(n4470), .Z(n4477) );
  IV U4831 ( .A(y[123]), .Z(n4471) );
  NOR U4832 ( .A(n6209), .B(n4471), .Z(n4474) );
  IV U4833 ( .A(y[283]), .Z(n4472) );
  NOR U4834 ( .A(n4472), .B(n6197), .Z(n4473) );
  NOR U4835 ( .A(n4474), .B(n4473), .Z(n4475) );
  IV U4836 ( .A(n4475), .Z(n4476) );
  NOR U4837 ( .A(n4477), .B(n4476), .Z(n4478) );
  IV U4838 ( .A(n4478), .Z(n4479) );
  NOR U4839 ( .A(n4480), .B(n4479), .Z(n4481) );
  IV U4840 ( .A(n4481), .Z(n4482) );
  NOR U4841 ( .A(n4483), .B(n4482), .Z(n4484) );
  IV U4842 ( .A(n4484), .Z(n4485) );
  NOR U4843 ( .A(n4486), .B(n4485), .Z(n4487) );
  IV U4844 ( .A(n4487), .Z(n4488) );
  NOR U4845 ( .A(n4489), .B(n4488), .Z(n4490) );
  IV U4846 ( .A(n4490), .Z(n4491) );
  NOR U4847 ( .A(n4492), .B(n4491), .Z(n6579) );
  IV U4848 ( .A(x[162]), .Z(n4493) );
  NOR U4849 ( .A(n6048), .B(n4493), .Z(n4524) );
  IV U4850 ( .A(x[130]), .Z(n4494) );
  NOR U4851 ( .A(n6051), .B(n4494), .Z(n4521) );
  IV U4852 ( .A(x[194]), .Z(n4495) );
  NOR U4853 ( .A(n6055), .B(n4495), .Z(n4518) );
  IV U4854 ( .A(x[66]), .Z(n4496) );
  NOR U4855 ( .A(n6059), .B(n4496), .Z(n4515) );
  IV U4856 ( .A(x[226]), .Z(n4497) );
  NOR U4857 ( .A(n6057), .B(n4497), .Z(n4512) );
  IV U4858 ( .A(x[34]), .Z(n4498) );
  NOR U4859 ( .A(n6067), .B(n4498), .Z(n4501) );
  IV U4860 ( .A(x[98]), .Z(n4499) );
  NOR U4861 ( .A(n6061), .B(n4499), .Z(n4500) );
  NOR U4862 ( .A(n4501), .B(n4500), .Z(n4502) );
  IV U4863 ( .A(n4502), .Z(n4509) );
  IV U4864 ( .A(x[258]), .Z(n4503) );
  NOR U4865 ( .A(n6065), .B(n4503), .Z(n4506) );
  IV U4866 ( .A(x[2]), .Z(n4504) );
  NOR U4867 ( .A(n6052), .B(n4504), .Z(n4505) );
  NOR U4868 ( .A(n4506), .B(n4505), .Z(n4507) );
  IV U4869 ( .A(n4507), .Z(n4508) );
  NOR U4870 ( .A(n4509), .B(n4508), .Z(n4510) );
  IV U4871 ( .A(n4510), .Z(n4511) );
  NOR U4872 ( .A(n4512), .B(n4511), .Z(n4513) );
  IV U4873 ( .A(n4513), .Z(n4514) );
  NOR U4874 ( .A(n4515), .B(n4514), .Z(n4516) );
  IV U4875 ( .A(n4516), .Z(n4517) );
  NOR U4876 ( .A(n4518), .B(n4517), .Z(n4519) );
  IV U4877 ( .A(n4519), .Z(n4520) );
  NOR U4878 ( .A(n4521), .B(n4520), .Z(n4522) );
  IV U4879 ( .A(n4522), .Z(n4523) );
  NOR U4880 ( .A(n4524), .B(n4523), .Z(n9584) );
  NOR U4881 ( .A(n6579), .B(n9584), .Z(n6345) );
  XOR U4882 ( .A(n6346), .B(n6345), .Z(n4525) );
  IV U4883 ( .A(n4525), .Z(n6347) );
  XOR U4884 ( .A(n6348), .B(n6347), .Z(n4693) );
  NOR U4885 ( .A(n4694), .B(n4693), .Z(n4697) );
  IV U4886 ( .A(y[244]), .Z(n4526) );
  NOR U4887 ( .A(n4526), .B(n6205), .Z(n4557) );
  IV U4888 ( .A(y[276]), .Z(n4527) );
  NOR U4889 ( .A(n6197), .B(n4527), .Z(n4554) );
  IV U4890 ( .A(y[20]), .Z(n4528) );
  NOR U4891 ( .A(n4528), .B(n6200), .Z(n4551) );
  IV U4892 ( .A(y[84]), .Z(n4529) );
  NOR U4893 ( .A(n6216), .B(n4529), .Z(n4548) );
  IV U4894 ( .A(y[180]), .Z(n4530) );
  NOR U4895 ( .A(n4530), .B(n6199), .Z(n4545) );
  IV U4896 ( .A(y[52]), .Z(n4531) );
  NOR U4897 ( .A(n6207), .B(n4531), .Z(n4534) );
  IV U4898 ( .A(y[116]), .Z(n4532) );
  NOR U4899 ( .A(n6209), .B(n4532), .Z(n4533) );
  NOR U4900 ( .A(n4534), .B(n4533), .Z(n4535) );
  IV U4901 ( .A(n4535), .Z(n4542) );
  IV U4902 ( .A(y[212]), .Z(n4536) );
  NOR U4903 ( .A(n6203), .B(n4536), .Z(n4539) );
  IV U4904 ( .A(y[148]), .Z(n4537) );
  NOR U4905 ( .A(n4537), .B(n6214), .Z(n4538) );
  NOR U4906 ( .A(n4539), .B(n4538), .Z(n4540) );
  IV U4907 ( .A(n4540), .Z(n4541) );
  NOR U4908 ( .A(n4542), .B(n4541), .Z(n4543) );
  IV U4909 ( .A(n4543), .Z(n4544) );
  NOR U4910 ( .A(n4545), .B(n4544), .Z(n4546) );
  IV U4911 ( .A(n4546), .Z(n4547) );
  NOR U4912 ( .A(n4548), .B(n4547), .Z(n4549) );
  IV U4913 ( .A(n4549), .Z(n4550) );
  NOR U4914 ( .A(n4551), .B(n4550), .Z(n4552) );
  IV U4915 ( .A(n4552), .Z(n4553) );
  NOR U4916 ( .A(n4554), .B(n4553), .Z(n4555) );
  IV U4917 ( .A(n4555), .Z(n4556) );
  NOR U4918 ( .A(n4557), .B(n4556), .Z(n7891) );
  IV U4919 ( .A(x[232]), .Z(n4558) );
  NOR U4920 ( .A(n6057), .B(n4558), .Z(n4589) );
  IV U4921 ( .A(x[168]), .Z(n4559) );
  NOR U4922 ( .A(n6048), .B(n4559), .Z(n4586) );
  IV U4923 ( .A(x[104]), .Z(n4560) );
  NOR U4924 ( .A(n4560), .B(n6061), .Z(n4583) );
  IV U4925 ( .A(x[72]), .Z(n4561) );
  NOR U4926 ( .A(n6059), .B(n4561), .Z(n4580) );
  IV U4927 ( .A(x[264]), .Z(n4562) );
  NOR U4928 ( .A(n6065), .B(n4562), .Z(n4577) );
  IV U4929 ( .A(x[200]), .Z(n4563) );
  NOR U4930 ( .A(n6055), .B(n4563), .Z(n4566) );
  IV U4931 ( .A(x[40]), .Z(n4564) );
  NOR U4932 ( .A(n6067), .B(n4564), .Z(n4565) );
  NOR U4933 ( .A(n4566), .B(n4565), .Z(n4567) );
  IV U4934 ( .A(n4567), .Z(n4574) );
  IV U4935 ( .A(x[136]), .Z(n4568) );
  NOR U4936 ( .A(n6051), .B(n4568), .Z(n4571) );
  IV U4937 ( .A(x[8]), .Z(n4569) );
  NOR U4938 ( .A(n6052), .B(n4569), .Z(n4570) );
  NOR U4939 ( .A(n4571), .B(n4570), .Z(n4572) );
  IV U4940 ( .A(n4572), .Z(n4573) );
  NOR U4941 ( .A(n4574), .B(n4573), .Z(n4575) );
  IV U4942 ( .A(n4575), .Z(n4576) );
  NOR U4943 ( .A(n4577), .B(n4576), .Z(n4578) );
  IV U4944 ( .A(n4578), .Z(n4579) );
  NOR U4945 ( .A(n4580), .B(n4579), .Z(n4581) );
  IV U4946 ( .A(n4581), .Z(n4582) );
  NOR U4947 ( .A(n4583), .B(n4582), .Z(n4584) );
  IV U4948 ( .A(n4584), .Z(n4585) );
  NOR U4949 ( .A(n4586), .B(n4585), .Z(n4587) );
  IV U4950 ( .A(n4587), .Z(n4588) );
  NOR U4951 ( .A(n4589), .B(n4588), .Z(n9316) );
  NOR U4952 ( .A(n7891), .B(n9316), .Z(n4590) );
  IV U4953 ( .A(n4590), .Z(n4625) );
  IV U4954 ( .A(x[246]), .Z(n4591) );
  NOR U4955 ( .A(n6057), .B(n4591), .Z(n4622) );
  IV U4956 ( .A(x[182]), .Z(n4592) );
  NOR U4957 ( .A(n6048), .B(n4592), .Z(n4619) );
  IV U4958 ( .A(x[118]), .Z(n4593) );
  NOR U4959 ( .A(n4593), .B(n6061), .Z(n4616) );
  IV U4960 ( .A(x[214]), .Z(n4594) );
  NOR U4961 ( .A(n6055), .B(n4594), .Z(n4613) );
  IV U4962 ( .A(x[278]), .Z(n4595) );
  NOR U4963 ( .A(n6065), .B(n4595), .Z(n4610) );
  IV U4964 ( .A(x[86]), .Z(n4596) );
  NOR U4965 ( .A(n6059), .B(n4596), .Z(n4599) );
  IV U4966 ( .A(x[54]), .Z(n4597) );
  NOR U4967 ( .A(n4597), .B(n6067), .Z(n4598) );
  NOR U4968 ( .A(n4599), .B(n4598), .Z(n4600) );
  IV U4969 ( .A(n4600), .Z(n4607) );
  IV U4970 ( .A(x[150]), .Z(n4601) );
  NOR U4971 ( .A(n6051), .B(n4601), .Z(n4604) );
  IV U4972 ( .A(x[22]), .Z(n4602) );
  NOR U4973 ( .A(n6052), .B(n4602), .Z(n4603) );
  NOR U4974 ( .A(n4604), .B(n4603), .Z(n4605) );
  IV U4975 ( .A(n4605), .Z(n4606) );
  NOR U4976 ( .A(n4607), .B(n4606), .Z(n4608) );
  IV U4977 ( .A(n4608), .Z(n4609) );
  NOR U4978 ( .A(n4610), .B(n4609), .Z(n4611) );
  IV U4979 ( .A(n4611), .Z(n4612) );
  NOR U4980 ( .A(n4613), .B(n4612), .Z(n4614) );
  IV U4981 ( .A(n4614), .Z(n4615) );
  NOR U4982 ( .A(n4616), .B(n4615), .Z(n4617) );
  IV U4983 ( .A(n4617), .Z(n4618) );
  NOR U4984 ( .A(n4619), .B(n4618), .Z(n4620) );
  IV U4985 ( .A(n4620), .Z(n4621) );
  NOR U4986 ( .A(n4622), .B(n4621), .Z(n7531) );
  NOR U4987 ( .A(n9429), .B(n7531), .Z(n4624) );
  IV U4988 ( .A(n4624), .Z(n4623) );
  NOR U4989 ( .A(n4625), .B(n4623), .Z(n4692) );
  XOR U4990 ( .A(n4625), .B(n4624), .Z(n5849) );
  IV U4991 ( .A(y[265]), .Z(n4626) );
  NOR U4992 ( .A(n6197), .B(n4626), .Z(n4657) );
  IV U4993 ( .A(y[137]), .Z(n4627) );
  NOR U4994 ( .A(n6214), .B(n4627), .Z(n4654) );
  IV U4995 ( .A(y[9]), .Z(n4628) );
  NOR U4996 ( .A(n4628), .B(n6200), .Z(n4651) );
  IV U4997 ( .A(y[73]), .Z(n4629) );
  NOR U4998 ( .A(n6216), .B(n4629), .Z(n4648) );
  IV U4999 ( .A(y[233]), .Z(n4630) );
  NOR U5000 ( .A(n6205), .B(n4630), .Z(n4645) );
  IV U5001 ( .A(y[41]), .Z(n4631) );
  NOR U5002 ( .A(n6207), .B(n4631), .Z(n4634) );
  IV U5003 ( .A(y[105]), .Z(n4632) );
  NOR U5004 ( .A(n6209), .B(n4632), .Z(n4633) );
  NOR U5005 ( .A(n4634), .B(n4633), .Z(n4635) );
  IV U5006 ( .A(n4635), .Z(n4642) );
  IV U5007 ( .A(y[201]), .Z(n4636) );
  NOR U5008 ( .A(n6203), .B(n4636), .Z(n4639) );
  IV U5009 ( .A(y[169]), .Z(n4637) );
  NOR U5010 ( .A(n4637), .B(n6199), .Z(n4638) );
  NOR U5011 ( .A(n4639), .B(n4638), .Z(n4640) );
  IV U5012 ( .A(n4640), .Z(n4641) );
  NOR U5013 ( .A(n4642), .B(n4641), .Z(n4643) );
  IV U5014 ( .A(n4643), .Z(n4644) );
  NOR U5015 ( .A(n4645), .B(n4644), .Z(n4646) );
  IV U5016 ( .A(n4646), .Z(n4647) );
  NOR U5017 ( .A(n4648), .B(n4647), .Z(n4649) );
  IV U5018 ( .A(n4649), .Z(n4650) );
  NOR U5019 ( .A(n4651), .B(n4650), .Z(n4652) );
  IV U5020 ( .A(n4652), .Z(n4653) );
  NOR U5021 ( .A(n4654), .B(n4653), .Z(n4655) );
  IV U5022 ( .A(n4655), .Z(n4656) );
  NOR U5023 ( .A(n4657), .B(n4656), .Z(n9237) );
  IV U5024 ( .A(x[179]), .Z(n4658) );
  NOR U5025 ( .A(n6048), .B(n4658), .Z(n4689) );
  IV U5026 ( .A(x[275]), .Z(n4659) );
  NOR U5027 ( .A(n6065), .B(n4659), .Z(n4686) );
  IV U5028 ( .A(x[19]), .Z(n4660) );
  NOR U5029 ( .A(n4660), .B(n6052), .Z(n4683) );
  IV U5030 ( .A(x[83]), .Z(n4661) );
  NOR U5031 ( .A(n6059), .B(n4661), .Z(n4680) );
  IV U5032 ( .A(x[243]), .Z(n4662) );
  NOR U5033 ( .A(n6057), .B(n4662), .Z(n4677) );
  IV U5034 ( .A(x[211]), .Z(n4663) );
  NOR U5035 ( .A(n6055), .B(n4663), .Z(n4666) );
  IV U5036 ( .A(x[51]), .Z(n4664) );
  NOR U5037 ( .A(n6067), .B(n4664), .Z(n4665) );
  NOR U5038 ( .A(n4666), .B(n4665), .Z(n4667) );
  IV U5039 ( .A(n4667), .Z(n4674) );
  IV U5040 ( .A(x[147]), .Z(n4668) );
  NOR U5041 ( .A(n6051), .B(n4668), .Z(n4671) );
  IV U5042 ( .A(x[115]), .Z(n4669) );
  NOR U5043 ( .A(n6061), .B(n4669), .Z(n4670) );
  NOR U5044 ( .A(n4671), .B(n4670), .Z(n4672) );
  IV U5045 ( .A(n4672), .Z(n4673) );
  NOR U5046 ( .A(n4674), .B(n4673), .Z(n4675) );
  IV U5047 ( .A(n4675), .Z(n4676) );
  NOR U5048 ( .A(n4677), .B(n4676), .Z(n4678) );
  IV U5049 ( .A(n4678), .Z(n4679) );
  NOR U5050 ( .A(n4680), .B(n4679), .Z(n4681) );
  IV U5051 ( .A(n4681), .Z(n4682) );
  NOR U5052 ( .A(n4683), .B(n4682), .Z(n4684) );
  IV U5053 ( .A(n4684), .Z(n4685) );
  NOR U5054 ( .A(n4686), .B(n4685), .Z(n4687) );
  IV U5055 ( .A(n4687), .Z(n4688) );
  NOR U5056 ( .A(n4689), .B(n4688), .Z(n8068) );
  NOR U5057 ( .A(n9237), .B(n8068), .Z(n4690) );
  IV U5058 ( .A(n4690), .Z(n5850) );
  NOR U5059 ( .A(n5849), .B(n5850), .Z(n4691) );
  NOR U5060 ( .A(n4692), .B(n4691), .Z(n5844) );
  XOR U5061 ( .A(n4694), .B(n4693), .Z(n5843) );
  IV U5062 ( .A(n5843), .Z(n4695) );
  NOR U5063 ( .A(n5844), .B(n4695), .Z(n4696) );
  NOR U5064 ( .A(n4697), .B(n4696), .Z(n5861) );
  IV U5065 ( .A(x[180]), .Z(n4698) );
  NOR U5066 ( .A(n4698), .B(n6048), .Z(n4729) );
  IV U5067 ( .A(x[148]), .Z(n4699) );
  NOR U5068 ( .A(n6051), .B(n4699), .Z(n4726) );
  IV U5069 ( .A(x[212]), .Z(n4700) );
  NOR U5070 ( .A(n4700), .B(n6055), .Z(n4723) );
  IV U5071 ( .A(x[84]), .Z(n4701) );
  NOR U5072 ( .A(n6059), .B(n4701), .Z(n4720) );
  IV U5073 ( .A(x[244]), .Z(n4702) );
  NOR U5074 ( .A(n6057), .B(n4702), .Z(n4717) );
  IV U5075 ( .A(x[20]), .Z(n4703) );
  NOR U5076 ( .A(n6052), .B(n4703), .Z(n4706) );
  IV U5077 ( .A(x[116]), .Z(n4704) );
  NOR U5078 ( .A(n6061), .B(n4704), .Z(n4705) );
  NOR U5079 ( .A(n4706), .B(n4705), .Z(n4707) );
  IV U5080 ( .A(n4707), .Z(n4714) );
  IV U5081 ( .A(x[276]), .Z(n4708) );
  NOR U5082 ( .A(n4708), .B(n6065), .Z(n4711) );
  IV U5083 ( .A(x[52]), .Z(n4709) );
  NOR U5084 ( .A(n4709), .B(n6067), .Z(n4710) );
  NOR U5085 ( .A(n4711), .B(n4710), .Z(n4712) );
  IV U5086 ( .A(n4712), .Z(n4713) );
  NOR U5087 ( .A(n4714), .B(n4713), .Z(n4715) );
  IV U5088 ( .A(n4715), .Z(n4716) );
  NOR U5089 ( .A(n4717), .B(n4716), .Z(n4718) );
  IV U5090 ( .A(n4718), .Z(n4719) );
  NOR U5091 ( .A(n4720), .B(n4719), .Z(n4721) );
  IV U5092 ( .A(n4721), .Z(n4722) );
  NOR U5093 ( .A(n4723), .B(n4722), .Z(n4724) );
  IV U5094 ( .A(n4724), .Z(n4725) );
  NOR U5095 ( .A(n4726), .B(n4725), .Z(n4727) );
  IV U5096 ( .A(n4727), .Z(n4728) );
  NOR U5097 ( .A(n4729), .B(n4728), .Z(n7851) );
  NOR U5098 ( .A(n9237), .B(n7851), .Z(n5942) );
  IV U5099 ( .A(y[250]), .Z(n4730) );
  NOR U5100 ( .A(n6205), .B(n4730), .Z(n4761) );
  IV U5101 ( .A(y[282]), .Z(n4731) );
  NOR U5102 ( .A(n6197), .B(n4731), .Z(n4758) );
  IV U5103 ( .A(y[122]), .Z(n4732) );
  NOR U5104 ( .A(n4732), .B(n6209), .Z(n4755) );
  IV U5105 ( .A(y[90]), .Z(n4733) );
  NOR U5106 ( .A(n6216), .B(n4733), .Z(n4752) );
  IV U5107 ( .A(y[186]), .Z(n4734) );
  NOR U5108 ( .A(n6199), .B(n4734), .Z(n4749) );
  IV U5109 ( .A(y[218]), .Z(n4735) );
  NOR U5110 ( .A(n6203), .B(n4735), .Z(n4738) );
  IV U5111 ( .A(y[58]), .Z(n4736) );
  NOR U5112 ( .A(n6207), .B(n4736), .Z(n4737) );
  NOR U5113 ( .A(n4738), .B(n4737), .Z(n4739) );
  IV U5114 ( .A(n4739), .Z(n4746) );
  IV U5115 ( .A(y[154]), .Z(n4740) );
  NOR U5116 ( .A(n6214), .B(n4740), .Z(n4743) );
  IV U5117 ( .A(y[26]), .Z(n4741) );
  NOR U5118 ( .A(n6200), .B(n4741), .Z(n4742) );
  NOR U5119 ( .A(n4743), .B(n4742), .Z(n4744) );
  IV U5120 ( .A(n4744), .Z(n4745) );
  NOR U5121 ( .A(n4746), .B(n4745), .Z(n4747) );
  IV U5122 ( .A(n4747), .Z(n4748) );
  NOR U5123 ( .A(n4749), .B(n4748), .Z(n4750) );
  IV U5124 ( .A(n4750), .Z(n4751) );
  NOR U5125 ( .A(n4752), .B(n4751), .Z(n4753) );
  IV U5126 ( .A(n4753), .Z(n4754) );
  NOR U5127 ( .A(n4755), .B(n4754), .Z(n4756) );
  IV U5128 ( .A(n4756), .Z(n4757) );
  NOR U5129 ( .A(n4758), .B(n4757), .Z(n4759) );
  IV U5130 ( .A(n4759), .Z(n4760) );
  NOR U5131 ( .A(n4761), .B(n4760), .Z(n6731) );
  IV U5132 ( .A(x[259]), .Z(n4762) );
  NOR U5133 ( .A(n4762), .B(n6065), .Z(n4793) );
  IV U5134 ( .A(x[131]), .Z(n4763) );
  NOR U5135 ( .A(n6051), .B(n4763), .Z(n4790) );
  IV U5136 ( .A(x[3]), .Z(n4764) );
  NOR U5137 ( .A(n6052), .B(n4764), .Z(n4787) );
  IV U5138 ( .A(x[195]), .Z(n4765) );
  NOR U5139 ( .A(n6055), .B(n4765), .Z(n4784) );
  IV U5140 ( .A(x[227]), .Z(n4766) );
  NOR U5141 ( .A(n6057), .B(n4766), .Z(n4781) );
  IV U5142 ( .A(x[67]), .Z(n4767) );
  NOR U5143 ( .A(n6059), .B(n4767), .Z(n4770) );
  IV U5144 ( .A(x[35]), .Z(n4768) );
  NOR U5145 ( .A(n4768), .B(n6067), .Z(n4769) );
  NOR U5146 ( .A(n4770), .B(n4769), .Z(n4771) );
  IV U5147 ( .A(n4771), .Z(n4778) );
  IV U5148 ( .A(x[99]), .Z(n4772) );
  NOR U5149 ( .A(n6061), .B(n4772), .Z(n4775) );
  IV U5150 ( .A(x[163]), .Z(n4773) );
  NOR U5151 ( .A(n6048), .B(n4773), .Z(n4774) );
  NOR U5152 ( .A(n4775), .B(n4774), .Z(n4776) );
  IV U5153 ( .A(n4776), .Z(n4777) );
  NOR U5154 ( .A(n4778), .B(n4777), .Z(n4779) );
  IV U5155 ( .A(n4779), .Z(n4780) );
  NOR U5156 ( .A(n4781), .B(n4780), .Z(n4782) );
  IV U5157 ( .A(n4782), .Z(n4783) );
  NOR U5158 ( .A(n4784), .B(n4783), .Z(n4785) );
  IV U5159 ( .A(n4785), .Z(n4786) );
  NOR U5160 ( .A(n4787), .B(n4786), .Z(n4788) );
  IV U5161 ( .A(n4788), .Z(n4789) );
  NOR U5162 ( .A(n4790), .B(n4789), .Z(n4791) );
  IV U5163 ( .A(n4791), .Z(n4792) );
  NOR U5164 ( .A(n4793), .B(n4792), .Z(n9493) );
  NOR U5165 ( .A(n6731), .B(n9493), .Z(n4794) );
  IV U5166 ( .A(n4794), .Z(n5943) );
  XOR U5167 ( .A(n5942), .B(n5943), .Z(n5945) );
  IV U5168 ( .A(y[281]), .Z(n4795) );
  NOR U5169 ( .A(n4795), .B(n6197), .Z(n4826) );
  IV U5170 ( .A(y[153]), .Z(n4796) );
  NOR U5171 ( .A(n6214), .B(n4796), .Z(n4823) );
  IV U5172 ( .A(y[57]), .Z(n4797) );
  NOR U5173 ( .A(n6207), .B(n4797), .Z(n4820) );
  IV U5174 ( .A(y[217]), .Z(n4798) );
  NOR U5175 ( .A(n6203), .B(n4798), .Z(n4817) );
  IV U5176 ( .A(y[249]), .Z(n4799) );
  NOR U5177 ( .A(n6205), .B(n4799), .Z(n4814) );
  IV U5178 ( .A(y[89]), .Z(n4800) );
  NOR U5179 ( .A(n6216), .B(n4800), .Z(n4803) );
  IV U5180 ( .A(y[121]), .Z(n4801) );
  NOR U5181 ( .A(n6209), .B(n4801), .Z(n4802) );
  NOR U5182 ( .A(n4803), .B(n4802), .Z(n4804) );
  IV U5183 ( .A(n4804), .Z(n4811) );
  IV U5184 ( .A(y[185]), .Z(n4805) );
  NOR U5185 ( .A(n6199), .B(n4805), .Z(n4808) );
  IV U5186 ( .A(y[25]), .Z(n4806) );
  NOR U5187 ( .A(n6200), .B(n4806), .Z(n4807) );
  NOR U5188 ( .A(n4808), .B(n4807), .Z(n4809) );
  IV U5189 ( .A(n4809), .Z(n4810) );
  NOR U5190 ( .A(n4811), .B(n4810), .Z(n4812) );
  IV U5191 ( .A(n4812), .Z(n4813) );
  NOR U5192 ( .A(n4814), .B(n4813), .Z(n4815) );
  IV U5193 ( .A(n4815), .Z(n4816) );
  NOR U5194 ( .A(n4817), .B(n4816), .Z(n4818) );
  IV U5195 ( .A(n4818), .Z(n4819) );
  NOR U5196 ( .A(n4820), .B(n4819), .Z(n4821) );
  IV U5197 ( .A(n4821), .Z(n4822) );
  NOR U5198 ( .A(n4823), .B(n4822), .Z(n4824) );
  IV U5199 ( .A(n4824), .Z(n4825) );
  NOR U5200 ( .A(n4826), .B(n4825), .Z(n6784) );
  IV U5201 ( .A(x[260]), .Z(n4827) );
  NOR U5202 ( .A(n4827), .B(n6065), .Z(n4858) );
  IV U5203 ( .A(x[132]), .Z(n4828) );
  NOR U5204 ( .A(n6051), .B(n4828), .Z(n4855) );
  IV U5205 ( .A(x[4]), .Z(n4829) );
  NOR U5206 ( .A(n4829), .B(n6052), .Z(n4852) );
  IV U5207 ( .A(x[68]), .Z(n4830) );
  NOR U5208 ( .A(n6059), .B(n4830), .Z(n4849) );
  IV U5209 ( .A(x[228]), .Z(n4831) );
  NOR U5210 ( .A(n6057), .B(n4831), .Z(n4846) );
  IV U5211 ( .A(x[196]), .Z(n4832) );
  NOR U5212 ( .A(n6055), .B(n4832), .Z(n4835) );
  IV U5213 ( .A(x[100]), .Z(n4833) );
  NOR U5214 ( .A(n6061), .B(n4833), .Z(n4834) );
  NOR U5215 ( .A(n4835), .B(n4834), .Z(n4836) );
  IV U5216 ( .A(n4836), .Z(n4843) );
  IV U5217 ( .A(x[36]), .Z(n4837) );
  NOR U5218 ( .A(n6067), .B(n4837), .Z(n4840) );
  IV U5219 ( .A(x[164]), .Z(n4838) );
  NOR U5220 ( .A(n4838), .B(n6048), .Z(n4839) );
  NOR U5221 ( .A(n4840), .B(n4839), .Z(n4841) );
  IV U5222 ( .A(n4841), .Z(n4842) );
  NOR U5223 ( .A(n4843), .B(n4842), .Z(n4844) );
  IV U5224 ( .A(n4844), .Z(n4845) );
  NOR U5225 ( .A(n4846), .B(n4845), .Z(n4847) );
  IV U5226 ( .A(n4847), .Z(n4848) );
  NOR U5227 ( .A(n4849), .B(n4848), .Z(n4850) );
  IV U5228 ( .A(n4850), .Z(n4851) );
  NOR U5229 ( .A(n4852), .B(n4851), .Z(n4853) );
  IV U5230 ( .A(n4853), .Z(n4854) );
  NOR U5231 ( .A(n4855), .B(n4854), .Z(n4856) );
  IV U5232 ( .A(n4856), .Z(n4857) );
  NOR U5233 ( .A(n4858), .B(n4857), .Z(n9526) );
  NOR U5234 ( .A(n6784), .B(n9526), .Z(n4859) );
  IV U5235 ( .A(n4859), .Z(n5944) );
  XOR U5236 ( .A(n5945), .B(n5944), .Z(n6342) );
  IV U5237 ( .A(y[231]), .Z(n4860) );
  NOR U5238 ( .A(n4860), .B(n6205), .Z(n4891) );
  IV U5239 ( .A(y[263]), .Z(n4861) );
  NOR U5240 ( .A(n6197), .B(n4861), .Z(n4888) );
  IV U5241 ( .A(y[103]), .Z(n4862) );
  NOR U5242 ( .A(n6209), .B(n4862), .Z(n4885) );
  IV U5243 ( .A(y[39]), .Z(n4863) );
  NOR U5244 ( .A(n6207), .B(n4863), .Z(n4882) );
  IV U5245 ( .A(y[167]), .Z(n4864) );
  NOR U5246 ( .A(n6199), .B(n4864), .Z(n4879) );
  IV U5247 ( .A(y[199]), .Z(n4865) );
  NOR U5248 ( .A(n6203), .B(n4865), .Z(n4868) );
  IV U5249 ( .A(y[71]), .Z(n4866) );
  NOR U5250 ( .A(n6216), .B(n4866), .Z(n4867) );
  NOR U5251 ( .A(n4868), .B(n4867), .Z(n4869) );
  IV U5252 ( .A(n4869), .Z(n4876) );
  IV U5253 ( .A(y[135]), .Z(n4870) );
  NOR U5254 ( .A(n6214), .B(n4870), .Z(n4873) );
  IV U5255 ( .A(y[7]), .Z(n4871) );
  NOR U5256 ( .A(n6200), .B(n4871), .Z(n4872) );
  NOR U5257 ( .A(n4873), .B(n4872), .Z(n4874) );
  IV U5258 ( .A(n4874), .Z(n4875) );
  NOR U5259 ( .A(n4876), .B(n4875), .Z(n4877) );
  IV U5260 ( .A(n4877), .Z(n4878) );
  NOR U5261 ( .A(n4879), .B(n4878), .Z(n4880) );
  IV U5262 ( .A(n4880), .Z(n4881) );
  NOR U5263 ( .A(n4882), .B(n4881), .Z(n4883) );
  IV U5264 ( .A(n4883), .Z(n4884) );
  NOR U5265 ( .A(n4885), .B(n4884), .Z(n4886) );
  IV U5266 ( .A(n4886), .Z(n4887) );
  NOR U5267 ( .A(n4888), .B(n4887), .Z(n4889) );
  IV U5268 ( .A(n4889), .Z(n4890) );
  NOR U5269 ( .A(n4891), .B(n4890), .Z(n9301) );
  NOR U5270 ( .A(n7531), .B(n9301), .Z(n6340) );
  IV U5271 ( .A(y[164]), .Z(n4892) );
  NOR U5272 ( .A(n6199), .B(n4892), .Z(n4923) );
  IV U5273 ( .A(y[132]), .Z(n4893) );
  NOR U5274 ( .A(n6214), .B(n4893), .Z(n4920) );
  IV U5275 ( .A(y[36]), .Z(n4894) );
  NOR U5276 ( .A(n6207), .B(n4894), .Z(n4917) );
  IV U5277 ( .A(y[196]), .Z(n4895) );
  NOR U5278 ( .A(n6203), .B(n4895), .Z(n4914) );
  IV U5279 ( .A(y[228]), .Z(n4896) );
  NOR U5280 ( .A(n6205), .B(n4896), .Z(n4911) );
  IV U5281 ( .A(y[68]), .Z(n4897) );
  NOR U5282 ( .A(n6216), .B(n4897), .Z(n4900) );
  IV U5283 ( .A(y[100]), .Z(n4898) );
  NOR U5284 ( .A(n6209), .B(n4898), .Z(n4899) );
  NOR U5285 ( .A(n4900), .B(n4899), .Z(n4901) );
  IV U5286 ( .A(n4901), .Z(n4908) );
  IV U5287 ( .A(y[4]), .Z(n4902) );
  NOR U5288 ( .A(n6200), .B(n4902), .Z(n4905) );
  IV U5289 ( .A(y[260]), .Z(n4903) );
  NOR U5290 ( .A(n6197), .B(n4903), .Z(n4904) );
  NOR U5291 ( .A(n4905), .B(n4904), .Z(n4906) );
  IV U5292 ( .A(n4906), .Z(n4907) );
  NOR U5293 ( .A(n4908), .B(n4907), .Z(n4909) );
  IV U5294 ( .A(n4909), .Z(n4910) );
  NOR U5295 ( .A(n4911), .B(n4910), .Z(n4912) );
  IV U5296 ( .A(n4912), .Z(n4913) );
  NOR U5297 ( .A(n4914), .B(n4913), .Z(n4915) );
  IV U5298 ( .A(n4915), .Z(n4916) );
  NOR U5299 ( .A(n4917), .B(n4916), .Z(n4918) );
  IV U5300 ( .A(n4918), .Z(n4919) );
  NOR U5301 ( .A(n4920), .B(n4919), .Z(n4921) );
  IV U5302 ( .A(n4921), .Z(n4922) );
  NOR U5303 ( .A(n4923), .B(n4922), .Z(n9472) );
  IV U5304 ( .A(x[249]), .Z(n4924) );
  NOR U5305 ( .A(n4924), .B(n6057), .Z(n4955) );
  IV U5306 ( .A(x[185]), .Z(n4925) );
  NOR U5307 ( .A(n6048), .B(n4925), .Z(n4952) );
  IV U5308 ( .A(x[25]), .Z(n4926) );
  NOR U5309 ( .A(n4926), .B(n6052), .Z(n4949) );
  IV U5310 ( .A(x[217]), .Z(n4927) );
  NOR U5311 ( .A(n6055), .B(n4927), .Z(n4946) );
  IV U5312 ( .A(x[121]), .Z(n4928) );
  NOR U5313 ( .A(n6061), .B(n4928), .Z(n4943) );
  IV U5314 ( .A(x[89]), .Z(n4929) );
  NOR U5315 ( .A(n6059), .B(n4929), .Z(n4932) );
  IV U5316 ( .A(x[57]), .Z(n4930) );
  NOR U5317 ( .A(n4930), .B(n6067), .Z(n4931) );
  NOR U5318 ( .A(n4932), .B(n4931), .Z(n4933) );
  IV U5319 ( .A(n4933), .Z(n4940) );
  IV U5320 ( .A(x[153]), .Z(n4934) );
  NOR U5321 ( .A(n6051), .B(n4934), .Z(n4937) );
  IV U5322 ( .A(x[281]), .Z(n4935) );
  NOR U5323 ( .A(n6065), .B(n4935), .Z(n4936) );
  NOR U5324 ( .A(n4937), .B(n4936), .Z(n4938) );
  IV U5325 ( .A(n4938), .Z(n4939) );
  NOR U5326 ( .A(n4940), .B(n4939), .Z(n4941) );
  IV U5327 ( .A(n4941), .Z(n4942) );
  NOR U5328 ( .A(n4943), .B(n4942), .Z(n4944) );
  IV U5329 ( .A(n4944), .Z(n4945) );
  NOR U5330 ( .A(n4946), .B(n4945), .Z(n4947) );
  IV U5331 ( .A(n4947), .Z(n4948) );
  NOR U5332 ( .A(n4949), .B(n4948), .Z(n4950) );
  IV U5333 ( .A(n4950), .Z(n4951) );
  NOR U5334 ( .A(n4952), .B(n4951), .Z(n4953) );
  IV U5335 ( .A(n4953), .Z(n4954) );
  NOR U5336 ( .A(n4955), .B(n4954), .Z(n6957) );
  NOR U5337 ( .A(n9472), .B(n6957), .Z(n6339) );
  XOR U5338 ( .A(n6340), .B(n6339), .Z(n4956) );
  IV U5339 ( .A(n4956), .Z(n6341) );
  XOR U5340 ( .A(n6342), .B(n6341), .Z(n5832) );
  IV U5341 ( .A(y[268]), .Z(n4957) );
  NOR U5342 ( .A(n4957), .B(n6197), .Z(n4988) );
  IV U5343 ( .A(y[172]), .Z(n4958) );
  NOR U5344 ( .A(n6199), .B(n4958), .Z(n4985) );
  IV U5345 ( .A(y[108]), .Z(n4959) );
  NOR U5346 ( .A(n4959), .B(n6209), .Z(n4982) );
  IV U5347 ( .A(y[204]), .Z(n4960) );
  NOR U5348 ( .A(n6203), .B(n4960), .Z(n4979) );
  IV U5349 ( .A(y[236]), .Z(n4961) );
  NOR U5350 ( .A(n6205), .B(n4961), .Z(n4976) );
  IV U5351 ( .A(y[12]), .Z(n4962) );
  NOR U5352 ( .A(n6200), .B(n4962), .Z(n4965) );
  IV U5353 ( .A(y[44]), .Z(n4963) );
  NOR U5354 ( .A(n6207), .B(n4963), .Z(n4964) );
  NOR U5355 ( .A(n4965), .B(n4964), .Z(n4966) );
  IV U5356 ( .A(n4966), .Z(n4973) );
  IV U5357 ( .A(y[140]), .Z(n4967) );
  NOR U5358 ( .A(n6214), .B(n4967), .Z(n4970) );
  IV U5359 ( .A(y[76]), .Z(n4968) );
  NOR U5360 ( .A(n6216), .B(n4968), .Z(n4969) );
  NOR U5361 ( .A(n4970), .B(n4969), .Z(n4971) );
  IV U5362 ( .A(n4971), .Z(n4972) );
  NOR U5363 ( .A(n4973), .B(n4972), .Z(n4974) );
  IV U5364 ( .A(n4974), .Z(n4975) );
  NOR U5365 ( .A(n4976), .B(n4975), .Z(n4977) );
  IV U5366 ( .A(n4977), .Z(n4978) );
  NOR U5367 ( .A(n4979), .B(n4978), .Z(n4980) );
  IV U5368 ( .A(n4980), .Z(n4981) );
  NOR U5369 ( .A(n4982), .B(n4981), .Z(n4983) );
  IV U5370 ( .A(n4983), .Z(n4984) );
  NOR U5371 ( .A(n4985), .B(n4984), .Z(n4986) );
  IV U5372 ( .A(n4986), .Z(n4987) );
  NOR U5373 ( .A(n4988), .B(n4987), .Z(n8948) );
  IV U5374 ( .A(x[241]), .Z(n4989) );
  NOR U5375 ( .A(n4989), .B(n6057), .Z(n5020) );
  IV U5376 ( .A(x[145]), .Z(n4990) );
  NOR U5377 ( .A(n6051), .B(n4990), .Z(n5017) );
  IV U5378 ( .A(x[17]), .Z(n4991) );
  NOR U5379 ( .A(n4991), .B(n6052), .Z(n5014) );
  IV U5380 ( .A(x[81]), .Z(n4992) );
  NOR U5381 ( .A(n6059), .B(n4992), .Z(n5011) );
  IV U5382 ( .A(x[177]), .Z(n4993) );
  NOR U5383 ( .A(n6048), .B(n4993), .Z(n5008) );
  IV U5384 ( .A(x[209]), .Z(n4994) );
  NOR U5385 ( .A(n6055), .B(n4994), .Z(n4997) );
  IV U5386 ( .A(x[49]), .Z(n4995) );
  NOR U5387 ( .A(n6067), .B(n4995), .Z(n4996) );
  NOR U5388 ( .A(n4997), .B(n4996), .Z(n4998) );
  IV U5389 ( .A(n4998), .Z(n5005) );
  IV U5390 ( .A(x[273]), .Z(n4999) );
  NOR U5391 ( .A(n6065), .B(n4999), .Z(n5002) );
  IV U5392 ( .A(x[113]), .Z(n5000) );
  NOR U5393 ( .A(n6061), .B(n5000), .Z(n5001) );
  NOR U5394 ( .A(n5002), .B(n5001), .Z(n5003) );
  IV U5395 ( .A(n5003), .Z(n5004) );
  NOR U5396 ( .A(n5005), .B(n5004), .Z(n5006) );
  IV U5397 ( .A(n5006), .Z(n5007) );
  NOR U5398 ( .A(n5008), .B(n5007), .Z(n5009) );
  IV U5399 ( .A(n5009), .Z(n5010) );
  NOR U5400 ( .A(n5011), .B(n5010), .Z(n5012) );
  IV U5401 ( .A(n5012), .Z(n5013) );
  NOR U5402 ( .A(n5014), .B(n5013), .Z(n5015) );
  IV U5403 ( .A(n5015), .Z(n5016) );
  NOR U5404 ( .A(n5017), .B(n5016), .Z(n5018) );
  IV U5405 ( .A(n5018), .Z(n5019) );
  NOR U5406 ( .A(n5020), .B(n5019), .Z(n8311) );
  NOR U5407 ( .A(n8948), .B(n8311), .Z(n6306) );
  IV U5408 ( .A(y[273]), .Z(n5021) );
  NOR U5409 ( .A(n6197), .B(n5021), .Z(n5052) );
  IV U5410 ( .A(y[145]), .Z(n5022) );
  NOR U5411 ( .A(n6214), .B(n5022), .Z(n5049) );
  IV U5412 ( .A(y[17]), .Z(n5023) );
  NOR U5413 ( .A(n5023), .B(n6200), .Z(n5046) );
  IV U5414 ( .A(y[81]), .Z(n5024) );
  NOR U5415 ( .A(n6216), .B(n5024), .Z(n5043) );
  IV U5416 ( .A(y[241]), .Z(n5025) );
  NOR U5417 ( .A(n6205), .B(n5025), .Z(n5040) );
  IV U5418 ( .A(y[49]), .Z(n5026) );
  NOR U5419 ( .A(n6207), .B(n5026), .Z(n5029) );
  IV U5420 ( .A(y[113]), .Z(n5027) );
  NOR U5421 ( .A(n6209), .B(n5027), .Z(n5028) );
  NOR U5422 ( .A(n5029), .B(n5028), .Z(n5030) );
  IV U5423 ( .A(n5030), .Z(n5037) );
  IV U5424 ( .A(y[209]), .Z(n5031) );
  NOR U5425 ( .A(n6203), .B(n5031), .Z(n5034) );
  IV U5426 ( .A(y[177]), .Z(n5032) );
  NOR U5427 ( .A(n5032), .B(n6199), .Z(n5033) );
  NOR U5428 ( .A(n5034), .B(n5033), .Z(n5035) );
  IV U5429 ( .A(n5035), .Z(n5036) );
  NOR U5430 ( .A(n5037), .B(n5036), .Z(n5038) );
  IV U5431 ( .A(n5038), .Z(n5039) );
  NOR U5432 ( .A(n5040), .B(n5039), .Z(n5041) );
  IV U5433 ( .A(n5041), .Z(n5042) );
  NOR U5434 ( .A(n5043), .B(n5042), .Z(n5044) );
  IV U5435 ( .A(n5044), .Z(n5045) );
  NOR U5436 ( .A(n5046), .B(n5045), .Z(n5047) );
  IV U5437 ( .A(n5047), .Z(n5048) );
  NOR U5438 ( .A(n5049), .B(n5048), .Z(n5050) );
  IV U5439 ( .A(n5050), .Z(n5051) );
  NOR U5440 ( .A(n5052), .B(n5051), .Z(n8290) );
  IV U5441 ( .A(x[172]), .Z(n5053) );
  NOR U5442 ( .A(n5053), .B(n6048), .Z(n5084) );
  IV U5443 ( .A(x[268]), .Z(n5054) );
  NOR U5444 ( .A(n6065), .B(n5054), .Z(n5081) );
  IV U5445 ( .A(x[108]), .Z(n5055) );
  NOR U5446 ( .A(n6061), .B(n5055), .Z(n5078) );
  IV U5447 ( .A(x[12]), .Z(n5056) );
  NOR U5448 ( .A(n6052), .B(n5056), .Z(n5075) );
  IV U5449 ( .A(x[236]), .Z(n5057) );
  NOR U5450 ( .A(n6057), .B(n5057), .Z(n5072) );
  IV U5451 ( .A(x[76]), .Z(n5058) );
  NOR U5452 ( .A(n6059), .B(n5058), .Z(n5061) );
  IV U5453 ( .A(x[44]), .Z(n5059) );
  NOR U5454 ( .A(n5059), .B(n6067), .Z(n5060) );
  NOR U5455 ( .A(n5061), .B(n5060), .Z(n5062) );
  IV U5456 ( .A(n5062), .Z(n5069) );
  IV U5457 ( .A(x[140]), .Z(n5063) );
  NOR U5458 ( .A(n6051), .B(n5063), .Z(n5066) );
  IV U5459 ( .A(x[204]), .Z(n5064) );
  NOR U5460 ( .A(n6055), .B(n5064), .Z(n5065) );
  NOR U5461 ( .A(n5066), .B(n5065), .Z(n5067) );
  IV U5462 ( .A(n5067), .Z(n5068) );
  NOR U5463 ( .A(n5069), .B(n5068), .Z(n5070) );
  IV U5464 ( .A(n5070), .Z(n5071) );
  NOR U5465 ( .A(n5072), .B(n5071), .Z(n5073) );
  IV U5466 ( .A(n5073), .Z(n5074) );
  NOR U5467 ( .A(n5075), .B(n5074), .Z(n5076) );
  IV U5468 ( .A(n5076), .Z(n5077) );
  NOR U5469 ( .A(n5078), .B(n5077), .Z(n5079) );
  IV U5470 ( .A(n5079), .Z(n5080) );
  NOR U5471 ( .A(n5081), .B(n5080), .Z(n5082) );
  IV U5472 ( .A(n5082), .Z(n5083) );
  NOR U5473 ( .A(n5084), .B(n5083), .Z(n8754) );
  NOR U5474 ( .A(n8290), .B(n8754), .Z(n6303) );
  IV U5475 ( .A(y[234]), .Z(n5085) );
  NOR U5476 ( .A(n5085), .B(n6205), .Z(n5116) );
  IV U5477 ( .A(y[266]), .Z(n5086) );
  NOR U5478 ( .A(n6197), .B(n5086), .Z(n5113) );
  IV U5479 ( .A(y[106]), .Z(n5087) );
  NOR U5480 ( .A(n6209), .B(n5087), .Z(n5110) );
  IV U5481 ( .A(y[10]), .Z(n5088) );
  NOR U5482 ( .A(n6200), .B(n5088), .Z(n5107) );
  IV U5483 ( .A(y[170]), .Z(n5089) );
  NOR U5484 ( .A(n6199), .B(n5089), .Z(n5104) );
  IV U5485 ( .A(y[74]), .Z(n5090) );
  NOR U5486 ( .A(n6216), .B(n5090), .Z(n5093) );
  IV U5487 ( .A(y[42]), .Z(n5091) );
  NOR U5488 ( .A(n6207), .B(n5091), .Z(n5092) );
  NOR U5489 ( .A(n5093), .B(n5092), .Z(n5094) );
  IV U5490 ( .A(n5094), .Z(n5101) );
  IV U5491 ( .A(y[202]), .Z(n5095) );
  NOR U5492 ( .A(n6203), .B(n5095), .Z(n5098) );
  IV U5493 ( .A(y[138]), .Z(n5096) );
  NOR U5494 ( .A(n5096), .B(n6214), .Z(n5097) );
  NOR U5495 ( .A(n5098), .B(n5097), .Z(n5099) );
  IV U5496 ( .A(n5099), .Z(n5100) );
  NOR U5497 ( .A(n5101), .B(n5100), .Z(n5102) );
  IV U5498 ( .A(n5102), .Z(n5103) );
  NOR U5499 ( .A(n5104), .B(n5103), .Z(n5105) );
  IV U5500 ( .A(n5105), .Z(n5106) );
  NOR U5501 ( .A(n5107), .B(n5106), .Z(n5108) );
  IV U5502 ( .A(n5108), .Z(n5109) );
  NOR U5503 ( .A(n5110), .B(n5109), .Z(n5111) );
  IV U5504 ( .A(n5111), .Z(n5112) );
  NOR U5505 ( .A(n5113), .B(n5112), .Z(n5114) );
  IV U5506 ( .A(n5114), .Z(n5115) );
  NOR U5507 ( .A(n5116), .B(n5115), .Z(n9113) );
  NOR U5508 ( .A(n8068), .B(n9113), .Z(n5117) );
  IV U5509 ( .A(n5117), .Z(n6304) );
  XOR U5510 ( .A(n6303), .B(n6304), .Z(n6307) );
  XOR U5511 ( .A(n6306), .B(n6307), .Z(n5939) );
  IV U5512 ( .A(x[234]), .Z(n5118) );
  NOR U5513 ( .A(n6057), .B(n5118), .Z(n5149) );
  IV U5514 ( .A(x[266]), .Z(n5119) );
  NOR U5515 ( .A(n6065), .B(n5119), .Z(n5146) );
  IV U5516 ( .A(x[202]), .Z(n5120) );
  NOR U5517 ( .A(n6055), .B(n5120), .Z(n5143) );
  IV U5518 ( .A(x[74]), .Z(n5121) );
  NOR U5519 ( .A(n6059), .B(n5121), .Z(n5140) );
  IV U5520 ( .A(x[170]), .Z(n5122) );
  NOR U5521 ( .A(n6048), .B(n5122), .Z(n5137) );
  IV U5522 ( .A(x[10]), .Z(n5123) );
  NOR U5523 ( .A(n6052), .B(n5123), .Z(n5126) );
  IV U5524 ( .A(x[106]), .Z(n5124) );
  NOR U5525 ( .A(n6061), .B(n5124), .Z(n5125) );
  NOR U5526 ( .A(n5126), .B(n5125), .Z(n5127) );
  IV U5527 ( .A(n5127), .Z(n5134) );
  IV U5528 ( .A(x[138]), .Z(n5128) );
  NOR U5529 ( .A(n5128), .B(n6051), .Z(n5131) );
  IV U5530 ( .A(x[42]), .Z(n5129) );
  NOR U5531 ( .A(n5129), .B(n6067), .Z(n5130) );
  NOR U5532 ( .A(n5131), .B(n5130), .Z(n5132) );
  IV U5533 ( .A(n5132), .Z(n5133) );
  NOR U5534 ( .A(n5134), .B(n5133), .Z(n5135) );
  IV U5535 ( .A(n5135), .Z(n5136) );
  NOR U5536 ( .A(n5137), .B(n5136), .Z(n5138) );
  IV U5537 ( .A(n5138), .Z(n5139) );
  NOR U5538 ( .A(n5140), .B(n5139), .Z(n5141) );
  IV U5539 ( .A(n5141), .Z(n5142) );
  NOR U5540 ( .A(n5143), .B(n5142), .Z(n5144) );
  IV U5541 ( .A(n5144), .Z(n5145) );
  NOR U5542 ( .A(n5146), .B(n5145), .Z(n5147) );
  IV U5543 ( .A(n5147), .Z(n5148) );
  NOR U5544 ( .A(n5149), .B(n5148), .Z(n9115) );
  IV U5545 ( .A(y[275]), .Z(n5150) );
  NOR U5546 ( .A(n6197), .B(n5150), .Z(n5181) );
  IV U5547 ( .A(y[147]), .Z(n5151) );
  NOR U5548 ( .A(n6214), .B(n5151), .Z(n5178) );
  IV U5549 ( .A(y[115]), .Z(n5152) );
  NOR U5550 ( .A(n5152), .B(n6209), .Z(n5175) );
  IV U5551 ( .A(y[211]), .Z(n5153) );
  NOR U5552 ( .A(n6203), .B(n5153), .Z(n5172) );
  IV U5553 ( .A(y[243]), .Z(n5154) );
  NOR U5554 ( .A(n6205), .B(n5154), .Z(n5169) );
  IV U5555 ( .A(y[19]), .Z(n5155) );
  NOR U5556 ( .A(n6200), .B(n5155), .Z(n5158) );
  IV U5557 ( .A(y[51]), .Z(n5156) );
  NOR U5558 ( .A(n6207), .B(n5156), .Z(n5157) );
  NOR U5559 ( .A(n5158), .B(n5157), .Z(n5159) );
  IV U5560 ( .A(n5159), .Z(n5166) );
  IV U5561 ( .A(y[179]), .Z(n5160) );
  NOR U5562 ( .A(n6199), .B(n5160), .Z(n5163) );
  IV U5563 ( .A(y[83]), .Z(n5161) );
  NOR U5564 ( .A(n6216), .B(n5161), .Z(n5162) );
  NOR U5565 ( .A(n5163), .B(n5162), .Z(n5164) );
  IV U5566 ( .A(n5164), .Z(n5165) );
  NOR U5567 ( .A(n5166), .B(n5165), .Z(n5167) );
  IV U5568 ( .A(n5167), .Z(n5168) );
  NOR U5569 ( .A(n5169), .B(n5168), .Z(n5170) );
  IV U5570 ( .A(n5170), .Z(n5171) );
  NOR U5571 ( .A(n5172), .B(n5171), .Z(n5173) );
  IV U5572 ( .A(n5173), .Z(n5174) );
  NOR U5573 ( .A(n5175), .B(n5174), .Z(n5176) );
  IV U5574 ( .A(n5176), .Z(n5177) );
  NOR U5575 ( .A(n5178), .B(n5177), .Z(n5179) );
  IV U5576 ( .A(n5179), .Z(n5180) );
  NOR U5577 ( .A(n5181), .B(n5180), .Z(n8069) );
  NOR U5578 ( .A(n9115), .B(n8069), .Z(n5845) );
  IV U5579 ( .A(x[265]), .Z(n5182) );
  NOR U5580 ( .A(n5182), .B(n6065), .Z(n5213) );
  IV U5581 ( .A(x[137]), .Z(n5183) );
  NOR U5582 ( .A(n6051), .B(n5183), .Z(n5210) );
  IV U5583 ( .A(x[9]), .Z(n5184) );
  NOR U5584 ( .A(n6052), .B(n5184), .Z(n5207) );
  IV U5585 ( .A(x[201]), .Z(n5185) );
  NOR U5586 ( .A(n6055), .B(n5185), .Z(n5204) );
  IV U5587 ( .A(x[233]), .Z(n5186) );
  NOR U5588 ( .A(n6057), .B(n5186), .Z(n5201) );
  IV U5589 ( .A(x[73]), .Z(n5187) );
  NOR U5590 ( .A(n6059), .B(n5187), .Z(n5190) );
  IV U5591 ( .A(x[41]), .Z(n5188) );
  NOR U5592 ( .A(n5188), .B(n6067), .Z(n5189) );
  NOR U5593 ( .A(n5190), .B(n5189), .Z(n5191) );
  IV U5594 ( .A(n5191), .Z(n5198) );
  IV U5595 ( .A(x[105]), .Z(n5192) );
  NOR U5596 ( .A(n6061), .B(n5192), .Z(n5195) );
  IV U5597 ( .A(x[169]), .Z(n5193) );
  NOR U5598 ( .A(n6048), .B(n5193), .Z(n5194) );
  NOR U5599 ( .A(n5195), .B(n5194), .Z(n5196) );
  IV U5600 ( .A(n5196), .Z(n5197) );
  NOR U5601 ( .A(n5198), .B(n5197), .Z(n5199) );
  IV U5602 ( .A(n5199), .Z(n5200) );
  NOR U5603 ( .A(n5201), .B(n5200), .Z(n5202) );
  IV U5604 ( .A(n5202), .Z(n5203) );
  NOR U5605 ( .A(n5204), .B(n5203), .Z(n5205) );
  IV U5606 ( .A(n5205), .Z(n5206) );
  NOR U5607 ( .A(n5207), .B(n5206), .Z(n5208) );
  IV U5608 ( .A(n5208), .Z(n5209) );
  NOR U5609 ( .A(n5210), .B(n5209), .Z(n5211) );
  IV U5610 ( .A(n5211), .Z(n5212) );
  NOR U5611 ( .A(n5213), .B(n5212), .Z(n9241) );
  NOR U5612 ( .A(n7891), .B(n9241), .Z(n5214) );
  XOR U5613 ( .A(n5845), .B(n5214), .Z(n5937) );
  XOR U5614 ( .A(n5939), .B(n5937), .Z(n5833) );
  NOR U5615 ( .A(n5832), .B(n5833), .Z(n5836) );
  IV U5616 ( .A(sum[28]), .Z(n5280) );
  IV U5617 ( .A(y[225]), .Z(n5215) );
  NOR U5618 ( .A(n6205), .B(n5215), .Z(n5246) );
  IV U5619 ( .A(y[161]), .Z(n5216) );
  NOR U5620 ( .A(n6199), .B(n5216), .Z(n5243) );
  IV U5621 ( .A(y[1]), .Z(n5217) );
  NOR U5622 ( .A(n5217), .B(n6200), .Z(n5240) );
  IV U5623 ( .A(y[65]), .Z(n5218) );
  NOR U5624 ( .A(n6216), .B(n5218), .Z(n5237) );
  IV U5625 ( .A(y[257]), .Z(n5219) );
  NOR U5626 ( .A(n6197), .B(n5219), .Z(n5234) );
  IV U5627 ( .A(y[193]), .Z(n5220) );
  NOR U5628 ( .A(n6203), .B(n5220), .Z(n5223) );
  IV U5629 ( .A(y[33]), .Z(n5221) );
  NOR U5630 ( .A(n6207), .B(n5221), .Z(n5222) );
  NOR U5631 ( .A(n5223), .B(n5222), .Z(n5224) );
  IV U5632 ( .A(n5224), .Z(n5231) );
  IV U5633 ( .A(y[129]), .Z(n5225) );
  NOR U5634 ( .A(n5225), .B(n6214), .Z(n5228) );
  IV U5635 ( .A(y[97]), .Z(n5226) );
  NOR U5636 ( .A(n5226), .B(n6209), .Z(n5227) );
  NOR U5637 ( .A(n5228), .B(n5227), .Z(n5229) );
  IV U5638 ( .A(n5229), .Z(n5230) );
  NOR U5639 ( .A(n5231), .B(n5230), .Z(n5232) );
  IV U5640 ( .A(n5232), .Z(n5233) );
  NOR U5641 ( .A(n5234), .B(n5233), .Z(n5235) );
  IV U5642 ( .A(n5235), .Z(n5236) );
  NOR U5643 ( .A(n5237), .B(n5236), .Z(n5238) );
  IV U5644 ( .A(n5238), .Z(n5239) );
  NOR U5645 ( .A(n5240), .B(n5239), .Z(n5241) );
  IV U5646 ( .A(n5241), .Z(n5242) );
  NOR U5647 ( .A(n5243), .B(n5242), .Z(n5244) );
  IV U5648 ( .A(n5244), .Z(n5245) );
  NOR U5649 ( .A(n5246), .B(n5245), .Z(n9593) );
  IV U5650 ( .A(x[187]), .Z(n5247) );
  NOR U5651 ( .A(n5247), .B(n6048), .Z(n5278) );
  IV U5652 ( .A(x[283]), .Z(n5248) );
  NOR U5653 ( .A(n6065), .B(n5248), .Z(n5275) );
  IV U5654 ( .A(x[27]), .Z(n5249) );
  NOR U5655 ( .A(n6052), .B(n5249), .Z(n5272) );
  IV U5656 ( .A(x[219]), .Z(n5250) );
  NOR U5657 ( .A(n6055), .B(n5250), .Z(n5269) );
  IV U5658 ( .A(x[251]), .Z(n5251) );
  NOR U5659 ( .A(n6057), .B(n5251), .Z(n5266) );
  IV U5660 ( .A(x[59]), .Z(n5252) );
  NOR U5661 ( .A(n6067), .B(n5252), .Z(n5255) );
  IV U5662 ( .A(x[123]), .Z(n5253) );
  NOR U5663 ( .A(n6061), .B(n5253), .Z(n5254) );
  NOR U5664 ( .A(n5255), .B(n5254), .Z(n5256) );
  IV U5665 ( .A(n5256), .Z(n5263) );
  IV U5666 ( .A(x[91]), .Z(n5257) );
  NOR U5667 ( .A(n6059), .B(n5257), .Z(n5260) );
  IV U5668 ( .A(x[155]), .Z(n5258) );
  NOR U5669 ( .A(n5258), .B(n6051), .Z(n5259) );
  NOR U5670 ( .A(n5260), .B(n5259), .Z(n5261) );
  IV U5671 ( .A(n5261), .Z(n5262) );
  NOR U5672 ( .A(n5263), .B(n5262), .Z(n5264) );
  IV U5673 ( .A(n5264), .Z(n5265) );
  NOR U5674 ( .A(n5266), .B(n5265), .Z(n5267) );
  IV U5675 ( .A(n5267), .Z(n5268) );
  NOR U5676 ( .A(n5269), .B(n5268), .Z(n5270) );
  IV U5677 ( .A(n5270), .Z(n5271) );
  NOR U5678 ( .A(n5272), .B(n5271), .Z(n5273) );
  IV U5679 ( .A(n5273), .Z(n5274) );
  NOR U5680 ( .A(n5275), .B(n5274), .Z(n5276) );
  IV U5681 ( .A(n5276), .Z(n5277) );
  NOR U5682 ( .A(n5278), .B(n5277), .Z(n6581) );
  NOR U5683 ( .A(n9593), .B(n6581), .Z(n5279) );
  IV U5684 ( .A(n5279), .Z(n6359) );
  NOR U5685 ( .A(n5280), .B(n6359), .Z(n5912) );
  IV U5686 ( .A(y[272]), .Z(n5281) );
  NOR U5687 ( .A(n5281), .B(n6197), .Z(n5312) );
  IV U5688 ( .A(y[176]), .Z(n5282) );
  NOR U5689 ( .A(n6199), .B(n5282), .Z(n5309) );
  IV U5690 ( .A(y[16]), .Z(n5283) );
  NOR U5691 ( .A(n5283), .B(n6200), .Z(n5306) );
  IV U5692 ( .A(y[80]), .Z(n5284) );
  NOR U5693 ( .A(n6216), .B(n5284), .Z(n5303) );
  IV U5694 ( .A(y[240]), .Z(n5285) );
  NOR U5695 ( .A(n6205), .B(n5285), .Z(n5300) );
  IV U5696 ( .A(y[208]), .Z(n5286) );
  NOR U5697 ( .A(n6203), .B(n5286), .Z(n5289) );
  IV U5698 ( .A(y[48]), .Z(n5287) );
  NOR U5699 ( .A(n6207), .B(n5287), .Z(n5288) );
  NOR U5700 ( .A(n5289), .B(n5288), .Z(n5290) );
  IV U5701 ( .A(n5290), .Z(n5297) );
  IV U5702 ( .A(y[144]), .Z(n5291) );
  NOR U5703 ( .A(n5291), .B(n6214), .Z(n5294) );
  IV U5704 ( .A(y[112]), .Z(n5292) );
  NOR U5705 ( .A(n5292), .B(n6209), .Z(n5293) );
  NOR U5706 ( .A(n5294), .B(n5293), .Z(n5295) );
  IV U5707 ( .A(n5295), .Z(n5296) );
  NOR U5708 ( .A(n5297), .B(n5296), .Z(n5298) );
  IV U5709 ( .A(n5298), .Z(n5299) );
  NOR U5710 ( .A(n5300), .B(n5299), .Z(n5301) );
  IV U5711 ( .A(n5301), .Z(n5302) );
  NOR U5712 ( .A(n5303), .B(n5302), .Z(n5304) );
  IV U5713 ( .A(n5304), .Z(n5305) );
  NOR U5714 ( .A(n5306), .B(n5305), .Z(n5307) );
  IV U5715 ( .A(n5307), .Z(n5308) );
  NOR U5716 ( .A(n5309), .B(n5308), .Z(n5310) );
  IV U5717 ( .A(n5310), .Z(n5311) );
  NOR U5718 ( .A(n5312), .B(n5311), .Z(n8501) );
  IV U5719 ( .A(x[269]), .Z(n5313) );
  NOR U5720 ( .A(n5313), .B(n6065), .Z(n5344) );
  IV U5721 ( .A(x[141]), .Z(n5314) );
  NOR U5722 ( .A(n6051), .B(n5314), .Z(n5341) );
  IV U5723 ( .A(x[13]), .Z(n5315) );
  NOR U5724 ( .A(n5315), .B(n6052), .Z(n5338) );
  IV U5725 ( .A(x[205]), .Z(n5316) );
  NOR U5726 ( .A(n6055), .B(n5316), .Z(n5335) );
  IV U5727 ( .A(x[237]), .Z(n5317) );
  NOR U5728 ( .A(n6057), .B(n5317), .Z(n5332) );
  IV U5729 ( .A(x[77]), .Z(n5318) );
  NOR U5730 ( .A(n5318), .B(n6059), .Z(n5321) );
  IV U5731 ( .A(x[45]), .Z(n5319) );
  NOR U5732 ( .A(n5319), .B(n6067), .Z(n5320) );
  NOR U5733 ( .A(n5321), .B(n5320), .Z(n5322) );
  IV U5734 ( .A(n5322), .Z(n5329) );
  IV U5735 ( .A(x[109]), .Z(n5323) );
  NOR U5736 ( .A(n6061), .B(n5323), .Z(n5326) );
  IV U5737 ( .A(x[173]), .Z(n5324) );
  NOR U5738 ( .A(n6048), .B(n5324), .Z(n5325) );
  NOR U5739 ( .A(n5326), .B(n5325), .Z(n5327) );
  IV U5740 ( .A(n5327), .Z(n5328) );
  NOR U5741 ( .A(n5329), .B(n5328), .Z(n5330) );
  IV U5742 ( .A(n5330), .Z(n5331) );
  NOR U5743 ( .A(n5332), .B(n5331), .Z(n5333) );
  IV U5744 ( .A(n5333), .Z(n5334) );
  NOR U5745 ( .A(n5335), .B(n5334), .Z(n5336) );
  IV U5746 ( .A(n5336), .Z(n5337) );
  NOR U5747 ( .A(n5338), .B(n5337), .Z(n5339) );
  IV U5748 ( .A(n5339), .Z(n5340) );
  NOR U5749 ( .A(n5341), .B(n5340), .Z(n5342) );
  IV U5750 ( .A(n5342), .Z(n5343) );
  NOR U5751 ( .A(n5344), .B(n5343), .Z(n8656) );
  NOR U5752 ( .A(n8501), .B(n8656), .Z(n5910) );
  IV U5753 ( .A(x[284]), .Z(n5345) );
  NOR U5754 ( .A(n5345), .B(n6065), .Z(n5376) );
  IV U5755 ( .A(x[156]), .Z(n5346) );
  NOR U5756 ( .A(n6051), .B(n5346), .Z(n5373) );
  IV U5757 ( .A(x[28]), .Z(n5347) );
  NOR U5758 ( .A(n5347), .B(n6052), .Z(n5370) );
  IV U5759 ( .A(x[60]), .Z(n5348) );
  NOR U5760 ( .A(n6067), .B(n5348), .Z(n5367) );
  IV U5761 ( .A(x[252]), .Z(n5349) );
  NOR U5762 ( .A(n6057), .B(n5349), .Z(n5364) );
  IV U5763 ( .A(x[92]), .Z(n5350) );
  NOR U5764 ( .A(n6059), .B(n5350), .Z(n5353) );
  IV U5765 ( .A(x[124]), .Z(n5351) );
  NOR U5766 ( .A(n6061), .B(n5351), .Z(n5352) );
  NOR U5767 ( .A(n5353), .B(n5352), .Z(n5354) );
  IV U5768 ( .A(n5354), .Z(n5361) );
  IV U5769 ( .A(x[220]), .Z(n5355) );
  NOR U5770 ( .A(n6055), .B(n5355), .Z(n5358) );
  IV U5771 ( .A(x[188]), .Z(n5356) );
  NOR U5772 ( .A(n6048), .B(n5356), .Z(n5357) );
  NOR U5773 ( .A(n5358), .B(n5357), .Z(n5359) );
  IV U5774 ( .A(n5359), .Z(n5360) );
  NOR U5775 ( .A(n5361), .B(n5360), .Z(n5362) );
  IV U5776 ( .A(n5362), .Z(n5363) );
  NOR U5777 ( .A(n5364), .B(n5363), .Z(n5365) );
  IV U5778 ( .A(n5365), .Z(n5366) );
  NOR U5779 ( .A(n5367), .B(n5366), .Z(n5368) );
  IV U5780 ( .A(n5368), .Z(n5369) );
  NOR U5781 ( .A(n5370), .B(n5369), .Z(n5371) );
  IV U5782 ( .A(n5371), .Z(n5372) );
  NOR U5783 ( .A(n5373), .B(n5372), .Z(n5374) );
  IV U5784 ( .A(n5374), .Z(n5375) );
  NOR U5785 ( .A(n5376), .B(n5375), .Z(n6450) );
  NOR U5786 ( .A(n9593), .B(n6450), .Z(n5377) );
  IV U5787 ( .A(n5377), .Z(n6269) );
  XOR U5788 ( .A(n6269), .B(sum[29]), .Z(n5911) );
  XOR U5789 ( .A(n5910), .B(n5911), .Z(n5913) );
  XOR U5790 ( .A(n5912), .B(n5913), .Z(n5957) );
  IV U5791 ( .A(x[166]), .Z(n5378) );
  NOR U5792 ( .A(n6048), .B(n5378), .Z(n5409) );
  IV U5793 ( .A(x[262]), .Z(n5379) );
  NOR U5794 ( .A(n6065), .B(n5379), .Z(n5406) );
  IV U5795 ( .A(x[38]), .Z(n5380) );
  NOR U5796 ( .A(n6067), .B(n5380), .Z(n5403) );
  IV U5797 ( .A(x[198]), .Z(n5381) );
  NOR U5798 ( .A(n6055), .B(n5381), .Z(n5400) );
  IV U5799 ( .A(x[230]), .Z(n5382) );
  NOR U5800 ( .A(n6057), .B(n5382), .Z(n5397) );
  IV U5801 ( .A(x[70]), .Z(n5383) );
  NOR U5802 ( .A(n6059), .B(n5383), .Z(n5386) );
  IV U5803 ( .A(x[102]), .Z(n5384) );
  NOR U5804 ( .A(n6061), .B(n5384), .Z(n5385) );
  NOR U5805 ( .A(n5386), .B(n5385), .Z(n5387) );
  IV U5806 ( .A(n5387), .Z(n5394) );
  IV U5807 ( .A(x[134]), .Z(n5388) );
  NOR U5808 ( .A(n6051), .B(n5388), .Z(n5391) );
  IV U5809 ( .A(x[6]), .Z(n5389) );
  NOR U5810 ( .A(n6052), .B(n5389), .Z(n5390) );
  NOR U5811 ( .A(n5391), .B(n5390), .Z(n5392) );
  IV U5812 ( .A(n5392), .Z(n5393) );
  NOR U5813 ( .A(n5394), .B(n5393), .Z(n5395) );
  IV U5814 ( .A(n5395), .Z(n5396) );
  NOR U5815 ( .A(n5397), .B(n5396), .Z(n5398) );
  IV U5816 ( .A(n5398), .Z(n5399) );
  NOR U5817 ( .A(n5400), .B(n5399), .Z(n5401) );
  IV U5818 ( .A(n5401), .Z(n5402) );
  NOR U5819 ( .A(n5403), .B(n5402), .Z(n5404) );
  IV U5820 ( .A(n5404), .Z(n5405) );
  NOR U5821 ( .A(n5406), .B(n5405), .Z(n5407) );
  IV U5822 ( .A(n5407), .Z(n5408) );
  NOR U5823 ( .A(n5409), .B(n5408), .Z(n9336) );
  IV U5824 ( .A(y[247]), .Z(n5410) );
  NOR U5825 ( .A(n6205), .B(n5410), .Z(n5441) );
  IV U5826 ( .A(y[279]), .Z(n5411) );
  NOR U5827 ( .A(n6197), .B(n5411), .Z(n5438) );
  IV U5828 ( .A(y[55]), .Z(n5412) );
  NOR U5829 ( .A(n5412), .B(n6207), .Z(n5435) );
  IV U5830 ( .A(y[215]), .Z(n5413) );
  NOR U5831 ( .A(n6203), .B(n5413), .Z(n5432) );
  IV U5832 ( .A(y[183]), .Z(n5414) );
  NOR U5833 ( .A(n6199), .B(n5414), .Z(n5429) );
  IV U5834 ( .A(y[87]), .Z(n5415) );
  NOR U5835 ( .A(n6216), .B(n5415), .Z(n5418) );
  IV U5836 ( .A(y[119]), .Z(n5416) );
  NOR U5837 ( .A(n6209), .B(n5416), .Z(n5417) );
  NOR U5838 ( .A(n5418), .B(n5417), .Z(n5419) );
  IV U5839 ( .A(n5419), .Z(n5426) );
  IV U5840 ( .A(y[151]), .Z(n5420) );
  NOR U5841 ( .A(n6214), .B(n5420), .Z(n5423) );
  IV U5842 ( .A(y[23]), .Z(n5421) );
  NOR U5843 ( .A(n6200), .B(n5421), .Z(n5422) );
  NOR U5844 ( .A(n5423), .B(n5422), .Z(n5424) );
  IV U5845 ( .A(n5424), .Z(n5425) );
  NOR U5846 ( .A(n5426), .B(n5425), .Z(n5427) );
  IV U5847 ( .A(n5427), .Z(n5428) );
  NOR U5848 ( .A(n5429), .B(n5428), .Z(n5430) );
  IV U5849 ( .A(n5430), .Z(n5431) );
  NOR U5850 ( .A(n5432), .B(n5431), .Z(n5433) );
  IV U5851 ( .A(n5433), .Z(n5434) );
  NOR U5852 ( .A(n5435), .B(n5434), .Z(n5436) );
  IV U5853 ( .A(n5436), .Z(n5437) );
  NOR U5854 ( .A(n5438), .B(n5437), .Z(n5439) );
  IV U5855 ( .A(n5439), .Z(n5440) );
  NOR U5856 ( .A(n5441), .B(n5440), .Z(n7321) );
  NOR U5857 ( .A(n9336), .B(n7321), .Z(n5507) );
  IV U5858 ( .A(x[231]), .Z(n5442) );
  NOR U5859 ( .A(n5442), .B(n6057), .Z(n5473) );
  IV U5860 ( .A(x[167]), .Z(n5443) );
  NOR U5861 ( .A(n6048), .B(n5443), .Z(n5470) );
  IV U5862 ( .A(x[103]), .Z(n5444) );
  NOR U5863 ( .A(n5444), .B(n6061), .Z(n5467) );
  IV U5864 ( .A(x[7]), .Z(n5445) );
  NOR U5865 ( .A(n6052), .B(n5445), .Z(n5464) );
  IV U5866 ( .A(x[263]), .Z(n5446) );
  NOR U5867 ( .A(n5446), .B(n6065), .Z(n5461) );
  IV U5868 ( .A(x[199]), .Z(n5447) );
  NOR U5869 ( .A(n6055), .B(n5447), .Z(n5450) );
  IV U5870 ( .A(x[39]), .Z(n5448) );
  NOR U5871 ( .A(n6067), .B(n5448), .Z(n5449) );
  NOR U5872 ( .A(n5450), .B(n5449), .Z(n5451) );
  IV U5873 ( .A(n5451), .Z(n5458) );
  IV U5874 ( .A(x[71]), .Z(n5452) );
  NOR U5875 ( .A(n6059), .B(n5452), .Z(n5455) );
  IV U5876 ( .A(x[135]), .Z(n5453) );
  NOR U5877 ( .A(n5453), .B(n6051), .Z(n5454) );
  NOR U5878 ( .A(n5455), .B(n5454), .Z(n5456) );
  IV U5879 ( .A(n5456), .Z(n5457) );
  NOR U5880 ( .A(n5458), .B(n5457), .Z(n5459) );
  IV U5881 ( .A(n5459), .Z(n5460) );
  NOR U5882 ( .A(n5461), .B(n5460), .Z(n5462) );
  IV U5883 ( .A(n5462), .Z(n5463) );
  NOR U5884 ( .A(n5464), .B(n5463), .Z(n5465) );
  IV U5885 ( .A(n5465), .Z(n5466) );
  NOR U5886 ( .A(n5467), .B(n5466), .Z(n5468) );
  IV U5887 ( .A(n5468), .Z(n5469) );
  NOR U5888 ( .A(n5470), .B(n5469), .Z(n5471) );
  IV U5889 ( .A(n5471), .Z(n5472) );
  NOR U5890 ( .A(n5473), .B(n5472), .Z(n9260) );
  IV U5891 ( .A(y[246]), .Z(n5474) );
  NOR U5892 ( .A(n5474), .B(n6205), .Z(n5505) );
  IV U5893 ( .A(y[150]), .Z(n5475) );
  NOR U5894 ( .A(n6214), .B(n5475), .Z(n5502) );
  IV U5895 ( .A(y[54]), .Z(n5476) );
  NOR U5896 ( .A(n5476), .B(n6207), .Z(n5499) );
  IV U5897 ( .A(y[22]), .Z(n5477) );
  NOR U5898 ( .A(n6200), .B(n5477), .Z(n5496) );
  IV U5899 ( .A(y[278]), .Z(n5478) );
  NOR U5900 ( .A(n6197), .B(n5478), .Z(n5493) );
  IV U5901 ( .A(y[214]), .Z(n5479) );
  NOR U5902 ( .A(n5479), .B(n6203), .Z(n5482) );
  IV U5903 ( .A(y[118]), .Z(n5480) );
  NOR U5904 ( .A(n5480), .B(n6209), .Z(n5481) );
  NOR U5905 ( .A(n5482), .B(n5481), .Z(n5483) );
  IV U5906 ( .A(n5483), .Z(n5490) );
  IV U5907 ( .A(y[182]), .Z(n5484) );
  NOR U5908 ( .A(n6199), .B(n5484), .Z(n5487) );
  IV U5909 ( .A(y[86]), .Z(n5485) );
  NOR U5910 ( .A(n6216), .B(n5485), .Z(n5486) );
  NOR U5911 ( .A(n5487), .B(n5486), .Z(n5488) );
  IV U5912 ( .A(n5488), .Z(n5489) );
  NOR U5913 ( .A(n5490), .B(n5489), .Z(n5491) );
  IV U5914 ( .A(n5491), .Z(n5492) );
  NOR U5915 ( .A(n5493), .B(n5492), .Z(n5494) );
  IV U5916 ( .A(n5494), .Z(n5495) );
  NOR U5917 ( .A(n5496), .B(n5495), .Z(n5497) );
  IV U5918 ( .A(n5497), .Z(n5498) );
  NOR U5919 ( .A(n5499), .B(n5498), .Z(n5500) );
  IV U5920 ( .A(n5500), .Z(n5501) );
  NOR U5921 ( .A(n5502), .B(n5501), .Z(n5503) );
  IV U5922 ( .A(n5503), .Z(n5504) );
  NOR U5923 ( .A(n5505), .B(n5504), .Z(n7529) );
  NOR U5924 ( .A(n9260), .B(n7529), .Z(n5506) );
  XOR U5925 ( .A(n5507), .B(n5506), .Z(n5866) );
  IV U5926 ( .A(y[181]), .Z(n5508) );
  NOR U5927 ( .A(n6199), .B(n5508), .Z(n5539) );
  IV U5928 ( .A(y[149]), .Z(n5509) );
  NOR U5929 ( .A(n6214), .B(n5509), .Z(n5536) );
  IV U5930 ( .A(y[21]), .Z(n5510) );
  NOR U5931 ( .A(n6200), .B(n5510), .Z(n5533) );
  IV U5932 ( .A(y[213]), .Z(n5511) );
  NOR U5933 ( .A(n6203), .B(n5511), .Z(n5530) );
  IV U5934 ( .A(y[245]), .Z(n5512) );
  NOR U5935 ( .A(n6205), .B(n5512), .Z(n5527) );
  IV U5936 ( .A(y[85]), .Z(n5513) );
  NOR U5937 ( .A(n6216), .B(n5513), .Z(n5516) );
  IV U5938 ( .A(y[53]), .Z(n5514) );
  NOR U5939 ( .A(n6207), .B(n5514), .Z(n5515) );
  NOR U5940 ( .A(n5516), .B(n5515), .Z(n5517) );
  IV U5941 ( .A(n5517), .Z(n5524) );
  IV U5942 ( .A(y[117]), .Z(n5518) );
  NOR U5943 ( .A(n6209), .B(n5518), .Z(n5521) );
  IV U5944 ( .A(y[277]), .Z(n5519) );
  NOR U5945 ( .A(n5519), .B(n6197), .Z(n5520) );
  NOR U5946 ( .A(n5521), .B(n5520), .Z(n5522) );
  IV U5947 ( .A(n5522), .Z(n5523) );
  NOR U5948 ( .A(n5524), .B(n5523), .Z(n5525) );
  IV U5949 ( .A(n5525), .Z(n5526) );
  NOR U5950 ( .A(n5527), .B(n5526), .Z(n5528) );
  IV U5951 ( .A(n5528), .Z(n5529) );
  NOR U5952 ( .A(n5530), .B(n5529), .Z(n5531) );
  IV U5953 ( .A(n5531), .Z(n5532) );
  NOR U5954 ( .A(n5533), .B(n5532), .Z(n5534) );
  IV U5955 ( .A(n5534), .Z(n5535) );
  NOR U5956 ( .A(n5536), .B(n5535), .Z(n5537) );
  IV U5957 ( .A(n5537), .Z(n5538) );
  NOR U5958 ( .A(n5539), .B(n5538), .Z(n7714) );
  NOR U5959 ( .A(n9316), .B(n7714), .Z(n5540) );
  IV U5960 ( .A(n5540), .Z(n5867) );
  XOR U5961 ( .A(n5866), .B(n5867), .Z(n5956) );
  XOR U5962 ( .A(n5957), .B(n5956), .Z(n5958) );
  IV U5963 ( .A(x[271]), .Z(n5541) );
  NOR U5964 ( .A(n6065), .B(n5541), .Z(n5572) );
  IV U5965 ( .A(x[143]), .Z(n5542) );
  NOR U5966 ( .A(n6051), .B(n5542), .Z(n5569) );
  IV U5967 ( .A(x[111]), .Z(n5543) );
  NOR U5968 ( .A(n6061), .B(n5543), .Z(n5566) );
  IV U5969 ( .A(x[47]), .Z(n5544) );
  NOR U5970 ( .A(n6067), .B(n5544), .Z(n5563) );
  IV U5971 ( .A(x[239]), .Z(n5545) );
  NOR U5972 ( .A(n6057), .B(n5545), .Z(n5560) );
  IV U5973 ( .A(x[79]), .Z(n5546) );
  NOR U5974 ( .A(n6059), .B(n5546), .Z(n5549) );
  IV U5975 ( .A(x[207]), .Z(n5547) );
  NOR U5976 ( .A(n6055), .B(n5547), .Z(n5548) );
  NOR U5977 ( .A(n5549), .B(n5548), .Z(n5550) );
  IV U5978 ( .A(n5550), .Z(n5557) );
  IV U5979 ( .A(x[15]), .Z(n5551) );
  NOR U5980 ( .A(n6052), .B(n5551), .Z(n5554) );
  IV U5981 ( .A(x[175]), .Z(n5552) );
  NOR U5982 ( .A(n6048), .B(n5552), .Z(n5553) );
  NOR U5983 ( .A(n5554), .B(n5553), .Z(n5555) );
  IV U5984 ( .A(n5555), .Z(n5556) );
  NOR U5985 ( .A(n5557), .B(n5556), .Z(n5558) );
  IV U5986 ( .A(n5558), .Z(n5559) );
  NOR U5987 ( .A(n5560), .B(n5559), .Z(n5561) );
  IV U5988 ( .A(n5561), .Z(n5562) );
  NOR U5989 ( .A(n5563), .B(n5562), .Z(n5564) );
  IV U5990 ( .A(n5564), .Z(n5565) );
  NOR U5991 ( .A(n5566), .B(n5565), .Z(n5567) );
  IV U5992 ( .A(n5567), .Z(n5568) );
  NOR U5993 ( .A(n5569), .B(n5568), .Z(n5570) );
  IV U5994 ( .A(n5570), .Z(n5571) );
  NOR U5995 ( .A(n5572), .B(n5571), .Z(n8422) );
  IV U5996 ( .A(y[238]), .Z(n5573) );
  NOR U5997 ( .A(n6205), .B(n5573), .Z(n5604) );
  IV U5998 ( .A(y[142]), .Z(n5574) );
  NOR U5999 ( .A(n6214), .B(n5574), .Z(n5601) );
  IV U6000 ( .A(y[46]), .Z(n5575) );
  NOR U6001 ( .A(n5575), .B(n6207), .Z(n5598) );
  IV U6002 ( .A(y[14]), .Z(n5576) );
  NOR U6003 ( .A(n6200), .B(n5576), .Z(n5595) );
  IV U6004 ( .A(y[270]), .Z(n5577) );
  NOR U6005 ( .A(n6197), .B(n5577), .Z(n5592) );
  IV U6006 ( .A(y[78]), .Z(n5578) );
  NOR U6007 ( .A(n6216), .B(n5578), .Z(n5581) );
  IV U6008 ( .A(y[110]), .Z(n5579) );
  NOR U6009 ( .A(n6209), .B(n5579), .Z(n5580) );
  NOR U6010 ( .A(n5581), .B(n5580), .Z(n5582) );
  IV U6011 ( .A(n5582), .Z(n5589) );
  IV U6012 ( .A(y[206]), .Z(n5583) );
  NOR U6013 ( .A(n6203), .B(n5583), .Z(n5586) );
  IV U6014 ( .A(y[174]), .Z(n5584) );
  NOR U6015 ( .A(n5584), .B(n6199), .Z(n5585) );
  NOR U6016 ( .A(n5586), .B(n5585), .Z(n5587) );
  IV U6017 ( .A(n5587), .Z(n5588) );
  NOR U6018 ( .A(n5589), .B(n5588), .Z(n5590) );
  IV U6019 ( .A(n5590), .Z(n5591) );
  NOR U6020 ( .A(n5592), .B(n5591), .Z(n5593) );
  IV U6021 ( .A(n5593), .Z(n5594) );
  NOR U6022 ( .A(n5595), .B(n5594), .Z(n5596) );
  IV U6023 ( .A(n5596), .Z(n5597) );
  NOR U6024 ( .A(n5598), .B(n5597), .Z(n5599) );
  IV U6025 ( .A(n5599), .Z(n5600) );
  NOR U6026 ( .A(n5601), .B(n5600), .Z(n5602) );
  IV U6027 ( .A(n5602), .Z(n5603) );
  NOR U6028 ( .A(n5604), .B(n5603), .Z(n8727) );
  NOR U6029 ( .A(n8422), .B(n8727), .Z(n6330) );
  IV U6030 ( .A(y[256]), .Z(n5605) );
  NOR U6031 ( .A(n5605), .B(n6197), .Z(n5636) );
  IV U6032 ( .A(y[160]), .Z(n5606) );
  NOR U6033 ( .A(n6199), .B(n5606), .Z(n5633) );
  IV U6034 ( .A(y[32]), .Z(n5607) );
  NOR U6035 ( .A(n6207), .B(n5607), .Z(n5630) );
  IV U6036 ( .A(y[64]), .Z(n5608) );
  NOR U6037 ( .A(n6216), .B(n5608), .Z(n5627) );
  IV U6038 ( .A(y[224]), .Z(n5609) );
  NOR U6039 ( .A(n6205), .B(n5609), .Z(n5624) );
  IV U6040 ( .A(y[192]), .Z(n5610) );
  NOR U6041 ( .A(n5610), .B(n6203), .Z(n5613) );
  IV U6042 ( .A(y[96]), .Z(n5611) );
  NOR U6043 ( .A(n5611), .B(n6209), .Z(n5612) );
  NOR U6044 ( .A(n5613), .B(n5612), .Z(n5614) );
  IV U6045 ( .A(n5614), .Z(n5621) );
  IV U6046 ( .A(y[128]), .Z(n5615) );
  NOR U6047 ( .A(n6214), .B(n5615), .Z(n5618) );
  IV U6048 ( .A(y[0]), .Z(n5616) );
  NOR U6049 ( .A(n6200), .B(n5616), .Z(n5617) );
  NOR U6050 ( .A(n5618), .B(n5617), .Z(n5619) );
  IV U6051 ( .A(n5619), .Z(n5620) );
  NOR U6052 ( .A(n5621), .B(n5620), .Z(n5622) );
  IV U6053 ( .A(n5622), .Z(n5623) );
  NOR U6054 ( .A(n5624), .B(n5623), .Z(n5625) );
  IV U6055 ( .A(n5625), .Z(n5626) );
  NOR U6056 ( .A(n5627), .B(n5626), .Z(n5628) );
  IV U6057 ( .A(n5628), .Z(n5629) );
  NOR U6058 ( .A(n5630), .B(n5629), .Z(n5631) );
  IV U6059 ( .A(n5631), .Z(n5632) );
  NOR U6060 ( .A(n5633), .B(n5632), .Z(n5634) );
  IV U6061 ( .A(n5634), .Z(n5635) );
  NOR U6062 ( .A(n5636), .B(n5635), .Z(n9600) );
  IV U6063 ( .A(x[253]), .Z(n5637) );
  NOR U6064 ( .A(n5637), .B(n6057), .Z(n5668) );
  IV U6065 ( .A(x[285]), .Z(n5638) );
  NOR U6066 ( .A(n6065), .B(n5638), .Z(n5665) );
  IV U6067 ( .A(x[221]), .Z(n5639) );
  NOR U6068 ( .A(n6055), .B(n5639), .Z(n5662) );
  IV U6069 ( .A(x[93]), .Z(n5640) );
  NOR U6070 ( .A(n6059), .B(n5640), .Z(n5659) );
  IV U6071 ( .A(x[189]), .Z(n5641) );
  NOR U6072 ( .A(n6048), .B(n5641), .Z(n5656) );
  IV U6073 ( .A(x[61]), .Z(n5642) );
  NOR U6074 ( .A(n6067), .B(n5642), .Z(n5645) );
  IV U6075 ( .A(x[125]), .Z(n5643) );
  NOR U6076 ( .A(n6061), .B(n5643), .Z(n5644) );
  NOR U6077 ( .A(n5645), .B(n5644), .Z(n5646) );
  IV U6078 ( .A(n5646), .Z(n5653) );
  IV U6079 ( .A(x[157]), .Z(n5647) );
  NOR U6080 ( .A(n6051), .B(n5647), .Z(n5650) );
  IV U6081 ( .A(x[29]), .Z(n5648) );
  NOR U6082 ( .A(n6052), .B(n5648), .Z(n5649) );
  NOR U6083 ( .A(n5650), .B(n5649), .Z(n5651) );
  IV U6084 ( .A(n5651), .Z(n5652) );
  NOR U6085 ( .A(n5653), .B(n5652), .Z(n5654) );
  IV U6086 ( .A(n5654), .Z(n5655) );
  NOR U6087 ( .A(n5656), .B(n5655), .Z(n5657) );
  IV U6088 ( .A(n5657), .Z(n5658) );
  NOR U6089 ( .A(n5659), .B(n5658), .Z(n5660) );
  IV U6090 ( .A(n5660), .Z(n5661) );
  NOR U6091 ( .A(n5662), .B(n5661), .Z(n5663) );
  IV U6092 ( .A(n5663), .Z(n5664) );
  NOR U6093 ( .A(n5665), .B(n5664), .Z(n5666) );
  IV U6094 ( .A(n5666), .Z(n5667) );
  NOR U6095 ( .A(n5668), .B(n5667), .Z(n6094) );
  NOR U6096 ( .A(n9600), .B(n6094), .Z(n5669) );
  IV U6097 ( .A(n5669), .Z(n6331) );
  XOR U6098 ( .A(n6330), .B(n6331), .Z(n6334) );
  IV U6099 ( .A(x[224]), .Z(n5670) );
  NOR U6100 ( .A(n5670), .B(n6057), .Z(n5701) );
  IV U6101 ( .A(x[160]), .Z(n5671) );
  NOR U6102 ( .A(n6048), .B(n5671), .Z(n5698) );
  IV U6103 ( .A(x[0]), .Z(n5672) );
  NOR U6104 ( .A(n5672), .B(n6052), .Z(n5695) );
  IV U6105 ( .A(x[32]), .Z(n5673) );
  NOR U6106 ( .A(n6067), .B(n5673), .Z(n5692) );
  IV U6107 ( .A(x[192]), .Z(n5674) );
  NOR U6108 ( .A(n6055), .B(n5674), .Z(n5689) );
  IV U6109 ( .A(x[64]), .Z(n5675) );
  NOR U6110 ( .A(n6059), .B(n5675), .Z(n5678) );
  IV U6111 ( .A(x[96]), .Z(n5676) );
  NOR U6112 ( .A(n6061), .B(n5676), .Z(n5677) );
  NOR U6113 ( .A(n5678), .B(n5677), .Z(n5679) );
  IV U6114 ( .A(n5679), .Z(n5686) );
  IV U6115 ( .A(x[128]), .Z(n5680) );
  NOR U6116 ( .A(n6051), .B(n5680), .Z(n5683) );
  IV U6117 ( .A(x[256]), .Z(n5681) );
  NOR U6118 ( .A(n6065), .B(n5681), .Z(n5682) );
  NOR U6119 ( .A(n5683), .B(n5682), .Z(n5684) );
  IV U6120 ( .A(n5684), .Z(n5685) );
  NOR U6121 ( .A(n5686), .B(n5685), .Z(n5687) );
  IV U6122 ( .A(n5687), .Z(n5688) );
  NOR U6123 ( .A(n5689), .B(n5688), .Z(n5690) );
  IV U6124 ( .A(n5690), .Z(n5691) );
  NOR U6125 ( .A(n5692), .B(n5691), .Z(n5693) );
  IV U6126 ( .A(n5693), .Z(n5694) );
  NOR U6127 ( .A(n5695), .B(n5694), .Z(n5696) );
  IV U6128 ( .A(n5696), .Z(n5697) );
  NOR U6129 ( .A(n5698), .B(n5697), .Z(n5699) );
  IV U6130 ( .A(n5699), .Z(n5700) );
  NOR U6131 ( .A(n5701), .B(n5700), .Z(n9592) );
  IV U6132 ( .A(y[253]), .Z(n5702) );
  NOR U6133 ( .A(n6205), .B(n5702), .Z(n5733) );
  IV U6134 ( .A(y[189]), .Z(n5703) );
  NOR U6135 ( .A(n6199), .B(n5703), .Z(n5730) );
  IV U6136 ( .A(y[29]), .Z(n5704) );
  NOR U6137 ( .A(n6200), .B(n5704), .Z(n5727) );
  IV U6138 ( .A(y[221]), .Z(n5705) );
  NOR U6139 ( .A(n6203), .B(n5705), .Z(n5724) );
  IV U6140 ( .A(y[285]), .Z(n5706) );
  NOR U6141 ( .A(n6197), .B(n5706), .Z(n5721) );
  IV U6142 ( .A(y[93]), .Z(n5707) );
  NOR U6143 ( .A(n6216), .B(n5707), .Z(n5710) );
  IV U6144 ( .A(y[61]), .Z(n5708) );
  NOR U6145 ( .A(n6207), .B(n5708), .Z(n5709) );
  NOR U6146 ( .A(n5710), .B(n5709), .Z(n5711) );
  IV U6147 ( .A(n5711), .Z(n5718) );
  IV U6148 ( .A(y[157]), .Z(n5712) );
  NOR U6149 ( .A(n5712), .B(n6214), .Z(n5715) );
  IV U6150 ( .A(y[125]), .Z(n5713) );
  NOR U6151 ( .A(n5713), .B(n6209), .Z(n5714) );
  NOR U6152 ( .A(n5715), .B(n5714), .Z(n5716) );
  IV U6153 ( .A(n5716), .Z(n5717) );
  NOR U6154 ( .A(n5718), .B(n5717), .Z(n5719) );
  IV U6155 ( .A(n5719), .Z(n5720) );
  NOR U6156 ( .A(n5721), .B(n5720), .Z(n5722) );
  IV U6157 ( .A(n5722), .Z(n5723) );
  NOR U6158 ( .A(n5724), .B(n5723), .Z(n5725) );
  IV U6159 ( .A(n5725), .Z(n5726) );
  NOR U6160 ( .A(n5727), .B(n5726), .Z(n5728) );
  IV U6161 ( .A(n5728), .Z(n5729) );
  NOR U6162 ( .A(n5730), .B(n5729), .Z(n5731) );
  IV U6163 ( .A(n5731), .Z(n5732) );
  NOR U6164 ( .A(n5733), .B(n5732), .Z(n6187) );
  NOR U6165 ( .A(n9592), .B(n6187), .Z(n5734) );
  IV U6166 ( .A(n5734), .Z(n6333) );
  XOR U6167 ( .A(n6334), .B(n6333), .Z(n5951) );
  IV U6168 ( .A(y[235]), .Z(n5735) );
  NOR U6169 ( .A(n6205), .B(n5735), .Z(n5766) );
  IV U6170 ( .A(y[267]), .Z(n5736) );
  NOR U6171 ( .A(n6197), .B(n5736), .Z(n5763) );
  IV U6172 ( .A(y[107]), .Z(n5737) );
  NOR U6173 ( .A(n5737), .B(n6209), .Z(n5760) );
  IV U6174 ( .A(y[75]), .Z(n5738) );
  NOR U6175 ( .A(n6216), .B(n5738), .Z(n5757) );
  IV U6176 ( .A(y[171]), .Z(n5739) );
  NOR U6177 ( .A(n6199), .B(n5739), .Z(n5754) );
  IV U6178 ( .A(y[203]), .Z(n5740) );
  NOR U6179 ( .A(n6203), .B(n5740), .Z(n5743) );
  IV U6180 ( .A(y[43]), .Z(n5741) );
  NOR U6181 ( .A(n6207), .B(n5741), .Z(n5742) );
  NOR U6182 ( .A(n5743), .B(n5742), .Z(n5744) );
  IV U6183 ( .A(n5744), .Z(n5751) );
  IV U6184 ( .A(y[139]), .Z(n5745) );
  NOR U6185 ( .A(n6214), .B(n5745), .Z(n5748) );
  IV U6186 ( .A(y[11]), .Z(n5746) );
  NOR U6187 ( .A(n6200), .B(n5746), .Z(n5747) );
  NOR U6188 ( .A(n5748), .B(n5747), .Z(n5749) );
  IV U6189 ( .A(n5749), .Z(n5750) );
  NOR U6190 ( .A(n5751), .B(n5750), .Z(n5752) );
  IV U6191 ( .A(n5752), .Z(n5753) );
  NOR U6192 ( .A(n5754), .B(n5753), .Z(n5755) );
  IV U6193 ( .A(n5755), .Z(n5756) );
  NOR U6194 ( .A(n5757), .B(n5756), .Z(n5758) );
  IV U6195 ( .A(n5758), .Z(n5759) );
  NOR U6196 ( .A(n5760), .B(n5759), .Z(n5761) );
  IV U6197 ( .A(n5761), .Z(n5762) );
  NOR U6198 ( .A(n5763), .B(n5762), .Z(n5764) );
  IV U6199 ( .A(n5764), .Z(n5765) );
  NOR U6200 ( .A(n5766), .B(n5765), .Z(n9080) );
  IV U6201 ( .A(x[274]), .Z(n5767) );
  NOR U6202 ( .A(n6065), .B(n5767), .Z(n5798) );
  IV U6203 ( .A(x[146]), .Z(n5768) );
  NOR U6204 ( .A(n6051), .B(n5768), .Z(n5795) );
  IV U6205 ( .A(x[50]), .Z(n5769) );
  NOR U6206 ( .A(n5769), .B(n6067), .Z(n5792) );
  IV U6207 ( .A(x[210]), .Z(n5770) );
  NOR U6208 ( .A(n6055), .B(n5770), .Z(n5789) );
  IV U6209 ( .A(x[242]), .Z(n5771) );
  NOR U6210 ( .A(n6057), .B(n5771), .Z(n5786) );
  IV U6211 ( .A(x[82]), .Z(n5772) );
  NOR U6212 ( .A(n6059), .B(n5772), .Z(n5775) );
  IV U6213 ( .A(x[114]), .Z(n5773) );
  NOR U6214 ( .A(n6061), .B(n5773), .Z(n5774) );
  NOR U6215 ( .A(n5775), .B(n5774), .Z(n5776) );
  IV U6216 ( .A(n5776), .Z(n5783) );
  IV U6217 ( .A(x[18]), .Z(n5777) );
  NOR U6218 ( .A(n6052), .B(n5777), .Z(n5780) );
  IV U6219 ( .A(x[178]), .Z(n5778) );
  NOR U6220 ( .A(n6048), .B(n5778), .Z(n5779) );
  NOR U6221 ( .A(n5780), .B(n5779), .Z(n5781) );
  IV U6222 ( .A(n5781), .Z(n5782) );
  NOR U6223 ( .A(n5783), .B(n5782), .Z(n5784) );
  IV U6224 ( .A(n5784), .Z(n5785) );
  NOR U6225 ( .A(n5786), .B(n5785), .Z(n5787) );
  IV U6226 ( .A(n5787), .Z(n5788) );
  NOR U6227 ( .A(n5789), .B(n5788), .Z(n5790) );
  IV U6228 ( .A(n5790), .Z(n5791) );
  NOR U6229 ( .A(n5792), .B(n5791), .Z(n5793) );
  IV U6230 ( .A(n5793), .Z(n5794) );
  NOR U6231 ( .A(n5795), .B(n5794), .Z(n5796) );
  IV U6232 ( .A(n5796), .Z(n5797) );
  NOR U6233 ( .A(n5798), .B(n5797), .Z(n8235) );
  NOR U6234 ( .A(n9080), .B(n8235), .Z(n5949) );
  IV U6235 ( .A(y[226]), .Z(n5799) );
  NOR U6236 ( .A(n6205), .B(n5799), .Z(n5830) );
  IV U6237 ( .A(y[130]), .Z(n5800) );
  NOR U6238 ( .A(n6214), .B(n5800), .Z(n5827) );
  IV U6239 ( .A(y[34]), .Z(n5801) );
  NOR U6240 ( .A(n5801), .B(n6207), .Z(n5824) );
  IV U6241 ( .A(y[66]), .Z(n5802) );
  NOR U6242 ( .A(n6216), .B(n5802), .Z(n5821) );
  IV U6243 ( .A(y[258]), .Z(n5803) );
  NOR U6244 ( .A(n6197), .B(n5803), .Z(n5818) );
  IV U6245 ( .A(y[2]), .Z(n5804) );
  NOR U6246 ( .A(n6200), .B(n5804), .Z(n5807) );
  IV U6247 ( .A(y[98]), .Z(n5805) );
  NOR U6248 ( .A(n6209), .B(n5805), .Z(n5806) );
  NOR U6249 ( .A(n5807), .B(n5806), .Z(n5808) );
  IV U6250 ( .A(n5808), .Z(n5815) );
  IV U6251 ( .A(y[194]), .Z(n5809) );
  NOR U6252 ( .A(n6203), .B(n5809), .Z(n5812) );
  IV U6253 ( .A(y[162]), .Z(n5810) );
  NOR U6254 ( .A(n5810), .B(n6199), .Z(n5811) );
  NOR U6255 ( .A(n5812), .B(n5811), .Z(n5813) );
  IV U6256 ( .A(n5813), .Z(n5814) );
  NOR U6257 ( .A(n5815), .B(n5814), .Z(n5816) );
  IV U6258 ( .A(n5816), .Z(n5817) );
  NOR U6259 ( .A(n5818), .B(n5817), .Z(n5819) );
  IV U6260 ( .A(n5819), .Z(n5820) );
  NOR U6261 ( .A(n5821), .B(n5820), .Z(n5822) );
  IV U6262 ( .A(n5822), .Z(n5823) );
  NOR U6263 ( .A(n5824), .B(n5823), .Z(n5825) );
  IV U6264 ( .A(n5825), .Z(n5826) );
  NOR U6265 ( .A(n5827), .B(n5826), .Z(n5828) );
  IV U6266 ( .A(n5828), .Z(n5829) );
  NOR U6267 ( .A(n5830), .B(n5829), .Z(n9571) );
  NOR U6268 ( .A(n6581), .B(n9571), .Z(n5948) );
  XOR U6269 ( .A(n5949), .B(n5948), .Z(n5831) );
  IV U6270 ( .A(n5831), .Z(n5950) );
  XOR U6271 ( .A(n5951), .B(n5950), .Z(n5960) );
  XOR U6272 ( .A(n5958), .B(n5960), .Z(n6377) );
  XOR U6273 ( .A(n5833), .B(n5832), .Z(n6376) );
  IV U6274 ( .A(n6376), .Z(n5834) );
  NOR U6275 ( .A(n6377), .B(n5834), .Z(n5835) );
  NOR U6276 ( .A(n5836), .B(n5835), .Z(n5860) );
  NOR U6277 ( .A(n5861), .B(n5860), .Z(n5864) );
  NOR U6278 ( .A(n9414), .B(n7314), .Z(n5837) );
  IV U6279 ( .A(n5837), .Z(n5839) );
  NOR U6280 ( .A(n9336), .B(n7529), .Z(n5838) );
  IV U6281 ( .A(n5838), .Z(n5865) );
  NOR U6282 ( .A(n5839), .B(n5865), .Z(n5842) );
  XOR U6283 ( .A(n5839), .B(n5838), .Z(n6393) );
  NOR U6284 ( .A(n7225), .B(n9472), .Z(n5840) );
  IV U6285 ( .A(n5840), .Z(n6392) );
  NOR U6286 ( .A(n6393), .B(n6392), .Z(n5841) );
  NOR U6287 ( .A(n5842), .B(n5841), .Z(n5856) );
  XOR U6288 ( .A(n5844), .B(n5843), .Z(n5855) );
  NOR U6289 ( .A(n5856), .B(n5855), .Z(n5859) );
  NOR U6290 ( .A(n9241), .B(n8228), .Z(n6629) );
  IV U6291 ( .A(n6629), .Z(n5847) );
  IV U6292 ( .A(n5845), .Z(n5846) );
  NOR U6293 ( .A(n5847), .B(n5846), .Z(n5854) );
  NOR U6294 ( .A(n9034), .B(n8290), .Z(n6405) );
  IV U6295 ( .A(n6405), .Z(n5848) );
  NOR U6296 ( .A(n9080), .B(n8311), .Z(n6404) );
  XOR U6297 ( .A(n5848), .B(n6404), .Z(n6406) );
  XOR U6298 ( .A(n5850), .B(n5849), .Z(n6407) );
  XOR U6299 ( .A(n6406), .B(n6407), .Z(n6511) );
  NOR U6300 ( .A(n8228), .B(n9115), .Z(n5851) );
  NOR U6301 ( .A(n9241), .B(n8069), .Z(n5936) );
  XOR U6302 ( .A(n5851), .B(n5936), .Z(n5852) );
  IV U6303 ( .A(n5852), .Z(n6512) );
  NOR U6304 ( .A(n6511), .B(n6512), .Z(n5853) );
  NOR U6305 ( .A(n5854), .B(n5853), .Z(n6412) );
  XOR U6306 ( .A(n5856), .B(n5855), .Z(n6411) );
  IV U6307 ( .A(n6411), .Z(n5857) );
  NOR U6308 ( .A(n6412), .B(n5857), .Z(n5858) );
  NOR U6309 ( .A(n5859), .B(n5858), .Z(n6384) );
  XOR U6310 ( .A(n5861), .B(n5860), .Z(n6383) );
  IV U6311 ( .A(n6383), .Z(n5862) );
  NOR U6312 ( .A(n6384), .B(n5862), .Z(n5863) );
  NOR U6313 ( .A(n5864), .B(n5863), .Z(n6427) );
  NOR U6314 ( .A(n9260), .B(n7321), .Z(n6150) );
  IV U6315 ( .A(n6150), .Z(n6255) );
  NOR U6316 ( .A(n5865), .B(n6255), .Z(n5870) );
  IV U6317 ( .A(n5866), .Z(n5868) );
  NOR U6318 ( .A(n5868), .B(n5867), .Z(n5869) );
  NOR U6319 ( .A(n5870), .B(n5869), .Z(n6295) );
  NOR U6320 ( .A(n7851), .B(n9113), .Z(n6115) );
  NOR U6321 ( .A(n6579), .B(n9493), .Z(n5871) );
  IV U6322 ( .A(n5871), .Z(n6116) );
  XOR U6323 ( .A(n6115), .B(n6116), .Z(n6119) );
  NOR U6324 ( .A(n7314), .B(n9301), .Z(n5872) );
  IV U6325 ( .A(n5872), .Z(n6118) );
  XOR U6326 ( .A(n6119), .B(n6118), .Z(n6162) );
  NOR U6327 ( .A(n7531), .B(n9202), .Z(n6160) );
  NOR U6328 ( .A(n6731), .B(n9526), .Z(n6159) );
  XOR U6329 ( .A(n6160), .B(n6159), .Z(n5873) );
  IV U6330 ( .A(n5873), .Z(n6161) );
  XOR U6331 ( .A(n6162), .B(n6161), .Z(n6293) );
  NOR U6332 ( .A(n8499), .B(n8727), .Z(n6248) );
  IV U6333 ( .A(x[190]), .Z(n5874) );
  NOR U6334 ( .A(n5874), .B(n6048), .Z(n5905) );
  IV U6335 ( .A(x[286]), .Z(n5875) );
  NOR U6336 ( .A(n6065), .B(n5875), .Z(n5902) );
  IV U6337 ( .A(x[30]), .Z(n5876) );
  NOR U6338 ( .A(n5876), .B(n6052), .Z(n5899) );
  IV U6339 ( .A(x[94]), .Z(n5877) );
  NOR U6340 ( .A(n6059), .B(n5877), .Z(n5896) );
  IV U6341 ( .A(x[254]), .Z(n5878) );
  NOR U6342 ( .A(n6057), .B(n5878), .Z(n5893) );
  IV U6343 ( .A(x[222]), .Z(n5879) );
  NOR U6344 ( .A(n6055), .B(n5879), .Z(n5882) );
  IV U6345 ( .A(x[126]), .Z(n5880) );
  NOR U6346 ( .A(n6061), .B(n5880), .Z(n5881) );
  NOR U6347 ( .A(n5882), .B(n5881), .Z(n5883) );
  IV U6348 ( .A(n5883), .Z(n5890) );
  IV U6349 ( .A(x[158]), .Z(n5884) );
  NOR U6350 ( .A(n5884), .B(n6051), .Z(n5887) );
  IV U6351 ( .A(x[62]), .Z(n5885) );
  NOR U6352 ( .A(n5885), .B(n6067), .Z(n5886) );
  NOR U6353 ( .A(n5887), .B(n5886), .Z(n5888) );
  IV U6354 ( .A(n5888), .Z(n5889) );
  NOR U6355 ( .A(n5890), .B(n5889), .Z(n5891) );
  IV U6356 ( .A(n5891), .Z(n5892) );
  NOR U6357 ( .A(n5893), .B(n5892), .Z(n5894) );
  IV U6358 ( .A(n5894), .Z(n5895) );
  NOR U6359 ( .A(n5896), .B(n5895), .Z(n5897) );
  IV U6360 ( .A(n5897), .Z(n5898) );
  NOR U6361 ( .A(n5899), .B(n5898), .Z(n5900) );
  IV U6362 ( .A(n5900), .Z(n5901) );
  NOR U6363 ( .A(n5902), .B(n5901), .Z(n5903) );
  IV U6364 ( .A(n5903), .Z(n5904) );
  NOR U6365 ( .A(n5905), .B(n5904), .Z(n6171) );
  NOR U6366 ( .A(n9600), .B(n6171), .Z(n5906) );
  IV U6367 ( .A(n5906), .Z(n6249) );
  XOR U6368 ( .A(n6248), .B(n6249), .Z(n6252) );
  NOR U6369 ( .A(n6450), .B(n9571), .Z(n5907) );
  IV U6370 ( .A(n5907), .Z(n6251) );
  XOR U6371 ( .A(n6252), .B(n6251), .Z(n6027) );
  NOR U6372 ( .A(n8422), .B(n8582), .Z(n6025) );
  NOR U6373 ( .A(n6581), .B(n9490), .Z(n6024) );
  XOR U6374 ( .A(n6025), .B(n6024), .Z(n5908) );
  IV U6375 ( .A(n5908), .Z(n6026) );
  XOR U6376 ( .A(n6027), .B(n6026), .Z(n6292) );
  XOR U6377 ( .A(n6293), .B(n6292), .Z(n5909) );
  IV U6378 ( .A(n5909), .Z(n6294) );
  XOR U6379 ( .A(n6295), .B(n6294), .Z(n5918) );
  IV U6380 ( .A(n5910), .Z(n8248) );
  NOR U6381 ( .A(n8248), .B(n5911), .Z(n5916) );
  IV U6382 ( .A(n5912), .Z(n5914) );
  NOR U6383 ( .A(n5914), .B(n5913), .Z(n5915) );
  NOR U6384 ( .A(n5916), .B(n5915), .Z(n5919) );
  IV U6385 ( .A(n5919), .Z(n5917) );
  NOR U6386 ( .A(n5918), .B(n5917), .Z(n5929) );
  XOR U6387 ( .A(n5919), .B(n5918), .Z(n6338) );
  IV U6388 ( .A(n5920), .Z(n5922) );
  NOR U6389 ( .A(n5922), .B(n5921), .Z(n5926) );
  NOR U6390 ( .A(n5924), .B(n5923), .Z(n5925) );
  NOR U6391 ( .A(n5926), .B(n5925), .Z(n5927) );
  IV U6392 ( .A(n5927), .Z(n6337) );
  NOR U6393 ( .A(n6338), .B(n6337), .Z(n5928) );
  NOR U6394 ( .A(n5929), .B(n5928), .Z(n6325) );
  NOR U6395 ( .A(n5931), .B(n5930), .Z(n5935) );
  NOR U6396 ( .A(n5933), .B(n5932), .Z(n5934) );
  NOR U6397 ( .A(n5935), .B(n5934), .Z(n5964) );
  IV U6398 ( .A(n5964), .Z(n5955) );
  IV U6399 ( .A(n5936), .Z(n7123) );
  NOR U6400 ( .A(n7891), .B(n9115), .Z(n6033) );
  IV U6401 ( .A(n6033), .Z(n6031) );
  NOR U6402 ( .A(n7123), .B(n6031), .Z(n5941) );
  IV U6403 ( .A(n5937), .Z(n5938) );
  NOR U6404 ( .A(n5939), .B(n5938), .Z(n5940) );
  NOR U6405 ( .A(n5941), .B(n5940), .Z(n5971) );
  IV U6406 ( .A(n5942), .Z(n7456) );
  NOR U6407 ( .A(n7456), .B(n5943), .Z(n5947) );
  NOR U6408 ( .A(n5945), .B(n5944), .Z(n5946) );
  NOR U6409 ( .A(n5947), .B(n5946), .Z(n5969) );
  NOR U6410 ( .A(n5949), .B(n5948), .Z(n5953) );
  NOR U6411 ( .A(n5951), .B(n5950), .Z(n5952) );
  NOR U6412 ( .A(n5953), .B(n5952), .Z(n5967) );
  XOR U6413 ( .A(n5969), .B(n5967), .Z(n5970) );
  XOR U6414 ( .A(n5971), .B(n5970), .Z(n5954) );
  IV U6415 ( .A(n5954), .Z(n5963) );
  NOR U6416 ( .A(n5955), .B(n5963), .Z(n5966) );
  NOR U6417 ( .A(n5957), .B(n5956), .Z(n5962) );
  IV U6418 ( .A(n5958), .Z(n5959) );
  NOR U6419 ( .A(n5960), .B(n5959), .Z(n5961) );
  NOR U6420 ( .A(n5962), .B(n5961), .Z(n6353) );
  XOR U6421 ( .A(n5964), .B(n5963), .Z(n6352) );
  NOR U6422 ( .A(n6353), .B(n6352), .Z(n5965) );
  NOR U6423 ( .A(n5966), .B(n5965), .Z(n6323) );
  IV U6424 ( .A(n5967), .Z(n5968) );
  NOR U6425 ( .A(n5969), .B(n5968), .Z(n5973) );
  NOR U6426 ( .A(n5971), .B(n5970), .Z(n5972) );
  NOR U6427 ( .A(n5973), .B(n5972), .Z(n6321) );
  NOR U6428 ( .A(n8290), .B(n8656), .Z(n6122) );
  IV U6429 ( .A(y[286]), .Z(n5974) );
  NOR U6430 ( .A(n5974), .B(n6197), .Z(n6005) );
  IV U6431 ( .A(y[158]), .Z(n5975) );
  NOR U6432 ( .A(n6214), .B(n5975), .Z(n6002) );
  IV U6433 ( .A(y[94]), .Z(n5976) );
  NOR U6434 ( .A(n6216), .B(n5976), .Z(n5999) );
  IV U6435 ( .A(y[222]), .Z(n5977) );
  NOR U6436 ( .A(n6203), .B(n5977), .Z(n5996) );
  IV U6437 ( .A(y[254]), .Z(n5978) );
  NOR U6438 ( .A(n6205), .B(n5978), .Z(n5993) );
  IV U6439 ( .A(y[30]), .Z(n5979) );
  NOR U6440 ( .A(n6200), .B(n5979), .Z(n5982) );
  IV U6441 ( .A(y[62]), .Z(n5980) );
  NOR U6442 ( .A(n6207), .B(n5980), .Z(n5981) );
  NOR U6443 ( .A(n5982), .B(n5981), .Z(n5983) );
  IV U6444 ( .A(n5983), .Z(n5990) );
  IV U6445 ( .A(y[190]), .Z(n5984) );
  NOR U6446 ( .A(n5984), .B(n6199), .Z(n5987) );
  IV U6447 ( .A(y[126]), .Z(n5985) );
  NOR U6448 ( .A(n5985), .B(n6209), .Z(n5986) );
  NOR U6449 ( .A(n5987), .B(n5986), .Z(n5988) );
  IV U6450 ( .A(n5988), .Z(n5989) );
  NOR U6451 ( .A(n5990), .B(n5989), .Z(n5991) );
  IV U6452 ( .A(n5991), .Z(n5992) );
  NOR U6453 ( .A(n5993), .B(n5992), .Z(n5994) );
  IV U6454 ( .A(n5994), .Z(n5995) );
  NOR U6455 ( .A(n5996), .B(n5995), .Z(n5997) );
  IV U6456 ( .A(n5997), .Z(n5998) );
  NOR U6457 ( .A(n5999), .B(n5998), .Z(n6000) );
  IV U6458 ( .A(n6000), .Z(n6001) );
  NOR U6459 ( .A(n6002), .B(n6001), .Z(n6003) );
  IV U6460 ( .A(n6003), .Z(n6004) );
  NOR U6461 ( .A(n6005), .B(n6004), .Z(n6180) );
  NOR U6462 ( .A(n9592), .B(n6180), .Z(n6006) );
  IV U6463 ( .A(n6006), .Z(n6123) );
  XOR U6464 ( .A(n6122), .B(n6123), .Z(n6126) );
  NOR U6465 ( .A(n6728), .B(n9472), .Z(n6007) );
  IV U6466 ( .A(n6007), .Z(n6125) );
  XOR U6467 ( .A(n6126), .B(n6125), .Z(n6144) );
  NOR U6468 ( .A(n8228), .B(n8754), .Z(n6142) );
  NOR U6469 ( .A(n9414), .B(n6957), .Z(n6141) );
  XOR U6470 ( .A(n6142), .B(n6141), .Z(n6008) );
  IV U6471 ( .A(n6008), .Z(n6143) );
  XOR U6472 ( .A(n6144), .B(n6143), .Z(n6020) );
  NOR U6473 ( .A(n9429), .B(n7225), .Z(n6165) );
  NOR U6474 ( .A(n8068), .B(n9080), .Z(n6009) );
  IV U6475 ( .A(n6009), .Z(n6166) );
  XOR U6476 ( .A(n6165), .B(n6166), .Z(n6168) );
  NOR U6477 ( .A(n9599), .B(n6187), .Z(n6010) );
  IV U6478 ( .A(n6010), .Z(n6167) );
  XOR U6479 ( .A(n6168), .B(n6167), .Z(n6138) );
  NOR U6480 ( .A(n8948), .B(n8235), .Z(n6136) );
  NOR U6481 ( .A(n6368), .B(n9584), .Z(n6135) );
  XOR U6482 ( .A(n6136), .B(n6135), .Z(n6011) );
  IV U6483 ( .A(n6011), .Z(n6137) );
  XOR U6484 ( .A(n6138), .B(n6137), .Z(n6019) );
  NOR U6485 ( .A(n6020), .B(n6019), .Z(n6023) );
  IV U6486 ( .A(n6012), .Z(n6014) );
  NOR U6487 ( .A(n6014), .B(n6013), .Z(n6018) );
  NOR U6488 ( .A(n6016), .B(n6015), .Z(n6017) );
  NOR U6489 ( .A(n6018), .B(n6017), .Z(n6327) );
  XOR U6490 ( .A(n6020), .B(n6019), .Z(n6326) );
  IV U6491 ( .A(n6326), .Z(n6021) );
  NOR U6492 ( .A(n6327), .B(n6021), .Z(n6022) );
  NOR U6493 ( .A(n6023), .B(n6022), .Z(n6319) );
  NOR U6494 ( .A(n6025), .B(n6024), .Z(n6029) );
  NOR U6495 ( .A(n6027), .B(n6026), .Z(n6028) );
  NOR U6496 ( .A(n6029), .B(n6028), .Z(n6134) );
  NOR U6497 ( .A(n6784), .B(n9388), .Z(n6030) );
  IV U6498 ( .A(n6030), .Z(n6032) );
  NOR U6499 ( .A(n6031), .B(n6032), .Z(n6036) );
  XOR U6500 ( .A(n6033), .B(n6032), .Z(n6153) );
  NOR U6501 ( .A(n9237), .B(n7772), .Z(n6034) );
  IV U6502 ( .A(n6034), .Z(n6152) );
  NOR U6503 ( .A(n6153), .B(n6152), .Z(n6035) );
  NOR U6504 ( .A(n6036), .B(n6035), .Z(n6114) );
  NOR U6505 ( .A(n8422), .B(n8501), .Z(n7698) );
  NOR U6506 ( .A(n6731), .B(n9388), .Z(n6043) );
  NOR U6507 ( .A(n8311), .B(n8727), .Z(n7365) );
  NOR U6508 ( .A(n9571), .B(n6094), .Z(n6040) );
  NOR U6509 ( .A(n7314), .B(n9202), .Z(n6037) );
  IV U6510 ( .A(n6037), .Z(n7312) );
  NOR U6511 ( .A(n8069), .B(n8754), .Z(n6038) );
  IV U6512 ( .A(n6038), .Z(n7682) );
  XOR U6513 ( .A(n7312), .B(n7682), .Z(n6039) );
  XOR U6514 ( .A(n6040), .B(n6039), .Z(n6041) );
  XOR U6515 ( .A(n7365), .B(n6041), .Z(n6042) );
  XOR U6516 ( .A(n6043), .B(n6042), .Z(n6044) );
  XOR U6517 ( .A(n7698), .B(n6044), .Z(n6045) );
  XOR U6518 ( .A(sum[31]), .B(n6045), .Z(n6112) );
  NOR U6519 ( .A(n8228), .B(n8656), .Z(n6047) );
  NOR U6520 ( .A(n9429), .B(n6957), .Z(n6046) );
  XOR U6521 ( .A(n6047), .B(n6046), .Z(n6093) );
  IV U6522 ( .A(x[191]), .Z(n6049) );
  NOR U6523 ( .A(n6049), .B(n6048), .Z(n6088) );
  IV U6524 ( .A(x[159]), .Z(n6050) );
  NOR U6525 ( .A(n6051), .B(n6050), .Z(n6085) );
  IV U6526 ( .A(x[31]), .Z(n6053) );
  NOR U6527 ( .A(n6053), .B(n6052), .Z(n6082) );
  IV U6528 ( .A(x[223]), .Z(n6054) );
  NOR U6529 ( .A(n6055), .B(n6054), .Z(n6079) );
  IV U6530 ( .A(x[255]), .Z(n6056) );
  NOR U6531 ( .A(n6057), .B(n6056), .Z(n6076) );
  IV U6532 ( .A(x[95]), .Z(n6058) );
  NOR U6533 ( .A(n6059), .B(n6058), .Z(n6063) );
  IV U6534 ( .A(x[127]), .Z(n6060) );
  NOR U6535 ( .A(n6061), .B(n6060), .Z(n6062) );
  NOR U6536 ( .A(n6063), .B(n6062), .Z(n6064) );
  IV U6537 ( .A(n6064), .Z(n6073) );
  IV U6538 ( .A(x[287]), .Z(n6066) );
  NOR U6539 ( .A(n6066), .B(n6065), .Z(n6070) );
  IV U6540 ( .A(x[63]), .Z(n6068) );
  NOR U6541 ( .A(n6068), .B(n6067), .Z(n6069) );
  NOR U6542 ( .A(n6070), .B(n6069), .Z(n6071) );
  IV U6543 ( .A(n6071), .Z(n6072) );
  NOR U6544 ( .A(n6073), .B(n6072), .Z(n6074) );
  IV U6545 ( .A(n6074), .Z(n6075) );
  NOR U6546 ( .A(n6076), .B(n6075), .Z(n6077) );
  IV U6547 ( .A(n6077), .Z(n6078) );
  NOR U6548 ( .A(n6079), .B(n6078), .Z(n6080) );
  IV U6549 ( .A(n6080), .Z(n6081) );
  NOR U6550 ( .A(n6082), .B(n6081), .Z(n6083) );
  IV U6551 ( .A(n6083), .Z(n6084) );
  NOR U6552 ( .A(n6085), .B(n6084), .Z(n6086) );
  IV U6553 ( .A(n6086), .Z(n6087) );
  NOR U6554 ( .A(n6088), .B(n6087), .Z(n6089) );
  NOR U6555 ( .A(n9600), .B(n6089), .Z(n6091) );
  NOR U6556 ( .A(n8582), .B(n8499), .Z(n6090) );
  XOR U6557 ( .A(n6091), .B(n6090), .Z(n6092) );
  XOR U6558 ( .A(n6093), .B(n6092), .Z(n6102) );
  IV U6559 ( .A(sum[30]), .Z(n6096) );
  NOR U6560 ( .A(n9593), .B(n6094), .Z(n6095) );
  IV U6561 ( .A(n6095), .Z(n6267) );
  NOR U6562 ( .A(n6096), .B(n6267), .Z(n6100) );
  NOR U6563 ( .A(n9336), .B(n6784), .Z(n6098) );
  NOR U6564 ( .A(n7225), .B(n9301), .Z(n6097) );
  XOR U6565 ( .A(n6098), .B(n6097), .Z(n6099) );
  XOR U6566 ( .A(n6100), .B(n6099), .Z(n6101) );
  XOR U6567 ( .A(n6102), .B(n6101), .Z(n6110) );
  NOR U6568 ( .A(n6728), .B(n9414), .Z(n6104) );
  NOR U6569 ( .A(n9260), .B(n7167), .Z(n6103) );
  XOR U6570 ( .A(n6104), .B(n6103), .Z(n6108) );
  NOR U6571 ( .A(n7772), .B(n9113), .Z(n6106) );
  NOR U6572 ( .A(n6581), .B(n9472), .Z(n6105) );
  XOR U6573 ( .A(n6106), .B(n6105), .Z(n6107) );
  XOR U6574 ( .A(n6108), .B(n6107), .Z(n6109) );
  XOR U6575 ( .A(n6110), .B(n6109), .Z(n6111) );
  XOR U6576 ( .A(n6112), .B(n6111), .Z(n6113) );
  XOR U6577 ( .A(n6114), .B(n6113), .Z(n6132) );
  IV U6578 ( .A(n6115), .Z(n6117) );
  NOR U6579 ( .A(n6117), .B(n6116), .Z(n6121) );
  NOR U6580 ( .A(n6119), .B(n6118), .Z(n6120) );
  NOR U6581 ( .A(n6121), .B(n6120), .Z(n6130) );
  IV U6582 ( .A(n6122), .Z(n6124) );
  NOR U6583 ( .A(n6124), .B(n6123), .Z(n6128) );
  NOR U6584 ( .A(n6126), .B(n6125), .Z(n6127) );
  NOR U6585 ( .A(n6128), .B(n6127), .Z(n6129) );
  XOR U6586 ( .A(n6130), .B(n6129), .Z(n6131) );
  XOR U6587 ( .A(n6132), .B(n6131), .Z(n6133) );
  XOR U6588 ( .A(n6134), .B(n6133), .Z(n6291) );
  NOR U6589 ( .A(n6136), .B(n6135), .Z(n6140) );
  NOR U6590 ( .A(n6138), .B(n6137), .Z(n6139) );
  NOR U6591 ( .A(n6140), .B(n6139), .Z(n6148) );
  NOR U6592 ( .A(n6142), .B(n6141), .Z(n6146) );
  NOR U6593 ( .A(n6144), .B(n6143), .Z(n6145) );
  NOR U6594 ( .A(n6146), .B(n6145), .Z(n6147) );
  XOR U6595 ( .A(n6148), .B(n6147), .Z(n6289) );
  NOR U6596 ( .A(n9316), .B(n7529), .Z(n6156) );
  IV U6597 ( .A(n6156), .Z(n6151) );
  NOR U6598 ( .A(n9034), .B(n8069), .Z(n6149) );
  IV U6599 ( .A(n6149), .Z(n8067) );
  XOR U6600 ( .A(n6150), .B(n8067), .Z(n6258) );
  NOR U6601 ( .A(n9241), .B(n7714), .Z(n6256) );
  XOR U6602 ( .A(n6258), .B(n6256), .Z(n6155) );
  NOR U6603 ( .A(n6151), .B(n6155), .Z(n6158) );
  XOR U6604 ( .A(n6153), .B(n6152), .Z(n6279) );
  NOR U6605 ( .A(n8311), .B(n8862), .Z(n6277) );
  NOR U6606 ( .A(n9336), .B(n7167), .Z(n6276) );
  XOR U6607 ( .A(n6277), .B(n6276), .Z(n6154) );
  IV U6608 ( .A(n6154), .Z(n6278) );
  XOR U6609 ( .A(n6279), .B(n6278), .Z(n6298) );
  XOR U6610 ( .A(n6156), .B(n6155), .Z(n6299) );
  NOR U6611 ( .A(n6298), .B(n6299), .Z(n6157) );
  NOR U6612 ( .A(n6158), .B(n6157), .Z(n6287) );
  NOR U6613 ( .A(n6160), .B(n6159), .Z(n6164) );
  NOR U6614 ( .A(n6162), .B(n6161), .Z(n6163) );
  NOR U6615 ( .A(n6164), .B(n6163), .Z(n6266) );
  IV U6616 ( .A(n6165), .Z(n6773) );
  NOR U6617 ( .A(n6773), .B(n6166), .Z(n6170) );
  NOR U6618 ( .A(n6168), .B(n6167), .Z(n6169) );
  NOR U6619 ( .A(n6170), .B(n6169), .Z(n6247) );
  NOR U6620 ( .A(n9593), .B(n6171), .Z(n6173) );
  NOR U6621 ( .A(n9316), .B(n7321), .Z(n6172) );
  XOR U6622 ( .A(n6173), .B(n6172), .Z(n6177) );
  NOR U6623 ( .A(n8290), .B(n8729), .Z(n6175) );
  NOR U6624 ( .A(n7891), .B(n9034), .Z(n6174) );
  XOR U6625 ( .A(n6175), .B(n6174), .Z(n6176) );
  XOR U6626 ( .A(n6177), .B(n6176), .Z(n6186) );
  NOR U6627 ( .A(n9493), .B(n6368), .Z(n6179) );
  NOR U6628 ( .A(n9241), .B(n7529), .Z(n6178) );
  XOR U6629 ( .A(n6179), .B(n6178), .Z(n6184) );
  NOR U6630 ( .A(n9599), .B(n6180), .Z(n6182) );
  NOR U6631 ( .A(n9080), .B(n7851), .Z(n6181) );
  XOR U6632 ( .A(n6182), .B(n6181), .Z(n6183) );
  XOR U6633 ( .A(n6184), .B(n6183), .Z(n6185) );
  XOR U6634 ( .A(n6186), .B(n6185), .Z(n6245) );
  NOR U6635 ( .A(n9584), .B(n6187), .Z(n6189) );
  NOR U6636 ( .A(n9490), .B(n6450), .Z(n6188) );
  XOR U6637 ( .A(n6189), .B(n6188), .Z(n6193) );
  NOR U6638 ( .A(n8862), .B(n8235), .Z(n6191) );
  NOR U6639 ( .A(n9115), .B(n7714), .Z(n6190) );
  XOR U6640 ( .A(n6191), .B(n6190), .Z(n6192) );
  XOR U6641 ( .A(n6193), .B(n6192), .Z(n6243) );
  NOR U6642 ( .A(n6579), .B(n9526), .Z(n6195) );
  NOR U6643 ( .A(n7531), .B(n9237), .Z(n6194) );
  XOR U6644 ( .A(n6195), .B(n6194), .Z(n6241) );
  IV U6645 ( .A(y[287]), .Z(n6196) );
  NOR U6646 ( .A(n6197), .B(n6196), .Z(n6236) );
  IV U6647 ( .A(y[191]), .Z(n6198) );
  NOR U6648 ( .A(n6199), .B(n6198), .Z(n6233) );
  IV U6649 ( .A(y[31]), .Z(n6201) );
  NOR U6650 ( .A(n6201), .B(n6200), .Z(n6230) );
  IV U6651 ( .A(y[223]), .Z(n6202) );
  NOR U6652 ( .A(n6203), .B(n6202), .Z(n6227) );
  IV U6653 ( .A(y[255]), .Z(n6204) );
  NOR U6654 ( .A(n6205), .B(n6204), .Z(n6224) );
  IV U6655 ( .A(y[63]), .Z(n6206) );
  NOR U6656 ( .A(n6207), .B(n6206), .Z(n6211) );
  IV U6657 ( .A(y[127]), .Z(n6208) );
  NOR U6658 ( .A(n6209), .B(n6208), .Z(n6210) );
  NOR U6659 ( .A(n6211), .B(n6210), .Z(n6212) );
  IV U6660 ( .A(n6212), .Z(n6221) );
  IV U6661 ( .A(y[159]), .Z(n6213) );
  NOR U6662 ( .A(n6214), .B(n6213), .Z(n6218) );
  IV U6663 ( .A(y[95]), .Z(n6215) );
  NOR U6664 ( .A(n6216), .B(n6215), .Z(n6217) );
  NOR U6665 ( .A(n6218), .B(n6217), .Z(n6219) );
  IV U6666 ( .A(n6219), .Z(n6220) );
  NOR U6667 ( .A(n6221), .B(n6220), .Z(n6222) );
  IV U6668 ( .A(n6222), .Z(n6223) );
  NOR U6669 ( .A(n6224), .B(n6223), .Z(n6225) );
  IV U6670 ( .A(n6225), .Z(n6226) );
  NOR U6671 ( .A(n6227), .B(n6226), .Z(n6228) );
  IV U6672 ( .A(n6228), .Z(n6229) );
  NOR U6673 ( .A(n6230), .B(n6229), .Z(n6231) );
  IV U6674 ( .A(n6231), .Z(n6232) );
  NOR U6675 ( .A(n6233), .B(n6232), .Z(n6234) );
  IV U6676 ( .A(n6234), .Z(n6235) );
  NOR U6677 ( .A(n6236), .B(n6235), .Z(n6237) );
  NOR U6678 ( .A(n9592), .B(n6237), .Z(n6239) );
  NOR U6679 ( .A(n8948), .B(n8068), .Z(n6238) );
  XOR U6680 ( .A(n6239), .B(n6238), .Z(n6240) );
  XOR U6681 ( .A(n6241), .B(n6240), .Z(n6242) );
  XOR U6682 ( .A(n6243), .B(n6242), .Z(n6244) );
  XOR U6683 ( .A(n6245), .B(n6244), .Z(n6246) );
  XOR U6684 ( .A(n6247), .B(n6246), .Z(n6264) );
  IV U6685 ( .A(n6248), .Z(n6250) );
  NOR U6686 ( .A(n6250), .B(n6249), .Z(n6254) );
  NOR U6687 ( .A(n6252), .B(n6251), .Z(n6253) );
  NOR U6688 ( .A(n6254), .B(n6253), .Z(n6262) );
  NOR U6689 ( .A(n6255), .B(n8067), .Z(n6260) );
  IV U6690 ( .A(n6256), .Z(n6257) );
  NOR U6691 ( .A(n6258), .B(n6257), .Z(n6259) );
  NOR U6692 ( .A(n6260), .B(n6259), .Z(n6261) );
  XOR U6693 ( .A(n6262), .B(n6261), .Z(n6263) );
  XOR U6694 ( .A(n6264), .B(n6263), .Z(n6265) );
  XOR U6695 ( .A(n6266), .B(n6265), .Z(n6285) );
  NOR U6696 ( .A(n8501), .B(n8729), .Z(n6272) );
  IV U6697 ( .A(n6272), .Z(n6268) );
  XOR U6698 ( .A(sum[30]), .B(n6267), .Z(n6271) );
  NOR U6699 ( .A(n6268), .B(n6271), .Z(n6275) );
  IV U6700 ( .A(sum[29]), .Z(n6270) );
  NOR U6701 ( .A(n6270), .B(n6269), .Z(n6301) );
  IV U6702 ( .A(n6301), .Z(n6273) );
  XOR U6703 ( .A(n6272), .B(n6271), .Z(n6300) );
  NOR U6704 ( .A(n6273), .B(n6300), .Z(n6274) );
  NOR U6705 ( .A(n6275), .B(n6274), .Z(n6283) );
  NOR U6706 ( .A(n6277), .B(n6276), .Z(n6281) );
  NOR U6707 ( .A(n6279), .B(n6278), .Z(n6280) );
  NOR U6708 ( .A(n6281), .B(n6280), .Z(n6282) );
  XOR U6709 ( .A(n6283), .B(n6282), .Z(n6284) );
  XOR U6710 ( .A(n6285), .B(n6284), .Z(n6286) );
  XOR U6711 ( .A(n6287), .B(n6286), .Z(n6288) );
  XOR U6712 ( .A(n6289), .B(n6288), .Z(n6290) );
  XOR U6713 ( .A(n6291), .B(n6290), .Z(n6317) );
  NOR U6714 ( .A(n6293), .B(n6292), .Z(n6297) );
  NOR U6715 ( .A(n6295), .B(n6294), .Z(n6296) );
  NOR U6716 ( .A(n6297), .B(n6296), .Z(n6315) );
  XOR U6717 ( .A(n6299), .B(n6298), .Z(n6311) );
  IV U6718 ( .A(n6311), .Z(n6302) );
  XOR U6719 ( .A(n6301), .B(n6300), .Z(n6310) );
  NOR U6720 ( .A(n6302), .B(n6310), .Z(n6313) );
  IV U6721 ( .A(n6303), .Z(n6305) );
  NOR U6722 ( .A(n6305), .B(n6304), .Z(n6309) );
  IV U6723 ( .A(n6306), .Z(n7880) );
  NOR U6724 ( .A(n7880), .B(n6307), .Z(n6308) );
  NOR U6725 ( .A(n6309), .B(n6308), .Z(n6329) );
  XOR U6726 ( .A(n6311), .B(n6310), .Z(n6328) );
  NOR U6727 ( .A(n6329), .B(n6328), .Z(n6312) );
  NOR U6728 ( .A(n6313), .B(n6312), .Z(n6314) );
  XOR U6729 ( .A(n6315), .B(n6314), .Z(n6316) );
  XOR U6730 ( .A(n6317), .B(n6316), .Z(n6318) );
  XOR U6731 ( .A(n6319), .B(n6318), .Z(n6320) );
  XOR U6732 ( .A(n6321), .B(n6320), .Z(n6322) );
  XOR U6733 ( .A(n6323), .B(n6322), .Z(n6324) );
  XOR U6734 ( .A(n6325), .B(n6324), .Z(n6425) );
  XOR U6735 ( .A(n6327), .B(n6326), .Z(n6440) );
  XOR U6736 ( .A(n6329), .B(n6328), .Z(n6436) );
  IV U6737 ( .A(n6330), .Z(n6332) );
  NOR U6738 ( .A(n6332), .B(n6331), .Z(n6336) );
  NOR U6739 ( .A(n6334), .B(n6333), .Z(n6335) );
  NOR U6740 ( .A(n6336), .B(n6335), .Z(n6438) );
  XOR U6741 ( .A(n6436), .B(n6438), .Z(n6439) );
  XOR U6742 ( .A(n6440), .B(n6439), .Z(n6355) );
  XOR U6743 ( .A(n6338), .B(n6337), .Z(n6433) );
  NOR U6744 ( .A(n6340), .B(n6339), .Z(n6344) );
  NOR U6745 ( .A(n6342), .B(n6341), .Z(n6343) );
  NOR U6746 ( .A(n6344), .B(n6343), .Z(n6429) );
  NOR U6747 ( .A(n6346), .B(n6345), .Z(n6350) );
  NOR U6748 ( .A(n6348), .B(n6347), .Z(n6349) );
  NOR U6749 ( .A(n6350), .B(n6349), .Z(n6351) );
  IV U6750 ( .A(n6351), .Z(n6430) );
  XOR U6751 ( .A(n6429), .B(n6430), .Z(n6432) );
  XOR U6752 ( .A(n6433), .B(n6432), .Z(n6354) );
  NOR U6753 ( .A(n6355), .B(n6354), .Z(n6358) );
  XOR U6754 ( .A(n6353), .B(n6352), .Z(n6508) );
  XOR U6755 ( .A(n6355), .B(n6354), .Z(n6507) );
  IV U6756 ( .A(n6507), .Z(n6356) );
  NOR U6757 ( .A(n6508), .B(n6356), .Z(n6357) );
  NOR U6758 ( .A(n6358), .B(n6357), .Z(n6423) );
  NOR U6759 ( .A(n8656), .B(n8582), .Z(n6364) );
  IV U6760 ( .A(n6364), .Z(n6360) );
  XOR U6761 ( .A(n6359), .B(sum[28]), .Z(n6363) );
  NOR U6762 ( .A(n6360), .B(n6363), .Z(n6367) );
  IV U6763 ( .A(sum[27]), .Z(n6362) );
  NOR U6764 ( .A(n9593), .B(n6728), .Z(n6361) );
  IV U6765 ( .A(n6361), .Z(n6591) );
  NOR U6766 ( .A(n6362), .B(n6591), .Z(n6514) );
  IV U6767 ( .A(n6514), .Z(n6365) );
  XOR U6768 ( .A(n6364), .B(n6363), .Z(n6513) );
  NOR U6769 ( .A(n6365), .B(n6513), .Z(n6366) );
  NOR U6770 ( .A(n6367), .B(n6366), .Z(n6379) );
  NOR U6771 ( .A(n8948), .B(n8499), .Z(n6372) );
  IV U6772 ( .A(n6372), .Z(n6370) );
  NOR U6773 ( .A(n9592), .B(n6368), .Z(n6369) );
  IV U6774 ( .A(n6369), .Z(n6371) );
  NOR U6775 ( .A(n6370), .B(n6371), .Z(n6375) );
  XOR U6776 ( .A(n6372), .B(n6371), .Z(n6480) );
  NOR U6777 ( .A(n6579), .B(n9599), .Z(n6373) );
  IV U6778 ( .A(n6373), .Z(n6479) );
  NOR U6779 ( .A(n6480), .B(n6479), .Z(n6374) );
  NOR U6780 ( .A(n6375), .B(n6374), .Z(n6378) );
  NOR U6781 ( .A(n6379), .B(n6378), .Z(n6382) );
  XOR U6782 ( .A(n6377), .B(n6376), .Z(n6463) );
  XOR U6783 ( .A(n6379), .B(n6378), .Z(n6462) );
  IV U6784 ( .A(n6462), .Z(n6380) );
  NOR U6785 ( .A(n6463), .B(n6380), .Z(n6381) );
  NOR U6786 ( .A(n6382), .B(n6381), .Z(n6418) );
  XOR U6787 ( .A(n6384), .B(n6383), .Z(n6417) );
  NOR U6788 ( .A(n6418), .B(n6417), .Z(n6421) );
  NOR U6789 ( .A(n7772), .B(n9301), .Z(n6388) );
  NOR U6790 ( .A(n7321), .B(n9388), .Z(n6387) );
  NOR U6791 ( .A(n6388), .B(n6387), .Z(n6391) );
  NOR U6792 ( .A(n9202), .B(n7851), .Z(n6398) );
  NOR U6793 ( .A(n9490), .B(n6957), .Z(n6385) );
  IV U6794 ( .A(n6385), .Z(n6399) );
  XOR U6795 ( .A(n6398), .B(n6399), .Z(n6401) );
  NOR U6796 ( .A(n9526), .B(n7167), .Z(n6386) );
  IV U6797 ( .A(n6386), .Z(n6400) );
  XOR U6798 ( .A(n6401), .B(n6400), .Z(n6532) );
  XOR U6799 ( .A(n6388), .B(n6387), .Z(n6389) );
  IV U6800 ( .A(n6389), .Z(n6533) );
  NOR U6801 ( .A(n6532), .B(n6533), .Z(n6390) );
  NOR U6802 ( .A(n6391), .B(n6390), .Z(n6414) );
  IV U6803 ( .A(n6414), .Z(n6410) );
  NOR U6804 ( .A(n8501), .B(n8754), .Z(n6394) );
  NOR U6805 ( .A(n9260), .B(n7714), .Z(n6395) );
  NOR U6806 ( .A(n6394), .B(n6395), .Z(n6397) );
  XOR U6807 ( .A(n6393), .B(n6392), .Z(n6445) );
  IV U6808 ( .A(n6394), .Z(n6750) );
  XOR U6809 ( .A(n6395), .B(n6750), .Z(n6446) );
  NOR U6810 ( .A(n6445), .B(n6446), .Z(n6396) );
  NOR U6811 ( .A(n6397), .B(n6396), .Z(n6502) );
  IV U6812 ( .A(n6398), .Z(n7849) );
  NOR U6813 ( .A(n7849), .B(n6399), .Z(n6403) );
  NOR U6814 ( .A(n6401), .B(n6400), .Z(n6402) );
  NOR U6815 ( .A(n6403), .B(n6402), .Z(n6501) );
  NOR U6816 ( .A(n6405), .B(n6404), .Z(n6409) );
  NOR U6817 ( .A(n6407), .B(n6406), .Z(n6408) );
  NOR U6818 ( .A(n6409), .B(n6408), .Z(n6499) );
  XOR U6819 ( .A(n6501), .B(n6499), .Z(n6503) );
  XOR U6820 ( .A(n6502), .B(n6503), .Z(n6413) );
  NOR U6821 ( .A(n6410), .B(n6413), .Z(n6416) );
  XOR U6822 ( .A(n6412), .B(n6411), .Z(n6467) );
  XOR U6823 ( .A(n6414), .B(n6413), .Z(n6466) );
  NOR U6824 ( .A(n6467), .B(n6466), .Z(n6415) );
  NOR U6825 ( .A(n6416), .B(n6415), .Z(n6660) );
  XOR U6826 ( .A(n6418), .B(n6417), .Z(n6419) );
  IV U6827 ( .A(n6419), .Z(n6659) );
  NOR U6828 ( .A(n6660), .B(n6659), .Z(n6420) );
  NOR U6829 ( .A(n6421), .B(n6420), .Z(n6422) );
  XOR U6830 ( .A(n6423), .B(n6422), .Z(n6424) );
  XOR U6831 ( .A(n6425), .B(n6424), .Z(n6426) );
  XOR U6832 ( .A(n6427), .B(n6426), .Z(n6428) );
  IV U6833 ( .A(n6428), .Z(n6673) );
  IV U6834 ( .A(n6429), .Z(n6431) );
  NOR U6835 ( .A(n6431), .B(n6430), .Z(n6435) );
  NOR U6836 ( .A(n6433), .B(n6432), .Z(n6434) );
  NOR U6837 ( .A(n6435), .B(n6434), .Z(n6444) );
  IV U6838 ( .A(n6436), .Z(n6437) );
  NOR U6839 ( .A(n6438), .B(n6437), .Z(n6442) );
  NOR U6840 ( .A(n6440), .B(n6439), .Z(n6441) );
  NOR U6841 ( .A(n6442), .B(n6441), .Z(n6443) );
  XOR U6842 ( .A(n6444), .B(n6443), .Z(n6671) );
  XOR U6843 ( .A(n6446), .B(n6445), .Z(n6457) );
  NOR U6844 ( .A(n8727), .B(n8729), .Z(n6488) );
  IV U6845 ( .A(n6488), .Z(n6447) );
  NOR U6846 ( .A(n9493), .B(n6784), .Z(n6487) );
  XOR U6847 ( .A(n6447), .B(n6487), .Z(n6489) );
  NOR U6848 ( .A(n6728), .B(n9571), .Z(n6448) );
  IV U6849 ( .A(n6448), .Z(n6475) );
  NOR U6850 ( .A(n8422), .B(n8862), .Z(n6449) );
  IV U6851 ( .A(n6449), .Z(n6474) );
  NOR U6852 ( .A(n9600), .B(n6450), .Z(n6472) );
  XOR U6853 ( .A(n6474), .B(n6472), .Z(n6476) );
  XOR U6854 ( .A(n6475), .B(n6476), .Z(n6490) );
  XOR U6855 ( .A(n6489), .B(n6490), .Z(n6458) );
  NOR U6856 ( .A(n6457), .B(n6458), .Z(n6461) );
  NOR U6857 ( .A(n8656), .B(n8727), .Z(n6451) );
  IV U6858 ( .A(n6451), .Z(n7118) );
  NOR U6859 ( .A(n9599), .B(n6731), .Z(n6454) );
  IV U6860 ( .A(n6454), .Z(n6452) );
  NOR U6861 ( .A(n7118), .B(n6452), .Z(n6456) );
  NOR U6862 ( .A(n9490), .B(n7225), .Z(n6453) );
  IV U6863 ( .A(n6453), .Z(n6569) );
  XOR U6864 ( .A(n6454), .B(n7118), .Z(n6568) );
  NOR U6865 ( .A(n6569), .B(n6568), .Z(n6455) );
  NOR U6866 ( .A(n6456), .B(n6455), .Z(n6615) );
  IV U6867 ( .A(n6457), .Z(n6459) );
  XOR U6868 ( .A(n6459), .B(n6458), .Z(n6614) );
  NOR U6869 ( .A(n6615), .B(n6614), .Z(n6460) );
  NOR U6870 ( .A(n6461), .B(n6460), .Z(n6465) );
  XOR U6871 ( .A(n6463), .B(n6462), .Z(n6464) );
  NOR U6872 ( .A(n6465), .B(n6464), .Z(n6471) );
  XOR U6873 ( .A(n6465), .B(n6464), .Z(n6564) );
  IV U6874 ( .A(n6564), .Z(n6469) );
  XOR U6875 ( .A(n6467), .B(n6466), .Z(n6468) );
  IV U6876 ( .A(n6468), .Z(n6565) );
  NOR U6877 ( .A(n6469), .B(n6565), .Z(n6470) );
  NOR U6878 ( .A(n6471), .B(n6470), .Z(n6551) );
  IV U6879 ( .A(n6472), .Z(n6473) );
  NOR U6880 ( .A(n6474), .B(n6473), .Z(n6478) );
  NOR U6881 ( .A(n6476), .B(n6475), .Z(n6477) );
  NOR U6882 ( .A(n6478), .B(n6477), .Z(n6495) );
  NOR U6883 ( .A(n9113), .B(n8235), .Z(n6482) );
  NOR U6884 ( .A(n6731), .B(n9584), .Z(n6481) );
  NOR U6885 ( .A(n6482), .B(n6481), .Z(n6485) );
  XOR U6886 ( .A(n6480), .B(n6479), .Z(n6531) );
  XOR U6887 ( .A(n6482), .B(n6481), .Z(n6483) );
  IV U6888 ( .A(n6483), .Z(n6530) );
  NOR U6889 ( .A(n6531), .B(n6530), .Z(n6484) );
  NOR U6890 ( .A(n6485), .B(n6484), .Z(n6494) );
  IV U6891 ( .A(n6494), .Z(n6486) );
  NOR U6892 ( .A(n6495), .B(n6486), .Z(n6497) );
  NOR U6893 ( .A(n6488), .B(n6487), .Z(n6492) );
  NOR U6894 ( .A(n6490), .B(n6489), .Z(n6491) );
  NOR U6895 ( .A(n6492), .B(n6491), .Z(n6493) );
  IV U6896 ( .A(n6493), .Z(n6510) );
  XOR U6897 ( .A(n6495), .B(n6494), .Z(n6509) );
  NOR U6898 ( .A(n6510), .B(n6509), .Z(n6496) );
  NOR U6899 ( .A(n6497), .B(n6496), .Z(n6498) );
  IV U6900 ( .A(n6498), .Z(n6559) );
  IV U6901 ( .A(n6499), .Z(n6500) );
  NOR U6902 ( .A(n6501), .B(n6500), .Z(n6506) );
  IV U6903 ( .A(n6502), .Z(n6504) );
  NOR U6904 ( .A(n6504), .B(n6503), .Z(n6505) );
  NOR U6905 ( .A(n6506), .B(n6505), .Z(n6555) );
  XOR U6906 ( .A(n6508), .B(n6507), .Z(n6557) );
  XOR U6907 ( .A(n6555), .B(n6557), .Z(n6558) );
  XOR U6908 ( .A(n6559), .B(n6558), .Z(n6550) );
  NOR U6909 ( .A(n6551), .B(n6550), .Z(n6554) );
  XOR U6910 ( .A(n6510), .B(n6509), .Z(n6529) );
  XOR U6911 ( .A(n6512), .B(n6511), .Z(n6524) );
  IV U6912 ( .A(n6524), .Z(n6515) );
  XOR U6913 ( .A(n6514), .B(n6513), .Z(n6523) );
  NOR U6914 ( .A(n6515), .B(n6523), .Z(n6526) );
  NOR U6915 ( .A(n9260), .B(n7891), .Z(n6516) );
  IV U6916 ( .A(n6516), .Z(n6519) );
  NOR U6917 ( .A(n8948), .B(n8422), .Z(n6518) );
  IV U6918 ( .A(n6518), .Z(n6517) );
  NOR U6919 ( .A(n6519), .B(n6517), .Z(n6522) );
  NOR U6920 ( .A(n9034), .B(n8501), .Z(n6631) );
  IV U6921 ( .A(n6631), .Z(n6520) );
  XOR U6922 ( .A(n6519), .B(n6518), .Z(n6630) );
  NOR U6923 ( .A(n6520), .B(n6630), .Z(n6521) );
  NOR U6924 ( .A(n6522), .B(n6521), .Z(n6617) );
  XOR U6925 ( .A(n6524), .B(n6523), .Z(n6616) );
  NOR U6926 ( .A(n6617), .B(n6616), .Z(n6525) );
  NOR U6927 ( .A(n6526), .B(n6525), .Z(n6528) );
  IV U6928 ( .A(n6528), .Z(n6527) );
  NOR U6929 ( .A(n6529), .B(n6527), .Z(n6548) );
  XOR U6930 ( .A(n6529), .B(n6528), .Z(n6920) );
  XOR U6931 ( .A(n6531), .B(n6530), .Z(n6542) );
  XOR U6932 ( .A(n6533), .B(n6532), .Z(n6541) );
  NOR U6933 ( .A(n6542), .B(n6541), .Z(n6545) );
  NOR U6934 ( .A(n8068), .B(n9202), .Z(n6538) );
  IV U6935 ( .A(n6538), .Z(n6535) );
  NOR U6936 ( .A(n9493), .B(n7167), .Z(n6534) );
  IV U6937 ( .A(n6534), .Z(n6537) );
  NOR U6938 ( .A(n6535), .B(n6537), .Z(n6540) );
  NOR U6939 ( .A(n9526), .B(n7321), .Z(n6536) );
  IV U6940 ( .A(n6536), .Z(n6644) );
  XOR U6941 ( .A(n6538), .B(n6537), .Z(n6643) );
  NOR U6942 ( .A(n6644), .B(n6643), .Z(n6539) );
  NOR U6943 ( .A(n6540), .B(n6539), .Z(n6567) );
  IV U6944 ( .A(n6541), .Z(n6543) );
  XOR U6945 ( .A(n6543), .B(n6542), .Z(n6566) );
  NOR U6946 ( .A(n6567), .B(n6566), .Z(n6544) );
  NOR U6947 ( .A(n6545), .B(n6544), .Z(n6546) );
  IV U6948 ( .A(n6546), .Z(n6919) );
  NOR U6949 ( .A(n6920), .B(n6919), .Z(n6547) );
  NOR U6950 ( .A(n6548), .B(n6547), .Z(n6549) );
  IV U6951 ( .A(n6549), .Z(n6665) );
  XOR U6952 ( .A(n6551), .B(n6550), .Z(n6664) );
  IV U6953 ( .A(n6664), .Z(n6552) );
  NOR U6954 ( .A(n6665), .B(n6552), .Z(n6553) );
  NOR U6955 ( .A(n6554), .B(n6553), .Z(n6563) );
  IV U6956 ( .A(n6555), .Z(n6556) );
  NOR U6957 ( .A(n6557), .B(n6556), .Z(n6561) );
  NOR U6958 ( .A(n6559), .B(n6558), .Z(n6560) );
  NOR U6959 ( .A(n6561), .B(n6560), .Z(n6562) );
  XOR U6960 ( .A(n6563), .B(n6562), .Z(n6669) );
  XOR U6961 ( .A(n6565), .B(n6564), .Z(n6654) );
  XOR U6962 ( .A(n6567), .B(n6566), .Z(n6601) );
  NOR U6963 ( .A(n9237), .B(n8235), .Z(n6570) );
  NOR U6964 ( .A(n6784), .B(n9584), .Z(n6571) );
  NOR U6965 ( .A(n6570), .B(n6571), .Z(n6574) );
  XOR U6966 ( .A(n6569), .B(n6568), .Z(n6737) );
  IV U6967 ( .A(n6570), .Z(n6572) );
  XOR U6968 ( .A(n6572), .B(n6571), .Z(n6738) );
  NOR U6969 ( .A(n6737), .B(n6738), .Z(n6573) );
  NOR U6970 ( .A(n6574), .B(n6573), .Z(n6602) );
  NOR U6971 ( .A(n6601), .B(n6602), .Z(n6605) );
  NOR U6972 ( .A(n8311), .B(n9113), .Z(n6575) );
  IV U6973 ( .A(n6575), .Z(n6578) );
  NOR U6974 ( .A(n9571), .B(n6957), .Z(n6577) );
  IV U6975 ( .A(n6577), .Z(n6576) );
  NOR U6976 ( .A(n6578), .B(n6576), .Z(n6583) );
  XOR U6977 ( .A(n6578), .B(n6577), .Z(n6709) );
  NOR U6978 ( .A(n9592), .B(n6579), .Z(n6621) );
  NOR U6979 ( .A(n9080), .B(n8499), .Z(n6580) );
  IV U6980 ( .A(n6580), .Z(n6620) );
  NOR U6981 ( .A(n6581), .B(n9600), .Z(n6618) );
  XOR U6982 ( .A(n6620), .B(n6618), .Z(n6622) );
  XOR U6983 ( .A(n6621), .B(n6622), .Z(n6708) );
  NOR U6984 ( .A(n6709), .B(n6708), .Z(n6582) );
  NOR U6985 ( .A(n6583), .B(n6582), .Z(n6938) );
  NOR U6986 ( .A(n9301), .B(n7851), .Z(n6584) );
  IV U6987 ( .A(n6584), .Z(n6587) );
  NOR U6988 ( .A(n7529), .B(n9388), .Z(n6586) );
  IV U6989 ( .A(n6586), .Z(n6585) );
  NOR U6990 ( .A(n6587), .B(n6585), .Z(n6590) );
  XOR U6991 ( .A(n6587), .B(n6586), .Z(n6608) );
  NOR U6992 ( .A(n9336), .B(n7714), .Z(n6588) );
  IV U6993 ( .A(n6588), .Z(n6607) );
  NOR U6994 ( .A(n6608), .B(n6607), .Z(n6589) );
  NOR U6995 ( .A(n6590), .B(n6589), .Z(n6936) );
  IV U6996 ( .A(n6936), .Z(n6600) );
  NOR U6997 ( .A(n8582), .B(n8754), .Z(n6596) );
  IV U6998 ( .A(n6596), .Z(n6592) );
  XOR U6999 ( .A(n6591), .B(sum[27]), .Z(n6595) );
  NOR U7000 ( .A(n6592), .B(n6595), .Z(n6599) );
  IV U7001 ( .A(sum[26]), .Z(n6594) );
  NOR U7002 ( .A(n9593), .B(n6957), .Z(n6593) );
  IV U7003 ( .A(n6593), .Z(n6712) );
  NOR U7004 ( .A(n6594), .B(n6712), .Z(n6740) );
  IV U7005 ( .A(n6740), .Z(n6597) );
  XOR U7006 ( .A(n6596), .B(n6595), .Z(n6739) );
  NOR U7007 ( .A(n6597), .B(n6739), .Z(n6598) );
  NOR U7008 ( .A(n6599), .B(n6598), .Z(n6935) );
  XOR U7009 ( .A(n6600), .B(n6935), .Z(n6937) );
  XOR U7010 ( .A(n6938), .B(n6937), .Z(n6856) );
  XOR U7011 ( .A(n6602), .B(n6601), .Z(n6603) );
  IV U7012 ( .A(n6603), .Z(n6857) );
  NOR U7013 ( .A(n6856), .B(n6857), .Z(n6604) );
  NOR U7014 ( .A(n6605), .B(n6604), .Z(n6655) );
  IV U7015 ( .A(n6655), .Z(n6606) );
  NOR U7016 ( .A(n6654), .B(n6606), .Z(n6658) );
  NOR U7017 ( .A(n8862), .B(n8729), .Z(n6609) );
  NOR U7018 ( .A(n7531), .B(n9414), .Z(n6610) );
  NOR U7019 ( .A(n6609), .B(n6610), .Z(n6613) );
  XOR U7020 ( .A(n6608), .B(n6607), .Z(n6632) );
  IV U7021 ( .A(n6609), .Z(n6611) );
  XOR U7022 ( .A(n6611), .B(n6610), .Z(n6633) );
  NOR U7023 ( .A(n6632), .B(n6633), .Z(n6612) );
  NOR U7024 ( .A(n6613), .B(n6612), .Z(n6650) );
  XOR U7025 ( .A(n6615), .B(n6614), .Z(n6925) );
  XOR U7026 ( .A(n6617), .B(n6616), .Z(n6923) );
  IV U7027 ( .A(n6618), .Z(n6619) );
  NOR U7028 ( .A(n6620), .B(n6619), .Z(n6625) );
  IV U7029 ( .A(n6621), .Z(n6623) );
  NOR U7030 ( .A(n6623), .B(n6622), .Z(n6624) );
  NOR U7031 ( .A(n6625), .B(n6624), .Z(n6921) );
  XOR U7032 ( .A(n6923), .B(n6921), .Z(n6924) );
  XOR U7033 ( .A(n6925), .B(n6924), .Z(n6651) );
  IV U7034 ( .A(n6651), .Z(n6626) );
  NOR U7035 ( .A(n6650), .B(n6626), .Z(n6653) );
  NOR U7036 ( .A(n8290), .B(n9115), .Z(n6627) );
  IV U7037 ( .A(n6627), .Z(n8288) );
  NOR U7038 ( .A(n9316), .B(n8069), .Z(n6628) );
  XOR U7039 ( .A(n6629), .B(n6628), .Z(n6638) );
  XOR U7040 ( .A(n6631), .B(n6630), .Z(n6639) );
  XOR U7041 ( .A(n6638), .B(n6639), .Z(n6634) );
  NOR U7042 ( .A(n8288), .B(n6634), .Z(n6637) );
  XOR U7043 ( .A(n6633), .B(n6632), .Z(n6706) );
  XOR U7044 ( .A(n8288), .B(n6634), .Z(n6707) );
  IV U7045 ( .A(n6707), .Z(n6635) );
  NOR U7046 ( .A(n6706), .B(n6635), .Z(n6636) );
  NOR U7047 ( .A(n6637), .B(n6636), .Z(n6932) );
  NOR U7048 ( .A(n9316), .B(n8228), .Z(n6692) );
  IV U7049 ( .A(n6692), .Z(n8003) );
  NOR U7050 ( .A(n7123), .B(n8003), .Z(n6642) );
  IV U7051 ( .A(n6638), .Z(n6640) );
  NOR U7052 ( .A(n6640), .B(n6639), .Z(n6641) );
  NOR U7053 ( .A(n6642), .B(n6641), .Z(n6930) );
  NOR U7054 ( .A(n7314), .B(n9472), .Z(n6646) );
  NOR U7055 ( .A(n9429), .B(n7772), .Z(n6645) );
  NOR U7056 ( .A(n6646), .B(n6645), .Z(n6649) );
  XOR U7057 ( .A(n6644), .B(n6643), .Z(n6711) );
  XOR U7058 ( .A(n6646), .B(n6645), .Z(n6647) );
  IV U7059 ( .A(n6647), .Z(n6710) );
  NOR U7060 ( .A(n6711), .B(n6710), .Z(n6648) );
  NOR U7061 ( .A(n6649), .B(n6648), .Z(n6928) );
  XOR U7062 ( .A(n6930), .B(n6928), .Z(n6931) );
  XOR U7063 ( .A(n6932), .B(n6931), .Z(n6882) );
  XOR U7064 ( .A(n6651), .B(n6650), .Z(n6881) );
  NOR U7065 ( .A(n6882), .B(n6881), .Z(n6652) );
  NOR U7066 ( .A(n6653), .B(n6652), .Z(n6918) );
  IV U7067 ( .A(n6918), .Z(n6656) );
  XOR U7068 ( .A(n6655), .B(n6654), .Z(n6917) );
  NOR U7069 ( .A(n6656), .B(n6917), .Z(n6657) );
  NOR U7070 ( .A(n6658), .B(n6657), .Z(n6662) );
  XOR U7071 ( .A(n6660), .B(n6659), .Z(n6663) );
  IV U7072 ( .A(n6663), .Z(n6661) );
  NOR U7073 ( .A(n6662), .B(n6661), .Z(n6667) );
  XOR U7074 ( .A(n6663), .B(n6662), .Z(n7087) );
  XOR U7075 ( .A(n6665), .B(n6664), .Z(n7086) );
  NOR U7076 ( .A(n7087), .B(n7086), .Z(n6666) );
  NOR U7077 ( .A(n6667), .B(n6666), .Z(n6668) );
  XOR U7078 ( .A(n6669), .B(n6668), .Z(n6670) );
  XOR U7079 ( .A(n6671), .B(n6670), .Z(n6672) );
  XOR U7080 ( .A(n6673), .B(n6672), .Z(n9749) );
  NOR U7081 ( .A(n8656), .B(n8862), .Z(n6778) );
  NOR U7082 ( .A(n9260), .B(n8069), .Z(n6779) );
  IV U7083 ( .A(n6779), .Z(n7971) );
  XOR U7084 ( .A(n6778), .B(n7971), .Z(n6780) );
  NOR U7085 ( .A(n7531), .B(n9472), .Z(n6674) );
  IV U7086 ( .A(n6674), .Z(n6725) );
  NOR U7087 ( .A(n9237), .B(n8311), .Z(n6721) );
  NOR U7088 ( .A(n9490), .B(n7314), .Z(n6675) );
  IV U7089 ( .A(n6675), .Z(n6722) );
  XOR U7090 ( .A(n6721), .B(n6722), .Z(n6724) );
  XOR U7091 ( .A(n6725), .B(n6724), .Z(n6781) );
  XOR U7092 ( .A(n6780), .B(n6781), .Z(n6687) );
  NOR U7093 ( .A(n8068), .B(n9301), .Z(n6803) );
  IV U7094 ( .A(n6803), .Z(n6676) );
  NOR U7095 ( .A(n7529), .B(n9526), .Z(n6802) );
  XOR U7096 ( .A(n6676), .B(n6802), .Z(n6804) );
  NOR U7097 ( .A(n9493), .B(n7321), .Z(n6677) );
  IV U7098 ( .A(n6677), .Z(n6703) );
  NOR U7099 ( .A(n8948), .B(n8729), .Z(n6699) );
  NOR U7100 ( .A(n7167), .B(n9584), .Z(n6678) );
  IV U7101 ( .A(n6678), .Z(n6700) );
  XOR U7102 ( .A(n6699), .B(n6700), .Z(n6702) );
  XOR U7103 ( .A(n6703), .B(n6702), .Z(n6805) );
  XOR U7104 ( .A(n6804), .B(n6805), .Z(n6686) );
  NOR U7105 ( .A(n6687), .B(n6686), .Z(n6690) );
  NOR U7106 ( .A(n9592), .B(n6784), .Z(n6683) );
  IV U7107 ( .A(n6683), .Z(n6680) );
  NOR U7108 ( .A(n8422), .B(n9113), .Z(n6679) );
  IV U7109 ( .A(n6679), .Z(n6682) );
  NOR U7110 ( .A(n6680), .B(n6682), .Z(n6685) );
  NOR U7111 ( .A(n9599), .B(n7167), .Z(n6681) );
  IV U7112 ( .A(n6681), .Z(n6959) );
  XOR U7113 ( .A(n6683), .B(n6682), .Z(n6958) );
  NOR U7114 ( .A(n6959), .B(n6958), .Z(n6684) );
  NOR U7115 ( .A(n6685), .B(n6684), .Z(n6974) );
  XOR U7116 ( .A(n6687), .B(n6686), .Z(n6688) );
  IV U7117 ( .A(n6688), .Z(n6973) );
  NOR U7118 ( .A(n6974), .B(n6973), .Z(n6689) );
  NOR U7119 ( .A(n6690), .B(n6689), .Z(n6742) );
  NOR U7120 ( .A(n8501), .B(n9115), .Z(n6694) );
  NOR U7121 ( .A(n8290), .B(n9241), .Z(n6695) );
  NOR U7122 ( .A(n6694), .B(n6695), .Z(n6698) );
  NOR U7123 ( .A(n9202), .B(n8235), .Z(n6691) );
  IV U7124 ( .A(n6691), .Z(n6808) );
  XOR U7125 ( .A(n6692), .B(n6808), .Z(n6810) );
  NOR U7126 ( .A(n9034), .B(n8582), .Z(n6693) );
  IV U7127 ( .A(n6693), .Z(n6809) );
  XOR U7128 ( .A(n6810), .B(n6809), .Z(n6746) );
  IV U7129 ( .A(n6694), .Z(n6696) );
  XOR U7130 ( .A(n6696), .B(n6695), .Z(n6747) );
  NOR U7131 ( .A(n6746), .B(n6747), .Z(n6697) );
  NOR U7132 ( .A(n6698), .B(n6697), .Z(n6845) );
  IV U7133 ( .A(n6699), .Z(n6701) );
  NOR U7134 ( .A(n6701), .B(n6700), .Z(n6705) );
  NOR U7135 ( .A(n6703), .B(n6702), .Z(n6704) );
  NOR U7136 ( .A(n6705), .B(n6704), .Z(n6841) );
  XOR U7137 ( .A(n6707), .B(n6706), .Z(n6853) );
  XOR U7138 ( .A(n6709), .B(n6708), .Z(n6849) );
  XOR U7139 ( .A(n6711), .B(n6710), .Z(n6851) );
  XOR U7140 ( .A(n6849), .B(n6851), .Z(n6852) );
  XOR U7141 ( .A(n6853), .B(n6852), .Z(n6843) );
  XOR U7142 ( .A(n6841), .B(n6843), .Z(n6844) );
  XOR U7143 ( .A(n6845), .B(n6844), .Z(n6741) );
  NOR U7144 ( .A(n6742), .B(n6741), .Z(n6745) );
  XOR U7145 ( .A(n6712), .B(sum[26]), .Z(n6716) );
  NOR U7146 ( .A(n8727), .B(n8754), .Z(n6717) );
  IV U7147 ( .A(n6717), .Z(n6713) );
  NOR U7148 ( .A(n6716), .B(n6713), .Z(n6720) );
  IV U7149 ( .A(sum[25]), .Z(n6715) );
  NOR U7150 ( .A(n9593), .B(n7225), .Z(n6714) );
  IV U7151 ( .A(n6714), .Z(n6948) );
  NOR U7152 ( .A(n6715), .B(n6948), .Z(n6749) );
  IV U7153 ( .A(n6749), .Z(n6718) );
  XOR U7154 ( .A(n6717), .B(n6716), .Z(n6748) );
  NOR U7155 ( .A(n6718), .B(n6748), .Z(n6719) );
  NOR U7156 ( .A(n6720), .B(n6719), .Z(n6860) );
  IV U7157 ( .A(n6721), .Z(n6723) );
  NOR U7158 ( .A(n6723), .B(n6722), .Z(n6727) );
  NOR U7159 ( .A(n6725), .B(n6724), .Z(n6726) );
  NOR U7160 ( .A(n6727), .B(n6726), .Z(n6859) );
  XOR U7161 ( .A(n6860), .B(n6859), .Z(n6861) );
  NOR U7162 ( .A(n6728), .B(n9600), .Z(n6734) );
  IV U7163 ( .A(n6734), .Z(n6730) );
  NOR U7164 ( .A(n8422), .B(n9080), .Z(n6729) );
  IV U7165 ( .A(n6729), .Z(n6733) );
  NOR U7166 ( .A(n6730), .B(n6733), .Z(n6736) );
  NOR U7167 ( .A(n9592), .B(n6731), .Z(n6732) );
  IV U7168 ( .A(n6732), .Z(n6787) );
  XOR U7169 ( .A(n6734), .B(n6733), .Z(n6786) );
  NOR U7170 ( .A(n6787), .B(n6786), .Z(n6735) );
  NOR U7171 ( .A(n6736), .B(n6735), .Z(n6877) );
  XOR U7172 ( .A(n6738), .B(n6737), .Z(n6874) );
  XOR U7173 ( .A(n6740), .B(n6739), .Z(n6873) );
  XOR U7174 ( .A(n6874), .B(n6873), .Z(n6875) );
  XOR U7175 ( .A(n6877), .B(n6875), .Z(n6863) );
  XOR U7176 ( .A(n6861), .B(n6863), .Z(n6822) );
  XOR U7177 ( .A(n6742), .B(n6741), .Z(n6821) );
  IV U7178 ( .A(n6821), .Z(n6743) );
  NOR U7179 ( .A(n6822), .B(n6743), .Z(n6744) );
  NOR U7180 ( .A(n6745), .B(n6744), .Z(n6885) );
  XOR U7181 ( .A(n6747), .B(n6746), .Z(n6757) );
  XOR U7182 ( .A(n6749), .B(n6748), .Z(n6756) );
  NOR U7183 ( .A(n6757), .B(n6756), .Z(n6760) );
  NOR U7184 ( .A(n9241), .B(n8862), .Z(n7618) );
  IV U7185 ( .A(n7618), .Z(n7621) );
  NOR U7186 ( .A(n6750), .B(n7621), .Z(n6755) );
  NOR U7187 ( .A(n9115), .B(n8582), .Z(n6992) );
  IV U7188 ( .A(n6992), .Z(n8445) );
  NOR U7189 ( .A(n8754), .B(n8862), .Z(n6752) );
  NOR U7190 ( .A(n8501), .B(n9241), .Z(n6751) );
  XOR U7191 ( .A(n6752), .B(n6751), .Z(n6753) );
  IV U7192 ( .A(n6753), .Z(n6993) );
  NOR U7193 ( .A(n8445), .B(n6993), .Z(n6754) );
  NOR U7194 ( .A(n6755), .B(n6754), .Z(n6976) );
  XOR U7195 ( .A(n6757), .B(n6756), .Z(n6758) );
  IV U7196 ( .A(n6758), .Z(n6975) );
  NOR U7197 ( .A(n6976), .B(n6975), .Z(n6759) );
  NOR U7198 ( .A(n6760), .B(n6759), .Z(n6761) );
  IV U7199 ( .A(n6761), .Z(n6830) );
  NOR U7200 ( .A(n9414), .B(n7772), .Z(n6766) );
  NOR U7201 ( .A(n7891), .B(n9336), .Z(n6767) );
  NOR U7202 ( .A(n6766), .B(n6767), .Z(n6770) );
  NOR U7203 ( .A(n7714), .B(n9388), .Z(n6762) );
  IV U7204 ( .A(n6762), .Z(n6775) );
  NOR U7205 ( .A(n7225), .B(n9571), .Z(n6764) );
  NOR U7206 ( .A(n9429), .B(n7851), .Z(n6763) );
  XOR U7207 ( .A(n6764), .B(n6763), .Z(n6765) );
  IV U7208 ( .A(n6765), .Z(n6774) );
  XOR U7209 ( .A(n6775), .B(n6774), .Z(n6789) );
  IV U7210 ( .A(n6766), .Z(n6768) );
  XOR U7211 ( .A(n6768), .B(n6767), .Z(n6788) );
  NOR U7212 ( .A(n6789), .B(n6788), .Z(n6769) );
  NOR U7213 ( .A(n6770), .B(n6769), .Z(n6771) );
  IV U7214 ( .A(n6771), .Z(n6870) );
  NOR U7215 ( .A(n9571), .B(n7851), .Z(n7459) );
  IV U7216 ( .A(n7459), .Z(n6772) );
  NOR U7217 ( .A(n6773), .B(n6772), .Z(n6777) );
  NOR U7218 ( .A(n6775), .B(n6774), .Z(n6776) );
  NOR U7219 ( .A(n6777), .B(n6776), .Z(n6868) );
  NOR U7220 ( .A(n6779), .B(n6778), .Z(n6783) );
  NOR U7221 ( .A(n6781), .B(n6780), .Z(n6782) );
  NOR U7222 ( .A(n6783), .B(n6782), .Z(n6866) );
  XOR U7223 ( .A(n6868), .B(n6866), .Z(n6869) );
  XOR U7224 ( .A(n6870), .B(n6869), .Z(n6828) );
  NOR U7225 ( .A(n9599), .B(n6784), .Z(n6814) );
  NOR U7226 ( .A(n8499), .B(n9113), .Z(n6813) );
  XOR U7227 ( .A(n6814), .B(n6813), .Z(n6785) );
  IV U7228 ( .A(n6785), .Z(n6815) );
  XOR U7229 ( .A(n6787), .B(n6786), .Z(n6816) );
  XOR U7230 ( .A(n6815), .B(n6816), .Z(n6797) );
  XOR U7231 ( .A(n6789), .B(n6788), .Z(n6798) );
  NOR U7232 ( .A(n6797), .B(n6798), .Z(n6801) );
  NOR U7233 ( .A(n7714), .B(n9526), .Z(n6790) );
  IV U7234 ( .A(n6790), .Z(n6793) );
  NOR U7235 ( .A(n9429), .B(n8068), .Z(n6792) );
  IV U7236 ( .A(n6792), .Z(n6791) );
  NOR U7237 ( .A(n6793), .B(n6791), .Z(n6796) );
  NOR U7238 ( .A(n7891), .B(n9388), .Z(n7017) );
  IV U7239 ( .A(n7017), .Z(n6794) );
  XOR U7240 ( .A(n6793), .B(n6792), .Z(n7016) );
  NOR U7241 ( .A(n6794), .B(n7016), .Z(n6795) );
  NOR U7242 ( .A(n6796), .B(n6795), .Z(n6982) );
  IV U7243 ( .A(n6797), .Z(n6799) );
  XOR U7244 ( .A(n6799), .B(n6798), .Z(n6981) );
  NOR U7245 ( .A(n6982), .B(n6981), .Z(n6800) );
  NOR U7246 ( .A(n6801), .B(n6800), .Z(n6826) );
  XOR U7247 ( .A(n6828), .B(n6826), .Z(n6829) );
  XOR U7248 ( .A(n6830), .B(n6829), .Z(n6820) );
  NOR U7249 ( .A(n6803), .B(n6802), .Z(n6807) );
  NOR U7250 ( .A(n6805), .B(n6804), .Z(n6806) );
  NOR U7251 ( .A(n6807), .B(n6806), .Z(n6836) );
  NOR U7252 ( .A(n8003), .B(n6808), .Z(n6812) );
  NOR U7253 ( .A(n6810), .B(n6809), .Z(n6811) );
  NOR U7254 ( .A(n6812), .B(n6811), .Z(n6835) );
  NOR U7255 ( .A(n6814), .B(n6813), .Z(n6818) );
  NOR U7256 ( .A(n6816), .B(n6815), .Z(n6817) );
  NOR U7257 ( .A(n6818), .B(n6817), .Z(n6833) );
  XOR U7258 ( .A(n6835), .B(n6833), .Z(n6837) );
  XOR U7259 ( .A(n6836), .B(n6837), .Z(n6819) );
  NOR U7260 ( .A(n6820), .B(n6819), .Z(n6825) );
  XOR U7261 ( .A(n6820), .B(n6819), .Z(n7006) );
  IV U7262 ( .A(n7006), .Z(n6823) );
  XOR U7263 ( .A(n6822), .B(n6821), .Z(n7005) );
  NOR U7264 ( .A(n6823), .B(n7005), .Z(n6824) );
  NOR U7265 ( .A(n6825), .B(n6824), .Z(n6884) );
  NOR U7266 ( .A(n6885), .B(n6884), .Z(n6888) );
  IV U7267 ( .A(n6826), .Z(n6827) );
  NOR U7268 ( .A(n6828), .B(n6827), .Z(n6832) );
  NOR U7269 ( .A(n6830), .B(n6829), .Z(n6831) );
  NOR U7270 ( .A(n6832), .B(n6831), .Z(n6893) );
  IV U7271 ( .A(n6833), .Z(n6834) );
  NOR U7272 ( .A(n6835), .B(n6834), .Z(n6840) );
  IV U7273 ( .A(n6836), .Z(n6838) );
  NOR U7274 ( .A(n6838), .B(n6837), .Z(n6839) );
  NOR U7275 ( .A(n6840), .B(n6839), .Z(n6889) );
  IV U7276 ( .A(n6841), .Z(n6842) );
  NOR U7277 ( .A(n6843), .B(n6842), .Z(n6847) );
  NOR U7278 ( .A(n6845), .B(n6844), .Z(n6846) );
  NOR U7279 ( .A(n6847), .B(n6846), .Z(n6848) );
  IV U7280 ( .A(n6848), .Z(n6899) );
  IV U7281 ( .A(n6849), .Z(n6850) );
  NOR U7282 ( .A(n6851), .B(n6850), .Z(n6855) );
  NOR U7283 ( .A(n6853), .B(n6852), .Z(n6854) );
  NOR U7284 ( .A(n6855), .B(n6854), .Z(n6897) );
  XOR U7285 ( .A(n6857), .B(n6856), .Z(n6896) );
  XOR U7286 ( .A(n6897), .B(n6896), .Z(n6858) );
  IV U7287 ( .A(n6858), .Z(n6898) );
  XOR U7288 ( .A(n6899), .B(n6898), .Z(n6906) );
  NOR U7289 ( .A(n6860), .B(n6859), .Z(n6865) );
  IV U7290 ( .A(n6861), .Z(n6862) );
  NOR U7291 ( .A(n6863), .B(n6862), .Z(n6864) );
  NOR U7292 ( .A(n6865), .B(n6864), .Z(n6902) );
  IV U7293 ( .A(n6866), .Z(n6867) );
  NOR U7294 ( .A(n6868), .B(n6867), .Z(n6872) );
  NOR U7295 ( .A(n6870), .B(n6869), .Z(n6871) );
  NOR U7296 ( .A(n6872), .B(n6871), .Z(n6912) );
  NOR U7297 ( .A(n6874), .B(n6873), .Z(n6879) );
  IV U7298 ( .A(n6875), .Z(n6876) );
  NOR U7299 ( .A(n6877), .B(n6876), .Z(n6878) );
  NOR U7300 ( .A(n6879), .B(n6878), .Z(n6880) );
  IV U7301 ( .A(n6880), .Z(n6910) );
  XOR U7302 ( .A(n6882), .B(n6881), .Z(n6909) );
  XOR U7303 ( .A(n6910), .B(n6909), .Z(n6914) );
  XOR U7304 ( .A(n6912), .B(n6914), .Z(n6904) );
  XOR U7305 ( .A(n6902), .B(n6904), .Z(n6905) );
  XOR U7306 ( .A(n6906), .B(n6905), .Z(n6883) );
  IV U7307 ( .A(n6883), .Z(n6890) );
  XOR U7308 ( .A(n6889), .B(n6890), .Z(n6892) );
  XOR U7309 ( .A(n6893), .B(n6892), .Z(n6946) );
  XOR U7310 ( .A(n6885), .B(n6884), .Z(n6886) );
  IV U7311 ( .A(n6886), .Z(n6947) );
  NOR U7312 ( .A(n6946), .B(n6947), .Z(n6887) );
  NOR U7313 ( .A(n6888), .B(n6887), .Z(n6943) );
  IV U7314 ( .A(n6889), .Z(n6891) );
  NOR U7315 ( .A(n6891), .B(n6890), .Z(n6895) );
  NOR U7316 ( .A(n6893), .B(n6892), .Z(n6894) );
  NOR U7317 ( .A(n6895), .B(n6894), .Z(n7058) );
  NOR U7318 ( .A(n6897), .B(n6896), .Z(n6901) );
  NOR U7319 ( .A(n6899), .B(n6898), .Z(n6900) );
  NOR U7320 ( .A(n6901), .B(n6900), .Z(n7057) );
  IV U7321 ( .A(n7057), .Z(n6942) );
  IV U7322 ( .A(n6902), .Z(n6903) );
  NOR U7323 ( .A(n6904), .B(n6903), .Z(n6908) );
  NOR U7324 ( .A(n6906), .B(n6905), .Z(n6907) );
  NOR U7325 ( .A(n6908), .B(n6907), .Z(n7066) );
  IV U7326 ( .A(n6909), .Z(n6911) );
  NOR U7327 ( .A(n6911), .B(n6910), .Z(n6916) );
  IV U7328 ( .A(n6912), .Z(n6913) );
  NOR U7329 ( .A(n6914), .B(n6913), .Z(n6915) );
  NOR U7330 ( .A(n6916), .B(n6915), .Z(n7063) );
  XOR U7331 ( .A(n6918), .B(n6917), .Z(n7074) );
  XOR U7332 ( .A(n6920), .B(n6919), .Z(n7072) );
  IV U7333 ( .A(n6921), .Z(n6922) );
  NOR U7334 ( .A(n6923), .B(n6922), .Z(n6927) );
  NOR U7335 ( .A(n6925), .B(n6924), .Z(n6926) );
  NOR U7336 ( .A(n6927), .B(n6926), .Z(n7081) );
  IV U7337 ( .A(n6928), .Z(n6929) );
  NOR U7338 ( .A(n6930), .B(n6929), .Z(n6934) );
  NOR U7339 ( .A(n6932), .B(n6931), .Z(n6933) );
  NOR U7340 ( .A(n6934), .B(n6933), .Z(n7079) );
  XOR U7341 ( .A(n7081), .B(n7079), .Z(n7083) );
  NOR U7342 ( .A(n6936), .B(n6935), .Z(n6940) );
  NOR U7343 ( .A(n6938), .B(n6937), .Z(n6939) );
  NOR U7344 ( .A(n6940), .B(n6939), .Z(n6941) );
  IV U7345 ( .A(n6941), .Z(n7082) );
  XOR U7346 ( .A(n7083), .B(n7082), .Z(n7071) );
  XOR U7347 ( .A(n7072), .B(n7071), .Z(n7073) );
  XOR U7348 ( .A(n7074), .B(n7073), .Z(n7064) );
  XOR U7349 ( .A(n7063), .B(n7064), .Z(n7067) );
  XOR U7350 ( .A(n7066), .B(n7067), .Z(n7056) );
  XOR U7351 ( .A(n6942), .B(n7056), .Z(n7060) );
  XOR U7352 ( .A(n7058), .B(n7060), .Z(n6944) );
  NOR U7353 ( .A(n6943), .B(n6944), .Z(n7055) );
  IV U7354 ( .A(n6943), .Z(n6945) );
  XOR U7355 ( .A(n6945), .B(n6944), .Z(n7091) );
  XOR U7356 ( .A(n6947), .B(n6946), .Z(n7013) );
  NOR U7357 ( .A(n9034), .B(n8727), .Z(n6953) );
  IV U7358 ( .A(n6953), .Z(n6949) );
  XOR U7359 ( .A(n6948), .B(sum[25]), .Z(n6952) );
  NOR U7360 ( .A(n6949), .B(n6952), .Z(n6956) );
  IV U7361 ( .A(sum[24]), .Z(n6951) );
  NOR U7362 ( .A(n9593), .B(n7314), .Z(n6950) );
  IV U7363 ( .A(n6950), .Z(n7222) );
  NOR U7364 ( .A(n6951), .B(n7222), .Z(n7148) );
  IV U7365 ( .A(n7148), .Z(n6954) );
  XOR U7366 ( .A(n6953), .B(n6952), .Z(n7147) );
  NOR U7367 ( .A(n6954), .B(n7147), .Z(n6955) );
  NOR U7368 ( .A(n6956), .B(n6955), .Z(n6978) );
  NOR U7369 ( .A(n9600), .B(n6957), .Z(n6961) );
  NOR U7370 ( .A(n9080), .B(n8729), .Z(n6960) );
  NOR U7371 ( .A(n6961), .B(n6960), .Z(n6964) );
  XOR U7372 ( .A(n6959), .B(n6958), .Z(n7162) );
  XOR U7373 ( .A(n6961), .B(n6960), .Z(n6962) );
  IV U7374 ( .A(n6962), .Z(n7163) );
  NOR U7375 ( .A(n7162), .B(n7163), .Z(n6963) );
  NOR U7376 ( .A(n6964), .B(n6963), .Z(n6977) );
  IV U7377 ( .A(n6977), .Z(n6965) );
  NOR U7378 ( .A(n6978), .B(n6965), .Z(n6980) );
  NOR U7379 ( .A(n9301), .B(n8235), .Z(n6966) );
  IV U7380 ( .A(n6966), .Z(n6969) );
  NOR U7381 ( .A(n9260), .B(n8228), .Z(n6968) );
  IV U7382 ( .A(n6968), .Z(n6967) );
  NOR U7383 ( .A(n6969), .B(n6967), .Z(n6972) );
  XOR U7384 ( .A(n6969), .B(n6968), .Z(n6995) );
  NOR U7385 ( .A(n7531), .B(n9490), .Z(n6970) );
  IV U7386 ( .A(n6970), .Z(n6996) );
  NOR U7387 ( .A(n6995), .B(n6996), .Z(n6971) );
  NOR U7388 ( .A(n6972), .B(n6971), .Z(n7035) );
  XOR U7389 ( .A(n6974), .B(n6973), .Z(n7037) );
  XOR U7390 ( .A(n7035), .B(n7037), .Z(n7038) );
  XOR U7391 ( .A(n6976), .B(n6975), .Z(n7039) );
  XOR U7392 ( .A(n7038), .B(n7039), .Z(n7102) );
  XOR U7393 ( .A(n6978), .B(n6977), .Z(n7103) );
  NOR U7394 ( .A(n7102), .B(n7103), .Z(n6979) );
  NOR U7395 ( .A(n6980), .B(n6979), .Z(n7007) );
  XOR U7396 ( .A(n6982), .B(n6981), .Z(n6991) );
  NOR U7397 ( .A(n8948), .B(n8656), .Z(n6983) );
  IV U7398 ( .A(n6983), .Z(n8459) );
  NOR U7399 ( .A(n7321), .B(n9584), .Z(n6986) );
  IV U7400 ( .A(n6986), .Z(n6984) );
  NOR U7401 ( .A(n8459), .B(n6984), .Z(n6988) );
  NOR U7402 ( .A(n7314), .B(n9571), .Z(n6985) );
  IV U7403 ( .A(n6985), .Z(n7096) );
  XOR U7404 ( .A(n6986), .B(n8459), .Z(n7095) );
  NOR U7405 ( .A(n7096), .B(n7095), .Z(n6987) );
  NOR U7406 ( .A(n6988), .B(n6987), .Z(n6990) );
  IV U7407 ( .A(n6990), .Z(n6989) );
  NOR U7408 ( .A(n6991), .B(n6989), .Z(n7003) );
  XOR U7409 ( .A(n6991), .B(n6990), .Z(n7030) );
  NOR U7410 ( .A(n9414), .B(n7851), .Z(n6998) );
  IV U7411 ( .A(n6998), .Z(n7279) );
  XOR U7412 ( .A(n6993), .B(n6992), .Z(n6997) );
  NOR U7413 ( .A(n7279), .B(n6997), .Z(n7000) );
  NOR U7414 ( .A(n9237), .B(n8499), .Z(n7023) );
  IV U7415 ( .A(n7023), .Z(n6994) );
  NOR U7416 ( .A(n9316), .B(n8290), .Z(n7022) );
  XOR U7417 ( .A(n6994), .B(n7022), .Z(n7024) );
  XOR U7418 ( .A(n6996), .B(n6995), .Z(n7025) );
  XOR U7419 ( .A(n7024), .B(n7025), .Z(n7129) );
  XOR U7420 ( .A(n6998), .B(n6997), .Z(n7130) );
  NOR U7421 ( .A(n7129), .B(n7130), .Z(n6999) );
  NOR U7422 ( .A(n7000), .B(n6999), .Z(n7001) );
  IV U7423 ( .A(n7001), .Z(n7029) );
  NOR U7424 ( .A(n7030), .B(n7029), .Z(n7002) );
  NOR U7425 ( .A(n7003), .B(n7002), .Z(n7008) );
  IV U7426 ( .A(n7008), .Z(n7004) );
  NOR U7427 ( .A(n7007), .B(n7004), .Z(n7010) );
  XOR U7428 ( .A(n7006), .B(n7005), .Z(n7044) );
  XOR U7429 ( .A(n7008), .B(n7007), .Z(n7043) );
  NOR U7430 ( .A(n7044), .B(n7043), .Z(n7009) );
  NOR U7431 ( .A(n7010), .B(n7009), .Z(n7012) );
  IV U7432 ( .A(n7012), .Z(n7011) );
  NOR U7433 ( .A(n7013), .B(n7011), .Z(n7052) );
  XOR U7434 ( .A(n7013), .B(n7012), .Z(n7093) );
  NOR U7435 ( .A(n8069), .B(n9336), .Z(n7019) );
  IV U7436 ( .A(n7019), .Z(n7015) );
  NOR U7437 ( .A(n9472), .B(n7772), .Z(n7014) );
  IV U7438 ( .A(n7014), .Z(n7018) );
  NOR U7439 ( .A(n7015), .B(n7018), .Z(n7021) );
  XOR U7440 ( .A(n7017), .B(n7016), .Z(n7164) );
  XOR U7441 ( .A(n7019), .B(n7018), .Z(n7165) );
  NOR U7442 ( .A(n7164), .B(n7165), .Z(n7020) );
  NOR U7443 ( .A(n7021), .B(n7020), .Z(n7032) );
  NOR U7444 ( .A(n7023), .B(n7022), .Z(n7027) );
  NOR U7445 ( .A(n7025), .B(n7024), .Z(n7026) );
  NOR U7446 ( .A(n7027), .B(n7026), .Z(n7031) );
  IV U7447 ( .A(n7031), .Z(n7028) );
  NOR U7448 ( .A(n7032), .B(n7028), .Z(n7034) );
  XOR U7449 ( .A(n7030), .B(n7029), .Z(n7109) );
  XOR U7450 ( .A(n7032), .B(n7031), .Z(n7108) );
  NOR U7451 ( .A(n7109), .B(n7108), .Z(n7033) );
  NOR U7452 ( .A(n7034), .B(n7033), .Z(n7045) );
  IV U7453 ( .A(n7035), .Z(n7036) );
  NOR U7454 ( .A(n7037), .B(n7036), .Z(n7041) );
  NOR U7455 ( .A(n7039), .B(n7038), .Z(n7040) );
  NOR U7456 ( .A(n7041), .B(n7040), .Z(n7046) );
  IV U7457 ( .A(n7046), .Z(n7042) );
  NOR U7458 ( .A(n7045), .B(n7042), .Z(n7049) );
  XOR U7459 ( .A(n7044), .B(n7043), .Z(n7114) );
  IV U7460 ( .A(n7114), .Z(n7047) );
  XOR U7461 ( .A(n7046), .B(n7045), .Z(n7113) );
  NOR U7462 ( .A(n7047), .B(n7113), .Z(n7048) );
  NOR U7463 ( .A(n7049), .B(n7048), .Z(n7094) );
  IV U7464 ( .A(n7094), .Z(n7050) );
  NOR U7465 ( .A(n7093), .B(n7050), .Z(n7051) );
  NOR U7466 ( .A(n7052), .B(n7051), .Z(n7092) );
  IV U7467 ( .A(n7092), .Z(n7053) );
  NOR U7468 ( .A(n7091), .B(n7053), .Z(n7054) );
  NOR U7469 ( .A(n7055), .B(n7054), .Z(n7090) );
  IV U7470 ( .A(n7090), .Z(n7088) );
  NOR U7471 ( .A(n7057), .B(n7056), .Z(n7062) );
  IV U7472 ( .A(n7058), .Z(n7059) );
  NOR U7473 ( .A(n7060), .B(n7059), .Z(n7061) );
  NOR U7474 ( .A(n7062), .B(n7061), .Z(n9741) );
  IV U7475 ( .A(n7063), .Z(n7065) );
  NOR U7476 ( .A(n7065), .B(n7064), .Z(n7070) );
  IV U7477 ( .A(n7066), .Z(n7068) );
  NOR U7478 ( .A(n7068), .B(n7067), .Z(n7069) );
  NOR U7479 ( .A(n7070), .B(n7069), .Z(n9738) );
  NOR U7480 ( .A(n7072), .B(n7071), .Z(n7077) );
  IV U7481 ( .A(n7073), .Z(n7075) );
  NOR U7482 ( .A(n7075), .B(n7074), .Z(n7076) );
  NOR U7483 ( .A(n7077), .B(n7076), .Z(n7078) );
  IV U7484 ( .A(n7078), .Z(n9732) );
  IV U7485 ( .A(n7079), .Z(n7080) );
  NOR U7486 ( .A(n7081), .B(n7080), .Z(n7085) );
  NOR U7487 ( .A(n7083), .B(n7082), .Z(n7084) );
  NOR U7488 ( .A(n7085), .B(n7084), .Z(n9730) );
  XOR U7489 ( .A(n7087), .B(n7086), .Z(n9729) );
  XOR U7490 ( .A(n9730), .B(n9729), .Z(n9731) );
  XOR U7491 ( .A(n9732), .B(n9731), .Z(n9740) );
  XOR U7492 ( .A(n9738), .B(n9740), .Z(n9743) );
  XOR U7493 ( .A(n9741), .B(n9743), .Z(n7089) );
  NOR U7494 ( .A(n7088), .B(n7089), .Z(n9728) );
  XOR U7495 ( .A(n7090), .B(n7089), .Z(n9754) );
  XOR U7496 ( .A(n7092), .B(n7091), .Z(n7274) );
  XOR U7497 ( .A(n7094), .B(n7093), .Z(n7195) );
  NOR U7498 ( .A(n7529), .B(n9493), .Z(n7098) );
  NOR U7499 ( .A(n8311), .B(n9202), .Z(n7097) );
  NOR U7500 ( .A(n7098), .B(n7097), .Z(n7101) );
  XOR U7501 ( .A(n7096), .B(n7095), .Z(n7132) );
  XOR U7502 ( .A(n7098), .B(n7097), .Z(n7099) );
  IV U7503 ( .A(n7099), .Z(n7131) );
  NOR U7504 ( .A(n7132), .B(n7131), .Z(n7100) );
  NOR U7505 ( .A(n7101), .B(n7100), .Z(n7107) );
  IV U7506 ( .A(n7107), .Z(n7105) );
  IV U7507 ( .A(n7102), .Z(n7104) );
  XOR U7508 ( .A(n7104), .B(n7103), .Z(n7106) );
  NOR U7509 ( .A(n7105), .B(n7106), .Z(n7112) );
  XOR U7510 ( .A(n7107), .B(n7106), .Z(n7179) );
  XOR U7511 ( .A(n7109), .B(n7108), .Z(n7110) );
  IV U7512 ( .A(n7110), .Z(n7178) );
  NOR U7513 ( .A(n7179), .B(n7178), .Z(n7111) );
  NOR U7514 ( .A(n7112), .B(n7111), .Z(n7116) );
  XOR U7515 ( .A(n7114), .B(n7113), .Z(n7115) );
  NOR U7516 ( .A(n7116), .B(n7115), .Z(n7193) );
  XOR U7517 ( .A(n7116), .B(n7115), .Z(n7117) );
  IV U7518 ( .A(n7117), .Z(n7205) );
  NOR U7519 ( .A(n9080), .B(n9115), .Z(n7753) );
  IV U7520 ( .A(n7753), .Z(n7749) );
  NOR U7521 ( .A(n7118), .B(n7749), .Z(n7122) );
  NOR U7522 ( .A(n8501), .B(n9316), .Z(n7223) );
  IV U7523 ( .A(n7223), .Z(n8498) );
  NOR U7524 ( .A(n9115), .B(n8727), .Z(n7119) );
  IV U7525 ( .A(n7119), .Z(n8054) );
  NOR U7526 ( .A(n9080), .B(n8656), .Z(n7120) );
  XOR U7527 ( .A(n8054), .B(n7120), .Z(n7224) );
  NOR U7528 ( .A(n8498), .B(n7224), .Z(n7121) );
  NOR U7529 ( .A(n7122), .B(n7121), .Z(n7150) );
  NOR U7530 ( .A(n8582), .B(n9388), .Z(n7958) );
  IV U7531 ( .A(n7958), .Z(n7953) );
  NOR U7532 ( .A(n7123), .B(n7953), .Z(n7128) );
  NOR U7533 ( .A(n8228), .B(n9336), .Z(n7124) );
  IV U7534 ( .A(n7124), .Z(n7212) );
  NOR U7535 ( .A(n8069), .B(n9388), .Z(n7125) );
  NOR U7536 ( .A(n9241), .B(n8582), .Z(n8120) );
  XOR U7537 ( .A(n7125), .B(n8120), .Z(n7211) );
  IV U7538 ( .A(n7211), .Z(n7126) );
  NOR U7539 ( .A(n7212), .B(n7126), .Z(n7127) );
  NOR U7540 ( .A(n7128), .B(n7127), .Z(n7157) );
  XOR U7541 ( .A(n7130), .B(n7129), .Z(n7153) );
  XOR U7542 ( .A(n7132), .B(n7131), .Z(n7155) );
  XOR U7543 ( .A(n7153), .B(n7155), .Z(n7156) );
  XOR U7544 ( .A(n7157), .B(n7156), .Z(n7149) );
  IV U7545 ( .A(n7149), .Z(n7133) );
  NOR U7546 ( .A(n7150), .B(n7133), .Z(n7152) );
  NOR U7547 ( .A(n8499), .B(n9472), .Z(n7972) );
  IV U7548 ( .A(n7972), .Z(n8016) );
  NOR U7549 ( .A(n7849), .B(n8016), .Z(n7139) );
  NOR U7550 ( .A(n7714), .B(n9493), .Z(n7134) );
  IV U7551 ( .A(n7134), .Z(n7249) );
  NOR U7552 ( .A(n9472), .B(n7851), .Z(n7136) );
  NOR U7553 ( .A(n8499), .B(n9202), .Z(n7135) );
  XOR U7554 ( .A(n7136), .B(n7135), .Z(n7137) );
  IV U7555 ( .A(n7137), .Z(n7248) );
  NOR U7556 ( .A(n7249), .B(n7248), .Z(n7138) );
  NOR U7557 ( .A(n7139), .B(n7138), .Z(n7184) );
  NOR U7558 ( .A(n7529), .B(n9584), .Z(n7144) );
  IV U7559 ( .A(n7144), .Z(n7141) );
  NOR U7560 ( .A(n8422), .B(n9237), .Z(n7140) );
  IV U7561 ( .A(n7140), .Z(n7143) );
  NOR U7562 ( .A(n7141), .B(n7143), .Z(n7146) );
  NOR U7563 ( .A(n7531), .B(n9571), .Z(n7142) );
  IV U7564 ( .A(n7142), .Z(n7243) );
  XOR U7565 ( .A(n7144), .B(n7143), .Z(n7242) );
  NOR U7566 ( .A(n7243), .B(n7242), .Z(n7145) );
  NOR U7567 ( .A(n7146), .B(n7145), .Z(n7181) );
  XOR U7568 ( .A(n7148), .B(n7147), .Z(n7180) );
  XOR U7569 ( .A(n7181), .B(n7180), .Z(n7182) );
  XOR U7570 ( .A(n7184), .B(n7182), .Z(n7296) );
  XOR U7571 ( .A(n7150), .B(n7149), .Z(n7295) );
  NOR U7572 ( .A(n7296), .B(n7295), .Z(n7151) );
  NOR U7573 ( .A(n7152), .B(n7151), .Z(n7188) );
  IV U7574 ( .A(n7188), .Z(n7161) );
  IV U7575 ( .A(n7153), .Z(n7154) );
  NOR U7576 ( .A(n7155), .B(n7154), .Z(n7159) );
  NOR U7577 ( .A(n7157), .B(n7156), .Z(n7158) );
  NOR U7578 ( .A(n7159), .B(n7158), .Z(n7160) );
  IV U7579 ( .A(n7160), .Z(n7187) );
  NOR U7580 ( .A(n7161), .B(n7187), .Z(n7190) );
  XOR U7581 ( .A(n7163), .B(n7162), .Z(n7175) );
  XOR U7582 ( .A(n7165), .B(n7164), .Z(n7174) );
  IV U7583 ( .A(n7174), .Z(n7166) );
  NOR U7584 ( .A(n7175), .B(n7166), .Z(n7177) );
  NOR U7585 ( .A(n8948), .B(n8754), .Z(n7170) );
  IV U7586 ( .A(n7170), .Z(n8615) );
  NOR U7587 ( .A(n9592), .B(n7167), .Z(n7168) );
  IV U7588 ( .A(n7168), .Z(n7171) );
  NOR U7589 ( .A(n8615), .B(n7171), .Z(n7173) );
  NOR U7590 ( .A(n9599), .B(n7321), .Z(n7169) );
  IV U7591 ( .A(n7169), .Z(n7228) );
  XOR U7592 ( .A(n7171), .B(n7170), .Z(n7227) );
  NOR U7593 ( .A(n7228), .B(n7227), .Z(n7172) );
  NOR U7594 ( .A(n7173), .B(n7172), .Z(n7209) );
  XOR U7595 ( .A(n7175), .B(n7174), .Z(n7208) );
  NOR U7596 ( .A(n7209), .B(n7208), .Z(n7176) );
  NOR U7597 ( .A(n7177), .B(n7176), .Z(n7200) );
  XOR U7598 ( .A(n7179), .B(n7178), .Z(n7199) );
  NOR U7599 ( .A(n7181), .B(n7180), .Z(n7186) );
  IV U7600 ( .A(n7182), .Z(n7183) );
  NOR U7601 ( .A(n7184), .B(n7183), .Z(n7185) );
  NOR U7602 ( .A(n7186), .B(n7185), .Z(n7197) );
  XOR U7603 ( .A(n7199), .B(n7197), .Z(n7202) );
  XOR U7604 ( .A(n7200), .B(n7202), .Z(n7237) );
  XOR U7605 ( .A(n7188), .B(n7187), .Z(n7238) );
  NOR U7606 ( .A(n7237), .B(n7238), .Z(n7189) );
  NOR U7607 ( .A(n7190), .B(n7189), .Z(n7206) );
  IV U7608 ( .A(n7206), .Z(n7191) );
  NOR U7609 ( .A(n7205), .B(n7191), .Z(n7192) );
  NOR U7610 ( .A(n7193), .B(n7192), .Z(n7196) );
  IV U7611 ( .A(n7196), .Z(n7194) );
  NOR U7612 ( .A(n7195), .B(n7194), .Z(n7272) );
  XOR U7613 ( .A(n7196), .B(n7195), .Z(n7503) );
  IV U7614 ( .A(n7197), .Z(n7198) );
  NOR U7615 ( .A(n7199), .B(n7198), .Z(n7204) );
  IV U7616 ( .A(n7200), .Z(n7201) );
  NOR U7617 ( .A(n7202), .B(n7201), .Z(n7203) );
  NOR U7618 ( .A(n7204), .B(n7203), .Z(n7266) );
  IV U7619 ( .A(n7266), .Z(n7207) );
  XOR U7620 ( .A(n7206), .B(n7205), .Z(n7265) );
  NOR U7621 ( .A(n7207), .B(n7265), .Z(n7269) );
  XOR U7622 ( .A(n7209), .B(n7208), .Z(n7219) );
  NOR U7623 ( .A(n9260), .B(n8290), .Z(n7213) );
  IV U7624 ( .A(n7213), .Z(n7329) );
  NOR U7625 ( .A(n8068), .B(n9414), .Z(n7210) );
  IV U7626 ( .A(n7210), .Z(n7214) );
  NOR U7627 ( .A(n7329), .B(n7214), .Z(n7216) );
  XOR U7628 ( .A(n7212), .B(n7211), .Z(n7363) );
  XOR U7629 ( .A(n7214), .B(n7213), .Z(n7362) );
  NOR U7630 ( .A(n7363), .B(n7362), .Z(n7215) );
  NOR U7631 ( .A(n7216), .B(n7215), .Z(n7218) );
  IV U7632 ( .A(n7218), .Z(n7217) );
  NOR U7633 ( .A(n7219), .B(n7217), .Z(n7236) );
  XOR U7634 ( .A(n7219), .B(n7218), .Z(n7257) );
  IV U7635 ( .A(sum[23]), .Z(n7221) );
  NOR U7636 ( .A(n7531), .B(n9593), .Z(n7220) );
  IV U7637 ( .A(n7220), .Z(n7383) );
  NOR U7638 ( .A(n7221), .B(n7383), .Z(n7300) );
  NOR U7639 ( .A(n9034), .B(n8862), .Z(n7297) );
  XOR U7640 ( .A(n7222), .B(sum[24]), .Z(n7298) );
  XOR U7641 ( .A(n7297), .B(n7298), .Z(n7301) );
  XOR U7642 ( .A(n7300), .B(n7301), .Z(n7229) );
  XOR U7643 ( .A(n7224), .B(n7223), .Z(n7230) );
  NOR U7644 ( .A(n7229), .B(n7230), .Z(n7233) );
  NOR U7645 ( .A(n8729), .B(n9113), .Z(n7306) );
  IV U7646 ( .A(n7306), .Z(n7226) );
  NOR U7647 ( .A(n9600), .B(n7225), .Z(n7305) );
  XOR U7648 ( .A(n7226), .B(n7305), .Z(n7307) );
  XOR U7649 ( .A(n7228), .B(n7227), .Z(n7308) );
  XOR U7650 ( .A(n7307), .B(n7308), .Z(n7289) );
  XOR U7651 ( .A(n7230), .B(n7229), .Z(n7288) );
  IV U7652 ( .A(n7288), .Z(n7231) );
  NOR U7653 ( .A(n7289), .B(n7231), .Z(n7232) );
  NOR U7654 ( .A(n7233), .B(n7232), .Z(n7234) );
  IV U7655 ( .A(n7234), .Z(n7256) );
  NOR U7656 ( .A(n7257), .B(n7256), .Z(n7235) );
  NOR U7657 ( .A(n7236), .B(n7235), .Z(n7241) );
  XOR U7658 ( .A(n7238), .B(n7237), .Z(n7240) );
  IV U7659 ( .A(n7240), .Z(n7239) );
  NOR U7660 ( .A(n7241), .B(n7239), .Z(n7264) );
  XOR U7661 ( .A(n7241), .B(n7240), .Z(n7409) );
  NOR U7662 ( .A(n8311), .B(n9301), .Z(n7244) );
  NOR U7663 ( .A(n9490), .B(n7772), .Z(n7245) );
  NOR U7664 ( .A(n7244), .B(n7245), .Z(n7247) );
  XOR U7665 ( .A(n7243), .B(n7242), .Z(n7360) );
  IV U7666 ( .A(n7244), .Z(n8079) );
  XOR U7667 ( .A(n7245), .B(n8079), .Z(n7361) );
  NOR U7668 ( .A(n7360), .B(n7361), .Z(n7246) );
  NOR U7669 ( .A(n7247), .B(n7246), .Z(n7259) );
  IV U7670 ( .A(n7259), .Z(n7255) );
  NOR U7671 ( .A(n9429), .B(n8235), .Z(n7250) );
  NOR U7672 ( .A(n7891), .B(n9526), .Z(n7251) );
  NOR U7673 ( .A(n7250), .B(n7251), .Z(n7253) );
  XOR U7674 ( .A(n7249), .B(n7248), .Z(n7287) );
  IV U7675 ( .A(n7250), .Z(n7519) );
  XOR U7676 ( .A(n7251), .B(n7519), .Z(n7286) );
  NOR U7677 ( .A(n7287), .B(n7286), .Z(n7252) );
  NOR U7678 ( .A(n7253), .B(n7252), .Z(n7254) );
  IV U7679 ( .A(n7254), .Z(n7258) );
  NOR U7680 ( .A(n7255), .B(n7258), .Z(n7261) );
  XOR U7681 ( .A(n7257), .B(n7256), .Z(n7358) );
  XOR U7682 ( .A(n7259), .B(n7258), .Z(n7359) );
  NOR U7683 ( .A(n7358), .B(n7359), .Z(n7260) );
  NOR U7684 ( .A(n7261), .B(n7260), .Z(n7410) );
  IV U7685 ( .A(n7410), .Z(n7262) );
  NOR U7686 ( .A(n7409), .B(n7262), .Z(n7263) );
  NOR U7687 ( .A(n7264), .B(n7263), .Z(n7277) );
  IV U7688 ( .A(n7277), .Z(n7267) );
  XOR U7689 ( .A(n7266), .B(n7265), .Z(n7276) );
  NOR U7690 ( .A(n7267), .B(n7276), .Z(n7268) );
  NOR U7691 ( .A(n7269), .B(n7268), .Z(n7504) );
  IV U7692 ( .A(n7504), .Z(n7270) );
  NOR U7693 ( .A(n7503), .B(n7270), .Z(n7271) );
  NOR U7694 ( .A(n7272), .B(n7271), .Z(n7275) );
  IV U7695 ( .A(n7275), .Z(n7273) );
  NOR U7696 ( .A(n7274), .B(n7273), .Z(n9725) );
  XOR U7697 ( .A(n7275), .B(n7274), .Z(n9759) );
  XOR U7698 ( .A(n7277), .B(n7276), .Z(n7498) );
  NOR U7699 ( .A(n9490), .B(n8235), .Z(n7278) );
  IV U7700 ( .A(n7278), .Z(n7723) );
  NOR U7701 ( .A(n7279), .B(n7723), .Z(n7285) );
  NOR U7702 ( .A(n8068), .B(n9472), .Z(n7280) );
  IV U7703 ( .A(n7280), .Z(n7451) );
  NOR U7704 ( .A(n9414), .B(n8235), .Z(n7282) );
  NOR U7705 ( .A(n9490), .B(n7851), .Z(n7281) );
  XOR U7706 ( .A(n7282), .B(n7281), .Z(n7283) );
  IV U7707 ( .A(n7283), .Z(n7450) );
  NOR U7708 ( .A(n7451), .B(n7450), .Z(n7284) );
  NOR U7709 ( .A(n7285), .B(n7284), .Z(n7290) );
  XOR U7710 ( .A(n7287), .B(n7286), .Z(n7291) );
  NOR U7711 ( .A(n7290), .B(n7291), .Z(n7294) );
  XOR U7712 ( .A(n7289), .B(n7288), .Z(n7395) );
  IV U7713 ( .A(n7290), .Z(n7292) );
  XOR U7714 ( .A(n7292), .B(n7291), .Z(n7394) );
  NOR U7715 ( .A(n7395), .B(n7394), .Z(n7293) );
  NOR U7716 ( .A(n7294), .B(n7293), .Z(n7344) );
  XOR U7717 ( .A(n7296), .B(n7295), .Z(n7352) );
  IV U7718 ( .A(n7297), .Z(n7299) );
  NOR U7719 ( .A(n7299), .B(n7298), .Z(n7304) );
  IV U7720 ( .A(n7300), .Z(n7302) );
  NOR U7721 ( .A(n7302), .B(n7301), .Z(n7303) );
  NOR U7722 ( .A(n7304), .B(n7303), .Z(n7351) );
  NOR U7723 ( .A(n7306), .B(n7305), .Z(n7310) );
  NOR U7724 ( .A(n7308), .B(n7307), .Z(n7309) );
  NOR U7725 ( .A(n7310), .B(n7309), .Z(n7349) );
  XOR U7726 ( .A(n7351), .B(n7349), .Z(n7354) );
  XOR U7727 ( .A(n7352), .B(n7354), .Z(n7343) );
  NOR U7728 ( .A(n7344), .B(n7343), .Z(n7347) );
  NOR U7729 ( .A(n8422), .B(n9600), .Z(n7311) );
  IV U7730 ( .A(n7311), .Z(n8626) );
  NOR U7731 ( .A(n8626), .B(n7312), .Z(n7319) );
  NOR U7732 ( .A(n7891), .B(n9493), .Z(n7313) );
  IV U7733 ( .A(n7313), .Z(n7419) );
  NOR U7734 ( .A(n9600), .B(n7314), .Z(n7316) );
  NOR U7735 ( .A(n8422), .B(n9202), .Z(n7315) );
  XOR U7736 ( .A(n7316), .B(n7315), .Z(n7317) );
  IV U7737 ( .A(n7317), .Z(n7418) );
  NOR U7738 ( .A(n7419), .B(n7418), .Z(n7318) );
  NOR U7739 ( .A(n7319), .B(n7318), .Z(n7340) );
  NOR U7740 ( .A(n7714), .B(n9584), .Z(n7323) );
  NOR U7741 ( .A(n9237), .B(n8729), .Z(n7324) );
  NOR U7742 ( .A(n7323), .B(n7324), .Z(n7327) );
  NOR U7743 ( .A(n9599), .B(n7529), .Z(n7320) );
  IV U7744 ( .A(n7320), .Z(n7380) );
  NOR U7745 ( .A(n9080), .B(n8754), .Z(n7376) );
  NOR U7746 ( .A(n9592), .B(n7321), .Z(n7322) );
  IV U7747 ( .A(n7322), .Z(n7377) );
  XOR U7748 ( .A(n7376), .B(n7377), .Z(n7379) );
  XOR U7749 ( .A(n7380), .B(n7379), .Z(n7526) );
  IV U7750 ( .A(n7323), .Z(n7325) );
  XOR U7751 ( .A(n7325), .B(n7324), .Z(n7527) );
  NOR U7752 ( .A(n7526), .B(n7527), .Z(n7326) );
  NOR U7753 ( .A(n7327), .B(n7326), .Z(n7339) );
  IV U7754 ( .A(n7339), .Z(n7328) );
  NOR U7755 ( .A(n7340), .B(n7328), .Z(n7342) );
  NOR U7756 ( .A(n8501), .B(n9336), .Z(n7649) );
  IV U7757 ( .A(n7649), .Z(n7589) );
  NOR U7758 ( .A(n7329), .B(n7589), .Z(n7338) );
  NOR U7759 ( .A(n9241), .B(n8727), .Z(n7331) );
  NOR U7760 ( .A(n9429), .B(n8311), .Z(n7330) );
  XOR U7761 ( .A(n7331), .B(n7330), .Z(n7332) );
  IV U7762 ( .A(n7332), .Z(n7368) );
  NOR U7763 ( .A(n8948), .B(n9034), .Z(n7333) );
  IV U7764 ( .A(n7333), .Z(n7367) );
  XOR U7765 ( .A(n7368), .B(n7367), .Z(n7478) );
  NOR U7766 ( .A(n8228), .B(n9388), .Z(n7475) );
  NOR U7767 ( .A(n9316), .B(n8582), .Z(n7476) );
  IV U7768 ( .A(n7476), .Z(n8580) );
  XOR U7769 ( .A(n7475), .B(n8580), .Z(n7477) );
  XOR U7770 ( .A(n7478), .B(n7477), .Z(n7436) );
  NOR U7771 ( .A(n8290), .B(n9336), .Z(n7335) );
  NOR U7772 ( .A(n9260), .B(n8501), .Z(n7334) );
  XOR U7773 ( .A(n7335), .B(n7334), .Z(n7435) );
  IV U7774 ( .A(n7435), .Z(n7336) );
  NOR U7775 ( .A(n7436), .B(n7336), .Z(n7337) );
  NOR U7776 ( .A(n7338), .B(n7337), .Z(n7482) );
  XOR U7777 ( .A(n7340), .B(n7339), .Z(n7483) );
  NOR U7778 ( .A(n7482), .B(n7483), .Z(n7341) );
  NOR U7779 ( .A(n7342), .B(n7341), .Z(n7415) );
  XOR U7780 ( .A(n7344), .B(n7343), .Z(n7345) );
  IV U7781 ( .A(n7345), .Z(n7414) );
  NOR U7782 ( .A(n7415), .B(n7414), .Z(n7346) );
  NOR U7783 ( .A(n7347), .B(n7346), .Z(n7348) );
  IV U7784 ( .A(n7348), .Z(n7405) );
  IV U7785 ( .A(n7349), .Z(n7350) );
  NOR U7786 ( .A(n7351), .B(n7350), .Z(n7356) );
  IV U7787 ( .A(n7352), .Z(n7353) );
  NOR U7788 ( .A(n7354), .B(n7353), .Z(n7355) );
  NOR U7789 ( .A(n7356), .B(n7355), .Z(n7404) );
  IV U7790 ( .A(n7404), .Z(n7357) );
  NOR U7791 ( .A(n7405), .B(n7357), .Z(n7407) );
  XOR U7792 ( .A(n7359), .B(n7358), .Z(n7401) );
  XOR U7793 ( .A(n7361), .B(n7360), .Z(n7372) );
  XOR U7794 ( .A(n7363), .B(n7362), .Z(n7371) );
  IV U7795 ( .A(n7371), .Z(n7364) );
  NOR U7796 ( .A(n7372), .B(n7364), .Z(n7374) );
  NOR U7797 ( .A(n9429), .B(n9241), .Z(n8680) );
  IV U7798 ( .A(n8680), .Z(n8627) );
  IV U7799 ( .A(n7365), .Z(n7366) );
  NOR U7800 ( .A(n8627), .B(n7366), .Z(n7370) );
  NOR U7801 ( .A(n7368), .B(n7367), .Z(n7369) );
  NOR U7802 ( .A(n7370), .B(n7369), .Z(n7417) );
  XOR U7803 ( .A(n7372), .B(n7371), .Z(n7416) );
  NOR U7804 ( .A(n7417), .B(n7416), .Z(n7373) );
  NOR U7805 ( .A(n7374), .B(n7373), .Z(n7400) );
  IV U7806 ( .A(n7400), .Z(n7375) );
  NOR U7807 ( .A(n7401), .B(n7375), .Z(n7403) );
  IV U7808 ( .A(n7376), .Z(n7378) );
  NOR U7809 ( .A(n7378), .B(n7377), .Z(n7382) );
  NOR U7810 ( .A(n7380), .B(n7379), .Z(n7381) );
  NOR U7811 ( .A(n7382), .B(n7381), .Z(n7397) );
  IV U7812 ( .A(n7397), .Z(n7393) );
  XOR U7813 ( .A(n7383), .B(sum[23]), .Z(n7387) );
  NOR U7814 ( .A(n9115), .B(n8862), .Z(n7388) );
  IV U7815 ( .A(n7388), .Z(n7384) );
  NOR U7816 ( .A(n7387), .B(n7384), .Z(n7391) );
  IV U7817 ( .A(sum[22]), .Z(n7386) );
  NOR U7818 ( .A(n9593), .B(n7772), .Z(n7385) );
  IV U7819 ( .A(n7385), .Z(n7578) );
  NOR U7820 ( .A(n7386), .B(n7578), .Z(n7453) );
  IV U7821 ( .A(n7453), .Z(n7389) );
  XOR U7822 ( .A(n7388), .B(n7387), .Z(n7452) );
  NOR U7823 ( .A(n7389), .B(n7452), .Z(n7390) );
  NOR U7824 ( .A(n7391), .B(n7390), .Z(n7392) );
  IV U7825 ( .A(n7392), .Z(n7396) );
  NOR U7826 ( .A(n7393), .B(n7396), .Z(n7399) );
  XOR U7827 ( .A(n7395), .B(n7394), .Z(n7427) );
  XOR U7828 ( .A(n7397), .B(n7396), .Z(n7428) );
  NOR U7829 ( .A(n7427), .B(n7428), .Z(n7398) );
  NOR U7830 ( .A(n7399), .B(n7398), .Z(n7515) );
  XOR U7831 ( .A(n7401), .B(n7400), .Z(n7516) );
  NOR U7832 ( .A(n7515), .B(n7516), .Z(n7402) );
  NOR U7833 ( .A(n7403), .B(n7402), .Z(n7411) );
  XOR U7834 ( .A(n7405), .B(n7404), .Z(n7412) );
  NOR U7835 ( .A(n7411), .B(n7412), .Z(n7406) );
  NOR U7836 ( .A(n7407), .B(n7406), .Z(n7499) );
  IV U7837 ( .A(n7499), .Z(n7408) );
  NOR U7838 ( .A(n7498), .B(n7408), .Z(n7502) );
  XOR U7839 ( .A(n7410), .B(n7409), .Z(n7495) );
  XOR U7840 ( .A(n7412), .B(n7411), .Z(n7494) );
  IV U7841 ( .A(n7494), .Z(n7413) );
  NOR U7842 ( .A(n7495), .B(n7413), .Z(n7497) );
  XOR U7843 ( .A(n7415), .B(n7414), .Z(n7489) );
  XOR U7844 ( .A(n7417), .B(n7416), .Z(n7425) );
  NOR U7845 ( .A(n8499), .B(n9301), .Z(n7421) );
  NOR U7846 ( .A(n9571), .B(n7772), .Z(n7420) );
  NOR U7847 ( .A(n7421), .B(n7420), .Z(n7424) );
  XOR U7848 ( .A(n7419), .B(n7418), .Z(n7434) );
  XOR U7849 ( .A(n7421), .B(n7420), .Z(n7433) );
  IV U7850 ( .A(n7433), .Z(n7422) );
  NOR U7851 ( .A(n7434), .B(n7422), .Z(n7423) );
  NOR U7852 ( .A(n7424), .B(n7423), .Z(n7426) );
  NOR U7853 ( .A(n7425), .B(n7426), .Z(n7432) );
  XOR U7854 ( .A(n7426), .B(n7425), .Z(n7541) );
  IV U7855 ( .A(n7541), .Z(n7430) );
  IV U7856 ( .A(n7427), .Z(n7429) );
  XOR U7857 ( .A(n7429), .B(n7428), .Z(n7542) );
  NOR U7858 ( .A(n7430), .B(n7542), .Z(n7431) );
  NOR U7859 ( .A(n7432), .B(n7431), .Z(n7490) );
  NOR U7860 ( .A(n7489), .B(n7490), .Z(n7493) );
  XOR U7861 ( .A(n7434), .B(n7433), .Z(n7446) );
  IV U7862 ( .A(n7446), .Z(n7437) );
  XOR U7863 ( .A(n7436), .B(n7435), .Z(n7445) );
  NOR U7864 ( .A(n7437), .B(n7445), .Z(n7448) );
  NOR U7865 ( .A(n8729), .B(n9202), .Z(n7438) );
  IV U7866 ( .A(n7438), .Z(n7442) );
  NOR U7867 ( .A(n8228), .B(n9526), .Z(n7441) );
  IV U7868 ( .A(n7441), .Z(n7439) );
  NOR U7869 ( .A(n7442), .B(n7439), .Z(n7444) );
  NOR U7870 ( .A(n9316), .B(n8727), .Z(n7440) );
  IV U7871 ( .A(n7440), .Z(n7591) );
  XOR U7872 ( .A(n7442), .B(n7441), .Z(n7590) );
  NOR U7873 ( .A(n7591), .B(n7590), .Z(n7443) );
  NOR U7874 ( .A(n7444), .B(n7443), .Z(n7545) );
  XOR U7875 ( .A(n7446), .B(n7445), .Z(n7544) );
  NOR U7876 ( .A(n7545), .B(n7544), .Z(n7447) );
  NOR U7877 ( .A(n7448), .B(n7447), .Z(n7449) );
  IV U7878 ( .A(n7449), .Z(n7486) );
  XOR U7879 ( .A(n7451), .B(n7450), .Z(n7472) );
  NOR U7880 ( .A(n8656), .B(n9113), .Z(n7469) );
  NOR U7881 ( .A(n8069), .B(n9526), .Z(n7468) );
  XOR U7882 ( .A(n7469), .B(n7468), .Z(n7470) );
  XOR U7883 ( .A(n7472), .B(n7470), .Z(n7464) );
  IV U7884 ( .A(n7464), .Z(n7454) );
  XOR U7885 ( .A(n7453), .B(n7452), .Z(n7463) );
  NOR U7886 ( .A(n7454), .B(n7463), .Z(n7466) );
  NOR U7887 ( .A(n8656), .B(n9571), .Z(n8679) );
  IV U7888 ( .A(n8679), .Z(n7455) );
  NOR U7889 ( .A(n7456), .B(n7455), .Z(n7462) );
  NOR U7890 ( .A(n8068), .B(n9490), .Z(n7457) );
  IV U7891 ( .A(n7457), .Z(n7620) );
  NOR U7892 ( .A(n9237), .B(n8656), .Z(n7458) );
  XOR U7893 ( .A(n7459), .B(n7458), .Z(n7460) );
  IV U7894 ( .A(n7460), .Z(n7619) );
  NOR U7895 ( .A(n7620), .B(n7619), .Z(n7461) );
  NOR U7896 ( .A(n7462), .B(n7461), .Z(n7554) );
  XOR U7897 ( .A(n7464), .B(n7463), .Z(n7553) );
  NOR U7898 ( .A(n7554), .B(n7553), .Z(n7465) );
  NOR U7899 ( .A(n7466), .B(n7465), .Z(n7485) );
  IV U7900 ( .A(n7485), .Z(n7467) );
  NOR U7901 ( .A(n7486), .B(n7467), .Z(n7488) );
  NOR U7902 ( .A(n7469), .B(n7468), .Z(n7474) );
  IV U7903 ( .A(n7470), .Z(n7471) );
  NOR U7904 ( .A(n7472), .B(n7471), .Z(n7473) );
  NOR U7905 ( .A(n7474), .B(n7473), .Z(n7508) );
  NOR U7906 ( .A(n7476), .B(n7475), .Z(n7480) );
  NOR U7907 ( .A(n7478), .B(n7477), .Z(n7479) );
  NOR U7908 ( .A(n7480), .B(n7479), .Z(n7481) );
  IV U7909 ( .A(n7481), .Z(n7509) );
  XOR U7910 ( .A(n7508), .B(n7509), .Z(n7512) );
  IV U7911 ( .A(n7482), .Z(n7484) );
  XOR U7912 ( .A(n7484), .B(n7483), .Z(n7511) );
  XOR U7913 ( .A(n7512), .B(n7511), .Z(n7606) );
  XOR U7914 ( .A(n7486), .B(n7485), .Z(n7605) );
  NOR U7915 ( .A(n7606), .B(n7605), .Z(n7487) );
  NOR U7916 ( .A(n7488), .B(n7487), .Z(n7574) );
  XOR U7917 ( .A(n7490), .B(n7489), .Z(n7573) );
  IV U7918 ( .A(n7573), .Z(n7491) );
  NOR U7919 ( .A(n7574), .B(n7491), .Z(n7492) );
  NOR U7920 ( .A(n7493), .B(n7492), .Z(n7569) );
  XOR U7921 ( .A(n7495), .B(n7494), .Z(n7568) );
  NOR U7922 ( .A(n7569), .B(n7568), .Z(n7496) );
  NOR U7923 ( .A(n7497), .B(n7496), .Z(n7507) );
  IV U7924 ( .A(n7507), .Z(n7500) );
  XOR U7925 ( .A(n7499), .B(n7498), .Z(n7506) );
  NOR U7926 ( .A(n7500), .B(n7506), .Z(n7501) );
  NOR U7927 ( .A(n7502), .B(n7501), .Z(n9719) );
  IV U7928 ( .A(n9719), .Z(n7505) );
  XOR U7929 ( .A(n7504), .B(n7503), .Z(n9718) );
  NOR U7930 ( .A(n7505), .B(n9718), .Z(n9722) );
  XOR U7931 ( .A(n7507), .B(n7506), .Z(n9714) );
  IV U7932 ( .A(n7508), .Z(n7510) );
  NOR U7933 ( .A(n7510), .B(n7509), .Z(n7514) );
  NOR U7934 ( .A(n7512), .B(n7511), .Z(n7513) );
  NOR U7935 ( .A(n7514), .B(n7513), .Z(n7565) );
  IV U7936 ( .A(n7565), .Z(n7518) );
  IV U7937 ( .A(n7515), .Z(n7517) );
  XOR U7938 ( .A(n7517), .B(n7516), .Z(n7564) );
  NOR U7939 ( .A(n7518), .B(n7564), .Z(n7567) );
  NOR U7940 ( .A(n8016), .B(n7519), .Z(n7525) );
  NOR U7941 ( .A(n8311), .B(n9414), .Z(n7520) );
  IV U7942 ( .A(n7520), .Z(n7594) );
  NOR U7943 ( .A(n9472), .B(n8235), .Z(n7522) );
  NOR U7944 ( .A(n9429), .B(n8499), .Z(n7521) );
  XOR U7945 ( .A(n7522), .B(n7521), .Z(n7523) );
  IV U7946 ( .A(n7523), .Z(n7593) );
  NOR U7947 ( .A(n7594), .B(n7593), .Z(n7524) );
  NOR U7948 ( .A(n7525), .B(n7524), .Z(n7537) );
  XOR U7949 ( .A(n7527), .B(n7526), .Z(n7536) );
  NOR U7950 ( .A(n7537), .B(n7536), .Z(n7540) );
  NOR U7951 ( .A(n9034), .B(n9080), .Z(n7528) );
  IV U7952 ( .A(n7528), .Z(n8558) );
  NOR U7953 ( .A(n9592), .B(n7529), .Z(n7533) );
  IV U7954 ( .A(n7533), .Z(n7530) );
  NOR U7955 ( .A(n8558), .B(n7530), .Z(n7535) );
  NOR U7956 ( .A(n7531), .B(n9600), .Z(n7532) );
  IV U7957 ( .A(n7532), .Z(n7547) );
  XOR U7958 ( .A(n7533), .B(n8558), .Z(n7546) );
  NOR U7959 ( .A(n7547), .B(n7546), .Z(n7534) );
  NOR U7960 ( .A(n7535), .B(n7534), .Z(n7587) );
  XOR U7961 ( .A(n7537), .B(n7536), .Z(n7588) );
  IV U7962 ( .A(n7588), .Z(n7538) );
  NOR U7963 ( .A(n7587), .B(n7538), .Z(n7539) );
  NOR U7964 ( .A(n7540), .B(n7539), .Z(n7561) );
  IV U7965 ( .A(n7561), .Z(n7543) );
  XOR U7966 ( .A(n7542), .B(n7541), .Z(n7560) );
  NOR U7967 ( .A(n7543), .B(n7560), .Z(n7563) );
  XOR U7968 ( .A(n7545), .B(n7544), .Z(n7556) );
  NOR U7969 ( .A(n9599), .B(n7714), .Z(n7548) );
  NOR U7970 ( .A(n8754), .B(n9113), .Z(n7549) );
  NOR U7971 ( .A(n7548), .B(n7549), .Z(n7552) );
  XOR U7972 ( .A(n7547), .B(n7546), .Z(n7679) );
  IV U7973 ( .A(n7548), .Z(n7550) );
  XOR U7974 ( .A(n7550), .B(n7549), .Z(n7680) );
  NOR U7975 ( .A(n7679), .B(n7680), .Z(n7551) );
  NOR U7976 ( .A(n7552), .B(n7551), .Z(n7555) );
  NOR U7977 ( .A(n7556), .B(n7555), .Z(n7559) );
  XOR U7978 ( .A(n7554), .B(n7553), .Z(n7627) );
  IV U7979 ( .A(n7555), .Z(n7557) );
  XOR U7980 ( .A(n7557), .B(n7556), .Z(n7626) );
  NOR U7981 ( .A(n7627), .B(n7626), .Z(n7558) );
  NOR U7982 ( .A(n7559), .B(n7558), .Z(n7647) );
  XOR U7983 ( .A(n7561), .B(n7560), .Z(n7646) );
  NOR U7984 ( .A(n7647), .B(n7646), .Z(n7562) );
  NOR U7985 ( .A(n7563), .B(n7562), .Z(n7576) );
  XOR U7986 ( .A(n7565), .B(n7564), .Z(n7575) );
  NOR U7987 ( .A(n7576), .B(n7575), .Z(n7566) );
  NOR U7988 ( .A(n7567), .B(n7566), .Z(n7572) );
  XOR U7989 ( .A(n7569), .B(n7568), .Z(n7571) );
  IV U7990 ( .A(n7571), .Z(n7570) );
  NOR U7991 ( .A(n7572), .B(n7570), .Z(n7642) );
  XOR U7992 ( .A(n7572), .B(n7571), .Z(n7803) );
  XOR U7993 ( .A(n7574), .B(n7573), .Z(n7636) );
  IV U7994 ( .A(n7636), .Z(n7577) );
  XOR U7995 ( .A(n7576), .B(n7575), .Z(n7635) );
  NOR U7996 ( .A(n7577), .B(n7635), .Z(n7639) );
  XOR U7997 ( .A(n7578), .B(sum[22]), .Z(n7582) );
  NOR U7998 ( .A(n8948), .B(n9115), .Z(n7583) );
  IV U7999 ( .A(n7583), .Z(n7579) );
  NOR U8000 ( .A(n7582), .B(n7579), .Z(n7586) );
  IV U8001 ( .A(sum[21]), .Z(n7581) );
  NOR U8002 ( .A(n9593), .B(n7851), .Z(n7580) );
  IV U8003 ( .A(n7580), .Z(n7748) );
  NOR U8004 ( .A(n7581), .B(n7748), .Z(n7697) );
  IV U8005 ( .A(n7697), .Z(n7584) );
  XOR U8006 ( .A(n7583), .B(n7582), .Z(n7696) );
  NOR U8007 ( .A(n7584), .B(n7696), .Z(n7585) );
  NOR U8008 ( .A(n7586), .B(n7585), .Z(n7601) );
  XOR U8009 ( .A(n7588), .B(n7587), .Z(n7600) );
  NOR U8010 ( .A(n7601), .B(n7600), .Z(n7604) );
  NOR U8011 ( .A(n9260), .B(n8582), .Z(n7648) );
  XOR U8012 ( .A(n7589), .B(n7648), .Z(n7650) );
  XOR U8013 ( .A(n7591), .B(n7590), .Z(n7651) );
  XOR U8014 ( .A(n7650), .B(n7651), .Z(n7597) );
  NOR U8015 ( .A(n8290), .B(n9388), .Z(n7596) );
  IV U8016 ( .A(n7596), .Z(n7592) );
  NOR U8017 ( .A(n7597), .B(n7592), .Z(n7599) );
  XOR U8018 ( .A(n7594), .B(n7593), .Z(n7614) );
  NOR U8019 ( .A(n8422), .B(n9301), .Z(n7612) );
  IV U8020 ( .A(n7612), .Z(n7595) );
  NOR U8021 ( .A(n8069), .B(n9493), .Z(n7611) );
  XOR U8022 ( .A(n7595), .B(n7611), .Z(n7613) );
  XOR U8023 ( .A(n7614), .B(n7613), .Z(n7759) );
  XOR U8024 ( .A(n7597), .B(n7596), .Z(n7760) );
  NOR U8025 ( .A(n7759), .B(n7760), .Z(n7598) );
  NOR U8026 ( .A(n7599), .B(n7598), .Z(n7660) );
  XOR U8027 ( .A(n7601), .B(n7600), .Z(n7661) );
  IV U8028 ( .A(n7661), .Z(n7602) );
  NOR U8029 ( .A(n7660), .B(n7602), .Z(n7603) );
  NOR U8030 ( .A(n7604), .B(n7603), .Z(n7610) );
  IV U8031 ( .A(n7610), .Z(n7608) );
  XOR U8032 ( .A(n7606), .B(n7605), .Z(n7607) );
  IV U8033 ( .A(n7607), .Z(n7609) );
  NOR U8034 ( .A(n7608), .B(n7609), .Z(n7634) );
  XOR U8035 ( .A(n7610), .B(n7609), .Z(n7668) );
  NOR U8036 ( .A(n7612), .B(n7611), .Z(n7616) );
  NOR U8037 ( .A(n7614), .B(n7613), .Z(n7615) );
  NOR U8038 ( .A(n7616), .B(n7615), .Z(n7617) );
  IV U8039 ( .A(n7617), .Z(n7629) );
  NOR U8040 ( .A(n7891), .B(n9584), .Z(n7622) );
  NOR U8041 ( .A(n7618), .B(n7622), .Z(n7624) );
  XOR U8042 ( .A(n7620), .B(n7619), .Z(n7695) );
  XOR U8043 ( .A(n7622), .B(n7621), .Z(n7694) );
  NOR U8044 ( .A(n7695), .B(n7694), .Z(n7623) );
  NOR U8045 ( .A(n7624), .B(n7623), .Z(n7628) );
  IV U8046 ( .A(n7628), .Z(n7625) );
  NOR U8047 ( .A(n7629), .B(n7625), .Z(n7631) );
  XOR U8048 ( .A(n7627), .B(n7626), .Z(n7655) );
  XOR U8049 ( .A(n7629), .B(n7628), .Z(n7654) );
  NOR U8050 ( .A(n7655), .B(n7654), .Z(n7630) );
  NOR U8051 ( .A(n7631), .B(n7630), .Z(n7669) );
  IV U8052 ( .A(n7669), .Z(n7632) );
  NOR U8053 ( .A(n7668), .B(n7632), .Z(n7633) );
  NOR U8054 ( .A(n7634), .B(n7633), .Z(n7645) );
  IV U8055 ( .A(n7645), .Z(n7637) );
  XOR U8056 ( .A(n7636), .B(n7635), .Z(n7644) );
  NOR U8057 ( .A(n7637), .B(n7644), .Z(n7638) );
  NOR U8058 ( .A(n7639), .B(n7638), .Z(n7804) );
  IV U8059 ( .A(n7804), .Z(n7640) );
  NOR U8060 ( .A(n7803), .B(n7640), .Z(n7641) );
  NOR U8061 ( .A(n7642), .B(n7641), .Z(n9715) );
  IV U8062 ( .A(n9715), .Z(n7643) );
  NOR U8063 ( .A(n9714), .B(n7643), .Z(n9717) );
  XOR U8064 ( .A(n7645), .B(n7644), .Z(n7798) );
  XOR U8065 ( .A(n7647), .B(n7646), .Z(n7666) );
  IV U8066 ( .A(n7666), .Z(n7665) );
  NOR U8067 ( .A(n7649), .B(n7648), .Z(n7653) );
  NOR U8068 ( .A(n7651), .B(n7650), .Z(n7652) );
  NOR U8069 ( .A(n7653), .B(n7652), .Z(n7659) );
  IV U8070 ( .A(n7659), .Z(n7657) );
  XOR U8071 ( .A(n7655), .B(n7654), .Z(n7656) );
  IV U8072 ( .A(n7656), .Z(n7658) );
  NOR U8073 ( .A(n7657), .B(n7658), .Z(n7663) );
  XOR U8074 ( .A(n7659), .B(n7658), .Z(n7745) );
  XOR U8075 ( .A(n7661), .B(n7660), .Z(n7746) );
  NOR U8076 ( .A(n7745), .B(n7746), .Z(n7662) );
  NOR U8077 ( .A(n7663), .B(n7662), .Z(n7664) );
  IV U8078 ( .A(n7664), .Z(n7667) );
  NOR U8079 ( .A(n7665), .B(n7667), .Z(n7671) );
  XOR U8080 ( .A(n7667), .B(n7666), .Z(n7739) );
  XOR U8081 ( .A(n7669), .B(n7668), .Z(n7738) );
  NOR U8082 ( .A(n7739), .B(n7738), .Z(n7670) );
  NOR U8083 ( .A(n7671), .B(n7670), .Z(n7799) );
  IV U8084 ( .A(n7799), .Z(n7672) );
  NOR U8085 ( .A(n7798), .B(n7672), .Z(n7802) );
  NOR U8086 ( .A(n8290), .B(n9526), .Z(n7676) );
  IV U8087 ( .A(n7676), .Z(n7674) );
  NOR U8088 ( .A(n8499), .B(n9414), .Z(n7673) );
  IV U8089 ( .A(n7673), .Z(n7675) );
  NOR U8090 ( .A(n7674), .B(n7675), .Z(n7678) );
  XOR U8091 ( .A(n7676), .B(n7675), .Z(n7722) );
  NOR U8092 ( .A(n7723), .B(n7722), .Z(n7677) );
  NOR U8093 ( .A(n7678), .B(n7677), .Z(n7690) );
  XOR U8094 ( .A(n7680), .B(n7679), .Z(n7689) );
  NOR U8095 ( .A(n7690), .B(n7689), .Z(n7693) );
  NOR U8096 ( .A(n9237), .B(n9584), .Z(n7681) );
  IV U8097 ( .A(n7681), .Z(n9082) );
  NOR U8098 ( .A(n9082), .B(n7682), .Z(n7688) );
  NOR U8099 ( .A(n8068), .B(n9571), .Z(n7683) );
  IV U8100 ( .A(n7683), .Z(n7763) );
  NOR U8101 ( .A(n8069), .B(n9584), .Z(n7685) );
  NOR U8102 ( .A(n9237), .B(n8754), .Z(n7684) );
  XOR U8103 ( .A(n7685), .B(n7684), .Z(n7686) );
  IV U8104 ( .A(n7686), .Z(n7762) );
  NOR U8105 ( .A(n7763), .B(n7762), .Z(n7687) );
  NOR U8106 ( .A(n7688), .B(n7687), .Z(n7731) );
  XOR U8107 ( .A(n7690), .B(n7689), .Z(n7732) );
  IV U8108 ( .A(n7732), .Z(n7691) );
  NOR U8109 ( .A(n7731), .B(n7691), .Z(n7692) );
  NOR U8110 ( .A(n7693), .B(n7692), .Z(n7713) );
  IV U8111 ( .A(n7713), .Z(n7711) );
  XOR U8112 ( .A(n7695), .B(n7694), .Z(n7706) );
  XOR U8113 ( .A(n7697), .B(n7696), .Z(n7705) );
  NOR U8114 ( .A(n7706), .B(n7705), .Z(n7709) );
  NOR U8115 ( .A(n9429), .B(n9388), .Z(n9045) );
  IV U8116 ( .A(n9045), .Z(n9041) );
  IV U8117 ( .A(n7698), .Z(n7699) );
  NOR U8118 ( .A(n9041), .B(n7699), .Z(n7704) );
  NOR U8119 ( .A(n9316), .B(n8862), .Z(n7700) );
  IV U8120 ( .A(n7700), .Z(n7780) );
  NOR U8121 ( .A(n8501), .B(n9388), .Z(n7701) );
  NOR U8122 ( .A(n8422), .B(n9429), .Z(n7838) );
  XOR U8123 ( .A(n7701), .B(n7838), .Z(n7702) );
  IV U8124 ( .A(n7702), .Z(n7779) );
  NOR U8125 ( .A(n7780), .B(n7779), .Z(n7703) );
  NOR U8126 ( .A(n7704), .B(n7703), .Z(n7758) );
  XOR U8127 ( .A(n7706), .B(n7705), .Z(n7757) );
  IV U8128 ( .A(n7757), .Z(n7707) );
  NOR U8129 ( .A(n7758), .B(n7707), .Z(n7708) );
  NOR U8130 ( .A(n7709), .B(n7708), .Z(n7710) );
  IV U8131 ( .A(n7710), .Z(n7712) );
  NOR U8132 ( .A(n7711), .B(n7712), .Z(n7737) );
  XOR U8133 ( .A(n7713), .B(n7712), .Z(n7744) );
  NOR U8134 ( .A(n9592), .B(n7714), .Z(n7719) );
  IV U8135 ( .A(n7719), .Z(n7716) );
  NOR U8136 ( .A(n9034), .B(n9113), .Z(n7715) );
  IV U8137 ( .A(n7715), .Z(n7718) );
  NOR U8138 ( .A(n7716), .B(n7718), .Z(n7721) );
  NOR U8139 ( .A(n7891), .B(n9599), .Z(n7717) );
  IV U8140 ( .A(n7717), .Z(n7774) );
  XOR U8141 ( .A(n7719), .B(n7718), .Z(n7773) );
  NOR U8142 ( .A(n7774), .B(n7773), .Z(n7720) );
  NOR U8143 ( .A(n7721), .B(n7720), .Z(n7730) );
  NOR U8144 ( .A(n8311), .B(n9472), .Z(n7724) );
  NOR U8145 ( .A(n8948), .B(n9241), .Z(n7725) );
  NOR U8146 ( .A(n7724), .B(n7725), .Z(n7727) );
  XOR U8147 ( .A(n7723), .B(n7722), .Z(n7886) );
  IV U8148 ( .A(n7724), .Z(n8309) );
  XOR U8149 ( .A(n7725), .B(n8309), .Z(n7887) );
  NOR U8150 ( .A(n7886), .B(n7887), .Z(n7726) );
  NOR U8151 ( .A(n7727), .B(n7726), .Z(n7729) );
  IV U8152 ( .A(n7729), .Z(n7728) );
  NOR U8153 ( .A(n7730), .B(n7728), .Z(n7734) );
  XOR U8154 ( .A(n7730), .B(n7729), .Z(n7787) );
  XOR U8155 ( .A(n7732), .B(n7731), .Z(n7788) );
  NOR U8156 ( .A(n7787), .B(n7788), .Z(n7733) );
  NOR U8157 ( .A(n7734), .B(n7733), .Z(n7735) );
  IV U8158 ( .A(n7735), .Z(n7743) );
  NOR U8159 ( .A(n7744), .B(n7743), .Z(n7736) );
  NOR U8160 ( .A(n7737), .B(n7736), .Z(n7742) );
  XOR U8161 ( .A(n7739), .B(n7738), .Z(n7741) );
  IV U8162 ( .A(n7741), .Z(n7740) );
  NOR U8163 ( .A(n7742), .B(n7740), .Z(n7797) );
  XOR U8164 ( .A(n7742), .B(n7741), .Z(n7810) );
  XOR U8165 ( .A(n7744), .B(n7743), .Z(n7792) );
  XOR U8166 ( .A(n7746), .B(n7745), .Z(n7791) );
  IV U8167 ( .A(n7791), .Z(n7747) );
  NOR U8168 ( .A(n7792), .B(n7747), .Z(n7794) );
  XOR U8169 ( .A(n7748), .B(sum[21]), .Z(n7752) );
  NOR U8170 ( .A(n7749), .B(n7752), .Z(n7756) );
  IV U8171 ( .A(sum[20]), .Z(n7751) );
  NOR U8172 ( .A(n8068), .B(n9593), .Z(n7750) );
  IV U8173 ( .A(n7750), .Z(n7942) );
  NOR U8174 ( .A(n7751), .B(n7942), .Z(n7864) );
  IV U8175 ( .A(n7864), .Z(n7754) );
  XOR U8176 ( .A(n7753), .B(n7752), .Z(n7863) );
  NOR U8177 ( .A(n7754), .B(n7863), .Z(n7755) );
  NOR U8178 ( .A(n7756), .B(n7755), .Z(n7816) );
  IV U8179 ( .A(n7816), .Z(n7761) );
  XOR U8180 ( .A(n7758), .B(n7757), .Z(n7814) );
  XOR U8181 ( .A(n7760), .B(n7759), .Z(n7812) );
  XOR U8182 ( .A(n7814), .B(n7812), .Z(n7815) );
  XOR U8183 ( .A(n7761), .B(n7815), .Z(n7770) );
  NOR U8184 ( .A(n8656), .B(n9202), .Z(n7764) );
  NOR U8185 ( .A(n8228), .B(n9493), .Z(n7765) );
  NOR U8186 ( .A(n7764), .B(n7765), .Z(n7768) );
  XOR U8187 ( .A(n7763), .B(n7762), .Z(n7847) );
  IV U8188 ( .A(n7764), .Z(n7766) );
  XOR U8189 ( .A(n7766), .B(n7765), .Z(n7846) );
  NOR U8190 ( .A(n7847), .B(n7846), .Z(n7767) );
  NOR U8191 ( .A(n7768), .B(n7767), .Z(n7771) );
  IV U8192 ( .A(n7771), .Z(n7769) );
  NOR U8193 ( .A(n7770), .B(n7769), .Z(n7790) );
  XOR U8194 ( .A(n7771), .B(n7770), .Z(n7912) );
  NOR U8195 ( .A(n8729), .B(n9301), .Z(n7775) );
  NOR U8196 ( .A(n9600), .B(n7772), .Z(n7776) );
  NOR U8197 ( .A(n7775), .B(n7776), .Z(n7778) );
  XOR U8198 ( .A(n7774), .B(n7773), .Z(n7889) );
  IV U8199 ( .A(n7775), .Z(n8770) );
  XOR U8200 ( .A(n7776), .B(n8770), .Z(n7888) );
  NOR U8201 ( .A(n7889), .B(n7888), .Z(n7777) );
  NOR U8202 ( .A(n7778), .B(n7777), .Z(n7819) );
  NOR U8203 ( .A(n8582), .B(n9336), .Z(n7782) );
  NOR U8204 ( .A(n9260), .B(n8727), .Z(n7781) );
  NOR U8205 ( .A(n7782), .B(n7781), .Z(n7785) );
  XOR U8206 ( .A(n7780), .B(n7779), .Z(n7862) );
  XOR U8207 ( .A(n7782), .B(n7781), .Z(n7861) );
  IV U8208 ( .A(n7861), .Z(n7783) );
  NOR U8209 ( .A(n7862), .B(n7783), .Z(n7784) );
  NOR U8210 ( .A(n7785), .B(n7784), .Z(n7786) );
  IV U8211 ( .A(n7786), .Z(n7820) );
  XOR U8212 ( .A(n7819), .B(n7820), .Z(n7824) );
  XOR U8213 ( .A(n7788), .B(n7787), .Z(n7822) );
  XOR U8214 ( .A(n7824), .B(n7822), .Z(n7911) );
  NOR U8215 ( .A(n7912), .B(n7911), .Z(n7789) );
  NOR U8216 ( .A(n7790), .B(n7789), .Z(n7830) );
  XOR U8217 ( .A(n7792), .B(n7791), .Z(n7829) );
  NOR U8218 ( .A(n7830), .B(n7829), .Z(n7793) );
  NOR U8219 ( .A(n7794), .B(n7793), .Z(n7811) );
  IV U8220 ( .A(n7811), .Z(n7795) );
  NOR U8221 ( .A(n7810), .B(n7795), .Z(n7796) );
  NOR U8222 ( .A(n7797), .B(n7796), .Z(n7809) );
  IV U8223 ( .A(n7809), .Z(n7800) );
  XOR U8224 ( .A(n7799), .B(n7798), .Z(n7808) );
  NOR U8225 ( .A(n7800), .B(n7808), .Z(n7801) );
  NOR U8226 ( .A(n7802), .B(n7801), .Z(n7807) );
  IV U8227 ( .A(n7807), .Z(n7805) );
  XOR U8228 ( .A(n7804), .B(n7803), .Z(n7806) );
  NOR U8229 ( .A(n7805), .B(n7806), .Z(n9712) );
  XOR U8230 ( .A(n7807), .B(n7806), .Z(n9774) );
  XOR U8231 ( .A(n7809), .B(n7808), .Z(n7935) );
  XOR U8232 ( .A(n7811), .B(n7810), .Z(n7836) );
  IV U8233 ( .A(n7812), .Z(n7813) );
  NOR U8234 ( .A(n7814), .B(n7813), .Z(n7818) );
  NOR U8235 ( .A(n7816), .B(n7815), .Z(n7817) );
  NOR U8236 ( .A(n7818), .B(n7817), .Z(n7828) );
  IV U8237 ( .A(n7819), .Z(n7821) );
  NOR U8238 ( .A(n7821), .B(n7820), .Z(n7826) );
  IV U8239 ( .A(n7822), .Z(n7823) );
  NOR U8240 ( .A(n7824), .B(n7823), .Z(n7825) );
  NOR U8241 ( .A(n7826), .B(n7825), .Z(n7827) );
  NOR U8242 ( .A(n7828), .B(n7827), .Z(n7834) );
  XOR U8243 ( .A(n7828), .B(n7827), .Z(n7928) );
  IV U8244 ( .A(n7928), .Z(n7832) );
  XOR U8245 ( .A(n7830), .B(n7829), .Z(n7831) );
  IV U8246 ( .A(n7831), .Z(n7927) );
  NOR U8247 ( .A(n7832), .B(n7927), .Z(n7833) );
  NOR U8248 ( .A(n7834), .B(n7833), .Z(n7837) );
  IV U8249 ( .A(n7837), .Z(n7835) );
  NOR U8250 ( .A(n7836), .B(n7835), .Z(n7933) );
  XOR U8251 ( .A(n7837), .B(n7836), .Z(n8101) );
  IV U8252 ( .A(n7838), .Z(n7839) );
  NOR U8253 ( .A(n9414), .B(n8729), .Z(n8137) );
  IV U8254 ( .A(n8137), .Z(n8119) );
  NOR U8255 ( .A(n7839), .B(n8119), .Z(n7845) );
  NOR U8256 ( .A(n8228), .B(n9584), .Z(n7840) );
  IV U8257 ( .A(n7840), .Z(n7955) );
  NOR U8258 ( .A(n9429), .B(n8729), .Z(n7842) );
  NOR U8259 ( .A(n8422), .B(n9414), .Z(n7841) );
  XOR U8260 ( .A(n7842), .B(n7841), .Z(n7843) );
  IV U8261 ( .A(n7843), .Z(n7954) );
  NOR U8262 ( .A(n7955), .B(n7954), .Z(n7844) );
  NOR U8263 ( .A(n7845), .B(n7844), .Z(n7857) );
  XOR U8264 ( .A(n7847), .B(n7846), .Z(n7856) );
  NOR U8265 ( .A(n7857), .B(n7856), .Z(n7860) );
  NOR U8266 ( .A(n9600), .B(n8754), .Z(n8951) );
  IV U8267 ( .A(n8951), .Z(n7848) );
  NOR U8268 ( .A(n7849), .B(n7848), .Z(n7855) );
  NOR U8269 ( .A(n9571), .B(n8235), .Z(n7850) );
  IV U8270 ( .A(n7850), .Z(n7893) );
  NOR U8271 ( .A(n8754), .B(n9202), .Z(n8356) );
  NOR U8272 ( .A(n9600), .B(n7851), .Z(n7852) );
  XOR U8273 ( .A(n8356), .B(n7852), .Z(n7853) );
  IV U8274 ( .A(n7853), .Z(n7892) );
  NOR U8275 ( .A(n7893), .B(n7892), .Z(n7854) );
  NOR U8276 ( .A(n7855), .B(n7854), .Z(n7963) );
  XOR U8277 ( .A(n7857), .B(n7856), .Z(n7964) );
  IV U8278 ( .A(n7964), .Z(n7858) );
  NOR U8279 ( .A(n7963), .B(n7858), .Z(n7859) );
  NOR U8280 ( .A(n7860), .B(n7859), .Z(n7879) );
  IV U8281 ( .A(n7879), .Z(n7877) );
  XOR U8282 ( .A(n7862), .B(n7861), .Z(n7873) );
  IV U8283 ( .A(n7873), .Z(n7865) );
  XOR U8284 ( .A(n7864), .B(n7863), .Z(n7872) );
  NOR U8285 ( .A(n7865), .B(n7872), .Z(n7875) );
  NOR U8286 ( .A(n9526), .B(n9301), .Z(n9058) );
  IV U8287 ( .A(n9058), .Z(n9362) );
  NOR U8288 ( .A(n8248), .B(n9362), .Z(n7871) );
  NOR U8289 ( .A(n8727), .B(n9336), .Z(n7952) );
  IV U8290 ( .A(n7952), .Z(n7869) );
  NOR U8291 ( .A(n8656), .B(n9301), .Z(n7866) );
  IV U8292 ( .A(n7866), .Z(n7868) );
  NOR U8293 ( .A(n8501), .B(n9526), .Z(n7867) );
  XOR U8294 ( .A(n7868), .B(n7867), .Z(n7951) );
  NOR U8295 ( .A(n7869), .B(n7951), .Z(n7870) );
  NOR U8296 ( .A(n7871), .B(n7870), .Z(n7899) );
  XOR U8297 ( .A(n7873), .B(n7872), .Z(n7898) );
  NOR U8298 ( .A(n7899), .B(n7898), .Z(n7874) );
  NOR U8299 ( .A(n7875), .B(n7874), .Z(n7876) );
  IV U8300 ( .A(n7876), .Z(n7878) );
  NOR U8301 ( .A(n7877), .B(n7878), .Z(n7915) );
  XOR U8302 ( .A(n7879), .B(n7878), .Z(n7941) );
  NOR U8303 ( .A(n9316), .B(n9490), .Z(n9074) );
  IV U8304 ( .A(n9074), .Z(n9313) );
  NOR U8305 ( .A(n7880), .B(n9313), .Z(n7885) );
  NOR U8306 ( .A(n8311), .B(n9490), .Z(n7882) );
  NOR U8307 ( .A(n8948), .B(n9316), .Z(n7881) );
  XOR U8308 ( .A(n7882), .B(n7881), .Z(n7883) );
  IV U8309 ( .A(n7883), .Z(n7973) );
  NOR U8310 ( .A(n8016), .B(n7973), .Z(n7884) );
  NOR U8311 ( .A(n7885), .B(n7884), .Z(n7908) );
  XOR U8312 ( .A(n7887), .B(n7886), .Z(n7906) );
  IV U8313 ( .A(n7906), .Z(n7890) );
  XOR U8314 ( .A(n7889), .B(n7888), .Z(n7905) );
  XOR U8315 ( .A(n7890), .B(n7905), .Z(n7907) );
  XOR U8316 ( .A(n7908), .B(n7907), .Z(n7901) );
  NOR U8317 ( .A(n9034), .B(n9237), .Z(n7894) );
  NOR U8318 ( .A(n7891), .B(n9592), .Z(n7895) );
  NOR U8319 ( .A(n7894), .B(n7895), .Z(n7897) );
  XOR U8320 ( .A(n7893), .B(n7892), .Z(n8051) );
  IV U8321 ( .A(n7894), .Z(n8712) );
  XOR U8322 ( .A(n7895), .B(n8712), .Z(n8050) );
  NOR U8323 ( .A(n8051), .B(n8050), .Z(n7896) );
  NOR U8324 ( .A(n7897), .B(n7896), .Z(n7900) );
  NOR U8325 ( .A(n7901), .B(n7900), .Z(n7904) );
  XOR U8326 ( .A(n7899), .B(n7898), .Z(n7987) );
  IV U8327 ( .A(n7900), .Z(n7902) );
  XOR U8328 ( .A(n7902), .B(n7901), .Z(n7986) );
  NOR U8329 ( .A(n7987), .B(n7986), .Z(n7903) );
  NOR U8330 ( .A(n7904), .B(n7903), .Z(n7921) );
  NOR U8331 ( .A(n7906), .B(n7905), .Z(n7910) );
  NOR U8332 ( .A(n7908), .B(n7907), .Z(n7909) );
  NOR U8333 ( .A(n7910), .B(n7909), .Z(n7917) );
  XOR U8334 ( .A(n7912), .B(n7911), .Z(n7919) );
  XOR U8335 ( .A(n7917), .B(n7919), .Z(n7920) );
  XOR U8336 ( .A(n7921), .B(n7920), .Z(n7940) );
  IV U8337 ( .A(n7940), .Z(n7913) );
  NOR U8338 ( .A(n7941), .B(n7913), .Z(n7914) );
  NOR U8339 ( .A(n7915), .B(n7914), .Z(n7916) );
  IV U8340 ( .A(n7916), .Z(n7926) );
  IV U8341 ( .A(n7917), .Z(n7918) );
  NOR U8342 ( .A(n7919), .B(n7918), .Z(n7923) );
  NOR U8343 ( .A(n7921), .B(n7920), .Z(n7922) );
  NOR U8344 ( .A(n7923), .B(n7922), .Z(n7925) );
  IV U8345 ( .A(n7925), .Z(n7924) );
  NOR U8346 ( .A(n7926), .B(n7924), .Z(n7930) );
  XOR U8347 ( .A(n7926), .B(n7925), .Z(n7938) );
  XOR U8348 ( .A(n7928), .B(n7927), .Z(n7937) );
  NOR U8349 ( .A(n7938), .B(n7937), .Z(n7929) );
  NOR U8350 ( .A(n7930), .B(n7929), .Z(n8102) );
  IV U8351 ( .A(n8102), .Z(n7931) );
  NOR U8352 ( .A(n8101), .B(n7931), .Z(n7932) );
  NOR U8353 ( .A(n7933), .B(n7932), .Z(n7936) );
  IV U8354 ( .A(n7936), .Z(n7934) );
  NOR U8355 ( .A(n7935), .B(n7934), .Z(n9709) );
  XOR U8356 ( .A(n7936), .B(n7935), .Z(n9779) );
  XOR U8357 ( .A(n7938), .B(n7937), .Z(n7939) );
  IV U8358 ( .A(n7939), .Z(n7996) );
  XOR U8359 ( .A(n7941), .B(n7940), .Z(n7969) );
  NOR U8360 ( .A(n9080), .B(n9241), .Z(n7947) );
  IV U8361 ( .A(n7947), .Z(n7943) );
  XOR U8362 ( .A(n7942), .B(sum[20]), .Z(n7946) );
  NOR U8363 ( .A(n7943), .B(n7946), .Z(n7950) );
  IV U8364 ( .A(sum[19]), .Z(n7945) );
  NOR U8365 ( .A(n9593), .B(n8235), .Z(n7944) );
  IV U8366 ( .A(n7944), .Z(n8023) );
  NOR U8367 ( .A(n7945), .B(n8023), .Z(n8001) );
  IV U8368 ( .A(n8001), .Z(n7948) );
  XOR U8369 ( .A(n7947), .B(n7946), .Z(n8000) );
  NOR U8370 ( .A(n7948), .B(n8000), .Z(n7949) );
  NOR U8371 ( .A(n7950), .B(n7949), .Z(n7962) );
  XOR U8372 ( .A(n7952), .B(n7951), .Z(n7957) );
  NOR U8373 ( .A(n7953), .B(n7957), .Z(n7960) );
  XOR U8374 ( .A(n7955), .B(n7954), .Z(n7982) );
  NOR U8375 ( .A(n8290), .B(n9493), .Z(n7980) );
  NOR U8376 ( .A(n9115), .B(n9113), .Z(n7979) );
  XOR U8377 ( .A(n7980), .B(n7979), .Z(n7956) );
  IV U8378 ( .A(n7956), .Z(n7981) );
  XOR U8379 ( .A(n7982), .B(n7981), .Z(n7998) );
  XOR U8380 ( .A(n7958), .B(n7957), .Z(n7999) );
  NOR U8381 ( .A(n7998), .B(n7999), .Z(n7959) );
  NOR U8382 ( .A(n7960), .B(n7959), .Z(n7961) );
  NOR U8383 ( .A(n7962), .B(n7961), .Z(n7967) );
  XOR U8384 ( .A(n7962), .B(n7961), .Z(n8015) );
  IV U8385 ( .A(n8015), .Z(n7965) );
  XOR U8386 ( .A(n7964), .B(n7963), .Z(n8014) );
  NOR U8387 ( .A(n7965), .B(n8014), .Z(n7966) );
  NOR U8388 ( .A(n7967), .B(n7966), .Z(n7970) );
  IV U8389 ( .A(n7970), .Z(n7968) );
  NOR U8390 ( .A(n7969), .B(n7968), .Z(n7994) );
  XOR U8391 ( .A(n7970), .B(n7969), .Z(n8045) );
  NOR U8392 ( .A(n9599), .B(n8862), .Z(n8737) );
  IV U8393 ( .A(n8737), .Z(n8739) );
  NOR U8394 ( .A(n7971), .B(n8739), .Z(n7978) );
  XOR U8395 ( .A(n7973), .B(n7972), .Z(n8052) );
  NOR U8396 ( .A(n8069), .B(n9599), .Z(n7975) );
  NOR U8397 ( .A(n9260), .B(n8862), .Z(n7974) );
  XOR U8398 ( .A(n7975), .B(n7974), .Z(n8053) );
  IV U8399 ( .A(n8053), .Z(n7976) );
  NOR U8400 ( .A(n8052), .B(n7976), .Z(n7977) );
  NOR U8401 ( .A(n7978), .B(n7977), .Z(n7989) );
  NOR U8402 ( .A(n7980), .B(n7979), .Z(n7984) );
  NOR U8403 ( .A(n7982), .B(n7981), .Z(n7983) );
  NOR U8404 ( .A(n7984), .B(n7983), .Z(n7988) );
  IV U8405 ( .A(n7988), .Z(n7985) );
  NOR U8406 ( .A(n7989), .B(n7985), .Z(n7991) );
  XOR U8407 ( .A(n7987), .B(n7986), .Z(n8049) );
  XOR U8408 ( .A(n7989), .B(n7988), .Z(n8048) );
  NOR U8409 ( .A(n8049), .B(n8048), .Z(n7990) );
  NOR U8410 ( .A(n7991), .B(n7990), .Z(n8046) );
  IV U8411 ( .A(n8046), .Z(n7992) );
  NOR U8412 ( .A(n8045), .B(n7992), .Z(n7993) );
  NOR U8413 ( .A(n7994), .B(n7993), .Z(n7997) );
  IV U8414 ( .A(n7997), .Z(n7995) );
  NOR U8415 ( .A(n7996), .B(n7995), .Z(n8100) );
  XOR U8416 ( .A(n7997), .B(n7996), .Z(n8104) );
  XOR U8417 ( .A(n7999), .B(n7998), .Z(n8011) );
  IV U8418 ( .A(n8011), .Z(n8002) );
  XOR U8419 ( .A(n8001), .B(n8000), .Z(n8010) );
  NOR U8420 ( .A(n8002), .B(n8010), .Z(n8013) );
  NOR U8421 ( .A(n9080), .B(n9599), .Z(n8971) );
  IV U8422 ( .A(n8971), .Z(n8930) );
  NOR U8423 ( .A(n8003), .B(n8930), .Z(n8009) );
  NOR U8424 ( .A(n8290), .B(n9584), .Z(n8004) );
  IV U8425 ( .A(n8004), .Z(n8118) );
  NOR U8426 ( .A(n8228), .B(n9599), .Z(n8006) );
  NOR U8427 ( .A(n9316), .B(n9080), .Z(n8005) );
  XOR U8428 ( .A(n8006), .B(n8005), .Z(n8007) );
  IV U8429 ( .A(n8007), .Z(n8117) );
  NOR U8430 ( .A(n8118), .B(n8117), .Z(n8008) );
  NOR U8431 ( .A(n8009), .B(n8008), .Z(n8036) );
  XOR U8432 ( .A(n8011), .B(n8010), .Z(n8035) );
  NOR U8433 ( .A(n8036), .B(n8035), .Z(n8012) );
  NOR U8434 ( .A(n8013), .B(n8012), .Z(n8041) );
  XOR U8435 ( .A(n8015), .B(n8014), .Z(n8040) );
  NOR U8436 ( .A(n8041), .B(n8040), .Z(n8044) );
  NOR U8437 ( .A(n8422), .B(n9490), .Z(n8262) );
  IV U8438 ( .A(n8262), .Z(n8265) );
  NOR U8439 ( .A(n8016), .B(n8265), .Z(n8022) );
  NOR U8440 ( .A(n9429), .B(n8656), .Z(n8017) );
  IV U8441 ( .A(n8017), .Z(n8116) );
  NOR U8442 ( .A(n8499), .B(n9490), .Z(n8019) );
  NOR U8443 ( .A(n8422), .B(n9472), .Z(n8018) );
  XOR U8444 ( .A(n8019), .B(n8018), .Z(n8020) );
  IV U8445 ( .A(n8020), .Z(n8115) );
  NOR U8446 ( .A(n8116), .B(n8115), .Z(n8021) );
  NOR U8447 ( .A(n8022), .B(n8021), .Z(n8033) );
  XOR U8448 ( .A(n8023), .B(sum[19]), .Z(n8027) );
  NOR U8449 ( .A(n9241), .B(n9113), .Z(n8028) );
  IV U8450 ( .A(n8028), .Z(n8024) );
  NOR U8451 ( .A(n8027), .B(n8024), .Z(n8031) );
  IV U8452 ( .A(sum[18]), .Z(n8026) );
  NOR U8453 ( .A(n8311), .B(n9593), .Z(n8025) );
  IV U8454 ( .A(n8025), .Z(n8184) );
  NOR U8455 ( .A(n8026), .B(n8184), .Z(n8172) );
  IV U8456 ( .A(n8172), .Z(n8029) );
  XOR U8457 ( .A(n8028), .B(n8027), .Z(n8171) );
  NOR U8458 ( .A(n8029), .B(n8171), .Z(n8030) );
  NOR U8459 ( .A(n8031), .B(n8030), .Z(n8032) );
  NOR U8460 ( .A(n8033), .B(n8032), .Z(n8039) );
  XOR U8461 ( .A(n8033), .B(n8032), .Z(n8034) );
  IV U8462 ( .A(n8034), .Z(n8135) );
  XOR U8463 ( .A(n8036), .B(n8035), .Z(n8134) );
  IV U8464 ( .A(n8134), .Z(n8037) );
  NOR U8465 ( .A(n8135), .B(n8037), .Z(n8038) );
  NOR U8466 ( .A(n8039), .B(n8038), .Z(n8112) );
  XOR U8467 ( .A(n8041), .B(n8040), .Z(n8111) );
  IV U8468 ( .A(n8111), .Z(n8042) );
  NOR U8469 ( .A(n8112), .B(n8042), .Z(n8043) );
  NOR U8470 ( .A(n8044), .B(n8043), .Z(n8095) );
  IV U8471 ( .A(n8095), .Z(n8047) );
  XOR U8472 ( .A(n8046), .B(n8045), .Z(n8094) );
  NOR U8473 ( .A(n8047), .B(n8094), .Z(n8097) );
  XOR U8474 ( .A(n8049), .B(n8048), .Z(n8091) );
  XOR U8475 ( .A(n8051), .B(n8050), .Z(n8060) );
  XOR U8476 ( .A(n8053), .B(n8052), .Z(n8059) );
  NOR U8477 ( .A(n8060), .B(n8059), .Z(n8063) );
  NOR U8478 ( .A(n9237), .B(n9388), .Z(n8715) );
  IV U8479 ( .A(n8715), .Z(n9236) );
  NOR U8480 ( .A(n8054), .B(n9236), .Z(n8058) );
  NOR U8481 ( .A(n9336), .B(n8862), .Z(n8173) );
  IV U8482 ( .A(n8173), .Z(n8195) );
  NOR U8483 ( .A(n8727), .B(n9388), .Z(n8055) );
  IV U8484 ( .A(n8055), .Z(n8056) );
  NOR U8485 ( .A(n9237), .B(n9115), .Z(n8868) );
  XOR U8486 ( .A(n8056), .B(n8868), .Z(n8174) );
  NOR U8487 ( .A(n8195), .B(n8174), .Z(n8057) );
  NOR U8488 ( .A(n8058), .B(n8057), .Z(n8066) );
  XOR U8489 ( .A(n8060), .B(n8059), .Z(n8061) );
  IV U8490 ( .A(n8061), .Z(n8065) );
  NOR U8491 ( .A(n8066), .B(n8065), .Z(n8062) );
  NOR U8492 ( .A(n8063), .B(n8062), .Z(n8090) );
  IV U8493 ( .A(n8090), .Z(n8064) );
  NOR U8494 ( .A(n8091), .B(n8064), .Z(n8093) );
  XOR U8495 ( .A(n8066), .B(n8065), .Z(n8078) );
  NOR U8496 ( .A(n9592), .B(n9202), .Z(n9303) );
  IV U8497 ( .A(n9303), .Z(n8861) );
  NOR U8498 ( .A(n8067), .B(n8861), .Z(n8075) );
  NOR U8499 ( .A(n8068), .B(n9600), .Z(n8081) );
  IV U8500 ( .A(n8081), .Z(n8073) );
  NOR U8501 ( .A(n8069), .B(n9592), .Z(n8070) );
  IV U8502 ( .A(n8070), .Z(n8072) );
  NOR U8503 ( .A(n9034), .B(n9202), .Z(n8071) );
  XOR U8504 ( .A(n8072), .B(n8071), .Z(n8080) );
  NOR U8505 ( .A(n8073), .B(n8080), .Z(n8074) );
  NOR U8506 ( .A(n8075), .B(n8074), .Z(n8077) );
  IV U8507 ( .A(n8077), .Z(n8076) );
  NOR U8508 ( .A(n8078), .B(n8076), .Z(n8089) );
  XOR U8509 ( .A(n8078), .B(n8077), .Z(n8113) );
  NOR U8510 ( .A(n8754), .B(n9571), .Z(n8726) );
  IV U8511 ( .A(n8726), .Z(n8734) );
  NOR U8512 ( .A(n8079), .B(n8734), .Z(n8086) );
  XOR U8513 ( .A(n8081), .B(n8080), .Z(n8177) );
  NOR U8514 ( .A(n8754), .B(n9301), .Z(n8083) );
  NOR U8515 ( .A(n8311), .B(n9571), .Z(n8082) );
  XOR U8516 ( .A(n8083), .B(n8082), .Z(n8178) );
  IV U8517 ( .A(n8178), .Z(n8084) );
  NOR U8518 ( .A(n8177), .B(n8084), .Z(n8085) );
  NOR U8519 ( .A(n8086), .B(n8085), .Z(n8114) );
  IV U8520 ( .A(n8114), .Z(n8087) );
  NOR U8521 ( .A(n8113), .B(n8087), .Z(n8088) );
  NOR U8522 ( .A(n8089), .B(n8088), .Z(n8110) );
  XOR U8523 ( .A(n8091), .B(n8090), .Z(n8109) );
  NOR U8524 ( .A(n8110), .B(n8109), .Z(n8092) );
  NOR U8525 ( .A(n8093), .B(n8092), .Z(n8106) );
  XOR U8526 ( .A(n8095), .B(n8094), .Z(n8107) );
  NOR U8527 ( .A(n8106), .B(n8107), .Z(n8096) );
  NOR U8528 ( .A(n8097), .B(n8096), .Z(n8105) );
  IV U8529 ( .A(n8105), .Z(n8098) );
  NOR U8530 ( .A(n8104), .B(n8098), .Z(n8099) );
  NOR U8531 ( .A(n8100), .B(n8099), .Z(n9703) );
  IV U8532 ( .A(n9703), .Z(n8103) );
  XOR U8533 ( .A(n8102), .B(n8101), .Z(n9702) );
  NOR U8534 ( .A(n8103), .B(n9702), .Z(n9706) );
  XOR U8535 ( .A(n8105), .B(n8104), .Z(n9698) );
  IV U8536 ( .A(n8106), .Z(n8108) );
  XOR U8537 ( .A(n8108), .B(n8107), .Z(n8160) );
  XOR U8538 ( .A(n8110), .B(n8109), .Z(n8154) );
  XOR U8539 ( .A(n8112), .B(n8111), .Z(n8153) );
  NOR U8540 ( .A(n8154), .B(n8153), .Z(n8158) );
  XOR U8541 ( .A(n8114), .B(n8113), .Z(n8149) );
  XOR U8542 ( .A(n8116), .B(n8115), .Z(n8145) );
  NOR U8543 ( .A(n8582), .B(n9526), .Z(n8142) );
  NOR U8544 ( .A(n9260), .B(n8948), .Z(n8143) );
  IV U8545 ( .A(n8143), .Z(n8830) );
  XOR U8546 ( .A(n8142), .B(n8830), .Z(n8144) );
  XOR U8547 ( .A(n8145), .B(n8144), .Z(n8129) );
  XOR U8548 ( .A(n8118), .B(n8117), .Z(n8139) );
  NOR U8549 ( .A(n8501), .B(n9493), .Z(n8136) );
  XOR U8550 ( .A(n8136), .B(n8119), .Z(n8138) );
  XOR U8551 ( .A(n8139), .B(n8138), .Z(n8128) );
  NOR U8552 ( .A(n8129), .B(n8128), .Z(n8132) );
  IV U8553 ( .A(n8120), .Z(n8121) );
  NOR U8554 ( .A(n9237), .B(n9493), .Z(n8985) );
  IV U8555 ( .A(n8985), .Z(n8980) );
  NOR U8556 ( .A(n8121), .B(n8980), .Z(n8127) );
  NOR U8557 ( .A(n9472), .B(n8729), .Z(n8122) );
  IV U8558 ( .A(n8122), .Z(n8197) );
  NOR U8559 ( .A(n8582), .B(n9493), .Z(n8124) );
  NOR U8560 ( .A(n9237), .B(n9241), .Z(n8123) );
  XOR U8561 ( .A(n8124), .B(n8123), .Z(n8125) );
  IV U8562 ( .A(n8125), .Z(n8196) );
  NOR U8563 ( .A(n8197), .B(n8196), .Z(n8126) );
  NOR U8564 ( .A(n8127), .B(n8126), .Z(n8225) );
  XOR U8565 ( .A(n8129), .B(n8128), .Z(n8130) );
  IV U8566 ( .A(n8130), .Z(n8224) );
  NOR U8567 ( .A(n8225), .B(n8224), .Z(n8131) );
  NOR U8568 ( .A(n8132), .B(n8131), .Z(n8150) );
  IV U8569 ( .A(n8150), .Z(n8133) );
  NOR U8570 ( .A(n8149), .B(n8133), .Z(n8152) );
  XOR U8571 ( .A(n8135), .B(n8134), .Z(n8166) );
  NOR U8572 ( .A(n8137), .B(n8136), .Z(n8141) );
  NOR U8573 ( .A(n8139), .B(n8138), .Z(n8140) );
  NOR U8574 ( .A(n8141), .B(n8140), .Z(n8162) );
  NOR U8575 ( .A(n8143), .B(n8142), .Z(n8147) );
  NOR U8576 ( .A(n8145), .B(n8144), .Z(n8146) );
  NOR U8577 ( .A(n8147), .B(n8146), .Z(n8148) );
  IV U8578 ( .A(n8148), .Z(n8163) );
  XOR U8579 ( .A(n8162), .B(n8163), .Z(n8165) );
  XOR U8580 ( .A(n8166), .B(n8165), .Z(n8183) );
  XOR U8581 ( .A(n8150), .B(n8149), .Z(n8182) );
  NOR U8582 ( .A(n8183), .B(n8182), .Z(n8151) );
  NOR U8583 ( .A(n8152), .B(n8151), .Z(n8170) );
  IV U8584 ( .A(n8170), .Z(n8156) );
  XOR U8585 ( .A(n8154), .B(n8153), .Z(n8155) );
  IV U8586 ( .A(n8155), .Z(n8169) );
  NOR U8587 ( .A(n8156), .B(n8169), .Z(n8157) );
  NOR U8588 ( .A(n8158), .B(n8157), .Z(n8161) );
  IV U8589 ( .A(n8161), .Z(n8159) );
  NOR U8590 ( .A(n8160), .B(n8159), .Z(n8220) );
  XOR U8591 ( .A(n8161), .B(n8160), .Z(n8349) );
  IV U8592 ( .A(n8162), .Z(n8164) );
  NOR U8593 ( .A(n8164), .B(n8163), .Z(n8168) );
  NOR U8594 ( .A(n8166), .B(n8165), .Z(n8167) );
  NOR U8595 ( .A(n8168), .B(n8167), .Z(n8214) );
  XOR U8596 ( .A(n8170), .B(n8169), .Z(n8213) );
  NOR U8597 ( .A(n8214), .B(n8213), .Z(n8217) );
  XOR U8598 ( .A(n8172), .B(n8171), .Z(n8175) );
  XOR U8599 ( .A(n8174), .B(n8173), .Z(n8176) );
  NOR U8600 ( .A(n8175), .B(n8176), .Z(n8181) );
  XOR U8601 ( .A(n8176), .B(n8175), .Z(n8193) );
  IV U8602 ( .A(n8193), .Z(n8179) );
  XOR U8603 ( .A(n8178), .B(n8177), .Z(n8194) );
  NOR U8604 ( .A(n8179), .B(n8194), .Z(n8180) );
  NOR U8605 ( .A(n8181), .B(n8180), .Z(n8208) );
  XOR U8606 ( .A(n8183), .B(n8182), .Z(n8209) );
  NOR U8607 ( .A(n8208), .B(n8209), .Z(n8212) );
  XOR U8608 ( .A(n8184), .B(sum[18]), .Z(n8188) );
  NOR U8609 ( .A(n9316), .B(n9113), .Z(n8189) );
  IV U8610 ( .A(n8189), .Z(n8185) );
  NOR U8611 ( .A(n8188), .B(n8185), .Z(n8192) );
  IV U8612 ( .A(sum[17]), .Z(n8187) );
  NOR U8613 ( .A(n9593), .B(n8499), .Z(n8186) );
  IV U8614 ( .A(n8186), .Z(n8420) );
  NOR U8615 ( .A(n8187), .B(n8420), .Z(n8305) );
  IV U8616 ( .A(n8305), .Z(n8190) );
  XOR U8617 ( .A(n8189), .B(n8188), .Z(n8304) );
  NOR U8618 ( .A(n8190), .B(n8304), .Z(n8191) );
  NOR U8619 ( .A(n8192), .B(n8191), .Z(n8204) );
  XOR U8620 ( .A(n8194), .B(n8193), .Z(n8203) );
  NOR U8621 ( .A(n8204), .B(n8203), .Z(n8207) );
  NOR U8622 ( .A(n8948), .B(n9388), .Z(n8379) );
  IV U8623 ( .A(n8379), .Z(n8382) );
  NOR U8624 ( .A(n8195), .B(n8382), .Z(n8202) );
  XOR U8625 ( .A(n8197), .B(n8196), .Z(n8258) );
  NOR U8626 ( .A(n8727), .B(n9526), .Z(n8256) );
  NOR U8627 ( .A(n9260), .B(n9080), .Z(n8255) );
  XOR U8628 ( .A(n8256), .B(n8255), .Z(n8198) );
  IV U8629 ( .A(n8198), .Z(n8257) );
  XOR U8630 ( .A(n8258), .B(n8257), .Z(n8307) );
  NOR U8631 ( .A(n8862), .B(n9388), .Z(n8859) );
  NOR U8632 ( .A(n8948), .B(n9336), .Z(n8199) );
  XOR U8633 ( .A(n8859), .B(n8199), .Z(n8306) );
  IV U8634 ( .A(n8306), .Z(n8200) );
  NOR U8635 ( .A(n8307), .B(n8200), .Z(n8201) );
  NOR U8636 ( .A(n8202), .B(n8201), .Z(n8328) );
  XOR U8637 ( .A(n8204), .B(n8203), .Z(n8327) );
  IV U8638 ( .A(n8327), .Z(n8205) );
  NOR U8639 ( .A(n8328), .B(n8205), .Z(n8206) );
  NOR U8640 ( .A(n8207), .B(n8206), .Z(n8276) );
  IV U8641 ( .A(n8208), .Z(n8210) );
  XOR U8642 ( .A(n8210), .B(n8209), .Z(n8275) );
  NOR U8643 ( .A(n8276), .B(n8275), .Z(n8211) );
  NOR U8644 ( .A(n8212), .B(n8211), .Z(n8223) );
  XOR U8645 ( .A(n8214), .B(n8213), .Z(n8222) );
  IV U8646 ( .A(n8222), .Z(n8215) );
  NOR U8647 ( .A(n8223), .B(n8215), .Z(n8216) );
  NOR U8648 ( .A(n8217), .B(n8216), .Z(n8350) );
  IV U8649 ( .A(n8350), .Z(n8218) );
  NOR U8650 ( .A(n8349), .B(n8218), .Z(n8219) );
  NOR U8651 ( .A(n8220), .B(n8219), .Z(n9699) );
  IV U8652 ( .A(n9699), .Z(n8221) );
  NOR U8653 ( .A(n9698), .B(n8221), .Z(n9701) );
  XOR U8654 ( .A(n8223), .B(n8222), .Z(n8344) );
  XOR U8655 ( .A(n8225), .B(n8224), .Z(n8244) );
  NOR U8656 ( .A(n9592), .B(n9301), .Z(n9364) );
  IV U8657 ( .A(n9364), .Z(n8579) );
  NOR U8658 ( .A(n8226), .B(n8579), .Z(n8233) );
  NOR U8659 ( .A(n8290), .B(n9599), .Z(n8227) );
  IV U8660 ( .A(n8227), .Z(n8237) );
  NOR U8661 ( .A(n8228), .B(n9592), .Z(n8230) );
  NOR U8662 ( .A(n9034), .B(n9301), .Z(n8229) );
  XOR U8663 ( .A(n8230), .B(n8229), .Z(n8231) );
  IV U8664 ( .A(n8231), .Z(n8236) );
  NOR U8665 ( .A(n8237), .B(n8236), .Z(n8232) );
  NOR U8666 ( .A(n8233), .B(n8232), .Z(n8243) );
  IV U8667 ( .A(n8243), .Z(n8234) );
  NOR U8668 ( .A(n8244), .B(n8234), .Z(n8246) );
  NOR U8669 ( .A(n9429), .B(n8754), .Z(n8238) );
  NOR U8670 ( .A(n9600), .B(n8235), .Z(n8239) );
  NOR U8671 ( .A(n8238), .B(n8239), .Z(n8242) );
  XOR U8672 ( .A(n8237), .B(n8236), .Z(n8287) );
  IV U8673 ( .A(n8238), .Z(n8240) );
  XOR U8674 ( .A(n8240), .B(n8239), .Z(n8286) );
  NOR U8675 ( .A(n8287), .B(n8286), .Z(n8241) );
  NOR U8676 ( .A(n8242), .B(n8241), .Z(n8326) );
  XOR U8677 ( .A(n8244), .B(n8243), .Z(n8325) );
  NOR U8678 ( .A(n8326), .B(n8325), .Z(n8245) );
  NOR U8679 ( .A(n8246), .B(n8245), .Z(n8278) );
  NOR U8680 ( .A(n9414), .B(n9584), .Z(n9390) );
  IV U8681 ( .A(n9390), .Z(n8247) );
  NOR U8682 ( .A(n8248), .B(n8247), .Z(n8254) );
  NOR U8683 ( .A(n8499), .B(n9571), .Z(n8249) );
  IV U8684 ( .A(n8249), .Z(n8264) );
  NOR U8685 ( .A(n8656), .B(n9414), .Z(n8251) );
  NOR U8686 ( .A(n8501), .B(n9584), .Z(n8250) );
  XOR U8687 ( .A(n8251), .B(n8250), .Z(n8252) );
  IV U8688 ( .A(n8252), .Z(n8263) );
  NOR U8689 ( .A(n8264), .B(n8263), .Z(n8253) );
  NOR U8690 ( .A(n8254), .B(n8253), .Z(n8271) );
  NOR U8691 ( .A(n8256), .B(n8255), .Z(n8260) );
  NOR U8692 ( .A(n8258), .B(n8257), .Z(n8259) );
  NOR U8693 ( .A(n8260), .B(n8259), .Z(n8270) );
  IV U8694 ( .A(n8270), .Z(n8261) );
  NOR U8695 ( .A(n8271), .B(n8261), .Z(n8273) );
  NOR U8696 ( .A(n9115), .B(n9202), .Z(n8266) );
  NOR U8697 ( .A(n8262), .B(n8266), .Z(n8268) );
  XOR U8698 ( .A(n8264), .B(n8263), .Z(n8285) );
  XOR U8699 ( .A(n8266), .B(n8265), .Z(n8284) );
  NOR U8700 ( .A(n8285), .B(n8284), .Z(n8267) );
  NOR U8701 ( .A(n8268), .B(n8267), .Z(n8269) );
  IV U8702 ( .A(n8269), .Z(n8283) );
  XOR U8703 ( .A(n8271), .B(n8270), .Z(n8282) );
  NOR U8704 ( .A(n8283), .B(n8282), .Z(n8272) );
  NOR U8705 ( .A(n8273), .B(n8272), .Z(n8277) );
  IV U8706 ( .A(n8277), .Z(n8274) );
  NOR U8707 ( .A(n8278), .B(n8274), .Z(n8280) );
  XOR U8708 ( .A(n8276), .B(n8275), .Z(n8338) );
  XOR U8709 ( .A(n8278), .B(n8277), .Z(n8337) );
  NOR U8710 ( .A(n8338), .B(n8337), .Z(n8279) );
  NOR U8711 ( .A(n8280), .B(n8279), .Z(n8345) );
  IV U8712 ( .A(n8345), .Z(n8281) );
  NOR U8713 ( .A(n8344), .B(n8281), .Z(n8348) );
  XOR U8714 ( .A(n8283), .B(n8282), .Z(n8303) );
  XOR U8715 ( .A(n8285), .B(n8284), .Z(n8297) );
  XOR U8716 ( .A(n8287), .B(n8286), .Z(n8296) );
  NOR U8717 ( .A(n8297), .B(n8296), .Z(n8300) );
  NOR U8718 ( .A(n8288), .B(n8579), .Z(n8295) );
  NOR U8719 ( .A(n8501), .B(n9599), .Z(n8289) );
  IV U8720 ( .A(n8289), .Z(n8364) );
  NOR U8721 ( .A(n9115), .B(n9301), .Z(n8292) );
  NOR U8722 ( .A(n8290), .B(n9592), .Z(n8291) );
  XOR U8723 ( .A(n8292), .B(n8291), .Z(n8293) );
  IV U8724 ( .A(n8293), .Z(n8363) );
  NOR U8725 ( .A(n8364), .B(n8363), .Z(n8294) );
  NOR U8726 ( .A(n8295), .B(n8294), .Z(n8372) );
  XOR U8727 ( .A(n8297), .B(n8296), .Z(n8371) );
  IV U8728 ( .A(n8371), .Z(n8298) );
  NOR U8729 ( .A(n8372), .B(n8298), .Z(n8299) );
  NOR U8730 ( .A(n8300), .B(n8299), .Z(n8302) );
  IV U8731 ( .A(n8302), .Z(n8301) );
  NOR U8732 ( .A(n8303), .B(n8301), .Z(n8324) );
  XOR U8733 ( .A(n8303), .B(n8302), .Z(n8330) );
  XOR U8734 ( .A(n8305), .B(n8304), .Z(n8317) );
  XOR U8735 ( .A(n8307), .B(n8306), .Z(n8318) );
  NOR U8736 ( .A(n8317), .B(n8318), .Z(n8321) );
  NOR U8737 ( .A(n8656), .B(n9600), .Z(n8308) );
  IV U8738 ( .A(n8308), .Z(n8886) );
  NOR U8739 ( .A(n8309), .B(n8886), .Z(n8316) );
  NOR U8740 ( .A(n8727), .B(n9493), .Z(n8310) );
  IV U8741 ( .A(n8310), .Z(n8388) );
  NOR U8742 ( .A(n8656), .B(n9472), .Z(n8313) );
  NOR U8743 ( .A(n8311), .B(n9600), .Z(n8312) );
  XOR U8744 ( .A(n8313), .B(n8312), .Z(n8314) );
  IV U8745 ( .A(n8314), .Z(n8387) );
  NOR U8746 ( .A(n8388), .B(n8387), .Z(n8315) );
  NOR U8747 ( .A(n8316), .B(n8315), .Z(n8419) );
  XOR U8748 ( .A(n8318), .B(n8317), .Z(n8319) );
  IV U8749 ( .A(n8319), .Z(n8418) );
  NOR U8750 ( .A(n8419), .B(n8418), .Z(n8320) );
  NOR U8751 ( .A(n8321), .B(n8320), .Z(n8322) );
  IV U8752 ( .A(n8322), .Z(n8329) );
  NOR U8753 ( .A(n8330), .B(n8329), .Z(n8323) );
  NOR U8754 ( .A(n8324), .B(n8323), .Z(n8339) );
  XOR U8755 ( .A(n8326), .B(n8325), .Z(n8332) );
  XOR U8756 ( .A(n8328), .B(n8327), .Z(n8331) );
  NOR U8757 ( .A(n8332), .B(n8331), .Z(n8335) );
  XOR U8758 ( .A(n8330), .B(n8329), .Z(n8378) );
  XOR U8759 ( .A(n8332), .B(n8331), .Z(n8377) );
  IV U8760 ( .A(n8377), .Z(n8333) );
  NOR U8761 ( .A(n8378), .B(n8333), .Z(n8334) );
  NOR U8762 ( .A(n8335), .B(n8334), .Z(n8340) );
  IV U8763 ( .A(n8340), .Z(n8336) );
  NOR U8764 ( .A(n8339), .B(n8336), .Z(n8343) );
  XOR U8765 ( .A(n8338), .B(n8337), .Z(n8355) );
  IV U8766 ( .A(n8355), .Z(n8341) );
  XOR U8767 ( .A(n8340), .B(n8339), .Z(n8354) );
  NOR U8768 ( .A(n8341), .B(n8354), .Z(n8342) );
  NOR U8769 ( .A(n8343), .B(n8342), .Z(n8353) );
  IV U8770 ( .A(n8353), .Z(n8346) );
  XOR U8771 ( .A(n8345), .B(n8344), .Z(n8352) );
  NOR U8772 ( .A(n8346), .B(n8352), .Z(n8347) );
  NOR U8773 ( .A(n8348), .B(n8347), .Z(n9693) );
  IV U8774 ( .A(n9693), .Z(n8351) );
  XOR U8775 ( .A(n8350), .B(n8349), .Z(n9692) );
  NOR U8776 ( .A(n8351), .B(n9692), .Z(n9696) );
  XOR U8777 ( .A(n8353), .B(n8352), .Z(n9688) );
  XOR U8778 ( .A(n8355), .B(n8354), .Z(n8414) );
  IV U8779 ( .A(n8356), .Z(n8358) );
  NOR U8780 ( .A(n9241), .B(n9414), .Z(n8733) );
  IV U8781 ( .A(n8733), .Z(n8357) );
  NOR U8782 ( .A(n8358), .B(n8357), .Z(n8362) );
  NOR U8783 ( .A(n9260), .B(n9113), .Z(n8359) );
  IV U8784 ( .A(n8359), .Z(n8381) );
  NOR U8785 ( .A(n9414), .B(n8754), .Z(n8946) );
  NOR U8786 ( .A(n9241), .B(n9202), .Z(n8925) );
  XOR U8787 ( .A(n8946), .B(n8925), .Z(n8360) );
  IV U8788 ( .A(n8360), .Z(n8380) );
  NOR U8789 ( .A(n8381), .B(n8380), .Z(n8361) );
  NOR U8790 ( .A(n8362), .B(n8361), .Z(n8373) );
  NOR U8791 ( .A(n9034), .B(n9429), .Z(n8366) );
  NOR U8792 ( .A(n8582), .B(n9584), .Z(n8365) );
  NOR U8793 ( .A(n8366), .B(n8365), .Z(n8369) );
  XOR U8794 ( .A(n8364), .B(n8363), .Z(n8441) );
  XOR U8795 ( .A(n8366), .B(n8365), .Z(n8440) );
  IV U8796 ( .A(n8440), .Z(n8367) );
  NOR U8797 ( .A(n8441), .B(n8367), .Z(n8368) );
  NOR U8798 ( .A(n8369), .B(n8368), .Z(n8374) );
  IV U8799 ( .A(n8374), .Z(n8370) );
  NOR U8800 ( .A(n8373), .B(n8370), .Z(n8376) );
  XOR U8801 ( .A(n8372), .B(n8371), .Z(n8432) );
  XOR U8802 ( .A(n8374), .B(n8373), .Z(n8431) );
  NOR U8803 ( .A(n8432), .B(n8431), .Z(n8375) );
  NOR U8804 ( .A(n8376), .B(n8375), .Z(n8409) );
  XOR U8805 ( .A(n8378), .B(n8377), .Z(n8408) );
  NOR U8806 ( .A(n8409), .B(n8408), .Z(n8412) );
  NOR U8807 ( .A(n9080), .B(n9336), .Z(n8383) );
  NOR U8808 ( .A(n8379), .B(n8383), .Z(n8385) );
  XOR U8809 ( .A(n8381), .B(n8380), .Z(n8396) );
  XOR U8810 ( .A(n8383), .B(n8382), .Z(n8395) );
  NOR U8811 ( .A(n8396), .B(n8395), .Z(n8384) );
  NOR U8812 ( .A(n8385), .B(n8384), .Z(n8386) );
  IV U8813 ( .A(n8386), .Z(n8405) );
  NOR U8814 ( .A(n9490), .B(n8729), .Z(n8389) );
  NOR U8815 ( .A(n8422), .B(n9571), .Z(n8390) );
  NOR U8816 ( .A(n8389), .B(n8390), .Z(n8393) );
  XOR U8817 ( .A(n8388), .B(n8387), .Z(n8399) );
  IV U8818 ( .A(n8389), .Z(n8391) );
  XOR U8819 ( .A(n8391), .B(n8390), .Z(n8398) );
  NOR U8820 ( .A(n8399), .B(n8398), .Z(n8392) );
  NOR U8821 ( .A(n8393), .B(n8392), .Z(n8404) );
  IV U8822 ( .A(n8404), .Z(n8394) );
  NOR U8823 ( .A(n8405), .B(n8394), .Z(n8407) );
  XOR U8824 ( .A(n8396), .B(n8395), .Z(n8401) );
  NOR U8825 ( .A(n8862), .B(n9526), .Z(n8400) );
  IV U8826 ( .A(n8400), .Z(n8397) );
  NOR U8827 ( .A(n8401), .B(n8397), .Z(n8403) );
  XOR U8828 ( .A(n8399), .B(n8398), .Z(n8536) );
  XOR U8829 ( .A(n8401), .B(n8400), .Z(n8537) );
  NOR U8830 ( .A(n8536), .B(n8537), .Z(n8402) );
  NOR U8831 ( .A(n8403), .B(n8402), .Z(n8439) );
  XOR U8832 ( .A(n8405), .B(n8404), .Z(n8438) );
  NOR U8833 ( .A(n8439), .B(n8438), .Z(n8406) );
  NOR U8834 ( .A(n8407), .B(n8406), .Z(n8417) );
  XOR U8835 ( .A(n8409), .B(n8408), .Z(n8416) );
  IV U8836 ( .A(n8416), .Z(n8410) );
  NOR U8837 ( .A(n8417), .B(n8410), .Z(n8411) );
  NOR U8838 ( .A(n8412), .B(n8411), .Z(n8415) );
  IV U8839 ( .A(n8415), .Z(n8413) );
  NOR U8840 ( .A(n8414), .B(n8413), .Z(n8492) );
  XOR U8841 ( .A(n8415), .B(n8414), .Z(n8605) );
  XOR U8842 ( .A(n8417), .B(n8416), .Z(n8485) );
  XOR U8843 ( .A(n8419), .B(n8418), .Z(n8434) );
  XOR U8844 ( .A(n8420), .B(sum[17]), .Z(n8425) );
  NOR U8845 ( .A(n9316), .B(n9237), .Z(n8426) );
  IV U8846 ( .A(n8426), .Z(n8421) );
  NOR U8847 ( .A(n8425), .B(n8421), .Z(n8429) );
  IV U8848 ( .A(sum[16]), .Z(n8424) );
  NOR U8849 ( .A(n8422), .B(n9593), .Z(n8423) );
  IV U8850 ( .A(n8423), .Z(n8469) );
  NOR U8851 ( .A(n8424), .B(n8469), .Z(n8443) );
  IV U8852 ( .A(n8443), .Z(n8427) );
  XOR U8853 ( .A(n8426), .B(n8425), .Z(n8442) );
  NOR U8854 ( .A(n8427), .B(n8442), .Z(n8428) );
  NOR U8855 ( .A(n8429), .B(n8428), .Z(n8433) );
  IV U8856 ( .A(n8433), .Z(n8430) );
  NOR U8857 ( .A(n8434), .B(n8430), .Z(n8436) );
  XOR U8858 ( .A(n8432), .B(n8431), .Z(n8497) );
  XOR U8859 ( .A(n8434), .B(n8433), .Z(n8496) );
  NOR U8860 ( .A(n8497), .B(n8496), .Z(n8435) );
  NOR U8861 ( .A(n8436), .B(n8435), .Z(n8486) );
  IV U8862 ( .A(n8486), .Z(n8437) );
  NOR U8863 ( .A(n8485), .B(n8437), .Z(n8489) );
  XOR U8864 ( .A(n8439), .B(n8438), .Z(n8482) );
  XOR U8865 ( .A(n8441), .B(n8440), .Z(n8453) );
  IV U8866 ( .A(n8453), .Z(n8444) );
  XOR U8867 ( .A(n8443), .B(n8442), .Z(n8452) );
  NOR U8868 ( .A(n8444), .B(n8452), .Z(n8455) );
  NOR U8869 ( .A(n9429), .B(n9599), .Z(n9389) );
  IV U8870 ( .A(n9389), .Z(n8829) );
  NOR U8871 ( .A(n8445), .B(n8829), .Z(n8451) );
  NOR U8872 ( .A(n8727), .B(n9584), .Z(n8446) );
  IV U8873 ( .A(n8446), .Z(n8513) );
  NOR U8874 ( .A(n8582), .B(n9599), .Z(n8448) );
  NOR U8875 ( .A(n9429), .B(n9115), .Z(n8447) );
  XOR U8876 ( .A(n8448), .B(n8447), .Z(n8449) );
  IV U8877 ( .A(n8449), .Z(n8512) );
  NOR U8878 ( .A(n8513), .B(n8512), .Z(n8450) );
  NOR U8879 ( .A(n8451), .B(n8450), .Z(n8458) );
  XOR U8880 ( .A(n8453), .B(n8452), .Z(n8457) );
  NOR U8881 ( .A(n8458), .B(n8457), .Z(n8454) );
  NOR U8882 ( .A(n8455), .B(n8454), .Z(n8481) );
  IV U8883 ( .A(n8481), .Z(n8456) );
  NOR U8884 ( .A(n8482), .B(n8456), .Z(n8484) );
  XOR U8885 ( .A(n8458), .B(n8457), .Z(n8468) );
  NOR U8886 ( .A(n9490), .B(n9526), .Z(n9363) );
  IV U8887 ( .A(n9363), .Z(n8926) );
  NOR U8888 ( .A(n8459), .B(n8926), .Z(n8465) );
  NOR U8889 ( .A(n9034), .B(n9414), .Z(n8460) );
  IV U8890 ( .A(n8460), .Z(n9033) );
  NOR U8891 ( .A(n8656), .B(n9490), .Z(n8462) );
  NOR U8892 ( .A(n8948), .B(n9526), .Z(n8461) );
  XOR U8893 ( .A(n8462), .B(n8461), .Z(n8463) );
  IV U8894 ( .A(n8463), .Z(n8506) );
  NOR U8895 ( .A(n9033), .B(n8506), .Z(n8464) );
  NOR U8896 ( .A(n8465), .B(n8464), .Z(n8467) );
  IV U8897 ( .A(n8467), .Z(n8466) );
  NOR U8898 ( .A(n8468), .B(n8466), .Z(n8480) );
  XOR U8899 ( .A(n8468), .B(n8467), .Z(n8570) );
  XOR U8900 ( .A(n8469), .B(sum[16]), .Z(n8473) );
  NOR U8901 ( .A(n9260), .B(n9237), .Z(n8474) );
  IV U8902 ( .A(n8474), .Z(n8470) );
  NOR U8903 ( .A(n8473), .B(n8470), .Z(n8477) );
  IV U8904 ( .A(sum[15]), .Z(n8472) );
  NOR U8905 ( .A(n9593), .B(n8729), .Z(n8471) );
  IV U8906 ( .A(n8471), .Z(n8654) );
  NOR U8907 ( .A(n8472), .B(n8654), .Z(n8557) );
  IV U8908 ( .A(n8557), .Z(n8475) );
  XOR U8909 ( .A(n8474), .B(n8473), .Z(n8556) );
  NOR U8910 ( .A(n8475), .B(n8556), .Z(n8476) );
  NOR U8911 ( .A(n8477), .B(n8476), .Z(n8571) );
  IV U8912 ( .A(n8571), .Z(n8478) );
  NOR U8913 ( .A(n8570), .B(n8478), .Z(n8479) );
  NOR U8914 ( .A(n8480), .B(n8479), .Z(n8550) );
  XOR U8915 ( .A(n8482), .B(n8481), .Z(n8549) );
  NOR U8916 ( .A(n8550), .B(n8549), .Z(n8483) );
  NOR U8917 ( .A(n8484), .B(n8483), .Z(n8495) );
  IV U8918 ( .A(n8495), .Z(n8487) );
  XOR U8919 ( .A(n8486), .B(n8485), .Z(n8494) );
  NOR U8920 ( .A(n8487), .B(n8494), .Z(n8488) );
  NOR U8921 ( .A(n8489), .B(n8488), .Z(n8606) );
  IV U8922 ( .A(n8606), .Z(n8490) );
  NOR U8923 ( .A(n8605), .B(n8490), .Z(n8491) );
  NOR U8924 ( .A(n8492), .B(n8491), .Z(n9689) );
  IV U8925 ( .A(n9689), .Z(n8493) );
  NOR U8926 ( .A(n9688), .B(n8493), .Z(n9691) );
  XOR U8927 ( .A(n8495), .B(n8494), .Z(n8601) );
  XOR U8928 ( .A(n8497), .B(n8496), .Z(n8526) );
  IV U8929 ( .A(n8526), .Z(n8525) );
  NOR U8930 ( .A(n8498), .B(n8861), .Z(n8505) );
  NOR U8931 ( .A(n8499), .B(n9600), .Z(n8530) );
  IV U8932 ( .A(n8530), .Z(n8503) );
  NOR U8933 ( .A(n9316), .B(n9202), .Z(n8500) );
  IV U8934 ( .A(n8500), .Z(n9123) );
  NOR U8935 ( .A(n8501), .B(n9592), .Z(n8502) );
  XOR U8936 ( .A(n9123), .B(n8502), .Z(n8529) );
  NOR U8937 ( .A(n8503), .B(n8529), .Z(n8504) );
  NOR U8938 ( .A(n8505), .B(n8504), .Z(n8520) );
  NOR U8939 ( .A(n9336), .B(n9113), .Z(n8507) );
  NOR U8940 ( .A(n9080), .B(n9388), .Z(n8508) );
  NOR U8941 ( .A(n8507), .B(n8508), .Z(n8510) );
  XOR U8942 ( .A(n9033), .B(n8506), .Z(n8555) );
  IV U8943 ( .A(n8507), .Z(n8968) );
  XOR U8944 ( .A(n8508), .B(n8968), .Z(n8554) );
  NOR U8945 ( .A(n8555), .B(n8554), .Z(n8509) );
  NOR U8946 ( .A(n8510), .B(n8509), .Z(n8519) );
  IV U8947 ( .A(n8519), .Z(n8511) );
  NOR U8948 ( .A(n8520), .B(n8511), .Z(n8523) );
  NOR U8949 ( .A(n9472), .B(n8754), .Z(n8514) );
  NOR U8950 ( .A(n8862), .B(n9493), .Z(n8515) );
  NOR U8951 ( .A(n8514), .B(n8515), .Z(n8518) );
  XOR U8952 ( .A(n8513), .B(n8512), .Z(n8576) );
  IV U8953 ( .A(n8514), .Z(n8516) );
  XOR U8954 ( .A(n8516), .B(n8515), .Z(n8575) );
  NOR U8955 ( .A(n8576), .B(n8575), .Z(n8517) );
  NOR U8956 ( .A(n8518), .B(n8517), .Z(n8542) );
  IV U8957 ( .A(n8542), .Z(n8521) );
  XOR U8958 ( .A(n8520), .B(n8519), .Z(n8541) );
  NOR U8959 ( .A(n8521), .B(n8541), .Z(n8522) );
  NOR U8960 ( .A(n8523), .B(n8522), .Z(n8524) );
  IV U8961 ( .A(n8524), .Z(n8527) );
  NOR U8962 ( .A(n8525), .B(n8527), .Z(n8547) );
  XOR U8963 ( .A(n8527), .B(n8526), .Z(n8552) );
  NOR U8964 ( .A(n9241), .B(n9571), .Z(n8528) );
  IV U8965 ( .A(n8528), .Z(n9076) );
  NOR U8966 ( .A(n8770), .B(n9076), .Z(n8535) );
  XOR U8967 ( .A(n8530), .B(n8529), .Z(n8577) );
  NOR U8968 ( .A(n9571), .B(n8729), .Z(n8532) );
  NOR U8969 ( .A(n9241), .B(n9301), .Z(n8531) );
  XOR U8970 ( .A(n8532), .B(n8531), .Z(n8578) );
  IV U8971 ( .A(n8578), .Z(n8533) );
  NOR U8972 ( .A(n8577), .B(n8533), .Z(n8534) );
  NOR U8973 ( .A(n8535), .B(n8534), .Z(n8540) );
  XOR U8974 ( .A(n8537), .B(n8536), .Z(n8539) );
  IV U8975 ( .A(n8539), .Z(n8538) );
  NOR U8976 ( .A(n8540), .B(n8538), .Z(n8544) );
  XOR U8977 ( .A(n8540), .B(n8539), .Z(n8638) );
  XOR U8978 ( .A(n8542), .B(n8541), .Z(n8637) );
  NOR U8979 ( .A(n8638), .B(n8637), .Z(n8543) );
  NOR U8980 ( .A(n8544), .B(n8543), .Z(n8551) );
  IV U8981 ( .A(n8551), .Z(n8545) );
  NOR U8982 ( .A(n8552), .B(n8545), .Z(n8546) );
  NOR U8983 ( .A(n8547), .B(n8546), .Z(n8602) );
  IV U8984 ( .A(n8602), .Z(n8548) );
  NOR U8985 ( .A(n8601), .B(n8548), .Z(n8604) );
  XOR U8986 ( .A(n8550), .B(n8549), .Z(n8597) );
  XOR U8987 ( .A(n8552), .B(n8551), .Z(n8598) );
  IV U8988 ( .A(n8598), .Z(n8553) );
  NOR U8989 ( .A(n8597), .B(n8553), .Z(n8600) );
  XOR U8990 ( .A(n8555), .B(n8554), .Z(n8566) );
  XOR U8991 ( .A(n8557), .B(n8556), .Z(n8565) );
  NOR U8992 ( .A(n8566), .B(n8565), .Z(n8569) );
  NOR U8993 ( .A(n9472), .B(n9526), .Z(n9340) );
  IV U8994 ( .A(n9340), .Z(n9525) );
  NOR U8995 ( .A(n8558), .B(n9525), .Z(n8564) );
  NOR U8996 ( .A(n9388), .B(n9113), .Z(n8623) );
  IV U8997 ( .A(n8623), .Z(n8562) );
  NOR U8998 ( .A(n9080), .B(n9526), .Z(n8559) );
  IV U8999 ( .A(n8559), .Z(n8561) );
  NOR U9000 ( .A(n9034), .B(n9472), .Z(n8560) );
  XOR U9001 ( .A(n8561), .B(n8560), .Z(n8622) );
  NOR U9002 ( .A(n8562), .B(n8622), .Z(n8563) );
  NOR U9003 ( .A(n8564), .B(n8563), .Z(n8653) );
  XOR U9004 ( .A(n8566), .B(n8565), .Z(n8567) );
  IV U9005 ( .A(n8567), .Z(n8652) );
  NOR U9006 ( .A(n8653), .B(n8652), .Z(n8568) );
  NOR U9007 ( .A(n8569), .B(n8568), .Z(n8574) );
  IV U9008 ( .A(n8574), .Z(n8572) );
  XOR U9009 ( .A(n8571), .B(n8570), .Z(n8573) );
  NOR U9010 ( .A(n8572), .B(n8573), .Z(n8595) );
  XOR U9011 ( .A(n8574), .B(n8573), .Z(n8641) );
  XOR U9012 ( .A(n8576), .B(n8575), .Z(n8589) );
  XOR U9013 ( .A(n8578), .B(n8577), .Z(n8588) );
  NOR U9014 ( .A(n8589), .B(n8588), .Z(n8592) );
  NOR U9015 ( .A(n8580), .B(n8579), .Z(n8587) );
  NOR U9016 ( .A(n8727), .B(n9599), .Z(n8581) );
  IV U9017 ( .A(n8581), .Z(n8673) );
  NOR U9018 ( .A(n8582), .B(n9592), .Z(n8584) );
  NOR U9019 ( .A(n9316), .B(n9301), .Z(n8583) );
  XOR U9020 ( .A(n8584), .B(n8583), .Z(n8585) );
  IV U9021 ( .A(n8585), .Z(n8672) );
  NOR U9022 ( .A(n8673), .B(n8672), .Z(n8586) );
  NOR U9023 ( .A(n8587), .B(n8586), .Z(n8621) );
  XOR U9024 ( .A(n8589), .B(n8588), .Z(n8620) );
  IV U9025 ( .A(n8620), .Z(n8590) );
  NOR U9026 ( .A(n8621), .B(n8590), .Z(n8591) );
  NOR U9027 ( .A(n8592), .B(n8591), .Z(n8640) );
  IV U9028 ( .A(n8640), .Z(n8593) );
  NOR U9029 ( .A(n8641), .B(n8593), .Z(n8594) );
  NOR U9030 ( .A(n8595), .B(n8594), .Z(n8596) );
  IV U9031 ( .A(n8596), .Z(n8614) );
  XOR U9032 ( .A(n8598), .B(n8597), .Z(n8613) );
  NOR U9033 ( .A(n8614), .B(n8613), .Z(n8599) );
  NOR U9034 ( .A(n8600), .B(n8599), .Z(n8610) );
  XOR U9035 ( .A(n8602), .B(n8601), .Z(n8611) );
  NOR U9036 ( .A(n8610), .B(n8611), .Z(n8603) );
  NOR U9037 ( .A(n8604), .B(n8603), .Z(n8609) );
  IV U9038 ( .A(n8609), .Z(n8607) );
  XOR U9039 ( .A(n8606), .B(n8605), .Z(n8608) );
  NOR U9040 ( .A(n8607), .B(n8608), .Z(n9686) );
  XOR U9041 ( .A(n8609), .B(n8608), .Z(n9804) );
  XOR U9042 ( .A(n8611), .B(n8610), .Z(n8612) );
  IV U9043 ( .A(n8612), .Z(n9680) );
  XOR U9044 ( .A(n8614), .B(n8613), .Z(n8649) );
  NOR U9045 ( .A(n9490), .B(n9493), .Z(n9442) );
  IV U9046 ( .A(n9442), .Z(n9438) );
  NOR U9047 ( .A(n8615), .B(n9438), .Z(n8619) );
  NOR U9048 ( .A(n9490), .B(n8754), .Z(n8616) );
  NOR U9049 ( .A(n8948), .B(n9493), .Z(n8762) );
  XOR U9050 ( .A(n8616), .B(n8762), .Z(n8617) );
  IV U9051 ( .A(n8617), .Z(n8625) );
  NOR U9052 ( .A(n8626), .B(n8625), .Z(n8618) );
  NOR U9053 ( .A(n8619), .B(n8618), .Z(n8632) );
  XOR U9054 ( .A(n8621), .B(n8620), .Z(n8633) );
  NOR U9055 ( .A(n8632), .B(n8633), .Z(n8636) );
  XOR U9056 ( .A(n8623), .B(n8622), .Z(n8628) );
  NOR U9057 ( .A(n9237), .B(n9336), .Z(n8629) );
  IV U9058 ( .A(n8629), .Z(n8624) );
  NOR U9059 ( .A(n8628), .B(n8624), .Z(n8631) );
  XOR U9060 ( .A(n8626), .B(n8625), .Z(n8682) );
  XOR U9061 ( .A(n8627), .B(n8679), .Z(n8681) );
  XOR U9062 ( .A(n8682), .B(n8681), .Z(n8708) );
  XOR U9063 ( .A(n8629), .B(n8628), .Z(n8709) );
  NOR U9064 ( .A(n8708), .B(n8709), .Z(n8630) );
  NOR U9065 ( .A(n8631), .B(n8630), .Z(n8666) );
  IV U9066 ( .A(n8632), .Z(n8634) );
  XOR U9067 ( .A(n8634), .B(n8633), .Z(n8665) );
  NOR U9068 ( .A(n8666), .B(n8665), .Z(n8635) );
  NOR U9069 ( .A(n8636), .B(n8635), .Z(n8643) );
  XOR U9070 ( .A(n8638), .B(n8637), .Z(n8642) );
  IV U9071 ( .A(n8642), .Z(n8639) );
  NOR U9072 ( .A(n8643), .B(n8639), .Z(n8646) );
  XOR U9073 ( .A(n8641), .B(n8640), .Z(n8651) );
  IV U9074 ( .A(n8651), .Z(n8644) );
  XOR U9075 ( .A(n8643), .B(n8642), .Z(n8650) );
  NOR U9076 ( .A(n8644), .B(n8650), .Z(n8645) );
  NOR U9077 ( .A(n8646), .B(n8645), .Z(n8648) );
  IV U9078 ( .A(n8648), .Z(n8647) );
  NOR U9079 ( .A(n8649), .B(n8647), .Z(n8699) );
  XOR U9080 ( .A(n8649), .B(n8648), .Z(n8814) );
  XOR U9081 ( .A(n8651), .B(n8650), .Z(n8693) );
  XOR U9082 ( .A(n8653), .B(n8652), .Z(n8668) );
  XOR U9083 ( .A(n8654), .B(sum[15]), .Z(n8659) );
  NOR U9084 ( .A(n9260), .B(n9202), .Z(n8660) );
  IV U9085 ( .A(n8660), .Z(n8655) );
  NOR U9086 ( .A(n8659), .B(n8655), .Z(n8663) );
  IV U9087 ( .A(sum[14]), .Z(n8658) );
  NOR U9088 ( .A(n9593), .B(n8656), .Z(n8657) );
  IV U9089 ( .A(n8657), .Z(n8753) );
  NOR U9090 ( .A(n8658), .B(n8753), .Z(n8776) );
  IV U9091 ( .A(n8776), .Z(n8661) );
  XOR U9092 ( .A(n8660), .B(n8659), .Z(n8775) );
  NOR U9093 ( .A(n8661), .B(n8775), .Z(n8662) );
  NOR U9094 ( .A(n8663), .B(n8662), .Z(n8667) );
  IV U9095 ( .A(n8667), .Z(n8664) );
  NOR U9096 ( .A(n8668), .B(n8664), .Z(n8670) );
  XOR U9097 ( .A(n8666), .B(n8665), .Z(n8687) );
  XOR U9098 ( .A(n8668), .B(n8667), .Z(n8688) );
  NOR U9099 ( .A(n8687), .B(n8688), .Z(n8669) );
  NOR U9100 ( .A(n8670), .B(n8669), .Z(n8694) );
  IV U9101 ( .A(n8694), .Z(n8671) );
  NOR U9102 ( .A(n8693), .B(n8671), .Z(n8696) );
  NOR U9103 ( .A(n9115), .B(n9414), .Z(n8674) );
  NOR U9104 ( .A(n8862), .B(n9584), .Z(n8675) );
  NOR U9105 ( .A(n8674), .B(n8675), .Z(n8678) );
  XOR U9106 ( .A(n8673), .B(n8672), .Z(n8707) );
  IV U9107 ( .A(n8674), .Z(n8676) );
  XOR U9108 ( .A(n8676), .B(n8675), .Z(n8706) );
  NOR U9109 ( .A(n8707), .B(n8706), .Z(n8677) );
  NOR U9110 ( .A(n8678), .B(n8677), .Z(n8690) );
  IV U9111 ( .A(n8690), .Z(n8686) );
  NOR U9112 ( .A(n8680), .B(n8679), .Z(n8684) );
  NOR U9113 ( .A(n8682), .B(n8681), .Z(n8683) );
  NOR U9114 ( .A(n8684), .B(n8683), .Z(n8685) );
  IV U9115 ( .A(n8685), .Z(n8689) );
  NOR U9116 ( .A(n8686), .B(n8689), .Z(n8692) );
  XOR U9117 ( .A(n8688), .B(n8687), .Z(n8704) );
  XOR U9118 ( .A(n8690), .B(n8689), .Z(n8705) );
  NOR U9119 ( .A(n8704), .B(n8705), .Z(n8691) );
  NOR U9120 ( .A(n8692), .B(n8691), .Z(n8701) );
  XOR U9121 ( .A(n8694), .B(n8693), .Z(n8702) );
  NOR U9122 ( .A(n8701), .B(n8702), .Z(n8695) );
  NOR U9123 ( .A(n8696), .B(n8695), .Z(n8815) );
  IV U9124 ( .A(n8815), .Z(n8697) );
  NOR U9125 ( .A(n8814), .B(n8697), .Z(n8698) );
  NOR U9126 ( .A(n8699), .B(n8698), .Z(n9681) );
  IV U9127 ( .A(n9681), .Z(n8700) );
  NOR U9128 ( .A(n9680), .B(n8700), .Z(n9683) );
  XOR U9129 ( .A(n8702), .B(n8701), .Z(n8703) );
  IV U9130 ( .A(n8703), .Z(n8809) );
  XOR U9131 ( .A(n8705), .B(n8704), .Z(n8749) );
  XOR U9132 ( .A(n8707), .B(n8706), .Z(n8720) );
  XOR U9133 ( .A(n8709), .B(n8708), .Z(n8719) );
  IV U9134 ( .A(n8719), .Z(n8710) );
  NOR U9135 ( .A(n8720), .B(n8710), .Z(n8722) );
  NOR U9136 ( .A(n9490), .B(n9388), .Z(n9318) );
  IV U9137 ( .A(n9318), .Z(n8711) );
  NOR U9138 ( .A(n8712), .B(n8711), .Z(n8718) );
  NOR U9139 ( .A(n9115), .B(n9472), .Z(n8713) );
  IV U9140 ( .A(n8713), .Z(n9112) );
  NOR U9141 ( .A(n9034), .B(n9490), .Z(n8714) );
  XOR U9142 ( .A(n8715), .B(n8714), .Z(n8716) );
  IV U9143 ( .A(n8716), .Z(n8738) );
  NOR U9144 ( .A(n9112), .B(n8738), .Z(n8717) );
  NOR U9145 ( .A(n8718), .B(n8717), .Z(n8725) );
  XOR U9146 ( .A(n8720), .B(n8719), .Z(n8724) );
  NOR U9147 ( .A(n8725), .B(n8724), .Z(n8721) );
  NOR U9148 ( .A(n8722), .B(n8721), .Z(n8748) );
  IV U9149 ( .A(n8748), .Z(n8723) );
  NOR U9150 ( .A(n8749), .B(n8723), .Z(n8751) );
  XOR U9151 ( .A(n8725), .B(n8724), .Z(n8743) );
  NOR U9152 ( .A(n8726), .B(n8733), .Z(n8736) );
  NOR U9153 ( .A(n9592), .B(n8727), .Z(n8728) );
  IV U9154 ( .A(n8728), .Z(n8772) );
  NOR U9155 ( .A(n9600), .B(n8729), .Z(n8731) );
  NOR U9156 ( .A(n9260), .B(n9301), .Z(n8730) );
  XOR U9157 ( .A(n8731), .B(n8730), .Z(n8732) );
  IV U9158 ( .A(n8732), .Z(n8771) );
  XOR U9159 ( .A(n8772), .B(n8771), .Z(n8782) );
  XOR U9160 ( .A(n8734), .B(n8733), .Z(n8781) );
  NOR U9161 ( .A(n8782), .B(n8781), .Z(n8735) );
  NOR U9162 ( .A(n8736), .B(n8735), .Z(n8744) );
  NOR U9163 ( .A(n8743), .B(n8744), .Z(n8747) );
  NOR U9164 ( .A(n9526), .B(n9113), .Z(n8740) );
  NOR U9165 ( .A(n8737), .B(n8740), .Z(n8742) );
  XOR U9166 ( .A(n9112), .B(n8738), .Z(n8826) );
  XOR U9167 ( .A(n8740), .B(n8739), .Z(n8825) );
  NOR U9168 ( .A(n8826), .B(n8825), .Z(n8741) );
  NOR U9169 ( .A(n8742), .B(n8741), .Z(n8822) );
  XOR U9170 ( .A(n8744), .B(n8743), .Z(n8745) );
  IV U9171 ( .A(n8745), .Z(n8821) );
  NOR U9172 ( .A(n8822), .B(n8821), .Z(n8746) );
  NOR U9173 ( .A(n8747), .B(n8746), .Z(n8805) );
  XOR U9174 ( .A(n8749), .B(n8748), .Z(n8804) );
  NOR U9175 ( .A(n8805), .B(n8804), .Z(n8750) );
  NOR U9176 ( .A(n8751), .B(n8750), .Z(n8810) );
  IV U9177 ( .A(n8810), .Z(n8752) );
  NOR U9178 ( .A(n8809), .B(n8752), .Z(n8813) );
  NOR U9179 ( .A(n9336), .B(n9202), .Z(n8758) );
  IV U9180 ( .A(n8758), .Z(n9200) );
  XOR U9181 ( .A(n8753), .B(sum[14]), .Z(n8757) );
  NOR U9182 ( .A(n9200), .B(n8757), .Z(n8761) );
  IV U9183 ( .A(sum[13]), .Z(n8756) );
  NOR U9184 ( .A(n9593), .B(n8754), .Z(n8755) );
  IV U9185 ( .A(n8755), .Z(n8850) );
  NOR U9186 ( .A(n8756), .B(n8850), .Z(n8780) );
  IV U9187 ( .A(n8780), .Z(n8759) );
  XOR U9188 ( .A(n8758), .B(n8757), .Z(n8779) );
  NOR U9189 ( .A(n8759), .B(n8779), .Z(n8760) );
  NOR U9190 ( .A(n8761), .B(n8760), .Z(n8789) );
  IV U9191 ( .A(n8762), .Z(n8763) );
  NOR U9192 ( .A(n9080), .B(n9584), .Z(n8871) );
  IV U9193 ( .A(n8871), .Z(n8834) );
  NOR U9194 ( .A(n8763), .B(n8834), .Z(n8769) );
  NOR U9195 ( .A(n9316), .B(n9429), .Z(n8778) );
  IV U9196 ( .A(n8778), .Z(n8767) );
  NOR U9197 ( .A(n9080), .B(n9493), .Z(n8764) );
  IV U9198 ( .A(n8764), .Z(n8766) );
  NOR U9199 ( .A(n8948), .B(n9584), .Z(n8765) );
  XOR U9200 ( .A(n8766), .B(n8765), .Z(n8777) );
  NOR U9201 ( .A(n8767), .B(n8777), .Z(n8768) );
  NOR U9202 ( .A(n8769), .B(n8768), .Z(n8798) );
  NOR U9203 ( .A(n9260), .B(n9600), .Z(n9391) );
  IV U9204 ( .A(n9391), .Z(n9367) );
  NOR U9205 ( .A(n8770), .B(n9367), .Z(n8774) );
  NOR U9206 ( .A(n8772), .B(n8771), .Z(n8773) );
  NOR U9207 ( .A(n8774), .B(n8773), .Z(n8795) );
  XOR U9208 ( .A(n8776), .B(n8775), .Z(n8794) );
  XOR U9209 ( .A(n8795), .B(n8794), .Z(n8796) );
  XOR U9210 ( .A(n8798), .B(n8796), .Z(n8788) );
  NOR U9211 ( .A(n8789), .B(n8788), .Z(n8792) );
  XOR U9212 ( .A(n8778), .B(n8777), .Z(n8784) );
  XOR U9213 ( .A(n8780), .B(n8779), .Z(n8783) );
  NOR U9214 ( .A(n8784), .B(n8783), .Z(n8787) );
  XOR U9215 ( .A(n8782), .B(n8781), .Z(n8827) );
  XOR U9216 ( .A(n8784), .B(n8783), .Z(n8828) );
  IV U9217 ( .A(n8828), .Z(n8785) );
  NOR U9218 ( .A(n8827), .B(n8785), .Z(n8786) );
  NOR U9219 ( .A(n8787), .B(n8786), .Z(n8824) );
  XOR U9220 ( .A(n8789), .B(n8788), .Z(n8823) );
  IV U9221 ( .A(n8823), .Z(n8790) );
  NOR U9222 ( .A(n8824), .B(n8790), .Z(n8791) );
  NOR U9223 ( .A(n8792), .B(n8791), .Z(n8793) );
  IV U9224 ( .A(n8793), .Z(n8803) );
  NOR U9225 ( .A(n8795), .B(n8794), .Z(n8800) );
  IV U9226 ( .A(n8796), .Z(n8797) );
  NOR U9227 ( .A(n8798), .B(n8797), .Z(n8799) );
  NOR U9228 ( .A(n8800), .B(n8799), .Z(n8802) );
  IV U9229 ( .A(n8802), .Z(n8801) );
  NOR U9230 ( .A(n8803), .B(n8801), .Z(n8808) );
  XOR U9231 ( .A(n8803), .B(n8802), .Z(n8820) );
  XOR U9232 ( .A(n8805), .B(n8804), .Z(n8819) );
  IV U9233 ( .A(n8819), .Z(n8806) );
  NOR U9234 ( .A(n8820), .B(n8806), .Z(n8807) );
  NOR U9235 ( .A(n8808), .B(n8807), .Z(n8818) );
  IV U9236 ( .A(n8818), .Z(n8811) );
  XOR U9237 ( .A(n8810), .B(n8809), .Z(n8817) );
  NOR U9238 ( .A(n8811), .B(n8817), .Z(n8812) );
  NOR U9239 ( .A(n8813), .B(n8812), .Z(n9675) );
  IV U9240 ( .A(n9675), .Z(n8816) );
  XOR U9241 ( .A(n8815), .B(n8814), .Z(n9674) );
  NOR U9242 ( .A(n8816), .B(n9674), .Z(n9678) );
  XOR U9243 ( .A(n8818), .B(n8817), .Z(n8910) );
  XOR U9244 ( .A(n8820), .B(n8819), .Z(n8848) );
  XOR U9245 ( .A(n8822), .B(n8821), .Z(n8842) );
  XOR U9246 ( .A(n8824), .B(n8823), .Z(n8843) );
  NOR U9247 ( .A(n8842), .B(n8843), .Z(n8846) );
  XOR U9248 ( .A(n8826), .B(n8825), .Z(n8837) );
  XOR U9249 ( .A(n8828), .B(n8827), .Z(n8838) );
  NOR U9250 ( .A(n8837), .B(n8838), .Z(n8841) );
  NOR U9251 ( .A(n8830), .B(n8829), .Z(n8836) );
  NOR U9252 ( .A(n8948), .B(n9599), .Z(n8832) );
  NOR U9253 ( .A(n9260), .B(n9429), .Z(n8831) );
  XOR U9254 ( .A(n8832), .B(n8831), .Z(n8872) );
  IV U9255 ( .A(n8872), .Z(n8833) );
  NOR U9256 ( .A(n8834), .B(n8833), .Z(n8835) );
  NOR U9257 ( .A(n8836), .B(n8835), .Z(n8884) );
  IV U9258 ( .A(n8837), .Z(n8839) );
  XOR U9259 ( .A(n8839), .B(n8838), .Z(n8883) );
  NOR U9260 ( .A(n8884), .B(n8883), .Z(n8840) );
  NOR U9261 ( .A(n8841), .B(n8840), .Z(n8901) );
  XOR U9262 ( .A(n8843), .B(n8842), .Z(n8900) );
  IV U9263 ( .A(n8900), .Z(n8844) );
  NOR U9264 ( .A(n8901), .B(n8844), .Z(n8845) );
  NOR U9265 ( .A(n8846), .B(n8845), .Z(n8849) );
  IV U9266 ( .A(n8849), .Z(n8847) );
  NOR U9267 ( .A(n8848), .B(n8847), .Z(n8908) );
  XOR U9268 ( .A(n8849), .B(n8848), .Z(n9003) );
  XOR U9269 ( .A(n8850), .B(sum[13]), .Z(n8854) );
  NOR U9270 ( .A(n9336), .B(n9301), .Z(n8855) );
  IV U9271 ( .A(n8855), .Z(n8851) );
  NOR U9272 ( .A(n8854), .B(n8851), .Z(n8858) );
  IV U9273 ( .A(sum[12]), .Z(n8853) );
  NOR U9274 ( .A(n9034), .B(n9593), .Z(n8852) );
  IV U9275 ( .A(n8852), .Z(n9008) );
  NOR U9276 ( .A(n8853), .B(n9008), .Z(n8956) );
  IV U9277 ( .A(n8956), .Z(n8856) );
  XOR U9278 ( .A(n8855), .B(n8854), .Z(n8955) );
  NOR U9279 ( .A(n8856), .B(n8955), .Z(n8857) );
  NOR U9280 ( .A(n8858), .B(n8857), .Z(n8878) );
  IV U9281 ( .A(n8859), .Z(n8860) );
  NOR U9282 ( .A(n8861), .B(n8860), .Z(n8867) );
  NOR U9283 ( .A(n9202), .B(n9388), .Z(n8864) );
  NOR U9284 ( .A(n9592), .B(n8862), .Z(n8863) );
  XOR U9285 ( .A(n8864), .B(n8863), .Z(n8865) );
  IV U9286 ( .A(n8865), .Z(n8885) );
  NOR U9287 ( .A(n8886), .B(n8885), .Z(n8866) );
  NOR U9288 ( .A(n8867), .B(n8866), .Z(n8879) );
  NOR U9289 ( .A(n8878), .B(n8879), .Z(n8882) );
  IV U9290 ( .A(n8868), .Z(n8869) );
  NOR U9291 ( .A(n8869), .B(n8926), .Z(n8877) );
  NOR U9292 ( .A(n9493), .B(n9113), .Z(n8916) );
  NOR U9293 ( .A(n9241), .B(n9472), .Z(n8915) );
  XOR U9294 ( .A(n8916), .B(n8915), .Z(n8870) );
  IV U9295 ( .A(n8870), .Z(n8917) );
  XOR U9296 ( .A(n8872), .B(n8871), .Z(n8918) );
  XOR U9297 ( .A(n8917), .B(n8918), .Z(n8924) );
  NOR U9298 ( .A(n9115), .B(n9490), .Z(n8874) );
  NOR U9299 ( .A(n9237), .B(n9526), .Z(n8873) );
  XOR U9300 ( .A(n8874), .B(n8873), .Z(n8923) );
  IV U9301 ( .A(n8923), .Z(n8875) );
  NOR U9302 ( .A(n8924), .B(n8875), .Z(n8876) );
  NOR U9303 ( .A(n8877), .B(n8876), .Z(n8893) );
  IV U9304 ( .A(n8878), .Z(n8880) );
  XOR U9305 ( .A(n8880), .B(n8879), .Z(n8892) );
  NOR U9306 ( .A(n8893), .B(n8892), .Z(n8881) );
  NOR U9307 ( .A(n8882), .B(n8881), .Z(n8903) );
  XOR U9308 ( .A(n8884), .B(n8883), .Z(n8894) );
  NOR U9309 ( .A(n9316), .B(n9414), .Z(n8887) );
  NOR U9310 ( .A(n9034), .B(n9571), .Z(n8888) );
  NOR U9311 ( .A(n8887), .B(n8888), .Z(n8891) );
  XOR U9312 ( .A(n8886), .B(n8885), .Z(n8921) );
  IV U9313 ( .A(n8887), .Z(n8889) );
  XOR U9314 ( .A(n8889), .B(n8888), .Z(n8922) );
  NOR U9315 ( .A(n8921), .B(n8922), .Z(n8890) );
  NOR U9316 ( .A(n8891), .B(n8890), .Z(n8895) );
  NOR U9317 ( .A(n8894), .B(n8895), .Z(n8898) );
  XOR U9318 ( .A(n8893), .B(n8892), .Z(n8940) );
  XOR U9319 ( .A(n8895), .B(n8894), .Z(n8939) );
  IV U9320 ( .A(n8939), .Z(n8896) );
  NOR U9321 ( .A(n8940), .B(n8896), .Z(n8897) );
  NOR U9322 ( .A(n8898), .B(n8897), .Z(n8902) );
  IV U9323 ( .A(n8902), .Z(n8899) );
  NOR U9324 ( .A(n8903), .B(n8899), .Z(n8905) );
  XOR U9325 ( .A(n8901), .B(n8900), .Z(n8912) );
  XOR U9326 ( .A(n8903), .B(n8902), .Z(n8913) );
  NOR U9327 ( .A(n8912), .B(n8913), .Z(n8904) );
  NOR U9328 ( .A(n8905), .B(n8904), .Z(n9004) );
  IV U9329 ( .A(n9004), .Z(n8906) );
  NOR U9330 ( .A(n9003), .B(n8906), .Z(n8907) );
  NOR U9331 ( .A(n8908), .B(n8907), .Z(n8911) );
  IV U9332 ( .A(n8911), .Z(n8909) );
  NOR U9333 ( .A(n8910), .B(n8909), .Z(n9673) );
  XOR U9334 ( .A(n8911), .B(n8910), .Z(n9819) );
  IV U9335 ( .A(n8912), .Z(n8914) );
  XOR U9336 ( .A(n8914), .B(n8913), .Z(n8998) );
  NOR U9337 ( .A(n8916), .B(n8915), .Z(n8920) );
  NOR U9338 ( .A(n8918), .B(n8917), .Z(n8919) );
  NOR U9339 ( .A(n8920), .B(n8919), .Z(n8942) );
  XOR U9340 ( .A(n8922), .B(n8921), .Z(n8934) );
  XOR U9341 ( .A(n8924), .B(n8923), .Z(n8933) );
  NOR U9342 ( .A(n8934), .B(n8933), .Z(n8937) );
  IV U9343 ( .A(n8925), .Z(n8927) );
  NOR U9344 ( .A(n8927), .B(n8926), .Z(n8932) );
  NOR U9345 ( .A(n9526), .B(n9202), .Z(n9056) );
  NOR U9346 ( .A(n9241), .B(n9490), .Z(n8928) );
  XOR U9347 ( .A(n9056), .B(n8928), .Z(n8929) );
  IV U9348 ( .A(n8929), .Z(n8972) );
  NOR U9349 ( .A(n8930), .B(n8972), .Z(n8931) );
  NOR U9350 ( .A(n8932), .B(n8931), .Z(n8958) );
  XOR U9351 ( .A(n8934), .B(n8933), .Z(n8957) );
  IV U9352 ( .A(n8957), .Z(n8935) );
  NOR U9353 ( .A(n8958), .B(n8935), .Z(n8936) );
  NOR U9354 ( .A(n8937), .B(n8936), .Z(n8941) );
  IV U9355 ( .A(n8941), .Z(n8938) );
  NOR U9356 ( .A(n8942), .B(n8938), .Z(n8944) );
  XOR U9357 ( .A(n8940), .B(n8939), .Z(n8966) );
  XOR U9358 ( .A(n8942), .B(n8941), .Z(n8965) );
  NOR U9359 ( .A(n8966), .B(n8965), .Z(n8943) );
  NOR U9360 ( .A(n8944), .B(n8943), .Z(n8999) );
  IV U9361 ( .A(n8999), .Z(n8945) );
  NOR U9362 ( .A(n8998), .B(n8945), .Z(n9002) );
  IV U9363 ( .A(n8946), .Z(n8947) );
  NOR U9364 ( .A(n8947), .B(n9367), .Z(n8954) );
  NOR U9365 ( .A(n8948), .B(n9592), .Z(n8949) );
  IV U9366 ( .A(n8949), .Z(n8982) );
  NOR U9367 ( .A(n9260), .B(n9414), .Z(n8950) );
  XOR U9368 ( .A(n8951), .B(n8950), .Z(n8952) );
  IV U9369 ( .A(n8952), .Z(n8981) );
  NOR U9370 ( .A(n8982), .B(n8981), .Z(n8953) );
  NOR U9371 ( .A(n8954), .B(n8953), .Z(n8960) );
  XOR U9372 ( .A(n8956), .B(n8955), .Z(n8959) );
  NOR U9373 ( .A(n8960), .B(n8959), .Z(n8963) );
  XOR U9374 ( .A(n8958), .B(n8957), .Z(n8976) );
  XOR U9375 ( .A(n8960), .B(n8959), .Z(n8977) );
  IV U9376 ( .A(n8977), .Z(n8961) );
  NOR U9377 ( .A(n8976), .B(n8961), .Z(n8962) );
  NOR U9378 ( .A(n8963), .B(n8962), .Z(n8964) );
  IV U9379 ( .A(n8964), .Z(n8994) );
  XOR U9380 ( .A(n8966), .B(n8965), .Z(n8993) );
  IV U9381 ( .A(n8993), .Z(n8967) );
  NOR U9382 ( .A(n8994), .B(n8967), .Z(n8997) );
  NOR U9383 ( .A(n9429), .B(n9584), .Z(n9300) );
  IV U9384 ( .A(n9300), .Z(n9460) );
  NOR U9385 ( .A(n8968), .B(n9460), .Z(n8975) );
  NOR U9386 ( .A(n9113), .B(n9584), .Z(n8970) );
  NOR U9387 ( .A(n9429), .B(n9336), .Z(n8969) );
  XOR U9388 ( .A(n8970), .B(n8969), .Z(n8979) );
  IV U9389 ( .A(n8979), .Z(n8973) );
  XOR U9390 ( .A(n8972), .B(n8971), .Z(n8978) );
  NOR U9391 ( .A(n8973), .B(n8978), .Z(n8974) );
  NOR U9392 ( .A(n8975), .B(n8974), .Z(n8989) );
  XOR U9393 ( .A(n8977), .B(n8976), .Z(n8988) );
  NOR U9394 ( .A(n8989), .B(n8988), .Z(n8992) );
  XOR U9395 ( .A(n8979), .B(n8978), .Z(n8984) );
  NOR U9396 ( .A(n8980), .B(n8984), .Z(n8987) );
  XOR U9397 ( .A(n8982), .B(n8981), .Z(n9020) );
  NOR U9398 ( .A(n9115), .B(n9571), .Z(n9018) );
  IV U9399 ( .A(n9018), .Z(n8983) );
  NOR U9400 ( .A(n9316), .B(n9472), .Z(n9017) );
  XOR U9401 ( .A(n8983), .B(n9017), .Z(n9019) );
  XOR U9402 ( .A(n9020), .B(n9019), .Z(n9052) );
  XOR U9403 ( .A(n8985), .B(n8984), .Z(n9053) );
  NOR U9404 ( .A(n9052), .B(n9053), .Z(n8986) );
  NOR U9405 ( .A(n8987), .B(n8986), .Z(n9027) );
  XOR U9406 ( .A(n8989), .B(n8988), .Z(n9026) );
  IV U9407 ( .A(n9026), .Z(n8990) );
  NOR U9408 ( .A(n9027), .B(n8990), .Z(n8991) );
  NOR U9409 ( .A(n8992), .B(n8991), .Z(n9031) );
  IV U9410 ( .A(n9031), .Z(n8995) );
  XOR U9411 ( .A(n8994), .B(n8993), .Z(n9030) );
  NOR U9412 ( .A(n8995), .B(n9030), .Z(n8996) );
  NOR U9413 ( .A(n8997), .B(n8996), .Z(n9007) );
  IV U9414 ( .A(n9007), .Z(n9000) );
  XOR U9415 ( .A(n8999), .B(n8998), .Z(n9006) );
  NOR U9416 ( .A(n9000), .B(n9006), .Z(n9001) );
  NOR U9417 ( .A(n9002), .B(n9001), .Z(n9667) );
  IV U9418 ( .A(n9667), .Z(n9005) );
  XOR U9419 ( .A(n9004), .B(n9003), .Z(n9666) );
  NOR U9420 ( .A(n9005), .B(n9666), .Z(n9670) );
  XOR U9421 ( .A(n9007), .B(n9006), .Z(n9662) );
  NOR U9422 ( .A(n9301), .B(n9388), .Z(n9013) );
  IV U9423 ( .A(n9013), .Z(n9009) );
  XOR U9424 ( .A(n9008), .B(sum[12]), .Z(n9012) );
  NOR U9425 ( .A(n9009), .B(n9012), .Z(n9016) );
  IV U9426 ( .A(sum[11]), .Z(n9011) );
  NOR U9427 ( .A(n9115), .B(n9593), .Z(n9010) );
  IV U9428 ( .A(n9010), .Z(n9040) );
  NOR U9429 ( .A(n9011), .B(n9040), .Z(n9055) );
  IV U9430 ( .A(n9055), .Z(n9014) );
  XOR U9431 ( .A(n9013), .B(n9012), .Z(n9054) );
  NOR U9432 ( .A(n9014), .B(n9054), .Z(n9015) );
  NOR U9433 ( .A(n9016), .B(n9015), .Z(n9024) );
  NOR U9434 ( .A(n9018), .B(n9017), .Z(n9022) );
  NOR U9435 ( .A(n9020), .B(n9019), .Z(n9021) );
  NOR U9436 ( .A(n9022), .B(n9021), .Z(n9025) );
  IV U9437 ( .A(n9025), .Z(n9023) );
  NOR U9438 ( .A(n9024), .B(n9023), .Z(n9029) );
  XOR U9439 ( .A(n9025), .B(n9024), .Z(n9109) );
  XOR U9440 ( .A(n9027), .B(n9026), .Z(n9110) );
  NOR U9441 ( .A(n9109), .B(n9110), .Z(n9028) );
  NOR U9442 ( .A(n9029), .B(n9028), .Z(n9100) );
  IV U9443 ( .A(n9100), .Z(n9032) );
  XOR U9444 ( .A(n9031), .B(n9030), .Z(n9099) );
  NOR U9445 ( .A(n9032), .B(n9099), .Z(n9102) );
  NOR U9446 ( .A(n9600), .B(n9336), .Z(n9428) );
  IV U9447 ( .A(n9428), .Z(n9433) );
  NOR U9448 ( .A(n9033), .B(n9433), .Z(n9039) );
  NOR U9449 ( .A(n9414), .B(n9336), .Z(n9036) );
  NOR U9450 ( .A(n9034), .B(n9600), .Z(n9035) );
  XOR U9451 ( .A(n9036), .B(n9035), .Z(n9037) );
  IV U9452 ( .A(n9037), .Z(n9075) );
  NOR U9453 ( .A(n9076), .B(n9075), .Z(n9038) );
  NOR U9454 ( .A(n9039), .B(n9038), .Z(n9050) );
  XOR U9455 ( .A(n9040), .B(sum[11]), .Z(n9044) );
  NOR U9456 ( .A(n9041), .B(n9044), .Z(n9048) );
  IV U9457 ( .A(sum[10]), .Z(n9043) );
  NOR U9458 ( .A(n9241), .B(n9593), .Z(n9042) );
  IV U9459 ( .A(n9042), .Z(n9165) );
  NOR U9460 ( .A(n9043), .B(n9165), .Z(n9131) );
  IV U9461 ( .A(n9131), .Z(n9046) );
  XOR U9462 ( .A(n9045), .B(n9044), .Z(n9130) );
  NOR U9463 ( .A(n9046), .B(n9130), .Z(n9047) );
  NOR U9464 ( .A(n9048), .B(n9047), .Z(n9049) );
  NOR U9465 ( .A(n9050), .B(n9049), .Z(n9064) );
  XOR U9466 ( .A(n9050), .B(n9049), .Z(n9051) );
  IV U9467 ( .A(n9051), .Z(n9089) );
  XOR U9468 ( .A(n9053), .B(n9052), .Z(n9066) );
  XOR U9469 ( .A(n9055), .B(n9054), .Z(n9067) );
  XOR U9470 ( .A(n9066), .B(n9067), .Z(n9069) );
  IV U9471 ( .A(n9069), .Z(n9062) );
  IV U9472 ( .A(n9056), .Z(n9057) );
  NOR U9473 ( .A(n9493), .B(n9301), .Z(n9181) );
  IV U9474 ( .A(n9181), .Z(n9176) );
  NOR U9475 ( .A(n9057), .B(n9176), .Z(n9061) );
  NOR U9476 ( .A(n9493), .B(n9202), .Z(n9329) );
  XOR U9477 ( .A(n9058), .B(n9329), .Z(n9059) );
  IV U9478 ( .A(n9059), .Z(n9081) );
  NOR U9479 ( .A(n9082), .B(n9081), .Z(n9060) );
  NOR U9480 ( .A(n9061), .B(n9060), .Z(n9070) );
  XOR U9481 ( .A(n9062), .B(n9070), .Z(n9088) );
  NOR U9482 ( .A(n9089), .B(n9088), .Z(n9063) );
  NOR U9483 ( .A(n9064), .B(n9063), .Z(n9065) );
  IV U9484 ( .A(n9065), .Z(n9096) );
  IV U9485 ( .A(n9066), .Z(n9068) );
  NOR U9486 ( .A(n9068), .B(n9067), .Z(n9072) );
  NOR U9487 ( .A(n9070), .B(n9069), .Z(n9071) );
  NOR U9488 ( .A(n9072), .B(n9071), .Z(n9095) );
  IV U9489 ( .A(n9095), .Z(n9073) );
  NOR U9490 ( .A(n9096), .B(n9073), .Z(n9098) );
  NOR U9491 ( .A(n9260), .B(n9472), .Z(n9077) );
  NOR U9492 ( .A(n9074), .B(n9077), .Z(n9079) );
  XOR U9493 ( .A(n9076), .B(n9075), .Z(n9122) );
  XOR U9494 ( .A(n9077), .B(n9313), .Z(n9121) );
  NOR U9495 ( .A(n9122), .B(n9121), .Z(n9078) );
  NOR U9496 ( .A(n9079), .B(n9078), .Z(n9091) );
  NOR U9497 ( .A(n9599), .B(n9113), .Z(n9084) );
  NOR U9498 ( .A(n9080), .B(n9592), .Z(n9083) );
  NOR U9499 ( .A(n9084), .B(n9083), .Z(n9087) );
  XOR U9500 ( .A(n9082), .B(n9081), .Z(n9133) );
  XOR U9501 ( .A(n9084), .B(n9083), .Z(n9085) );
  IV U9502 ( .A(n9085), .Z(n9132) );
  NOR U9503 ( .A(n9133), .B(n9132), .Z(n9086) );
  NOR U9504 ( .A(n9087), .B(n9086), .Z(n9090) );
  NOR U9505 ( .A(n9091), .B(n9090), .Z(n9094) );
  XOR U9506 ( .A(n9089), .B(n9088), .Z(n9150) );
  XOR U9507 ( .A(n9091), .B(n9090), .Z(n9151) );
  IV U9508 ( .A(n9151), .Z(n9092) );
  NOR U9509 ( .A(n9150), .B(n9092), .Z(n9093) );
  NOR U9510 ( .A(n9094), .B(n9093), .Z(n9108) );
  XOR U9511 ( .A(n9096), .B(n9095), .Z(n9107) );
  NOR U9512 ( .A(n9108), .B(n9107), .Z(n9097) );
  NOR U9513 ( .A(n9098), .B(n9097), .Z(n9104) );
  XOR U9514 ( .A(n9100), .B(n9099), .Z(n9105) );
  NOR U9515 ( .A(n9104), .B(n9105), .Z(n9101) );
  NOR U9516 ( .A(n9102), .B(n9101), .Z(n9663) );
  IV U9517 ( .A(n9663), .Z(n9103) );
  NOR U9518 ( .A(n9662), .B(n9103), .Z(n9665) );
  IV U9519 ( .A(n9104), .Z(n9106) );
  XOR U9520 ( .A(n9106), .B(n9105), .Z(n9656) );
  XOR U9521 ( .A(n9108), .B(n9107), .Z(n9155) );
  XOR U9522 ( .A(n9110), .B(n9109), .Z(n9154) );
  IV U9523 ( .A(n9154), .Z(n9111) );
  NOR U9524 ( .A(n9155), .B(n9111), .Z(n9158) );
  NOR U9525 ( .A(n9112), .B(n9433), .Z(n9120) );
  NOR U9526 ( .A(n9592), .B(n9113), .Z(n9114) );
  IV U9527 ( .A(n9114), .Z(n9178) );
  NOR U9528 ( .A(n9336), .B(n9472), .Z(n9117) );
  NOR U9529 ( .A(n9115), .B(n9600), .Z(n9116) );
  XOR U9530 ( .A(n9117), .B(n9116), .Z(n9118) );
  IV U9531 ( .A(n9118), .Z(n9177) );
  NOR U9532 ( .A(n9178), .B(n9177), .Z(n9119) );
  NOR U9533 ( .A(n9120), .B(n9119), .Z(n9135) );
  XOR U9534 ( .A(n9122), .B(n9121), .Z(n9134) );
  NOR U9535 ( .A(n9135), .B(n9134), .Z(n9138) );
  NOR U9536 ( .A(n9571), .B(n9584), .Z(n9539) );
  IV U9537 ( .A(n9539), .Z(n9535) );
  NOR U9538 ( .A(n9123), .B(n9535), .Z(n9129) );
  NOR U9539 ( .A(n9429), .B(n9526), .Z(n9175) );
  IV U9540 ( .A(n9175), .Z(n9127) );
  NOR U9541 ( .A(n9202), .B(n9584), .Z(n9124) );
  IV U9542 ( .A(n9124), .Z(n9126) );
  NOR U9543 ( .A(n9316), .B(n9571), .Z(n9125) );
  XOR U9544 ( .A(n9126), .B(n9125), .Z(n9174) );
  NOR U9545 ( .A(n9127), .B(n9174), .Z(n9128) );
  NOR U9546 ( .A(n9129), .B(n9128), .Z(n9144) );
  XOR U9547 ( .A(n9131), .B(n9130), .Z(n9140) );
  XOR U9548 ( .A(n9133), .B(n9132), .Z(n9141) );
  XOR U9549 ( .A(n9140), .B(n9141), .Z(n9142) );
  XOR U9550 ( .A(n9144), .B(n9142), .Z(n9187) );
  XOR U9551 ( .A(n9135), .B(n9134), .Z(n9186) );
  IV U9552 ( .A(n9186), .Z(n9136) );
  NOR U9553 ( .A(n9187), .B(n9136), .Z(n9137) );
  NOR U9554 ( .A(n9138), .B(n9137), .Z(n9139) );
  IV U9555 ( .A(n9139), .Z(n9149) );
  NOR U9556 ( .A(n9141), .B(n9140), .Z(n9146) );
  IV U9557 ( .A(n9142), .Z(n9143) );
  NOR U9558 ( .A(n9144), .B(n9143), .Z(n9145) );
  NOR U9559 ( .A(n9146), .B(n9145), .Z(n9148) );
  IV U9560 ( .A(n9148), .Z(n9147) );
  NOR U9561 ( .A(n9149), .B(n9147), .Z(n9153) );
  XOR U9562 ( .A(n9149), .B(n9148), .Z(n9163) );
  XOR U9563 ( .A(n9151), .B(n9150), .Z(n9162) );
  NOR U9564 ( .A(n9163), .B(n9162), .Z(n9152) );
  NOR U9565 ( .A(n9153), .B(n9152), .Z(n9161) );
  IV U9566 ( .A(n9161), .Z(n9156) );
  XOR U9567 ( .A(n9155), .B(n9154), .Z(n9160) );
  NOR U9568 ( .A(n9156), .B(n9160), .Z(n9157) );
  NOR U9569 ( .A(n9158), .B(n9157), .Z(n9657) );
  IV U9570 ( .A(n9657), .Z(n9159) );
  NOR U9571 ( .A(n9656), .B(n9159), .Z(n9660) );
  XOR U9572 ( .A(n9161), .B(n9160), .Z(n9229) );
  XOR U9573 ( .A(n9163), .B(n9162), .Z(n9164) );
  IV U9574 ( .A(n9164), .Z(n9192) );
  NOR U9575 ( .A(n9414), .B(n9388), .Z(n9170) );
  IV U9576 ( .A(n9170), .Z(n9166) );
  XOR U9577 ( .A(n9165), .B(sum[10]), .Z(n9169) );
  NOR U9578 ( .A(n9166), .B(n9169), .Z(n9173) );
  IV U9579 ( .A(sum[9]), .Z(n9168) );
  NOR U9580 ( .A(n9316), .B(n9593), .Z(n9167) );
  IV U9581 ( .A(n9167), .Z(n9258) );
  NOR U9582 ( .A(n9168), .B(n9258), .Z(n9195) );
  IV U9583 ( .A(n9195), .Z(n9171) );
  XOR U9584 ( .A(n9170), .B(n9169), .Z(n9194) );
  NOR U9585 ( .A(n9171), .B(n9194), .Z(n9172) );
  NOR U9586 ( .A(n9173), .B(n9172), .Z(n9185) );
  XOR U9587 ( .A(n9175), .B(n9174), .Z(n9180) );
  NOR U9588 ( .A(n9176), .B(n9180), .Z(n9183) );
  XOR U9589 ( .A(n9178), .B(n9177), .Z(n9215) );
  NOR U9590 ( .A(n9237), .B(n9599), .Z(n9213) );
  NOR U9591 ( .A(n9260), .B(n9490), .Z(n9212) );
  XOR U9592 ( .A(n9213), .B(n9212), .Z(n9179) );
  IV U9593 ( .A(n9179), .Z(n9214) );
  XOR U9594 ( .A(n9215), .B(n9214), .Z(n9196) );
  XOR U9595 ( .A(n9181), .B(n9180), .Z(n9197) );
  NOR U9596 ( .A(n9196), .B(n9197), .Z(n9182) );
  NOR U9597 ( .A(n9183), .B(n9182), .Z(n9184) );
  NOR U9598 ( .A(n9185), .B(n9184), .Z(n9190) );
  XOR U9599 ( .A(n9185), .B(n9184), .Z(n9222) );
  IV U9600 ( .A(n9222), .Z(n9188) );
  XOR U9601 ( .A(n9187), .B(n9186), .Z(n9221) );
  NOR U9602 ( .A(n9188), .B(n9221), .Z(n9189) );
  NOR U9603 ( .A(n9190), .B(n9189), .Z(n9193) );
  IV U9604 ( .A(n9193), .Z(n9191) );
  NOR U9605 ( .A(n9192), .B(n9191), .Z(n9227) );
  XOR U9606 ( .A(n9193), .B(n9192), .Z(n9290) );
  XOR U9607 ( .A(n9195), .B(n9194), .Z(n9208) );
  XOR U9608 ( .A(n9197), .B(n9196), .Z(n9209) );
  IV U9609 ( .A(n9209), .Z(n9198) );
  NOR U9610 ( .A(n9208), .B(n9198), .Z(n9211) );
  NOR U9611 ( .A(n9599), .B(n9490), .Z(n9199) );
  IV U9612 ( .A(n9199), .Z(n9553) );
  NOR U9613 ( .A(n9200), .B(n9553), .Z(n9207) );
  NOR U9614 ( .A(n9301), .B(n9584), .Z(n9271) );
  IV U9615 ( .A(n9271), .Z(n9205) );
  NOR U9616 ( .A(n9490), .B(n9336), .Z(n9201) );
  IV U9617 ( .A(n9201), .Z(n9204) );
  NOR U9618 ( .A(n9599), .B(n9202), .Z(n9203) );
  XOR U9619 ( .A(n9204), .B(n9203), .Z(n9270) );
  NOR U9620 ( .A(n9205), .B(n9270), .Z(n9206) );
  NOR U9621 ( .A(n9207), .B(n9206), .Z(n9235) );
  XOR U9622 ( .A(n9209), .B(n9208), .Z(n9234) );
  NOR U9623 ( .A(n9235), .B(n9234), .Z(n9210) );
  NOR U9624 ( .A(n9211), .B(n9210), .Z(n9220) );
  NOR U9625 ( .A(n9213), .B(n9212), .Z(n9217) );
  NOR U9626 ( .A(n9215), .B(n9214), .Z(n9216) );
  NOR U9627 ( .A(n9217), .B(n9216), .Z(n9219) );
  IV U9628 ( .A(n9219), .Z(n9218) );
  NOR U9629 ( .A(n9220), .B(n9218), .Z(n9224) );
  XOR U9630 ( .A(n9220), .B(n9219), .Z(n9231) );
  XOR U9631 ( .A(n9222), .B(n9221), .Z(n9232) );
  NOR U9632 ( .A(n9231), .B(n9232), .Z(n9223) );
  NOR U9633 ( .A(n9224), .B(n9223), .Z(n9291) );
  IV U9634 ( .A(n9291), .Z(n9225) );
  NOR U9635 ( .A(n9290), .B(n9225), .Z(n9226) );
  NOR U9636 ( .A(n9227), .B(n9226), .Z(n9230) );
  IV U9637 ( .A(n9230), .Z(n9228) );
  NOR U9638 ( .A(n9229), .B(n9228), .Z(n9655) );
  XOR U9639 ( .A(n9230), .B(n9229), .Z(n9839) );
  XOR U9640 ( .A(n9232), .B(n9231), .Z(n9233) );
  IV U9641 ( .A(n9233), .Z(n9286) );
  XOR U9642 ( .A(n9235), .B(n9234), .Z(n9254) );
  NOR U9643 ( .A(n9592), .B(n9472), .Z(n9528) );
  IV U9644 ( .A(n9528), .Z(n9459) );
  NOR U9645 ( .A(n9236), .B(n9459), .Z(n9244) );
  NOR U9646 ( .A(n9472), .B(n9388), .Z(n9239) );
  NOR U9647 ( .A(n9237), .B(n9592), .Z(n9238) );
  XOR U9648 ( .A(n9239), .B(n9238), .Z(n9240) );
  IV U9649 ( .A(n9240), .Z(n9247) );
  NOR U9650 ( .A(n9241), .B(n9600), .Z(n9242) );
  IV U9651 ( .A(n9242), .Z(n9246) );
  NOR U9652 ( .A(n9247), .B(n9246), .Z(n9243) );
  NOR U9653 ( .A(n9244), .B(n9243), .Z(n9253) );
  IV U9654 ( .A(n9253), .Z(n9245) );
  NOR U9655 ( .A(n9254), .B(n9245), .Z(n9256) );
  NOR U9656 ( .A(n9429), .B(n9493), .Z(n9248) );
  NOR U9657 ( .A(n9260), .B(n9571), .Z(n9249) );
  NOR U9658 ( .A(n9248), .B(n9249), .Z(n9252) );
  XOR U9659 ( .A(n9247), .B(n9246), .Z(n9273) );
  IV U9660 ( .A(n9248), .Z(n9250) );
  XOR U9661 ( .A(n9250), .B(n9249), .Z(n9272) );
  NOR U9662 ( .A(n9273), .B(n9272), .Z(n9251) );
  NOR U9663 ( .A(n9252), .B(n9251), .Z(n9280) );
  XOR U9664 ( .A(n9254), .B(n9253), .Z(n9279) );
  NOR U9665 ( .A(n9280), .B(n9279), .Z(n9255) );
  NOR U9666 ( .A(n9256), .B(n9255), .Z(n9287) );
  IV U9667 ( .A(n9287), .Z(n9257) );
  NOR U9668 ( .A(n9286), .B(n9257), .Z(n9289) );
  XOR U9669 ( .A(n9258), .B(sum[9]), .Z(n9263) );
  NOR U9670 ( .A(n9414), .B(n9526), .Z(n9264) );
  IV U9671 ( .A(n9264), .Z(n9259) );
  NOR U9672 ( .A(n9263), .B(n9259), .Z(n9267) );
  IV U9673 ( .A(sum[8]), .Z(n9262) );
  NOR U9674 ( .A(n9260), .B(n9593), .Z(n9261) );
  IV U9675 ( .A(n9261), .Z(n9335) );
  NOR U9676 ( .A(n9262), .B(n9335), .Z(n9269) );
  IV U9677 ( .A(n9269), .Z(n9265) );
  XOR U9678 ( .A(n9264), .B(n9263), .Z(n9268) );
  NOR U9679 ( .A(n9265), .B(n9268), .Z(n9266) );
  NOR U9680 ( .A(n9267), .B(n9266), .Z(n9282) );
  XOR U9681 ( .A(n9269), .B(n9268), .Z(n9274) );
  XOR U9682 ( .A(n9271), .B(n9270), .Z(n9275) );
  NOR U9683 ( .A(n9274), .B(n9275), .Z(n9278) );
  XOR U9684 ( .A(n9273), .B(n9272), .Z(n9310) );
  XOR U9685 ( .A(n9275), .B(n9274), .Z(n9309) );
  IV U9686 ( .A(n9309), .Z(n9276) );
  NOR U9687 ( .A(n9310), .B(n9276), .Z(n9277) );
  NOR U9688 ( .A(n9278), .B(n9277), .Z(n9281) );
  NOR U9689 ( .A(n9282), .B(n9281), .Z(n9285) );
  XOR U9690 ( .A(n9280), .B(n9279), .Z(n9298) );
  XOR U9691 ( .A(n9282), .B(n9281), .Z(n9283) );
  IV U9692 ( .A(n9283), .Z(n9299) );
  NOR U9693 ( .A(n9298), .B(n9299), .Z(n9284) );
  NOR U9694 ( .A(n9285), .B(n9284), .Z(n9295) );
  XOR U9695 ( .A(n9287), .B(n9286), .Z(n9296) );
  NOR U9696 ( .A(n9295), .B(n9296), .Z(n9288) );
  NOR U9697 ( .A(n9289), .B(n9288), .Z(n9294) );
  IV U9698 ( .A(n9294), .Z(n9292) );
  XOR U9699 ( .A(n9291), .B(n9290), .Z(n9293) );
  NOR U9700 ( .A(n9292), .B(n9293), .Z(n9652) );
  XOR U9701 ( .A(n9294), .B(n9293), .Z(n9844) );
  XOR U9702 ( .A(n9296), .B(n9295), .Z(n9297) );
  IV U9703 ( .A(n9297), .Z(n9356) );
  XOR U9704 ( .A(n9299), .B(n9298), .Z(n9328) );
  NOR U9705 ( .A(n9336), .B(n9571), .Z(n9306) );
  NOR U9706 ( .A(n9300), .B(n9306), .Z(n9308) );
  NOR U9707 ( .A(n9599), .B(n9301), .Z(n9302) );
  IV U9708 ( .A(n9302), .Z(n9332) );
  NOR U9709 ( .A(n9414), .B(n9493), .Z(n9304) );
  XOR U9710 ( .A(n9304), .B(n9303), .Z(n9305) );
  IV U9711 ( .A(n9305), .Z(n9331) );
  XOR U9712 ( .A(n9332), .B(n9331), .Z(n9315) );
  XOR U9713 ( .A(n9306), .B(n9460), .Z(n9314) );
  NOR U9714 ( .A(n9315), .B(n9314), .Z(n9307) );
  NOR U9715 ( .A(n9308), .B(n9307), .Z(n9323) );
  IV U9716 ( .A(n9323), .Z(n9311) );
  XOR U9717 ( .A(n9310), .B(n9309), .Z(n9322) );
  NOR U9718 ( .A(n9311), .B(n9322), .Z(n9325) );
  NOR U9719 ( .A(n9600), .B(n9388), .Z(n9474) );
  IV U9720 ( .A(n9474), .Z(n9312) );
  NOR U9721 ( .A(n9313), .B(n9312), .Z(n9321) );
  XOR U9722 ( .A(n9315), .B(n9314), .Z(n9359) );
  NOR U9723 ( .A(n9316), .B(n9600), .Z(n9317) );
  XOR U9724 ( .A(n9318), .B(n9317), .Z(n9358) );
  IV U9725 ( .A(n9358), .Z(n9319) );
  NOR U9726 ( .A(n9359), .B(n9319), .Z(n9320) );
  NOR U9727 ( .A(n9321), .B(n9320), .Z(n9347) );
  XOR U9728 ( .A(n9323), .B(n9322), .Z(n9346) );
  NOR U9729 ( .A(n9347), .B(n9346), .Z(n9324) );
  NOR U9730 ( .A(n9325), .B(n9324), .Z(n9327) );
  IV U9731 ( .A(n9327), .Z(n9326) );
  NOR U9732 ( .A(n9328), .B(n9326), .Z(n9354) );
  XOR U9733 ( .A(n9328), .B(n9327), .Z(n9409) );
  IV U9734 ( .A(n9329), .Z(n9330) );
  NOR U9735 ( .A(n9592), .B(n9414), .Z(n9503) );
  IV U9736 ( .A(n9503), .Z(n9507) );
  NOR U9737 ( .A(n9330), .B(n9507), .Z(n9334) );
  NOR U9738 ( .A(n9332), .B(n9331), .Z(n9333) );
  NOR U9739 ( .A(n9334), .B(n9333), .Z(n9345) );
  XOR U9740 ( .A(n9335), .B(sum[8]), .Z(n9339) );
  NOR U9741 ( .A(n9525), .B(n9339), .Z(n9343) );
  IV U9742 ( .A(sum[7]), .Z(n9338) );
  NOR U9743 ( .A(n9593), .B(n9336), .Z(n9337) );
  IV U9744 ( .A(n9337), .Z(n9377) );
  NOR U9745 ( .A(n9338), .B(n9377), .Z(n9361) );
  IV U9746 ( .A(n9361), .Z(n9341) );
  XOR U9747 ( .A(n9340), .B(n9339), .Z(n9360) );
  NOR U9748 ( .A(n9341), .B(n9360), .Z(n9342) );
  NOR U9749 ( .A(n9343), .B(n9342), .Z(n9344) );
  NOR U9750 ( .A(n9345), .B(n9344), .Z(n9351) );
  XOR U9751 ( .A(n9345), .B(n9344), .Z(n9376) );
  IV U9752 ( .A(n9376), .Z(n9349) );
  XOR U9753 ( .A(n9347), .B(n9346), .Z(n9348) );
  IV U9754 ( .A(n9348), .Z(n9375) );
  NOR U9755 ( .A(n9349), .B(n9375), .Z(n9350) );
  NOR U9756 ( .A(n9351), .B(n9350), .Z(n9410) );
  IV U9757 ( .A(n9410), .Z(n9352) );
  NOR U9758 ( .A(n9409), .B(n9352), .Z(n9353) );
  NOR U9759 ( .A(n9354), .B(n9353), .Z(n9357) );
  IV U9760 ( .A(n9357), .Z(n9355) );
  NOR U9761 ( .A(n9356), .B(n9355), .Z(n9649) );
  XOR U9762 ( .A(n9357), .B(n9356), .Z(n9849) );
  XOR U9763 ( .A(n9359), .B(n9358), .Z(n9371) );
  XOR U9764 ( .A(n9361), .B(n9360), .Z(n9370) );
  NOR U9765 ( .A(n9371), .B(n9370), .Z(n9374) );
  NOR U9766 ( .A(n9592), .B(n9490), .Z(n9561) );
  IV U9767 ( .A(n9561), .Z(n9556) );
  NOR U9768 ( .A(n9362), .B(n9556), .Z(n9369) );
  NOR U9769 ( .A(n9364), .B(n9363), .Z(n9365) );
  NOR U9770 ( .A(n9369), .B(n9365), .Z(n9366) );
  IV U9771 ( .A(n9366), .Z(n9392) );
  NOR U9772 ( .A(n9367), .B(n9392), .Z(n9368) );
  NOR U9773 ( .A(n9369), .B(n9368), .Z(n9387) );
  XOR U9774 ( .A(n9371), .B(n9370), .Z(n9386) );
  IV U9775 ( .A(n9386), .Z(n9372) );
  NOR U9776 ( .A(n9387), .B(n9372), .Z(n9373) );
  NOR U9777 ( .A(n9374), .B(n9373), .Z(n9405) );
  XOR U9778 ( .A(n9376), .B(n9375), .Z(n9404) );
  NOR U9779 ( .A(n9405), .B(n9404), .Z(n9408) );
  XOR U9780 ( .A(n9377), .B(sum[7]), .Z(n9381) );
  NOR U9781 ( .A(n9472), .B(n9493), .Z(n9382) );
  IV U9782 ( .A(n9382), .Z(n9378) );
  NOR U9783 ( .A(n9381), .B(n9378), .Z(n9385) );
  IV U9784 ( .A(sum[6]), .Z(n9380) );
  NOR U9785 ( .A(n9593), .B(n9388), .Z(n9379) );
  IV U9786 ( .A(n9379), .Z(n9437) );
  NOR U9787 ( .A(n9380), .B(n9437), .Z(n9394) );
  IV U9788 ( .A(n9394), .Z(n9383) );
  XOR U9789 ( .A(n9382), .B(n9381), .Z(n9393) );
  NOR U9790 ( .A(n9383), .B(n9393), .Z(n9384) );
  NOR U9791 ( .A(n9385), .B(n9384), .Z(n9400) );
  XOR U9792 ( .A(n9387), .B(n9386), .Z(n9399) );
  NOR U9793 ( .A(n9400), .B(n9399), .Z(n9403) );
  NOR U9794 ( .A(n9571), .B(n9388), .Z(n9396) );
  IV U9795 ( .A(n9396), .Z(n9471) );
  XOR U9796 ( .A(n9390), .B(n9389), .Z(n9416) );
  XOR U9797 ( .A(n9392), .B(n9391), .Z(n9417) );
  XOR U9798 ( .A(n9416), .B(n9417), .Z(n9395) );
  NOR U9799 ( .A(n9471), .B(n9395), .Z(n9398) );
  XOR U9800 ( .A(n9394), .B(n9393), .Z(n9427) );
  XOR U9801 ( .A(n9396), .B(n9395), .Z(n9426) );
  NOR U9802 ( .A(n9427), .B(n9426), .Z(n9397) );
  NOR U9803 ( .A(n9398), .B(n9397), .Z(n9422) );
  XOR U9804 ( .A(n9400), .B(n9399), .Z(n9421) );
  IV U9805 ( .A(n9421), .Z(n9401) );
  NOR U9806 ( .A(n9422), .B(n9401), .Z(n9402) );
  NOR U9807 ( .A(n9403), .B(n9402), .Z(n9456) );
  XOR U9808 ( .A(n9405), .B(n9404), .Z(n9455) );
  IV U9809 ( .A(n9455), .Z(n9406) );
  NOR U9810 ( .A(n9456), .B(n9406), .Z(n9407) );
  NOR U9811 ( .A(n9408), .B(n9407), .Z(n9413) );
  IV U9812 ( .A(n9413), .Z(n9411) );
  XOR U9813 ( .A(n9410), .B(n9409), .Z(n9412) );
  NOR U9814 ( .A(n9411), .B(n9412), .Z(n9646) );
  XOR U9815 ( .A(n9413), .B(n9412), .Z(n9854) );
  NOR U9816 ( .A(n9599), .B(n9414), .Z(n9415) );
  IV U9817 ( .A(n9415), .Z(n9462) );
  NOR U9818 ( .A(n9460), .B(n9462), .Z(n9420) );
  IV U9819 ( .A(n9416), .Z(n9418) );
  NOR U9820 ( .A(n9418), .B(n9417), .Z(n9419) );
  NOR U9821 ( .A(n9420), .B(n9419), .Z(n9423) );
  XOR U9822 ( .A(n9422), .B(n9421), .Z(n9424) );
  NOR U9823 ( .A(n9423), .B(n9424), .Z(n9454) );
  IV U9824 ( .A(n9423), .Z(n9425) );
  XOR U9825 ( .A(n9425), .B(n9424), .Z(n9458) );
  XOR U9826 ( .A(n9427), .B(n9426), .Z(n9447) );
  NOR U9827 ( .A(n9571), .B(n9526), .Z(n9434) );
  NOR U9828 ( .A(n9428), .B(n9434), .Z(n9436) );
  NOR U9829 ( .A(n9472), .B(n9584), .Z(n9431) );
  NOR U9830 ( .A(n9429), .B(n9592), .Z(n9430) );
  XOR U9831 ( .A(n9431), .B(n9430), .Z(n9432) );
  IV U9832 ( .A(n9432), .Z(n9461) );
  XOR U9833 ( .A(n9462), .B(n9461), .Z(n9468) );
  XOR U9834 ( .A(n9434), .B(n9433), .Z(n9467) );
  NOR U9835 ( .A(n9468), .B(n9467), .Z(n9435) );
  NOR U9836 ( .A(n9436), .B(n9435), .Z(n9448) );
  NOR U9837 ( .A(n9447), .B(n9448), .Z(n9451) );
  XOR U9838 ( .A(n9437), .B(sum[6]), .Z(n9441) );
  NOR U9839 ( .A(n9438), .B(n9441), .Z(n9445) );
  IV U9840 ( .A(sum[5]), .Z(n9440) );
  NOR U9841 ( .A(n9593), .B(n9526), .Z(n9439) );
  IV U9842 ( .A(n9439), .Z(n9491) );
  NOR U9843 ( .A(n9440), .B(n9491), .Z(n9470) );
  IV U9844 ( .A(n9470), .Z(n9443) );
  XOR U9845 ( .A(n9442), .B(n9441), .Z(n9469) );
  NOR U9846 ( .A(n9443), .B(n9469), .Z(n9444) );
  NOR U9847 ( .A(n9445), .B(n9444), .Z(n9446) );
  IV U9848 ( .A(n9446), .Z(n9466) );
  XOR U9849 ( .A(n9448), .B(n9447), .Z(n9449) );
  IV U9850 ( .A(n9449), .Z(n9465) );
  NOR U9851 ( .A(n9466), .B(n9465), .Z(n9450) );
  NOR U9852 ( .A(n9451), .B(n9450), .Z(n9452) );
  IV U9853 ( .A(n9452), .Z(n9457) );
  NOR U9854 ( .A(n9458), .B(n9457), .Z(n9453) );
  NOR U9855 ( .A(n9454), .B(n9453), .Z(n9640) );
  XOR U9856 ( .A(n9456), .B(n9455), .Z(n9639) );
  NOR U9857 ( .A(n9640), .B(n9639), .Z(n9643) );
  XOR U9858 ( .A(n9458), .B(n9457), .Z(n9634) );
  NOR U9859 ( .A(n9460), .B(n9459), .Z(n9464) );
  NOR U9860 ( .A(n9462), .B(n9461), .Z(n9463) );
  NOR U9861 ( .A(n9464), .B(n9463), .Z(n9485) );
  XOR U9862 ( .A(n9466), .B(n9465), .Z(n9484) );
  NOR U9863 ( .A(n9485), .B(n9484), .Z(n9488) );
  XOR U9864 ( .A(n9468), .B(n9467), .Z(n9480) );
  XOR U9865 ( .A(n9470), .B(n9469), .Z(n9479) );
  NOR U9866 ( .A(n9480), .B(n9479), .Z(n9483) );
  NOR U9867 ( .A(n9600), .B(n9493), .Z(n9572) );
  IV U9868 ( .A(n9572), .Z(n9575) );
  NOR U9869 ( .A(n9471), .B(n9575), .Z(n9478) );
  NOR U9870 ( .A(n9599), .B(n9472), .Z(n9473) );
  IV U9871 ( .A(n9473), .Z(n9502) );
  NOR U9872 ( .A(n9571), .B(n9493), .Z(n9475) );
  XOR U9873 ( .A(n9475), .B(n9474), .Z(n9476) );
  IV U9874 ( .A(n9476), .Z(n9501) );
  NOR U9875 ( .A(n9502), .B(n9501), .Z(n9477) );
  NOR U9876 ( .A(n9478), .B(n9477), .Z(n9513) );
  XOR U9877 ( .A(n9480), .B(n9479), .Z(n9514) );
  IV U9878 ( .A(n9514), .Z(n9481) );
  NOR U9879 ( .A(n9513), .B(n9481), .Z(n9482) );
  NOR U9880 ( .A(n9483), .B(n9482), .Z(n9518) );
  XOR U9881 ( .A(n9485), .B(n9484), .Z(n9517) );
  IV U9882 ( .A(n9517), .Z(n9486) );
  NOR U9883 ( .A(n9518), .B(n9486), .Z(n9487) );
  NOR U9884 ( .A(n9488), .B(n9487), .Z(n9633) );
  IV U9885 ( .A(n9633), .Z(n9489) );
  NOR U9886 ( .A(n9634), .B(n9489), .Z(n9637) );
  NOR U9887 ( .A(n9490), .B(n9584), .Z(n9498) );
  IV U9888 ( .A(n9498), .Z(n9492) );
  XOR U9889 ( .A(n9491), .B(sum[5]), .Z(n9497) );
  NOR U9890 ( .A(n9492), .B(n9497), .Z(n9500) );
  IV U9891 ( .A(sum[4]), .Z(n9495) );
  NOR U9892 ( .A(n9593), .B(n9493), .Z(n9494) );
  IV U9893 ( .A(n9494), .Z(n9534) );
  NOR U9894 ( .A(n9495), .B(n9534), .Z(n9496) );
  IV U9895 ( .A(n9496), .Z(n9505) );
  XOR U9896 ( .A(n9498), .B(n9497), .Z(n9504) );
  NOR U9897 ( .A(n9505), .B(n9504), .Z(n9499) );
  NOR U9898 ( .A(n9500), .B(n9499), .Z(n9512) );
  XOR U9899 ( .A(n9502), .B(n9501), .Z(n9506) );
  NOR U9900 ( .A(n9503), .B(n9506), .Z(n9509) );
  XOR U9901 ( .A(n9505), .B(n9504), .Z(n9532) );
  XOR U9902 ( .A(n9507), .B(n9506), .Z(n9533) );
  NOR U9903 ( .A(n9532), .B(n9533), .Z(n9508) );
  NOR U9904 ( .A(n9509), .B(n9508), .Z(n9511) );
  IV U9905 ( .A(n9511), .Z(n9510) );
  NOR U9906 ( .A(n9512), .B(n9510), .Z(n9516) );
  XOR U9907 ( .A(n9512), .B(n9511), .Z(n9523) );
  XOR U9908 ( .A(n9514), .B(n9513), .Z(n9522) );
  NOR U9909 ( .A(n9523), .B(n9522), .Z(n9515) );
  NOR U9910 ( .A(n9516), .B(n9515), .Z(n9520) );
  XOR U9911 ( .A(n9518), .B(n9517), .Z(n9519) );
  NOR U9912 ( .A(n9520), .B(n9519), .Z(n9632) );
  XOR U9913 ( .A(n9520), .B(n9519), .Z(n9521) );
  IV U9914 ( .A(n9521), .Z(n9869) );
  XOR U9915 ( .A(n9523), .B(n9522), .Z(n9550) );
  NOR U9916 ( .A(n9600), .B(n9592), .Z(n9524) );
  IV U9917 ( .A(n9524), .Z(n9903) );
  NOR U9918 ( .A(n9525), .B(n9903), .Z(n9531) );
  NOR U9919 ( .A(n9600), .B(n9526), .Z(n9527) );
  XOR U9920 ( .A(n9528), .B(n9527), .Z(n9554) );
  IV U9921 ( .A(n9554), .Z(n9529) );
  NOR U9922 ( .A(n9553), .B(n9529), .Z(n9530) );
  NOR U9923 ( .A(n9531), .B(n9530), .Z(n9544) );
  XOR U9924 ( .A(n9533), .B(n9532), .Z(n9543) );
  NOR U9925 ( .A(n9544), .B(n9543), .Z(n9547) );
  XOR U9926 ( .A(n9534), .B(sum[4]), .Z(n9538) );
  NOR U9927 ( .A(n9535), .B(n9538), .Z(n9542) );
  IV U9928 ( .A(sum[3]), .Z(n9537) );
  NOR U9929 ( .A(n9593), .B(n9584), .Z(n9536) );
  IV U9930 ( .A(n9536), .Z(n9555) );
  NOR U9931 ( .A(n9537), .B(n9555), .Z(n9552) );
  IV U9932 ( .A(n9552), .Z(n9540) );
  XOR U9933 ( .A(n9539), .B(n9538), .Z(n9551) );
  NOR U9934 ( .A(n9540), .B(n9551), .Z(n9541) );
  NOR U9935 ( .A(n9542), .B(n9541), .Z(n9570) );
  XOR U9936 ( .A(n9544), .B(n9543), .Z(n9569) );
  IV U9937 ( .A(n9569), .Z(n9545) );
  NOR U9938 ( .A(n9570), .B(n9545), .Z(n9546) );
  NOR U9939 ( .A(n9547), .B(n9546), .Z(n9549) );
  IV U9940 ( .A(n9549), .Z(n9548) );
  NOR U9941 ( .A(n9550), .B(n9548), .Z(n9629) );
  XOR U9942 ( .A(n9550), .B(n9549), .Z(n9874) );
  XOR U9943 ( .A(n9552), .B(n9551), .Z(n9564) );
  XOR U9944 ( .A(n9554), .B(n9553), .Z(n9565) );
  NOR U9945 ( .A(n9564), .B(n9565), .Z(n9568) );
  XOR U9946 ( .A(n9555), .B(sum[3]), .Z(n9560) );
  NOR U9947 ( .A(n9556), .B(n9560), .Z(n9563) );
  IV U9948 ( .A(sum[2]), .Z(n9558) );
  NOR U9949 ( .A(n9592), .B(n9571), .Z(n9557) );
  IV U9950 ( .A(n9557), .Z(n9582) );
  NOR U9951 ( .A(n9558), .B(n9582), .Z(n9559) );
  IV U9952 ( .A(n9559), .Z(n9574) );
  XOR U9953 ( .A(n9561), .B(n9560), .Z(n9573) );
  NOR U9954 ( .A(n9574), .B(n9573), .Z(n9562) );
  NOR U9955 ( .A(n9563), .B(n9562), .Z(n9580) );
  XOR U9956 ( .A(n9565), .B(n9564), .Z(n9579) );
  IV U9957 ( .A(n9579), .Z(n9566) );
  NOR U9958 ( .A(n9580), .B(n9566), .Z(n9567) );
  NOR U9959 ( .A(n9568), .B(n9567), .Z(n9623) );
  XOR U9960 ( .A(n9570), .B(n9569), .Z(n9622) );
  NOR U9961 ( .A(n9623), .B(n9622), .Z(n9626) );
  NOR U9962 ( .A(n9599), .B(n9571), .Z(n9576) );
  NOR U9963 ( .A(n9572), .B(n9576), .Z(n9578) );
  XOR U9964 ( .A(n9574), .B(n9573), .Z(n9590) );
  XOR U9965 ( .A(n9576), .B(n9575), .Z(n9591) );
  NOR U9966 ( .A(n9590), .B(n9591), .Z(n9577) );
  NOR U9967 ( .A(n9578), .B(n9577), .Z(n9619) );
  IV U9968 ( .A(n9619), .Z(n9581) );
  XOR U9969 ( .A(n9580), .B(n9579), .Z(n9618) );
  NOR U9970 ( .A(n9581), .B(n9618), .Z(n9621) );
  NOR U9971 ( .A(n9593), .B(n9599), .Z(n9586) );
  IV U9972 ( .A(n9586), .Z(n9583) );
  XOR U9973 ( .A(n9582), .B(sum[2]), .Z(n9585) );
  NOR U9974 ( .A(n9583), .B(n9585), .Z(n9589) );
  NOR U9975 ( .A(n9600), .B(n9584), .Z(n9597) );
  IV U9976 ( .A(n9597), .Z(n9587) );
  XOR U9977 ( .A(n9586), .B(n9585), .Z(n9596) );
  NOR U9978 ( .A(n9587), .B(n9596), .Z(n9588) );
  NOR U9979 ( .A(n9589), .B(n9588), .Z(n9613) );
  XOR U9980 ( .A(n9591), .B(n9590), .Z(n9614) );
  NOR U9981 ( .A(n9613), .B(n9614), .Z(n9617) );
  IV U9982 ( .A(sum[1]), .Z(n9595) );
  NOR U9983 ( .A(n9593), .B(n9592), .Z(n9594) );
  IV U9984 ( .A(n9594), .Z(n9601) );
  NOR U9985 ( .A(n9595), .B(n9601), .Z(n9610) );
  IV U9986 ( .A(n9610), .Z(n9598) );
  XOR U9987 ( .A(n9597), .B(n9596), .Z(n9609) );
  NOR U9988 ( .A(n9598), .B(n9609), .Z(n9612) );
  NOR U9989 ( .A(n9600), .B(n9599), .Z(n9606) );
  IV U9990 ( .A(n9606), .Z(n9602) );
  XOR U9991 ( .A(n9601), .B(sum[1]), .Z(n9605) );
  NOR U9992 ( .A(n9602), .B(n9605), .Z(n9608) );
  IV U9993 ( .A(sum[0]), .Z(n9603) );
  NOR U9994 ( .A(n9903), .B(n9603), .Z(n9604) );
  IV U9995 ( .A(n9604), .Z(n9899) );
  XOR U9996 ( .A(n9606), .B(n9605), .Z(n9898) );
  NOR U9997 ( .A(n9899), .B(n9898), .Z(n9607) );
  NOR U9998 ( .A(n9608), .B(n9607), .Z(n9893) );
  XOR U9999 ( .A(n9610), .B(n9609), .Z(n9894) );
  NOR U10000 ( .A(n9893), .B(n9894), .Z(n9611) );
  NOR U10001 ( .A(n9612), .B(n9611), .Z(n9889) );
  IV U10002 ( .A(n9613), .Z(n9615) );
  XOR U10003 ( .A(n9615), .B(n9614), .Z(n9888) );
  NOR U10004 ( .A(n9889), .B(n9888), .Z(n9616) );
  NOR U10005 ( .A(n9617), .B(n9616), .Z(n9883) );
  XOR U10006 ( .A(n9619), .B(n9618), .Z(n9884) );
  NOR U10007 ( .A(n9883), .B(n9884), .Z(n9620) );
  NOR U10008 ( .A(n9621), .B(n9620), .Z(n9878) );
  XOR U10009 ( .A(n9623), .B(n9622), .Z(n9624) );
  IV U10010 ( .A(n9624), .Z(n9879) );
  NOR U10011 ( .A(n9878), .B(n9879), .Z(n9625) );
  NOR U10012 ( .A(n9626), .B(n9625), .Z(n9873) );
  IV U10013 ( .A(n9873), .Z(n9627) );
  NOR U10014 ( .A(n9874), .B(n9627), .Z(n9628) );
  NOR U10015 ( .A(n9629), .B(n9628), .Z(n9630) );
  IV U10016 ( .A(n9630), .Z(n9868) );
  NOR U10017 ( .A(n9869), .B(n9868), .Z(n9631) );
  NOR U10018 ( .A(n9632), .B(n9631), .Z(n9864) );
  IV U10019 ( .A(n9864), .Z(n9635) );
  XOR U10020 ( .A(n9634), .B(n9633), .Z(n9863) );
  NOR U10021 ( .A(n9635), .B(n9863), .Z(n9636) );
  NOR U10022 ( .A(n9637), .B(n9636), .Z(n9638) );
  IV U10023 ( .A(n9638), .Z(n9859) );
  XOR U10024 ( .A(n9640), .B(n9639), .Z(n9641) );
  IV U10025 ( .A(n9641), .Z(n9858) );
  NOR U10026 ( .A(n9859), .B(n9858), .Z(n9642) );
  NOR U10027 ( .A(n9643), .B(n9642), .Z(n9853) );
  IV U10028 ( .A(n9853), .Z(n9644) );
  NOR U10029 ( .A(n9854), .B(n9644), .Z(n9645) );
  NOR U10030 ( .A(n9646), .B(n9645), .Z(n9647) );
  IV U10031 ( .A(n9647), .Z(n9848) );
  NOR U10032 ( .A(n9849), .B(n9848), .Z(n9648) );
  NOR U10033 ( .A(n9649), .B(n9648), .Z(n9843) );
  IV U10034 ( .A(n9843), .Z(n9650) );
  NOR U10035 ( .A(n9844), .B(n9650), .Z(n9651) );
  NOR U10036 ( .A(n9652), .B(n9651), .Z(n9653) );
  IV U10037 ( .A(n9653), .Z(n9838) );
  NOR U10038 ( .A(n9839), .B(n9838), .Z(n9654) );
  NOR U10039 ( .A(n9655), .B(n9654), .Z(n9834) );
  IV U10040 ( .A(n9834), .Z(n9658) );
  XOR U10041 ( .A(n9657), .B(n9656), .Z(n9833) );
  NOR U10042 ( .A(n9658), .B(n9833), .Z(n9659) );
  NOR U10043 ( .A(n9660), .B(n9659), .Z(n9661) );
  IV U10044 ( .A(n9661), .Z(n9829) );
  XOR U10045 ( .A(n9663), .B(n9662), .Z(n9828) );
  NOR U10046 ( .A(n9829), .B(n9828), .Z(n9664) );
  NOR U10047 ( .A(n9665), .B(n9664), .Z(n9824) );
  IV U10048 ( .A(n9824), .Z(n9668) );
  XOR U10049 ( .A(n9667), .B(n9666), .Z(n9823) );
  NOR U10050 ( .A(n9668), .B(n9823), .Z(n9669) );
  NOR U10051 ( .A(n9670), .B(n9669), .Z(n9671) );
  IV U10052 ( .A(n9671), .Z(n9818) );
  NOR U10053 ( .A(n9819), .B(n9818), .Z(n9672) );
  NOR U10054 ( .A(n9673), .B(n9672), .Z(n9814) );
  IV U10055 ( .A(n9814), .Z(n9676) );
  XOR U10056 ( .A(n9675), .B(n9674), .Z(n9813) );
  NOR U10057 ( .A(n9676), .B(n9813), .Z(n9677) );
  NOR U10058 ( .A(n9678), .B(n9677), .Z(n9679) );
  IV U10059 ( .A(n9679), .Z(n9809) );
  XOR U10060 ( .A(n9681), .B(n9680), .Z(n9808) );
  NOR U10061 ( .A(n9809), .B(n9808), .Z(n9682) );
  NOR U10062 ( .A(n9683), .B(n9682), .Z(n9803) );
  IV U10063 ( .A(n9803), .Z(n9684) );
  NOR U10064 ( .A(n9804), .B(n9684), .Z(n9685) );
  NOR U10065 ( .A(n9686), .B(n9685), .Z(n9687) );
  IV U10066 ( .A(n9687), .Z(n9799) );
  XOR U10067 ( .A(n9689), .B(n9688), .Z(n9798) );
  NOR U10068 ( .A(n9799), .B(n9798), .Z(n9690) );
  NOR U10069 ( .A(n9691), .B(n9690), .Z(n9794) );
  IV U10070 ( .A(n9794), .Z(n9694) );
  XOR U10071 ( .A(n9693), .B(n9692), .Z(n9793) );
  NOR U10072 ( .A(n9694), .B(n9793), .Z(n9695) );
  NOR U10073 ( .A(n9696), .B(n9695), .Z(n9697) );
  IV U10074 ( .A(n9697), .Z(n9789) );
  XOR U10075 ( .A(n9699), .B(n9698), .Z(n9788) );
  NOR U10076 ( .A(n9789), .B(n9788), .Z(n9700) );
  NOR U10077 ( .A(n9701), .B(n9700), .Z(n9784) );
  IV U10078 ( .A(n9784), .Z(n9704) );
  XOR U10079 ( .A(n9703), .B(n9702), .Z(n9783) );
  NOR U10080 ( .A(n9704), .B(n9783), .Z(n9705) );
  NOR U10081 ( .A(n9706), .B(n9705), .Z(n9707) );
  IV U10082 ( .A(n9707), .Z(n9778) );
  NOR U10083 ( .A(n9779), .B(n9778), .Z(n9708) );
  NOR U10084 ( .A(n9709), .B(n9708), .Z(n9773) );
  IV U10085 ( .A(n9773), .Z(n9710) );
  NOR U10086 ( .A(n9774), .B(n9710), .Z(n9711) );
  NOR U10087 ( .A(n9712), .B(n9711), .Z(n9713) );
  IV U10088 ( .A(n9713), .Z(n9769) );
  XOR U10089 ( .A(n9715), .B(n9714), .Z(n9768) );
  NOR U10090 ( .A(n9769), .B(n9768), .Z(n9716) );
  NOR U10091 ( .A(n9717), .B(n9716), .Z(n9764) );
  IV U10092 ( .A(n9764), .Z(n9720) );
  XOR U10093 ( .A(n9719), .B(n9718), .Z(n9763) );
  NOR U10094 ( .A(n9720), .B(n9763), .Z(n9721) );
  NOR U10095 ( .A(n9722), .B(n9721), .Z(n9723) );
  IV U10096 ( .A(n9723), .Z(n9758) );
  NOR U10097 ( .A(n9759), .B(n9758), .Z(n9724) );
  NOR U10098 ( .A(n9725), .B(n9724), .Z(n9753) );
  IV U10099 ( .A(n9753), .Z(n9726) );
  NOR U10100 ( .A(n9754), .B(n9726), .Z(n9727) );
  NOR U10101 ( .A(n9728), .B(n9727), .Z(n9737) );
  NOR U10102 ( .A(n9730), .B(n9729), .Z(n9735) );
  IV U10103 ( .A(n9731), .Z(n9733) );
  NOR U10104 ( .A(n9733), .B(n9732), .Z(n9734) );
  NOR U10105 ( .A(n9735), .B(n9734), .Z(n9736) );
  XOR U10106 ( .A(n9737), .B(n9736), .Z(n9747) );
  IV U10107 ( .A(n9738), .Z(n9739) );
  NOR U10108 ( .A(n9740), .B(n9739), .Z(n9745) );
  IV U10109 ( .A(n9741), .Z(n9742) );
  NOR U10110 ( .A(n9743), .B(n9742), .Z(n9744) );
  NOR U10111 ( .A(n9745), .B(n9744), .Z(n9746) );
  XOR U10112 ( .A(n9747), .B(n9746), .Z(n9748) );
  XOR U10113 ( .A(n9749), .B(n9748), .Z(n9750) );
  NOR U10114 ( .A(n9904), .B(n9750), .Z(n9751) );
  NOR U10115 ( .A(n9752), .B(n9751), .Z(n979) );
  NOR U10116 ( .A(sum[30]), .B(n3237), .Z(n9757) );
  XOR U10117 ( .A(n9754), .B(n9753), .Z(n9755) );
  NOR U10118 ( .A(n9904), .B(n9755), .Z(n9756) );
  NOR U10119 ( .A(n9757), .B(n9756), .Z(n980) );
  NOR U10120 ( .A(sum[29]), .B(n3237), .Z(n9762) );
  XOR U10121 ( .A(n9759), .B(n9758), .Z(n9760) );
  NOR U10122 ( .A(n9904), .B(n9760), .Z(n9761) );
  NOR U10123 ( .A(n9762), .B(n9761), .Z(n981) );
  NOR U10124 ( .A(sum[28]), .B(n3237), .Z(n9767) );
  XOR U10125 ( .A(n9764), .B(n9763), .Z(n9765) );
  NOR U10126 ( .A(n9904), .B(n9765), .Z(n9766) );
  NOR U10127 ( .A(n9767), .B(n9766), .Z(n982) );
  NOR U10128 ( .A(sum[27]), .B(n3237), .Z(n9772) );
  XOR U10129 ( .A(n9769), .B(n9768), .Z(n9770) );
  NOR U10130 ( .A(n9904), .B(n9770), .Z(n9771) );
  NOR U10131 ( .A(n9772), .B(n9771), .Z(n983) );
  NOR U10132 ( .A(sum[26]), .B(n3237), .Z(n9777) );
  XOR U10133 ( .A(n9774), .B(n9773), .Z(n9775) );
  NOR U10134 ( .A(n9904), .B(n9775), .Z(n9776) );
  NOR U10135 ( .A(n9777), .B(n9776), .Z(n984) );
  NOR U10136 ( .A(sum[25]), .B(n3237), .Z(n9782) );
  XOR U10137 ( .A(n9779), .B(n9778), .Z(n9780) );
  NOR U10138 ( .A(n9904), .B(n9780), .Z(n9781) );
  NOR U10139 ( .A(n9782), .B(n9781), .Z(n985) );
  NOR U10140 ( .A(sum[24]), .B(n3237), .Z(n9787) );
  XOR U10141 ( .A(n9784), .B(n9783), .Z(n9785) );
  NOR U10142 ( .A(n9904), .B(n9785), .Z(n9786) );
  NOR U10143 ( .A(n9787), .B(n9786), .Z(n986) );
  NOR U10144 ( .A(sum[23]), .B(n3237), .Z(n9792) );
  XOR U10145 ( .A(n9789), .B(n9788), .Z(n9790) );
  NOR U10146 ( .A(n9904), .B(n9790), .Z(n9791) );
  NOR U10147 ( .A(n9792), .B(n9791), .Z(n987) );
  NOR U10148 ( .A(sum[22]), .B(n3237), .Z(n9797) );
  XOR U10149 ( .A(n9794), .B(n9793), .Z(n9795) );
  NOR U10150 ( .A(n9904), .B(n9795), .Z(n9796) );
  NOR U10151 ( .A(n9797), .B(n9796), .Z(n988) );
  NOR U10152 ( .A(sum[21]), .B(n3237), .Z(n9802) );
  XOR U10153 ( .A(n9799), .B(n9798), .Z(n9800) );
  NOR U10154 ( .A(n9904), .B(n9800), .Z(n9801) );
  NOR U10155 ( .A(n9802), .B(n9801), .Z(n989) );
  NOR U10156 ( .A(sum[20]), .B(n3237), .Z(n9807) );
  XOR U10157 ( .A(n9804), .B(n9803), .Z(n9805) );
  NOR U10158 ( .A(n9904), .B(n9805), .Z(n9806) );
  NOR U10159 ( .A(n9807), .B(n9806), .Z(n990) );
  NOR U10160 ( .A(sum[19]), .B(n3237), .Z(n9812) );
  XOR U10161 ( .A(n9809), .B(n9808), .Z(n9810) );
  NOR U10162 ( .A(n9904), .B(n9810), .Z(n9811) );
  NOR U10163 ( .A(n9812), .B(n9811), .Z(n991) );
  NOR U10164 ( .A(sum[18]), .B(n3237), .Z(n9817) );
  XOR U10165 ( .A(n9814), .B(n9813), .Z(n9815) );
  NOR U10166 ( .A(n9904), .B(n9815), .Z(n9816) );
  NOR U10167 ( .A(n9817), .B(n9816), .Z(n992) );
  NOR U10168 ( .A(sum[17]), .B(n3237), .Z(n9822) );
  XOR U10169 ( .A(n9819), .B(n9818), .Z(n9820) );
  NOR U10170 ( .A(n9904), .B(n9820), .Z(n9821) );
  NOR U10171 ( .A(n9822), .B(n9821), .Z(n993) );
  NOR U10172 ( .A(sum[16]), .B(n3237), .Z(n9827) );
  XOR U10173 ( .A(n9824), .B(n9823), .Z(n9825) );
  NOR U10174 ( .A(n9904), .B(n9825), .Z(n9826) );
  NOR U10175 ( .A(n9827), .B(n9826), .Z(n994) );
  NOR U10176 ( .A(sum[15]), .B(n3237), .Z(n9832) );
  XOR U10177 ( .A(n9829), .B(n9828), .Z(n9830) );
  NOR U10178 ( .A(n9904), .B(n9830), .Z(n9831) );
  NOR U10179 ( .A(n9832), .B(n9831), .Z(n995) );
  NOR U10180 ( .A(sum[14]), .B(n3237), .Z(n9837) );
  XOR U10181 ( .A(n9834), .B(n9833), .Z(n9835) );
  NOR U10182 ( .A(n9904), .B(n9835), .Z(n9836) );
  NOR U10183 ( .A(n9837), .B(n9836), .Z(n996) );
  NOR U10184 ( .A(sum[13]), .B(n3237), .Z(n9842) );
  XOR U10185 ( .A(n9839), .B(n9838), .Z(n9840) );
  NOR U10186 ( .A(n9904), .B(n9840), .Z(n9841) );
  NOR U10187 ( .A(n9842), .B(n9841), .Z(n997) );
  NOR U10188 ( .A(sum[12]), .B(n3237), .Z(n9847) );
  XOR U10189 ( .A(n9844), .B(n9843), .Z(n9845) );
  NOR U10190 ( .A(n9904), .B(n9845), .Z(n9846) );
  NOR U10191 ( .A(n9847), .B(n9846), .Z(n998) );
  NOR U10192 ( .A(sum[11]), .B(n3237), .Z(n9852) );
  XOR U10193 ( .A(n9849), .B(n9848), .Z(n9850) );
  NOR U10194 ( .A(n9904), .B(n9850), .Z(n9851) );
  NOR U10195 ( .A(n9852), .B(n9851), .Z(n999) );
  NOR U10196 ( .A(sum[10]), .B(n3237), .Z(n9857) );
  XOR U10197 ( .A(n9854), .B(n9853), .Z(n9855) );
  NOR U10198 ( .A(n9904), .B(n9855), .Z(n9856) );
  NOR U10199 ( .A(n9857), .B(n9856), .Z(n1000) );
  NOR U10200 ( .A(sum[9]), .B(n3237), .Z(n9862) );
  XOR U10201 ( .A(n9859), .B(n9858), .Z(n9860) );
  NOR U10202 ( .A(n9904), .B(n9860), .Z(n9861) );
  NOR U10203 ( .A(n9862), .B(n9861), .Z(n1001) );
  NOR U10204 ( .A(sum[8]), .B(n3237), .Z(n9867) );
  XOR U10205 ( .A(n9864), .B(n9863), .Z(n9865) );
  NOR U10206 ( .A(n9904), .B(n9865), .Z(n9866) );
  NOR U10207 ( .A(n9867), .B(n9866), .Z(n1002) );
  NOR U10208 ( .A(sum[7]), .B(n3237), .Z(n9872) );
  XOR U10209 ( .A(n9869), .B(n9868), .Z(n9870) );
  NOR U10210 ( .A(n9904), .B(n9870), .Z(n9871) );
  NOR U10211 ( .A(n9872), .B(n9871), .Z(n1003) );
  NOR U10212 ( .A(sum[6]), .B(n3237), .Z(n9877) );
  XOR U10213 ( .A(n9874), .B(n9873), .Z(n9875) );
  NOR U10214 ( .A(n9904), .B(n9875), .Z(n9876) );
  NOR U10215 ( .A(n9877), .B(n9876), .Z(n1004) );
  NOR U10216 ( .A(sum[5]), .B(n3237), .Z(n9882) );
  XOR U10217 ( .A(n9879), .B(n9878), .Z(n9880) );
  NOR U10218 ( .A(n9904), .B(n9880), .Z(n9881) );
  NOR U10219 ( .A(n9882), .B(n9881), .Z(n1005) );
  NOR U10220 ( .A(sum[4]), .B(n3237), .Z(n9887) );
  XOR U10221 ( .A(n9884), .B(n9883), .Z(n9885) );
  NOR U10222 ( .A(n9904), .B(n9885), .Z(n9886) );
  NOR U10223 ( .A(n9887), .B(n9886), .Z(n1006) );
  NOR U10224 ( .A(sum[3]), .B(n3237), .Z(n9892) );
  XOR U10225 ( .A(n9889), .B(n9888), .Z(n9890) );
  NOR U10226 ( .A(n9904), .B(n9890), .Z(n9891) );
  NOR U10227 ( .A(n9892), .B(n9891), .Z(n1007) );
  NOR U10228 ( .A(sum[2]), .B(n3237), .Z(n9897) );
  XOR U10229 ( .A(n9894), .B(n9893), .Z(n9895) );
  NOR U10230 ( .A(n9904), .B(n9895), .Z(n9896) );
  NOR U10231 ( .A(n9897), .B(n9896), .Z(n1008) );
  NOR U10232 ( .A(sum[1]), .B(n3237), .Z(n9902) );
  XOR U10233 ( .A(n9899), .B(n9898), .Z(n9900) );
  NOR U10234 ( .A(n9904), .B(n9900), .Z(n9901) );
  NOR U10235 ( .A(n9902), .B(n9901), .Z(n1009) );
  NOR U10236 ( .A(n9904), .B(n9903), .Z(n9905) );
  XOR U10237 ( .A(sum[0]), .B(n9905), .Z(n1010) );
  XOR U10238 ( .A(i[0]), .B(n9906), .Z(n1011) );
endmodule

