
module mult_N128_CC128 ( clk, rst, a, b, c );
  input [127:0] a;
  input [0:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637;
  wire   [255:0] sreg;

  DFF \sreg_reg[254]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U4 ( .A(b[0]), .B(a[0]), .Z(n1) );
  XNOR U5 ( .A(n1), .B(sreg[127]), .Z(c[127]) );
  NAND U6 ( .A(b[0]), .B(a[1]), .Z(n2) );
  XOR U7 ( .A(sreg[128]), .B(n2), .Z(n4) );
  NANDN U8 ( .A(n1), .B(sreg[127]), .Z(n3) );
  XOR U9 ( .A(n4), .B(n3), .Z(c[128]) );
  NAND U10 ( .A(b[0]), .B(a[2]), .Z(n7) );
  XOR U11 ( .A(sreg[129]), .B(n7), .Z(n9) );
  NANDN U12 ( .A(n2), .B(sreg[128]), .Z(n6) );
  OR U13 ( .A(n4), .B(n3), .Z(n5) );
  AND U14 ( .A(n6), .B(n5), .Z(n8) );
  XOR U15 ( .A(n9), .B(n8), .Z(c[129]) );
  NAND U16 ( .A(b[0]), .B(a[3]), .Z(n12) );
  XOR U17 ( .A(sreg[130]), .B(n12), .Z(n14) );
  NANDN U18 ( .A(n7), .B(sreg[129]), .Z(n11) );
  OR U19 ( .A(n9), .B(n8), .Z(n10) );
  AND U20 ( .A(n11), .B(n10), .Z(n13) );
  XOR U21 ( .A(n14), .B(n13), .Z(c[130]) );
  NAND U22 ( .A(b[0]), .B(a[4]), .Z(n17) );
  XOR U23 ( .A(sreg[131]), .B(n17), .Z(n19) );
  NANDN U24 ( .A(n12), .B(sreg[130]), .Z(n16) );
  OR U25 ( .A(n14), .B(n13), .Z(n15) );
  AND U26 ( .A(n16), .B(n15), .Z(n18) );
  XOR U27 ( .A(n19), .B(n18), .Z(c[131]) );
  NAND U28 ( .A(b[0]), .B(a[5]), .Z(n22) );
  XOR U29 ( .A(sreg[132]), .B(n22), .Z(n24) );
  NANDN U30 ( .A(n17), .B(sreg[131]), .Z(n21) );
  OR U31 ( .A(n19), .B(n18), .Z(n20) );
  AND U32 ( .A(n21), .B(n20), .Z(n23) );
  XOR U33 ( .A(n24), .B(n23), .Z(c[132]) );
  NAND U34 ( .A(b[0]), .B(a[6]), .Z(n27) );
  XOR U35 ( .A(sreg[133]), .B(n27), .Z(n29) );
  NANDN U36 ( .A(n22), .B(sreg[132]), .Z(n26) );
  OR U37 ( .A(n24), .B(n23), .Z(n25) );
  AND U38 ( .A(n26), .B(n25), .Z(n28) );
  XOR U39 ( .A(n29), .B(n28), .Z(c[133]) );
  NAND U40 ( .A(b[0]), .B(a[7]), .Z(n32) );
  XOR U41 ( .A(sreg[134]), .B(n32), .Z(n34) );
  NANDN U42 ( .A(n27), .B(sreg[133]), .Z(n31) );
  OR U43 ( .A(n29), .B(n28), .Z(n30) );
  AND U44 ( .A(n31), .B(n30), .Z(n33) );
  XOR U45 ( .A(n34), .B(n33), .Z(c[134]) );
  NAND U46 ( .A(b[0]), .B(a[8]), .Z(n37) );
  XOR U47 ( .A(sreg[135]), .B(n37), .Z(n39) );
  NANDN U48 ( .A(n32), .B(sreg[134]), .Z(n36) );
  OR U49 ( .A(n34), .B(n33), .Z(n35) );
  AND U50 ( .A(n36), .B(n35), .Z(n38) );
  XOR U51 ( .A(n39), .B(n38), .Z(c[135]) );
  NAND U52 ( .A(b[0]), .B(a[9]), .Z(n42) );
  XOR U53 ( .A(sreg[136]), .B(n42), .Z(n44) );
  NANDN U54 ( .A(n37), .B(sreg[135]), .Z(n41) );
  OR U55 ( .A(n39), .B(n38), .Z(n40) );
  AND U56 ( .A(n41), .B(n40), .Z(n43) );
  XOR U57 ( .A(n44), .B(n43), .Z(c[136]) );
  NAND U58 ( .A(b[0]), .B(a[10]), .Z(n47) );
  XOR U59 ( .A(sreg[137]), .B(n47), .Z(n49) );
  NANDN U60 ( .A(n42), .B(sreg[136]), .Z(n46) );
  OR U61 ( .A(n44), .B(n43), .Z(n45) );
  AND U62 ( .A(n46), .B(n45), .Z(n48) );
  XOR U63 ( .A(n49), .B(n48), .Z(c[137]) );
  NAND U64 ( .A(b[0]), .B(a[11]), .Z(n52) );
  XOR U65 ( .A(sreg[138]), .B(n52), .Z(n54) );
  NANDN U66 ( .A(n47), .B(sreg[137]), .Z(n51) );
  OR U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XOR U69 ( .A(n54), .B(n53), .Z(c[138]) );
  NAND U70 ( .A(b[0]), .B(a[12]), .Z(n57) );
  XOR U71 ( .A(sreg[139]), .B(n57), .Z(n59) );
  NANDN U72 ( .A(n52), .B(sreg[138]), .Z(n56) );
  OR U73 ( .A(n54), .B(n53), .Z(n55) );
  AND U74 ( .A(n56), .B(n55), .Z(n58) );
  XOR U75 ( .A(n59), .B(n58), .Z(c[139]) );
  NAND U76 ( .A(b[0]), .B(a[13]), .Z(n62) );
  XOR U77 ( .A(sreg[140]), .B(n62), .Z(n64) );
  NANDN U78 ( .A(n57), .B(sreg[139]), .Z(n61) );
  OR U79 ( .A(n59), .B(n58), .Z(n60) );
  AND U80 ( .A(n61), .B(n60), .Z(n63) );
  XOR U81 ( .A(n64), .B(n63), .Z(c[140]) );
  NAND U82 ( .A(b[0]), .B(a[14]), .Z(n67) );
  XOR U83 ( .A(sreg[141]), .B(n67), .Z(n69) );
  NANDN U84 ( .A(n62), .B(sreg[140]), .Z(n66) );
  OR U85 ( .A(n64), .B(n63), .Z(n65) );
  AND U86 ( .A(n66), .B(n65), .Z(n68) );
  XOR U87 ( .A(n69), .B(n68), .Z(c[141]) );
  NAND U88 ( .A(b[0]), .B(a[15]), .Z(n72) );
  XOR U89 ( .A(sreg[142]), .B(n72), .Z(n74) );
  NANDN U90 ( .A(n67), .B(sreg[141]), .Z(n71) );
  OR U91 ( .A(n69), .B(n68), .Z(n70) );
  AND U92 ( .A(n71), .B(n70), .Z(n73) );
  XOR U93 ( .A(n74), .B(n73), .Z(c[142]) );
  NAND U94 ( .A(b[0]), .B(a[16]), .Z(n77) );
  XOR U95 ( .A(sreg[143]), .B(n77), .Z(n79) );
  NANDN U96 ( .A(n72), .B(sreg[142]), .Z(n76) );
  OR U97 ( .A(n74), .B(n73), .Z(n75) );
  AND U98 ( .A(n76), .B(n75), .Z(n78) );
  XOR U99 ( .A(n79), .B(n78), .Z(c[143]) );
  NAND U100 ( .A(b[0]), .B(a[17]), .Z(n82) );
  XOR U101 ( .A(sreg[144]), .B(n82), .Z(n84) );
  NANDN U102 ( .A(n77), .B(sreg[143]), .Z(n81) );
  OR U103 ( .A(n79), .B(n78), .Z(n80) );
  AND U104 ( .A(n81), .B(n80), .Z(n83) );
  XOR U105 ( .A(n84), .B(n83), .Z(c[144]) );
  NAND U106 ( .A(b[0]), .B(a[18]), .Z(n87) );
  XOR U107 ( .A(sreg[145]), .B(n87), .Z(n89) );
  NANDN U108 ( .A(n82), .B(sreg[144]), .Z(n86) );
  OR U109 ( .A(n84), .B(n83), .Z(n85) );
  AND U110 ( .A(n86), .B(n85), .Z(n88) );
  XOR U111 ( .A(n89), .B(n88), .Z(c[145]) );
  NAND U112 ( .A(b[0]), .B(a[19]), .Z(n92) );
  XOR U113 ( .A(sreg[146]), .B(n92), .Z(n94) );
  NANDN U114 ( .A(n87), .B(sreg[145]), .Z(n91) );
  OR U115 ( .A(n89), .B(n88), .Z(n90) );
  AND U116 ( .A(n91), .B(n90), .Z(n93) );
  XOR U117 ( .A(n94), .B(n93), .Z(c[146]) );
  NAND U118 ( .A(b[0]), .B(a[20]), .Z(n97) );
  XOR U119 ( .A(sreg[147]), .B(n97), .Z(n99) );
  NANDN U120 ( .A(n92), .B(sreg[146]), .Z(n96) );
  OR U121 ( .A(n94), .B(n93), .Z(n95) );
  AND U122 ( .A(n96), .B(n95), .Z(n98) );
  XOR U123 ( .A(n99), .B(n98), .Z(c[147]) );
  NAND U124 ( .A(b[0]), .B(a[21]), .Z(n102) );
  XOR U125 ( .A(sreg[148]), .B(n102), .Z(n104) );
  NANDN U126 ( .A(n97), .B(sreg[147]), .Z(n101) );
  OR U127 ( .A(n99), .B(n98), .Z(n100) );
  AND U128 ( .A(n101), .B(n100), .Z(n103) );
  XOR U129 ( .A(n104), .B(n103), .Z(c[148]) );
  NAND U130 ( .A(b[0]), .B(a[22]), .Z(n107) );
  XOR U131 ( .A(sreg[149]), .B(n107), .Z(n109) );
  NANDN U132 ( .A(n102), .B(sreg[148]), .Z(n106) );
  OR U133 ( .A(n104), .B(n103), .Z(n105) );
  AND U134 ( .A(n106), .B(n105), .Z(n108) );
  XOR U135 ( .A(n109), .B(n108), .Z(c[149]) );
  NAND U136 ( .A(b[0]), .B(a[23]), .Z(n112) );
  XOR U137 ( .A(sreg[150]), .B(n112), .Z(n114) );
  NANDN U138 ( .A(n107), .B(sreg[149]), .Z(n111) );
  OR U139 ( .A(n109), .B(n108), .Z(n110) );
  AND U140 ( .A(n111), .B(n110), .Z(n113) );
  XOR U141 ( .A(n114), .B(n113), .Z(c[150]) );
  NAND U142 ( .A(b[0]), .B(a[24]), .Z(n117) );
  XOR U143 ( .A(sreg[151]), .B(n117), .Z(n119) );
  NANDN U144 ( .A(n112), .B(sreg[150]), .Z(n116) );
  OR U145 ( .A(n114), .B(n113), .Z(n115) );
  AND U146 ( .A(n116), .B(n115), .Z(n118) );
  XOR U147 ( .A(n119), .B(n118), .Z(c[151]) );
  NAND U148 ( .A(b[0]), .B(a[25]), .Z(n122) );
  XOR U149 ( .A(sreg[152]), .B(n122), .Z(n124) );
  NANDN U150 ( .A(n117), .B(sreg[151]), .Z(n121) );
  OR U151 ( .A(n119), .B(n118), .Z(n120) );
  AND U152 ( .A(n121), .B(n120), .Z(n123) );
  XOR U153 ( .A(n124), .B(n123), .Z(c[152]) );
  NAND U154 ( .A(b[0]), .B(a[26]), .Z(n127) );
  XOR U155 ( .A(sreg[153]), .B(n127), .Z(n129) );
  NANDN U156 ( .A(n122), .B(sreg[152]), .Z(n126) );
  OR U157 ( .A(n124), .B(n123), .Z(n125) );
  AND U158 ( .A(n126), .B(n125), .Z(n128) );
  XOR U159 ( .A(n129), .B(n128), .Z(c[153]) );
  NAND U160 ( .A(b[0]), .B(a[27]), .Z(n132) );
  XOR U161 ( .A(sreg[154]), .B(n132), .Z(n134) );
  NANDN U162 ( .A(n127), .B(sreg[153]), .Z(n131) );
  OR U163 ( .A(n129), .B(n128), .Z(n130) );
  AND U164 ( .A(n131), .B(n130), .Z(n133) );
  XOR U165 ( .A(n134), .B(n133), .Z(c[154]) );
  NAND U166 ( .A(b[0]), .B(a[28]), .Z(n137) );
  XOR U167 ( .A(sreg[155]), .B(n137), .Z(n139) );
  NANDN U168 ( .A(n132), .B(sreg[154]), .Z(n136) );
  OR U169 ( .A(n134), .B(n133), .Z(n135) );
  AND U170 ( .A(n136), .B(n135), .Z(n138) );
  XOR U171 ( .A(n139), .B(n138), .Z(c[155]) );
  NAND U172 ( .A(b[0]), .B(a[29]), .Z(n142) );
  XOR U173 ( .A(sreg[156]), .B(n142), .Z(n144) );
  NANDN U174 ( .A(n137), .B(sreg[155]), .Z(n141) );
  OR U175 ( .A(n139), .B(n138), .Z(n140) );
  AND U176 ( .A(n141), .B(n140), .Z(n143) );
  XOR U177 ( .A(n144), .B(n143), .Z(c[156]) );
  NAND U178 ( .A(b[0]), .B(a[30]), .Z(n147) );
  XOR U179 ( .A(sreg[157]), .B(n147), .Z(n149) );
  NANDN U180 ( .A(n142), .B(sreg[156]), .Z(n146) );
  OR U181 ( .A(n144), .B(n143), .Z(n145) );
  AND U182 ( .A(n146), .B(n145), .Z(n148) );
  XOR U183 ( .A(n149), .B(n148), .Z(c[157]) );
  NAND U184 ( .A(b[0]), .B(a[31]), .Z(n152) );
  XOR U185 ( .A(sreg[158]), .B(n152), .Z(n154) );
  NANDN U186 ( .A(n147), .B(sreg[157]), .Z(n151) );
  OR U187 ( .A(n149), .B(n148), .Z(n150) );
  AND U188 ( .A(n151), .B(n150), .Z(n153) );
  XOR U189 ( .A(n154), .B(n153), .Z(c[158]) );
  NAND U190 ( .A(b[0]), .B(a[32]), .Z(n157) );
  XOR U191 ( .A(sreg[159]), .B(n157), .Z(n159) );
  NANDN U192 ( .A(n152), .B(sreg[158]), .Z(n156) );
  OR U193 ( .A(n154), .B(n153), .Z(n155) );
  AND U194 ( .A(n156), .B(n155), .Z(n158) );
  XOR U195 ( .A(n159), .B(n158), .Z(c[159]) );
  NAND U196 ( .A(b[0]), .B(a[33]), .Z(n162) );
  XOR U197 ( .A(sreg[160]), .B(n162), .Z(n164) );
  NANDN U198 ( .A(n157), .B(sreg[159]), .Z(n161) );
  OR U199 ( .A(n159), .B(n158), .Z(n160) );
  AND U200 ( .A(n161), .B(n160), .Z(n163) );
  XOR U201 ( .A(n164), .B(n163), .Z(c[160]) );
  NAND U202 ( .A(b[0]), .B(a[34]), .Z(n167) );
  XOR U203 ( .A(sreg[161]), .B(n167), .Z(n169) );
  NANDN U204 ( .A(n162), .B(sreg[160]), .Z(n166) );
  OR U205 ( .A(n164), .B(n163), .Z(n165) );
  AND U206 ( .A(n166), .B(n165), .Z(n168) );
  XOR U207 ( .A(n169), .B(n168), .Z(c[161]) );
  NAND U208 ( .A(b[0]), .B(a[35]), .Z(n172) );
  XOR U209 ( .A(sreg[162]), .B(n172), .Z(n174) );
  NANDN U210 ( .A(n167), .B(sreg[161]), .Z(n171) );
  OR U211 ( .A(n169), .B(n168), .Z(n170) );
  AND U212 ( .A(n171), .B(n170), .Z(n173) );
  XOR U213 ( .A(n174), .B(n173), .Z(c[162]) );
  NAND U214 ( .A(b[0]), .B(a[36]), .Z(n177) );
  XOR U215 ( .A(sreg[163]), .B(n177), .Z(n179) );
  NANDN U216 ( .A(n172), .B(sreg[162]), .Z(n176) );
  OR U217 ( .A(n174), .B(n173), .Z(n175) );
  AND U218 ( .A(n176), .B(n175), .Z(n178) );
  XOR U219 ( .A(n179), .B(n178), .Z(c[163]) );
  NAND U220 ( .A(b[0]), .B(a[37]), .Z(n182) );
  XOR U221 ( .A(sreg[164]), .B(n182), .Z(n184) );
  NANDN U222 ( .A(n177), .B(sreg[163]), .Z(n181) );
  OR U223 ( .A(n179), .B(n178), .Z(n180) );
  AND U224 ( .A(n181), .B(n180), .Z(n183) );
  XOR U225 ( .A(n184), .B(n183), .Z(c[164]) );
  NAND U226 ( .A(b[0]), .B(a[38]), .Z(n187) );
  XOR U227 ( .A(sreg[165]), .B(n187), .Z(n189) );
  NANDN U228 ( .A(n182), .B(sreg[164]), .Z(n186) );
  OR U229 ( .A(n184), .B(n183), .Z(n185) );
  AND U230 ( .A(n186), .B(n185), .Z(n188) );
  XOR U231 ( .A(n189), .B(n188), .Z(c[165]) );
  NAND U232 ( .A(b[0]), .B(a[39]), .Z(n192) );
  XOR U233 ( .A(sreg[166]), .B(n192), .Z(n194) );
  NANDN U234 ( .A(n187), .B(sreg[165]), .Z(n191) );
  OR U235 ( .A(n189), .B(n188), .Z(n190) );
  AND U236 ( .A(n191), .B(n190), .Z(n193) );
  XOR U237 ( .A(n194), .B(n193), .Z(c[166]) );
  NAND U238 ( .A(b[0]), .B(a[40]), .Z(n197) );
  XOR U239 ( .A(sreg[167]), .B(n197), .Z(n199) );
  NANDN U240 ( .A(n192), .B(sreg[166]), .Z(n196) );
  OR U241 ( .A(n194), .B(n193), .Z(n195) );
  AND U242 ( .A(n196), .B(n195), .Z(n198) );
  XOR U243 ( .A(n199), .B(n198), .Z(c[167]) );
  NAND U244 ( .A(b[0]), .B(a[41]), .Z(n202) );
  XOR U245 ( .A(sreg[168]), .B(n202), .Z(n204) );
  NANDN U246 ( .A(n197), .B(sreg[167]), .Z(n201) );
  OR U247 ( .A(n199), .B(n198), .Z(n200) );
  AND U248 ( .A(n201), .B(n200), .Z(n203) );
  XOR U249 ( .A(n204), .B(n203), .Z(c[168]) );
  NAND U250 ( .A(b[0]), .B(a[42]), .Z(n207) );
  XOR U251 ( .A(sreg[169]), .B(n207), .Z(n209) );
  NANDN U252 ( .A(n202), .B(sreg[168]), .Z(n206) );
  OR U253 ( .A(n204), .B(n203), .Z(n205) );
  AND U254 ( .A(n206), .B(n205), .Z(n208) );
  XOR U255 ( .A(n209), .B(n208), .Z(c[169]) );
  NAND U256 ( .A(b[0]), .B(a[43]), .Z(n212) );
  XOR U257 ( .A(sreg[170]), .B(n212), .Z(n214) );
  NANDN U258 ( .A(n207), .B(sreg[169]), .Z(n211) );
  OR U259 ( .A(n209), .B(n208), .Z(n210) );
  AND U260 ( .A(n211), .B(n210), .Z(n213) );
  XOR U261 ( .A(n214), .B(n213), .Z(c[170]) );
  NAND U262 ( .A(b[0]), .B(a[44]), .Z(n217) );
  XOR U263 ( .A(sreg[171]), .B(n217), .Z(n219) );
  NANDN U264 ( .A(n212), .B(sreg[170]), .Z(n216) );
  OR U265 ( .A(n214), .B(n213), .Z(n215) );
  AND U266 ( .A(n216), .B(n215), .Z(n218) );
  XOR U267 ( .A(n219), .B(n218), .Z(c[171]) );
  NAND U268 ( .A(b[0]), .B(a[45]), .Z(n222) );
  XOR U269 ( .A(sreg[172]), .B(n222), .Z(n224) );
  NANDN U270 ( .A(n217), .B(sreg[171]), .Z(n221) );
  OR U271 ( .A(n219), .B(n218), .Z(n220) );
  AND U272 ( .A(n221), .B(n220), .Z(n223) );
  XOR U273 ( .A(n224), .B(n223), .Z(c[172]) );
  NAND U274 ( .A(b[0]), .B(a[46]), .Z(n227) );
  XOR U275 ( .A(sreg[173]), .B(n227), .Z(n229) );
  NANDN U276 ( .A(n222), .B(sreg[172]), .Z(n226) );
  OR U277 ( .A(n224), .B(n223), .Z(n225) );
  AND U278 ( .A(n226), .B(n225), .Z(n228) );
  XOR U279 ( .A(n229), .B(n228), .Z(c[173]) );
  NAND U280 ( .A(b[0]), .B(a[47]), .Z(n232) );
  XOR U281 ( .A(sreg[174]), .B(n232), .Z(n234) );
  NANDN U282 ( .A(n227), .B(sreg[173]), .Z(n231) );
  OR U283 ( .A(n229), .B(n228), .Z(n230) );
  AND U284 ( .A(n231), .B(n230), .Z(n233) );
  XOR U285 ( .A(n234), .B(n233), .Z(c[174]) );
  NAND U286 ( .A(b[0]), .B(a[48]), .Z(n237) );
  XOR U287 ( .A(sreg[175]), .B(n237), .Z(n239) );
  NANDN U288 ( .A(n232), .B(sreg[174]), .Z(n236) );
  OR U289 ( .A(n234), .B(n233), .Z(n235) );
  AND U290 ( .A(n236), .B(n235), .Z(n238) );
  XOR U291 ( .A(n239), .B(n238), .Z(c[175]) );
  NAND U292 ( .A(b[0]), .B(a[49]), .Z(n242) );
  XOR U293 ( .A(sreg[176]), .B(n242), .Z(n244) );
  NANDN U294 ( .A(n237), .B(sreg[175]), .Z(n241) );
  OR U295 ( .A(n239), .B(n238), .Z(n240) );
  AND U296 ( .A(n241), .B(n240), .Z(n243) );
  XOR U297 ( .A(n244), .B(n243), .Z(c[176]) );
  NAND U298 ( .A(b[0]), .B(a[50]), .Z(n247) );
  XOR U299 ( .A(sreg[177]), .B(n247), .Z(n249) );
  NANDN U300 ( .A(n242), .B(sreg[176]), .Z(n246) );
  OR U301 ( .A(n244), .B(n243), .Z(n245) );
  AND U302 ( .A(n246), .B(n245), .Z(n248) );
  XOR U303 ( .A(n249), .B(n248), .Z(c[177]) );
  NAND U304 ( .A(b[0]), .B(a[51]), .Z(n252) );
  XOR U305 ( .A(sreg[178]), .B(n252), .Z(n254) );
  NANDN U306 ( .A(n247), .B(sreg[177]), .Z(n251) );
  OR U307 ( .A(n249), .B(n248), .Z(n250) );
  AND U308 ( .A(n251), .B(n250), .Z(n253) );
  XOR U309 ( .A(n254), .B(n253), .Z(c[178]) );
  NAND U310 ( .A(b[0]), .B(a[52]), .Z(n257) );
  XOR U311 ( .A(sreg[179]), .B(n257), .Z(n259) );
  NANDN U312 ( .A(n252), .B(sreg[178]), .Z(n256) );
  OR U313 ( .A(n254), .B(n253), .Z(n255) );
  AND U314 ( .A(n256), .B(n255), .Z(n258) );
  XOR U315 ( .A(n259), .B(n258), .Z(c[179]) );
  NAND U316 ( .A(b[0]), .B(a[53]), .Z(n262) );
  XOR U317 ( .A(sreg[180]), .B(n262), .Z(n264) );
  NANDN U318 ( .A(n257), .B(sreg[179]), .Z(n261) );
  OR U319 ( .A(n259), .B(n258), .Z(n260) );
  AND U320 ( .A(n261), .B(n260), .Z(n263) );
  XOR U321 ( .A(n264), .B(n263), .Z(c[180]) );
  NAND U322 ( .A(b[0]), .B(a[54]), .Z(n267) );
  XOR U323 ( .A(sreg[181]), .B(n267), .Z(n269) );
  NANDN U324 ( .A(n262), .B(sreg[180]), .Z(n266) );
  OR U325 ( .A(n264), .B(n263), .Z(n265) );
  AND U326 ( .A(n266), .B(n265), .Z(n268) );
  XOR U327 ( .A(n269), .B(n268), .Z(c[181]) );
  NAND U328 ( .A(b[0]), .B(a[55]), .Z(n272) );
  XOR U329 ( .A(sreg[182]), .B(n272), .Z(n274) );
  NANDN U330 ( .A(n267), .B(sreg[181]), .Z(n271) );
  OR U331 ( .A(n269), .B(n268), .Z(n270) );
  AND U332 ( .A(n271), .B(n270), .Z(n273) );
  XOR U333 ( .A(n274), .B(n273), .Z(c[182]) );
  NAND U334 ( .A(b[0]), .B(a[56]), .Z(n277) );
  XOR U335 ( .A(sreg[183]), .B(n277), .Z(n279) );
  NANDN U336 ( .A(n272), .B(sreg[182]), .Z(n276) );
  OR U337 ( .A(n274), .B(n273), .Z(n275) );
  AND U338 ( .A(n276), .B(n275), .Z(n278) );
  XOR U339 ( .A(n279), .B(n278), .Z(c[183]) );
  NAND U340 ( .A(b[0]), .B(a[57]), .Z(n282) );
  XOR U341 ( .A(sreg[184]), .B(n282), .Z(n284) );
  NANDN U342 ( .A(n277), .B(sreg[183]), .Z(n281) );
  OR U343 ( .A(n279), .B(n278), .Z(n280) );
  AND U344 ( .A(n281), .B(n280), .Z(n283) );
  XOR U345 ( .A(n284), .B(n283), .Z(c[184]) );
  NAND U346 ( .A(b[0]), .B(a[58]), .Z(n287) );
  XOR U347 ( .A(sreg[185]), .B(n287), .Z(n289) );
  NANDN U348 ( .A(n282), .B(sreg[184]), .Z(n286) );
  OR U349 ( .A(n284), .B(n283), .Z(n285) );
  AND U350 ( .A(n286), .B(n285), .Z(n288) );
  XOR U351 ( .A(n289), .B(n288), .Z(c[185]) );
  NAND U352 ( .A(b[0]), .B(a[59]), .Z(n292) );
  XOR U353 ( .A(sreg[186]), .B(n292), .Z(n294) );
  NANDN U354 ( .A(n287), .B(sreg[185]), .Z(n291) );
  OR U355 ( .A(n289), .B(n288), .Z(n290) );
  AND U356 ( .A(n291), .B(n290), .Z(n293) );
  XOR U357 ( .A(n294), .B(n293), .Z(c[186]) );
  NAND U358 ( .A(b[0]), .B(a[60]), .Z(n297) );
  XOR U359 ( .A(sreg[187]), .B(n297), .Z(n299) );
  NANDN U360 ( .A(n292), .B(sreg[186]), .Z(n296) );
  OR U361 ( .A(n294), .B(n293), .Z(n295) );
  AND U362 ( .A(n296), .B(n295), .Z(n298) );
  XOR U363 ( .A(n299), .B(n298), .Z(c[187]) );
  NAND U364 ( .A(b[0]), .B(a[61]), .Z(n302) );
  XOR U365 ( .A(sreg[188]), .B(n302), .Z(n304) );
  NANDN U366 ( .A(n297), .B(sreg[187]), .Z(n301) );
  OR U367 ( .A(n299), .B(n298), .Z(n300) );
  AND U368 ( .A(n301), .B(n300), .Z(n303) );
  XOR U369 ( .A(n304), .B(n303), .Z(c[188]) );
  NAND U370 ( .A(b[0]), .B(a[62]), .Z(n307) );
  XOR U371 ( .A(sreg[189]), .B(n307), .Z(n309) );
  NANDN U372 ( .A(n302), .B(sreg[188]), .Z(n306) );
  OR U373 ( .A(n304), .B(n303), .Z(n305) );
  AND U374 ( .A(n306), .B(n305), .Z(n308) );
  XOR U375 ( .A(n309), .B(n308), .Z(c[189]) );
  NAND U376 ( .A(b[0]), .B(a[63]), .Z(n312) );
  XOR U377 ( .A(sreg[190]), .B(n312), .Z(n314) );
  NANDN U378 ( .A(n307), .B(sreg[189]), .Z(n311) );
  OR U379 ( .A(n309), .B(n308), .Z(n310) );
  AND U380 ( .A(n311), .B(n310), .Z(n313) );
  XOR U381 ( .A(n314), .B(n313), .Z(c[190]) );
  NAND U382 ( .A(b[0]), .B(a[64]), .Z(n317) );
  XOR U383 ( .A(sreg[191]), .B(n317), .Z(n319) );
  NANDN U384 ( .A(n312), .B(sreg[190]), .Z(n316) );
  OR U385 ( .A(n314), .B(n313), .Z(n315) );
  AND U386 ( .A(n316), .B(n315), .Z(n318) );
  XOR U387 ( .A(n319), .B(n318), .Z(c[191]) );
  NAND U388 ( .A(b[0]), .B(a[65]), .Z(n322) );
  XOR U389 ( .A(sreg[192]), .B(n322), .Z(n324) );
  NANDN U390 ( .A(n317), .B(sreg[191]), .Z(n321) );
  OR U391 ( .A(n319), .B(n318), .Z(n320) );
  AND U392 ( .A(n321), .B(n320), .Z(n323) );
  XOR U393 ( .A(n324), .B(n323), .Z(c[192]) );
  NAND U394 ( .A(b[0]), .B(a[66]), .Z(n327) );
  XOR U395 ( .A(sreg[193]), .B(n327), .Z(n329) );
  NANDN U396 ( .A(n322), .B(sreg[192]), .Z(n326) );
  OR U397 ( .A(n324), .B(n323), .Z(n325) );
  AND U398 ( .A(n326), .B(n325), .Z(n328) );
  XOR U399 ( .A(n329), .B(n328), .Z(c[193]) );
  NAND U400 ( .A(b[0]), .B(a[67]), .Z(n332) );
  XOR U401 ( .A(sreg[194]), .B(n332), .Z(n334) );
  NANDN U402 ( .A(n327), .B(sreg[193]), .Z(n331) );
  OR U403 ( .A(n329), .B(n328), .Z(n330) );
  AND U404 ( .A(n331), .B(n330), .Z(n333) );
  XOR U405 ( .A(n334), .B(n333), .Z(c[194]) );
  NAND U406 ( .A(b[0]), .B(a[68]), .Z(n337) );
  XOR U407 ( .A(sreg[195]), .B(n337), .Z(n339) );
  NANDN U408 ( .A(n332), .B(sreg[194]), .Z(n336) );
  OR U409 ( .A(n334), .B(n333), .Z(n335) );
  AND U410 ( .A(n336), .B(n335), .Z(n338) );
  XOR U411 ( .A(n339), .B(n338), .Z(c[195]) );
  NAND U412 ( .A(b[0]), .B(a[69]), .Z(n342) );
  XOR U413 ( .A(sreg[196]), .B(n342), .Z(n344) );
  NANDN U414 ( .A(n337), .B(sreg[195]), .Z(n341) );
  OR U415 ( .A(n339), .B(n338), .Z(n340) );
  AND U416 ( .A(n341), .B(n340), .Z(n343) );
  XOR U417 ( .A(n344), .B(n343), .Z(c[196]) );
  NAND U418 ( .A(b[0]), .B(a[70]), .Z(n347) );
  XOR U419 ( .A(sreg[197]), .B(n347), .Z(n349) );
  NANDN U420 ( .A(n342), .B(sreg[196]), .Z(n346) );
  OR U421 ( .A(n344), .B(n343), .Z(n345) );
  AND U422 ( .A(n346), .B(n345), .Z(n348) );
  XOR U423 ( .A(n349), .B(n348), .Z(c[197]) );
  NAND U424 ( .A(b[0]), .B(a[71]), .Z(n352) );
  XOR U425 ( .A(sreg[198]), .B(n352), .Z(n354) );
  NANDN U426 ( .A(n347), .B(sreg[197]), .Z(n351) );
  OR U427 ( .A(n349), .B(n348), .Z(n350) );
  AND U428 ( .A(n351), .B(n350), .Z(n353) );
  XOR U429 ( .A(n354), .B(n353), .Z(c[198]) );
  NAND U430 ( .A(b[0]), .B(a[72]), .Z(n357) );
  XOR U431 ( .A(sreg[199]), .B(n357), .Z(n359) );
  NANDN U432 ( .A(n352), .B(sreg[198]), .Z(n356) );
  OR U433 ( .A(n354), .B(n353), .Z(n355) );
  AND U434 ( .A(n356), .B(n355), .Z(n358) );
  XOR U435 ( .A(n359), .B(n358), .Z(c[199]) );
  NAND U436 ( .A(b[0]), .B(a[73]), .Z(n362) );
  XOR U437 ( .A(sreg[200]), .B(n362), .Z(n364) );
  NANDN U438 ( .A(n357), .B(sreg[199]), .Z(n361) );
  OR U439 ( .A(n359), .B(n358), .Z(n360) );
  AND U440 ( .A(n361), .B(n360), .Z(n363) );
  XOR U441 ( .A(n364), .B(n363), .Z(c[200]) );
  NAND U442 ( .A(b[0]), .B(a[74]), .Z(n367) );
  XOR U443 ( .A(sreg[201]), .B(n367), .Z(n369) );
  NANDN U444 ( .A(n362), .B(sreg[200]), .Z(n366) );
  OR U445 ( .A(n364), .B(n363), .Z(n365) );
  AND U446 ( .A(n366), .B(n365), .Z(n368) );
  XOR U447 ( .A(n369), .B(n368), .Z(c[201]) );
  NAND U448 ( .A(b[0]), .B(a[75]), .Z(n372) );
  XOR U449 ( .A(sreg[202]), .B(n372), .Z(n374) );
  NANDN U450 ( .A(n367), .B(sreg[201]), .Z(n371) );
  OR U451 ( .A(n369), .B(n368), .Z(n370) );
  AND U452 ( .A(n371), .B(n370), .Z(n373) );
  XOR U453 ( .A(n374), .B(n373), .Z(c[202]) );
  NAND U454 ( .A(b[0]), .B(a[76]), .Z(n377) );
  XOR U455 ( .A(sreg[203]), .B(n377), .Z(n379) );
  NANDN U456 ( .A(n372), .B(sreg[202]), .Z(n376) );
  OR U457 ( .A(n374), .B(n373), .Z(n375) );
  AND U458 ( .A(n376), .B(n375), .Z(n378) );
  XOR U459 ( .A(n379), .B(n378), .Z(c[203]) );
  NAND U460 ( .A(b[0]), .B(a[77]), .Z(n382) );
  XOR U461 ( .A(sreg[204]), .B(n382), .Z(n384) );
  NANDN U462 ( .A(n377), .B(sreg[203]), .Z(n381) );
  OR U463 ( .A(n379), .B(n378), .Z(n380) );
  AND U464 ( .A(n381), .B(n380), .Z(n383) );
  XOR U465 ( .A(n384), .B(n383), .Z(c[204]) );
  NAND U466 ( .A(b[0]), .B(a[78]), .Z(n387) );
  XOR U467 ( .A(sreg[205]), .B(n387), .Z(n389) );
  NANDN U468 ( .A(n382), .B(sreg[204]), .Z(n386) );
  OR U469 ( .A(n384), .B(n383), .Z(n385) );
  AND U470 ( .A(n386), .B(n385), .Z(n388) );
  XOR U471 ( .A(n389), .B(n388), .Z(c[205]) );
  NAND U472 ( .A(b[0]), .B(a[79]), .Z(n392) );
  XOR U473 ( .A(sreg[206]), .B(n392), .Z(n394) );
  NANDN U474 ( .A(n387), .B(sreg[205]), .Z(n391) );
  OR U475 ( .A(n389), .B(n388), .Z(n390) );
  AND U476 ( .A(n391), .B(n390), .Z(n393) );
  XOR U477 ( .A(n394), .B(n393), .Z(c[206]) );
  NAND U478 ( .A(b[0]), .B(a[80]), .Z(n397) );
  XOR U479 ( .A(sreg[207]), .B(n397), .Z(n399) );
  NANDN U480 ( .A(n392), .B(sreg[206]), .Z(n396) );
  OR U481 ( .A(n394), .B(n393), .Z(n395) );
  AND U482 ( .A(n396), .B(n395), .Z(n398) );
  XOR U483 ( .A(n399), .B(n398), .Z(c[207]) );
  NAND U484 ( .A(b[0]), .B(a[81]), .Z(n402) );
  XOR U485 ( .A(sreg[208]), .B(n402), .Z(n404) );
  NANDN U486 ( .A(n397), .B(sreg[207]), .Z(n401) );
  OR U487 ( .A(n399), .B(n398), .Z(n400) );
  AND U488 ( .A(n401), .B(n400), .Z(n403) );
  XOR U489 ( .A(n404), .B(n403), .Z(c[208]) );
  NAND U490 ( .A(b[0]), .B(a[82]), .Z(n407) );
  XOR U491 ( .A(sreg[209]), .B(n407), .Z(n409) );
  NANDN U492 ( .A(n402), .B(sreg[208]), .Z(n406) );
  OR U493 ( .A(n404), .B(n403), .Z(n405) );
  AND U494 ( .A(n406), .B(n405), .Z(n408) );
  XOR U495 ( .A(n409), .B(n408), .Z(c[209]) );
  NAND U496 ( .A(b[0]), .B(a[83]), .Z(n412) );
  XOR U497 ( .A(sreg[210]), .B(n412), .Z(n414) );
  NANDN U498 ( .A(n407), .B(sreg[209]), .Z(n411) );
  OR U499 ( .A(n409), .B(n408), .Z(n410) );
  AND U500 ( .A(n411), .B(n410), .Z(n413) );
  XOR U501 ( .A(n414), .B(n413), .Z(c[210]) );
  NAND U502 ( .A(b[0]), .B(a[84]), .Z(n417) );
  XOR U503 ( .A(sreg[211]), .B(n417), .Z(n419) );
  NANDN U504 ( .A(n412), .B(sreg[210]), .Z(n416) );
  OR U505 ( .A(n414), .B(n413), .Z(n415) );
  AND U506 ( .A(n416), .B(n415), .Z(n418) );
  XOR U507 ( .A(n419), .B(n418), .Z(c[211]) );
  NAND U508 ( .A(b[0]), .B(a[85]), .Z(n422) );
  XOR U509 ( .A(sreg[212]), .B(n422), .Z(n424) );
  NANDN U510 ( .A(n417), .B(sreg[211]), .Z(n421) );
  OR U511 ( .A(n419), .B(n418), .Z(n420) );
  AND U512 ( .A(n421), .B(n420), .Z(n423) );
  XOR U513 ( .A(n424), .B(n423), .Z(c[212]) );
  NAND U514 ( .A(b[0]), .B(a[86]), .Z(n427) );
  XOR U515 ( .A(sreg[213]), .B(n427), .Z(n429) );
  NANDN U516 ( .A(n422), .B(sreg[212]), .Z(n426) );
  OR U517 ( .A(n424), .B(n423), .Z(n425) );
  AND U518 ( .A(n426), .B(n425), .Z(n428) );
  XOR U519 ( .A(n429), .B(n428), .Z(c[213]) );
  NAND U520 ( .A(b[0]), .B(a[87]), .Z(n432) );
  XOR U521 ( .A(sreg[214]), .B(n432), .Z(n434) );
  NANDN U522 ( .A(n427), .B(sreg[213]), .Z(n431) );
  OR U523 ( .A(n429), .B(n428), .Z(n430) );
  AND U524 ( .A(n431), .B(n430), .Z(n433) );
  XOR U525 ( .A(n434), .B(n433), .Z(c[214]) );
  NAND U526 ( .A(b[0]), .B(a[88]), .Z(n437) );
  XOR U527 ( .A(sreg[215]), .B(n437), .Z(n439) );
  NANDN U528 ( .A(n432), .B(sreg[214]), .Z(n436) );
  OR U529 ( .A(n434), .B(n433), .Z(n435) );
  AND U530 ( .A(n436), .B(n435), .Z(n438) );
  XOR U531 ( .A(n439), .B(n438), .Z(c[215]) );
  NAND U532 ( .A(b[0]), .B(a[89]), .Z(n442) );
  XOR U533 ( .A(sreg[216]), .B(n442), .Z(n444) );
  NANDN U534 ( .A(n437), .B(sreg[215]), .Z(n441) );
  OR U535 ( .A(n439), .B(n438), .Z(n440) );
  AND U536 ( .A(n441), .B(n440), .Z(n443) );
  XOR U537 ( .A(n444), .B(n443), .Z(c[216]) );
  NAND U538 ( .A(b[0]), .B(a[90]), .Z(n447) );
  XOR U539 ( .A(sreg[217]), .B(n447), .Z(n449) );
  NANDN U540 ( .A(n442), .B(sreg[216]), .Z(n446) );
  OR U541 ( .A(n444), .B(n443), .Z(n445) );
  AND U542 ( .A(n446), .B(n445), .Z(n448) );
  XOR U543 ( .A(n449), .B(n448), .Z(c[217]) );
  NAND U544 ( .A(b[0]), .B(a[91]), .Z(n452) );
  XOR U545 ( .A(sreg[218]), .B(n452), .Z(n454) );
  NANDN U546 ( .A(n447), .B(sreg[217]), .Z(n451) );
  OR U547 ( .A(n449), .B(n448), .Z(n450) );
  AND U548 ( .A(n451), .B(n450), .Z(n453) );
  XOR U549 ( .A(n454), .B(n453), .Z(c[218]) );
  NAND U550 ( .A(b[0]), .B(a[92]), .Z(n457) );
  XOR U551 ( .A(sreg[219]), .B(n457), .Z(n459) );
  NANDN U552 ( .A(n452), .B(sreg[218]), .Z(n456) );
  OR U553 ( .A(n454), .B(n453), .Z(n455) );
  AND U554 ( .A(n456), .B(n455), .Z(n458) );
  XOR U555 ( .A(n459), .B(n458), .Z(c[219]) );
  NAND U556 ( .A(b[0]), .B(a[93]), .Z(n462) );
  XOR U557 ( .A(sreg[220]), .B(n462), .Z(n464) );
  NANDN U558 ( .A(n457), .B(sreg[219]), .Z(n461) );
  OR U559 ( .A(n459), .B(n458), .Z(n460) );
  AND U560 ( .A(n461), .B(n460), .Z(n463) );
  XOR U561 ( .A(n464), .B(n463), .Z(c[220]) );
  NAND U562 ( .A(b[0]), .B(a[94]), .Z(n467) );
  XOR U563 ( .A(sreg[221]), .B(n467), .Z(n469) );
  NANDN U564 ( .A(n462), .B(sreg[220]), .Z(n466) );
  OR U565 ( .A(n464), .B(n463), .Z(n465) );
  AND U566 ( .A(n466), .B(n465), .Z(n468) );
  XOR U567 ( .A(n469), .B(n468), .Z(c[221]) );
  NAND U568 ( .A(b[0]), .B(a[95]), .Z(n472) );
  XOR U569 ( .A(sreg[222]), .B(n472), .Z(n474) );
  NANDN U570 ( .A(n467), .B(sreg[221]), .Z(n471) );
  OR U571 ( .A(n469), .B(n468), .Z(n470) );
  AND U572 ( .A(n471), .B(n470), .Z(n473) );
  XOR U573 ( .A(n474), .B(n473), .Z(c[222]) );
  NAND U574 ( .A(b[0]), .B(a[96]), .Z(n477) );
  XOR U575 ( .A(sreg[223]), .B(n477), .Z(n479) );
  NANDN U576 ( .A(n472), .B(sreg[222]), .Z(n476) );
  OR U577 ( .A(n474), .B(n473), .Z(n475) );
  AND U578 ( .A(n476), .B(n475), .Z(n478) );
  XOR U579 ( .A(n479), .B(n478), .Z(c[223]) );
  NAND U580 ( .A(b[0]), .B(a[97]), .Z(n482) );
  XOR U581 ( .A(sreg[224]), .B(n482), .Z(n484) );
  NANDN U582 ( .A(n477), .B(sreg[223]), .Z(n481) );
  OR U583 ( .A(n479), .B(n478), .Z(n480) );
  AND U584 ( .A(n481), .B(n480), .Z(n483) );
  XOR U585 ( .A(n484), .B(n483), .Z(c[224]) );
  NAND U586 ( .A(b[0]), .B(a[98]), .Z(n487) );
  XOR U587 ( .A(sreg[225]), .B(n487), .Z(n489) );
  NANDN U588 ( .A(n482), .B(sreg[224]), .Z(n486) );
  OR U589 ( .A(n484), .B(n483), .Z(n485) );
  AND U590 ( .A(n486), .B(n485), .Z(n488) );
  XOR U591 ( .A(n489), .B(n488), .Z(c[225]) );
  NAND U592 ( .A(b[0]), .B(a[99]), .Z(n492) );
  XOR U593 ( .A(sreg[226]), .B(n492), .Z(n494) );
  NANDN U594 ( .A(n487), .B(sreg[225]), .Z(n491) );
  OR U595 ( .A(n489), .B(n488), .Z(n490) );
  AND U596 ( .A(n491), .B(n490), .Z(n493) );
  XOR U597 ( .A(n494), .B(n493), .Z(c[226]) );
  NAND U598 ( .A(b[0]), .B(a[100]), .Z(n497) );
  XOR U599 ( .A(sreg[227]), .B(n497), .Z(n499) );
  NANDN U600 ( .A(n492), .B(sreg[226]), .Z(n496) );
  OR U601 ( .A(n494), .B(n493), .Z(n495) );
  AND U602 ( .A(n496), .B(n495), .Z(n498) );
  XOR U603 ( .A(n499), .B(n498), .Z(c[227]) );
  NAND U604 ( .A(b[0]), .B(a[101]), .Z(n502) );
  XOR U605 ( .A(sreg[228]), .B(n502), .Z(n504) );
  NANDN U606 ( .A(n497), .B(sreg[227]), .Z(n501) );
  OR U607 ( .A(n499), .B(n498), .Z(n500) );
  AND U608 ( .A(n501), .B(n500), .Z(n503) );
  XOR U609 ( .A(n504), .B(n503), .Z(c[228]) );
  NAND U610 ( .A(b[0]), .B(a[102]), .Z(n507) );
  XOR U611 ( .A(sreg[229]), .B(n507), .Z(n509) );
  NANDN U612 ( .A(n502), .B(sreg[228]), .Z(n506) );
  OR U613 ( .A(n504), .B(n503), .Z(n505) );
  AND U614 ( .A(n506), .B(n505), .Z(n508) );
  XOR U615 ( .A(n509), .B(n508), .Z(c[229]) );
  NAND U616 ( .A(b[0]), .B(a[103]), .Z(n512) );
  XOR U617 ( .A(sreg[230]), .B(n512), .Z(n514) );
  NANDN U618 ( .A(n507), .B(sreg[229]), .Z(n511) );
  OR U619 ( .A(n509), .B(n508), .Z(n510) );
  AND U620 ( .A(n511), .B(n510), .Z(n513) );
  XOR U621 ( .A(n514), .B(n513), .Z(c[230]) );
  NAND U622 ( .A(b[0]), .B(a[104]), .Z(n517) );
  XOR U623 ( .A(sreg[231]), .B(n517), .Z(n519) );
  NANDN U624 ( .A(n512), .B(sreg[230]), .Z(n516) );
  OR U625 ( .A(n514), .B(n513), .Z(n515) );
  AND U626 ( .A(n516), .B(n515), .Z(n518) );
  XOR U627 ( .A(n519), .B(n518), .Z(c[231]) );
  NAND U628 ( .A(b[0]), .B(a[105]), .Z(n522) );
  XOR U629 ( .A(sreg[232]), .B(n522), .Z(n524) );
  NANDN U630 ( .A(n517), .B(sreg[231]), .Z(n521) );
  OR U631 ( .A(n519), .B(n518), .Z(n520) );
  AND U632 ( .A(n521), .B(n520), .Z(n523) );
  XOR U633 ( .A(n524), .B(n523), .Z(c[232]) );
  NAND U634 ( .A(b[0]), .B(a[106]), .Z(n527) );
  XOR U635 ( .A(sreg[233]), .B(n527), .Z(n529) );
  NANDN U636 ( .A(n522), .B(sreg[232]), .Z(n526) );
  OR U637 ( .A(n524), .B(n523), .Z(n525) );
  AND U638 ( .A(n526), .B(n525), .Z(n528) );
  XOR U639 ( .A(n529), .B(n528), .Z(c[233]) );
  NAND U640 ( .A(b[0]), .B(a[107]), .Z(n532) );
  XOR U641 ( .A(sreg[234]), .B(n532), .Z(n534) );
  NANDN U642 ( .A(n527), .B(sreg[233]), .Z(n531) );
  OR U643 ( .A(n529), .B(n528), .Z(n530) );
  AND U644 ( .A(n531), .B(n530), .Z(n533) );
  XOR U645 ( .A(n534), .B(n533), .Z(c[234]) );
  NAND U646 ( .A(b[0]), .B(a[108]), .Z(n537) );
  XOR U647 ( .A(sreg[235]), .B(n537), .Z(n539) );
  NANDN U648 ( .A(n532), .B(sreg[234]), .Z(n536) );
  OR U649 ( .A(n534), .B(n533), .Z(n535) );
  AND U650 ( .A(n536), .B(n535), .Z(n538) );
  XOR U651 ( .A(n539), .B(n538), .Z(c[235]) );
  NAND U652 ( .A(b[0]), .B(a[109]), .Z(n542) );
  XOR U653 ( .A(sreg[236]), .B(n542), .Z(n544) );
  NANDN U654 ( .A(n537), .B(sreg[235]), .Z(n541) );
  OR U655 ( .A(n539), .B(n538), .Z(n540) );
  AND U656 ( .A(n541), .B(n540), .Z(n543) );
  XOR U657 ( .A(n544), .B(n543), .Z(c[236]) );
  NAND U658 ( .A(b[0]), .B(a[110]), .Z(n547) );
  XOR U659 ( .A(sreg[237]), .B(n547), .Z(n549) );
  NANDN U660 ( .A(n542), .B(sreg[236]), .Z(n546) );
  OR U661 ( .A(n544), .B(n543), .Z(n545) );
  AND U662 ( .A(n546), .B(n545), .Z(n548) );
  XOR U663 ( .A(n549), .B(n548), .Z(c[237]) );
  NAND U664 ( .A(b[0]), .B(a[111]), .Z(n552) );
  XOR U665 ( .A(sreg[238]), .B(n552), .Z(n554) );
  NANDN U666 ( .A(n547), .B(sreg[237]), .Z(n551) );
  OR U667 ( .A(n549), .B(n548), .Z(n550) );
  AND U668 ( .A(n551), .B(n550), .Z(n553) );
  XOR U669 ( .A(n554), .B(n553), .Z(c[238]) );
  NAND U670 ( .A(b[0]), .B(a[112]), .Z(n557) );
  XOR U671 ( .A(sreg[239]), .B(n557), .Z(n559) );
  NANDN U672 ( .A(n552), .B(sreg[238]), .Z(n556) );
  OR U673 ( .A(n554), .B(n553), .Z(n555) );
  AND U674 ( .A(n556), .B(n555), .Z(n558) );
  XOR U675 ( .A(n559), .B(n558), .Z(c[239]) );
  NAND U676 ( .A(b[0]), .B(a[113]), .Z(n562) );
  XOR U677 ( .A(sreg[240]), .B(n562), .Z(n564) );
  NANDN U678 ( .A(n557), .B(sreg[239]), .Z(n561) );
  OR U679 ( .A(n559), .B(n558), .Z(n560) );
  AND U680 ( .A(n561), .B(n560), .Z(n563) );
  XOR U681 ( .A(n564), .B(n563), .Z(c[240]) );
  NAND U682 ( .A(b[0]), .B(a[114]), .Z(n567) );
  XOR U683 ( .A(sreg[241]), .B(n567), .Z(n569) );
  NANDN U684 ( .A(n562), .B(sreg[240]), .Z(n566) );
  OR U685 ( .A(n564), .B(n563), .Z(n565) );
  AND U686 ( .A(n566), .B(n565), .Z(n568) );
  XOR U687 ( .A(n569), .B(n568), .Z(c[241]) );
  NAND U688 ( .A(b[0]), .B(a[115]), .Z(n572) );
  XOR U689 ( .A(sreg[242]), .B(n572), .Z(n574) );
  NANDN U690 ( .A(n567), .B(sreg[241]), .Z(n571) );
  OR U691 ( .A(n569), .B(n568), .Z(n570) );
  AND U692 ( .A(n571), .B(n570), .Z(n573) );
  XOR U693 ( .A(n574), .B(n573), .Z(c[242]) );
  NAND U694 ( .A(b[0]), .B(a[116]), .Z(n577) );
  XOR U695 ( .A(sreg[243]), .B(n577), .Z(n579) );
  NANDN U696 ( .A(n572), .B(sreg[242]), .Z(n576) );
  OR U697 ( .A(n574), .B(n573), .Z(n575) );
  AND U698 ( .A(n576), .B(n575), .Z(n578) );
  XOR U699 ( .A(n579), .B(n578), .Z(c[243]) );
  NAND U700 ( .A(b[0]), .B(a[117]), .Z(n582) );
  XOR U701 ( .A(sreg[244]), .B(n582), .Z(n584) );
  NANDN U702 ( .A(n577), .B(sreg[243]), .Z(n581) );
  OR U703 ( .A(n579), .B(n578), .Z(n580) );
  AND U704 ( .A(n581), .B(n580), .Z(n583) );
  XOR U705 ( .A(n584), .B(n583), .Z(c[244]) );
  NAND U706 ( .A(b[0]), .B(a[118]), .Z(n587) );
  XOR U707 ( .A(sreg[245]), .B(n587), .Z(n589) );
  NANDN U708 ( .A(n582), .B(sreg[244]), .Z(n586) );
  OR U709 ( .A(n584), .B(n583), .Z(n585) );
  AND U710 ( .A(n586), .B(n585), .Z(n588) );
  XOR U711 ( .A(n589), .B(n588), .Z(c[245]) );
  NAND U712 ( .A(b[0]), .B(a[119]), .Z(n592) );
  XOR U713 ( .A(sreg[246]), .B(n592), .Z(n594) );
  NANDN U714 ( .A(n587), .B(sreg[245]), .Z(n591) );
  OR U715 ( .A(n589), .B(n588), .Z(n590) );
  AND U716 ( .A(n591), .B(n590), .Z(n593) );
  XOR U717 ( .A(n594), .B(n593), .Z(c[246]) );
  NAND U718 ( .A(b[0]), .B(a[120]), .Z(n597) );
  XOR U719 ( .A(sreg[247]), .B(n597), .Z(n599) );
  NANDN U720 ( .A(n592), .B(sreg[246]), .Z(n596) );
  OR U721 ( .A(n594), .B(n593), .Z(n595) );
  AND U722 ( .A(n596), .B(n595), .Z(n598) );
  XOR U723 ( .A(n599), .B(n598), .Z(c[247]) );
  NAND U724 ( .A(b[0]), .B(a[121]), .Z(n602) );
  XOR U725 ( .A(sreg[248]), .B(n602), .Z(n604) );
  NANDN U726 ( .A(n597), .B(sreg[247]), .Z(n601) );
  OR U727 ( .A(n599), .B(n598), .Z(n600) );
  AND U728 ( .A(n601), .B(n600), .Z(n603) );
  XOR U729 ( .A(n604), .B(n603), .Z(c[248]) );
  NAND U730 ( .A(b[0]), .B(a[122]), .Z(n607) );
  XOR U731 ( .A(sreg[249]), .B(n607), .Z(n609) );
  NANDN U732 ( .A(n602), .B(sreg[248]), .Z(n606) );
  OR U733 ( .A(n604), .B(n603), .Z(n605) );
  AND U734 ( .A(n606), .B(n605), .Z(n608) );
  XOR U735 ( .A(n609), .B(n608), .Z(c[249]) );
  NAND U736 ( .A(b[0]), .B(a[123]), .Z(n612) );
  XOR U737 ( .A(sreg[250]), .B(n612), .Z(n614) );
  NANDN U738 ( .A(n607), .B(sreg[249]), .Z(n611) );
  OR U739 ( .A(n609), .B(n608), .Z(n610) );
  AND U740 ( .A(n611), .B(n610), .Z(n613) );
  XOR U741 ( .A(n614), .B(n613), .Z(c[250]) );
  NAND U742 ( .A(b[0]), .B(a[124]), .Z(n617) );
  XOR U743 ( .A(sreg[251]), .B(n617), .Z(n619) );
  NANDN U744 ( .A(n612), .B(sreg[250]), .Z(n616) );
  OR U745 ( .A(n614), .B(n613), .Z(n615) );
  AND U746 ( .A(n616), .B(n615), .Z(n618) );
  XOR U747 ( .A(n619), .B(n618), .Z(c[251]) );
  NAND U748 ( .A(b[0]), .B(a[125]), .Z(n622) );
  XOR U749 ( .A(sreg[252]), .B(n622), .Z(n624) );
  NANDN U750 ( .A(n617), .B(sreg[251]), .Z(n621) );
  OR U751 ( .A(n619), .B(n618), .Z(n620) );
  AND U752 ( .A(n621), .B(n620), .Z(n623) );
  XOR U753 ( .A(n624), .B(n623), .Z(c[252]) );
  NAND U754 ( .A(b[0]), .B(a[126]), .Z(n627) );
  XOR U755 ( .A(sreg[253]), .B(n627), .Z(n629) );
  NANDN U756 ( .A(n622), .B(sreg[252]), .Z(n626) );
  OR U757 ( .A(n624), .B(n623), .Z(n625) );
  AND U758 ( .A(n626), .B(n625), .Z(n628) );
  XOR U759 ( .A(n629), .B(n628), .Z(c[253]) );
  NANDN U760 ( .A(n627), .B(sreg[253]), .Z(n631) );
  OR U761 ( .A(n629), .B(n628), .Z(n630) );
  AND U762 ( .A(n631), .B(n630), .Z(n635) );
  AND U763 ( .A(a[127]), .B(b[0]), .Z(n633) );
  XNOR U764 ( .A(sreg[254]), .B(n633), .Z(n632) );
  XOR U765 ( .A(n635), .B(n632), .Z(c[254]) );
  NAND U766 ( .A(sreg[254]), .B(n633), .Z(n637) );
  XOR U767 ( .A(n633), .B(sreg[254]), .Z(n634) );
  NANDN U768 ( .A(n635), .B(n634), .Z(n636) );
  NAND U769 ( .A(n637), .B(n636), .Z(c[255]) );
endmodule

