
module hamming_N1600_CC1 ( clk, rst, x, y, o );
  input [1599:0] x;
  input [1599:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569;

  NANDN U1601 ( .A(n929), .B(n928), .Z(n1) );
  NANDN U1602 ( .A(n927), .B(n926), .Z(n2) );
  AND U1603 ( .A(n1), .B(n2), .Z(n5384) );
  NANDN U1604 ( .A(n3832), .B(n3831), .Z(n3) );
  NANDN U1605 ( .A(n3834), .B(n3833), .Z(n4) );
  NAND U1606 ( .A(n3), .B(n4), .Z(n6114) );
  NANDN U1607 ( .A(n3253), .B(n3252), .Z(n5) );
  NANDN U1608 ( .A(n3255), .B(n3254), .Z(n6) );
  NAND U1609 ( .A(n5), .B(n6), .Z(n5754) );
  NANDN U1610 ( .A(n3273), .B(n3272), .Z(n7) );
  NANDN U1611 ( .A(n3275), .B(n3274), .Z(n8) );
  NAND U1612 ( .A(n7), .B(n8), .Z(n5743) );
  NANDN U1613 ( .A(n1139), .B(n1138), .Z(n9) );
  NANDN U1614 ( .A(n1141), .B(n1140), .Z(n10) );
  NAND U1615 ( .A(n9), .B(n10), .Z(n6025) );
  NANDN U1616 ( .A(n853), .B(n852), .Z(n11) );
  NANDN U1617 ( .A(n855), .B(n854), .Z(n12) );
  NAND U1618 ( .A(n11), .B(n12), .Z(n6019) );
  NANDN U1619 ( .A(n2855), .B(n2854), .Z(n13) );
  NANDN U1620 ( .A(n2857), .B(n2856), .Z(n14) );
  NAND U1621 ( .A(n13), .B(n14), .Z(n7059) );
  NANDN U1622 ( .A(n2769), .B(n2768), .Z(n15) );
  NANDN U1623 ( .A(n2771), .B(n2770), .Z(n16) );
  NAND U1624 ( .A(n15), .B(n16), .Z(n7065) );
  NANDN U1625 ( .A(n3887), .B(n3886), .Z(n17) );
  NANDN U1626 ( .A(n3889), .B(n3888), .Z(n18) );
  NAND U1627 ( .A(n17), .B(n18), .Z(n7028) );
  NANDN U1628 ( .A(n3869), .B(n3868), .Z(n19) );
  NANDN U1629 ( .A(n3871), .B(n3870), .Z(n20) );
  NAND U1630 ( .A(n19), .B(n20), .Z(n6612) );
  NANDN U1631 ( .A(n891), .B(n890), .Z(n21) );
  NANDN U1632 ( .A(n893), .B(n892), .Z(n22) );
  NAND U1633 ( .A(n21), .B(n22), .Z(n5977) );
  NANDN U1634 ( .A(n3145), .B(n3144), .Z(n23) );
  NANDN U1635 ( .A(n3147), .B(n3146), .Z(n24) );
  NAND U1636 ( .A(n23), .B(n24), .Z(n5328) );
  NANDN U1637 ( .A(n1205), .B(n1204), .Z(n25) );
  NANDN U1638 ( .A(n1207), .B(n1206), .Z(n26) );
  NAND U1639 ( .A(n25), .B(n26), .Z(n6077) );
  NANDN U1640 ( .A(n2879), .B(n2878), .Z(n27) );
  NANDN U1641 ( .A(n2881), .B(n2880), .Z(n28) );
  NAND U1642 ( .A(n27), .B(n28), .Z(n6655) );
  NANDN U1643 ( .A(n4293), .B(n4292), .Z(n29) );
  NANDN U1644 ( .A(n4295), .B(n4294), .Z(n30) );
  NAND U1645 ( .A(n29), .B(n30), .Z(n6485) );
  NANDN U1646 ( .A(n5519), .B(n5518), .Z(n31) );
  NANDN U1647 ( .A(n5521), .B(n5520), .Z(n32) );
  NAND U1648 ( .A(n31), .B(n32), .Z(n8409) );
  XOR U1649 ( .A(n1010), .B(n1011), .Z(n1012) );
  XOR U1650 ( .A(n2076), .B(n2077), .Z(n2078) );
  NANDN U1651 ( .A(n3314), .B(n3313), .Z(n33) );
  NANDN U1652 ( .A(n3316), .B(n3315), .Z(n34) );
  NAND U1653 ( .A(n33), .B(n34), .Z(n6239) );
  NANDN U1654 ( .A(n1725), .B(n1724), .Z(n35) );
  NANDN U1655 ( .A(n1727), .B(n1726), .Z(n36) );
  NAND U1656 ( .A(n35), .B(n36), .Z(n5310) );
  NANDN U1657 ( .A(n4715), .B(n4714), .Z(n37) );
  NANDN U1658 ( .A(n4717), .B(n4716), .Z(n38) );
  NAND U1659 ( .A(n37), .B(n38), .Z(n5444) );
  NANDN U1660 ( .A(n933), .B(n932), .Z(n39) );
  NANDN U1661 ( .A(n931), .B(n930), .Z(n40) );
  AND U1662 ( .A(n39), .B(n40), .Z(n5385) );
  NANDN U1663 ( .A(n3843), .B(n3842), .Z(n41) );
  NANDN U1664 ( .A(n3845), .B(n3844), .Z(n42) );
  NAND U1665 ( .A(n41), .B(n42), .Z(n6116) );
  NANDN U1666 ( .A(n3249), .B(n3248), .Z(n43) );
  NANDN U1667 ( .A(n3251), .B(n3250), .Z(n44) );
  NAND U1668 ( .A(n43), .B(n44), .Z(n5755) );
  NANDN U1669 ( .A(n3284), .B(n3283), .Z(n45) );
  NANDN U1670 ( .A(n3286), .B(n3285), .Z(n46) );
  NAND U1671 ( .A(n45), .B(n46), .Z(n5745) );
  NANDN U1672 ( .A(n1135), .B(n1134), .Z(n47) );
  NANDN U1673 ( .A(n1137), .B(n1136), .Z(n48) );
  NAND U1674 ( .A(n47), .B(n48), .Z(n6026) );
  NANDN U1675 ( .A(n849), .B(n848), .Z(n49) );
  NANDN U1676 ( .A(n851), .B(n850), .Z(n50) );
  NAND U1677 ( .A(n49), .B(n50), .Z(n6020) );
  NANDN U1678 ( .A(n2851), .B(n2850), .Z(n51) );
  NANDN U1679 ( .A(n2853), .B(n2852), .Z(n52) );
  NAND U1680 ( .A(n51), .B(n52), .Z(n7060) );
  NANDN U1681 ( .A(n2765), .B(n2764), .Z(n53) );
  NANDN U1682 ( .A(n2767), .B(n2766), .Z(n54) );
  NAND U1683 ( .A(n53), .B(n54), .Z(n7066) );
  NANDN U1684 ( .A(n3883), .B(n3882), .Z(n55) );
  NANDN U1685 ( .A(n3885), .B(n3884), .Z(n56) );
  NAND U1686 ( .A(n55), .B(n56), .Z(n7029) );
  NANDN U1687 ( .A(n3865), .B(n3864), .Z(n57) );
  NANDN U1688 ( .A(n3867), .B(n3866), .Z(n58) );
  NAND U1689 ( .A(n57), .B(n58), .Z(n6613) );
  NANDN U1690 ( .A(n2891), .B(n2890), .Z(n59) );
  NANDN U1691 ( .A(n2893), .B(n2892), .Z(n60) );
  NAND U1692 ( .A(n59), .B(n60), .Z(n6570) );
  NANDN U1693 ( .A(n1005), .B(n1004), .Z(n61) );
  NANDN U1694 ( .A(n1003), .B(n1002), .Z(n62) );
  AND U1695 ( .A(n61), .B(n62), .Z(n5564) );
  NANDN U1696 ( .A(n1109), .B(n1108), .Z(n63) );
  NANDN U1697 ( .A(n1111), .B(n1110), .Z(n64) );
  NAND U1698 ( .A(n63), .B(n64), .Z(n5612) );
  NANDN U1699 ( .A(n903), .B(n902), .Z(n65) );
  NANDN U1700 ( .A(n905), .B(n904), .Z(n66) );
  NAND U1701 ( .A(n65), .B(n66), .Z(n5606) );
  NANDN U1702 ( .A(n915), .B(n914), .Z(n67) );
  NANDN U1703 ( .A(n917), .B(n916), .Z(n68) );
  NAND U1704 ( .A(n67), .B(n68), .Z(n5989) );
  NANDN U1705 ( .A(n887), .B(n886), .Z(n69) );
  NANDN U1706 ( .A(n889), .B(n888), .Z(n70) );
  NAND U1707 ( .A(n69), .B(n70), .Z(n5978) );
  NANDN U1708 ( .A(n3141), .B(n3140), .Z(n71) );
  NANDN U1709 ( .A(n3143), .B(n3142), .Z(n72) );
  NAND U1710 ( .A(n71), .B(n72), .Z(n5329) );
  NANDN U1711 ( .A(n1587), .B(n1586), .Z(n73) );
  NANDN U1712 ( .A(n1585), .B(n1584), .Z(n74) );
  AND U1713 ( .A(n73), .B(n74), .Z(n5334) );
  NANDN U1714 ( .A(n3512), .B(n3511), .Z(n75) );
  NANDN U1715 ( .A(n3514), .B(n3513), .Z(n76) );
  NAND U1716 ( .A(n75), .B(n76), .Z(n6126) );
  NANDN U1717 ( .A(n1201), .B(n1200), .Z(n77) );
  NANDN U1718 ( .A(n1203), .B(n1202), .Z(n78) );
  NAND U1719 ( .A(n77), .B(n78), .Z(n6078) );
  NANDN U1720 ( .A(n2947), .B(n2946), .Z(n79) );
  NANDN U1721 ( .A(n2949), .B(n2948), .Z(n80) );
  NAND U1722 ( .A(n79), .B(n80), .Z(n6667) );
  NANDN U1723 ( .A(n2883), .B(n2882), .Z(n81) );
  NANDN U1724 ( .A(n2885), .B(n2884), .Z(n82) );
  NAND U1725 ( .A(n81), .B(n82), .Z(n6658) );
  NANDN U1726 ( .A(n1777), .B(n1776), .Z(n83) );
  NANDN U1727 ( .A(n1775), .B(n1774), .Z(n84) );
  AND U1728 ( .A(n83), .B(n84), .Z(n5232) );
  XNOR U1729 ( .A(n5597), .B(n5596), .Z(n7146) );
  NANDN U1730 ( .A(n4217), .B(n4216), .Z(n85) );
  NANDN U1731 ( .A(n4219), .B(n4218), .Z(n86) );
  NAND U1732 ( .A(n85), .B(n86), .Z(n6185) );
  NANDN U1733 ( .A(n4687), .B(n4686), .Z(n87) );
  NANDN U1734 ( .A(n4685), .B(n4684), .Z(n88) );
  AND U1735 ( .A(n87), .B(n88), .Z(n6149) );
  NANDN U1736 ( .A(n4865), .B(n4864), .Z(n89) );
  NANDN U1737 ( .A(n4863), .B(n4862), .Z(n90) );
  AND U1738 ( .A(n89), .B(n90), .Z(n6155) );
  NANDN U1739 ( .A(n4281), .B(n4280), .Z(n91) );
  NANDN U1740 ( .A(n4283), .B(n4282), .Z(n92) );
  NAND U1741 ( .A(n91), .B(n92), .Z(n6491) );
  NANDN U1742 ( .A(n4289), .B(n4288), .Z(n93) );
  NANDN U1743 ( .A(n4291), .B(n4290), .Z(n94) );
  NAND U1744 ( .A(n93), .B(n94), .Z(n6486) );
  NANDN U1745 ( .A(n4229), .B(n4228), .Z(n95) );
  NANDN U1746 ( .A(n4231), .B(n4230), .Z(n96) );
  NAND U1747 ( .A(n95), .B(n96), .Z(n6063) );
  NANDN U1748 ( .A(n2255), .B(n2254), .Z(n97) );
  NANDN U1749 ( .A(n2253), .B(n2252), .Z(n98) );
  AND U1750 ( .A(n97), .B(n98), .Z(n6059) );
  NANDN U1751 ( .A(n2167), .B(n2166), .Z(n99) );
  NANDN U1752 ( .A(n2169), .B(n2168), .Z(n100) );
  NAND U1753 ( .A(n99), .B(n100), .Z(n6056) );
  NANDN U1754 ( .A(n2415), .B(n2414), .Z(n101) );
  NANDN U1755 ( .A(n2413), .B(n2412), .Z(n102) );
  AND U1756 ( .A(n101), .B(n102), .Z(n5510) );
  NANDN U1757 ( .A(n5515), .B(n5514), .Z(n103) );
  NANDN U1758 ( .A(n5517), .B(n5516), .Z(n104) );
  NAND U1759 ( .A(n103), .B(n104), .Z(n8408) );
  XNOR U1760 ( .A(n9004), .B(n9005), .Z(n9007) );
  NAND U1761 ( .A(n7895), .B(n7894), .Z(n105) );
  NANDN U1762 ( .A(n7897), .B(n7896), .Z(n106) );
  NAND U1763 ( .A(n105), .B(n106), .Z(n8739) );
  XNOR U1764 ( .A(n9353), .B(n9354), .Z(n9356) );
  NAND U1765 ( .A(n9537), .B(n9538), .Z(n107) );
  NANDN U1766 ( .A(n9536), .B(n9535), .Z(n108) );
  NAND U1767 ( .A(n107), .B(n108), .Z(n9558) );
  XNOR U1768 ( .A(n2829), .B(n2828), .Z(n1482) );
  XNOR U1769 ( .A(n4042), .B(n4043), .Z(n4045) );
  XNOR U1770 ( .A(n3922), .B(n3923), .Z(n3925) );
  NANDN U1771 ( .A(n4925), .B(n4924), .Z(n109) );
  NANDN U1772 ( .A(n4927), .B(n4926), .Z(n110) );
  NAND U1773 ( .A(n109), .B(n110), .Z(n6254) );
  NANDN U1774 ( .A(n3310), .B(n3309), .Z(n111) );
  NANDN U1775 ( .A(n3312), .B(n3311), .Z(n112) );
  NAND U1776 ( .A(n111), .B(n112), .Z(n6240) );
  NANDN U1777 ( .A(n1721), .B(n1720), .Z(n113) );
  NANDN U1778 ( .A(n1723), .B(n1722), .Z(n114) );
  NAND U1779 ( .A(n113), .B(n114), .Z(n5311) );
  NANDN U1780 ( .A(n4711), .B(n4710), .Z(n115) );
  NANDN U1781 ( .A(n4713), .B(n4712), .Z(n116) );
  NAND U1782 ( .A(n115), .B(n116), .Z(n5445) );
  NANDN U1783 ( .A(n3025), .B(n3024), .Z(n117) );
  NANDN U1784 ( .A(n3023), .B(n3022), .Z(n118) );
  AND U1785 ( .A(n117), .B(n118), .Z(n5450) );
  NANDN U1786 ( .A(n1877), .B(n1876), .Z(n119) );
  NANDN U1787 ( .A(n1875), .B(n1874), .Z(n120) );
  AND U1788 ( .A(n119), .B(n120), .Z(n5396) );
  NAND U1789 ( .A(n924), .B(n925), .Z(n121) );
  NANDN U1790 ( .A(n923), .B(n922), .Z(n122) );
  NAND U1791 ( .A(n121), .B(n122), .Z(n5387) );
  NANDN U1792 ( .A(n879), .B(n878), .Z(n123) );
  NANDN U1793 ( .A(n881), .B(n880), .Z(n124) );
  NAND U1794 ( .A(n123), .B(n124), .Z(n5492) );
  NANDN U1795 ( .A(n3215), .B(n3214), .Z(n125) );
  NANDN U1796 ( .A(n3217), .B(n3216), .Z(n126) );
  NAND U1797 ( .A(n125), .B(n126), .Z(n5486) );
  XOR U1798 ( .A(n6113), .B(n6114), .Z(n6115) );
  NANDN U1799 ( .A(n3772), .B(n3771), .Z(n127) );
  NANDN U1800 ( .A(n3774), .B(n3773), .Z(n128) );
  NAND U1801 ( .A(n127), .B(n128), .Z(n6546) );
  NANDN U1802 ( .A(n1381), .B(n1380), .Z(n129) );
  NANDN U1803 ( .A(n1383), .B(n1382), .Z(n130) );
  NAND U1804 ( .A(n129), .B(n130), .Z(n6540) );
  NANDN U1805 ( .A(n1715), .B(n1714), .Z(n131) );
  NANDN U1806 ( .A(n1713), .B(n1712), .Z(n132) );
  AND U1807 ( .A(n131), .B(n132), .Z(n6293) );
  NANDN U1808 ( .A(n4129), .B(n4128), .Z(n133) );
  NANDN U1809 ( .A(n4127), .B(n4126), .Z(n134) );
  AND U1810 ( .A(n133), .B(n134), .Z(n6287) );
  NANDN U1811 ( .A(n3338), .B(n3337), .Z(n135) );
  NANDN U1812 ( .A(n3340), .B(n3339), .Z(n136) );
  NAND U1813 ( .A(n135), .B(n136), .Z(n5346) );
  NANDN U1814 ( .A(n3257), .B(n3256), .Z(n137) );
  NANDN U1815 ( .A(n3259), .B(n3258), .Z(n138) );
  NAND U1816 ( .A(n137), .B(n138), .Z(n5757) );
  XOR U1817 ( .A(n5742), .B(n5743), .Z(n5744) );
  NANDN U1818 ( .A(n1143), .B(n1142), .Z(n139) );
  NANDN U1819 ( .A(n1145), .B(n1144), .Z(n140) );
  NAND U1820 ( .A(n139), .B(n140), .Z(n6028) );
  NANDN U1821 ( .A(n857), .B(n856), .Z(n141) );
  NANDN U1822 ( .A(n859), .B(n858), .Z(n142) );
  NAND U1823 ( .A(n141), .B(n142), .Z(n6022) );
  XOR U1824 ( .A(n7059), .B(n7060), .Z(n7061) );
  NANDN U1825 ( .A(n2773), .B(n2772), .Z(n143) );
  NANDN U1826 ( .A(n2775), .B(n2774), .Z(n144) );
  NAND U1827 ( .A(n143), .B(n144), .Z(n7068) );
  NANDN U1828 ( .A(n3622), .B(n3621), .Z(n145) );
  NANDN U1829 ( .A(n3624), .B(n3623), .Z(n146) );
  NAND U1830 ( .A(n145), .B(n146), .Z(n7017) );
  NANDN U1831 ( .A(n3891), .B(n3890), .Z(n147) );
  NANDN U1832 ( .A(n3893), .B(n3892), .Z(n148) );
  NAND U1833 ( .A(n147), .B(n148), .Z(n7031) );
  NANDN U1834 ( .A(n3941), .B(n3940), .Z(n149) );
  NANDN U1835 ( .A(n3939), .B(n3938), .Z(n150) );
  AND U1836 ( .A(n149), .B(n150), .Z(n7053) );
  NANDN U1837 ( .A(n3107), .B(n3106), .Z(n151) );
  NANDN U1838 ( .A(n3109), .B(n3108), .Z(n152) );
  NAND U1839 ( .A(n151), .B(n152), .Z(n5293) );
  NANDN U1840 ( .A(n1573), .B(n1572), .Z(n153) );
  NANDN U1841 ( .A(n1571), .B(n1570), .Z(n154) );
  AND U1842 ( .A(n153), .B(n154), .Z(n5298) );
  NANDN U1843 ( .A(n3873), .B(n3872), .Z(n155) );
  NANDN U1844 ( .A(n3875), .B(n3874), .Z(n156) );
  NAND U1845 ( .A(n155), .B(n156), .Z(n6615) );
  NANDN U1846 ( .A(n2887), .B(n2886), .Z(n157) );
  NANDN U1847 ( .A(n2889), .B(n2888), .Z(n158) );
  NAND U1848 ( .A(n157), .B(n158), .Z(n6571) );
  NANDN U1849 ( .A(n2025), .B(n2024), .Z(n159) );
  NANDN U1850 ( .A(n2023), .B(n2022), .Z(n160) );
  AND U1851 ( .A(n159), .B(n160), .Z(n6377) );
  NANDN U1852 ( .A(n3786), .B(n3785), .Z(n161) );
  NANDN U1853 ( .A(n3784), .B(n3783), .Z(n162) );
  AND U1854 ( .A(n161), .B(n162), .Z(n6365) );
  NANDN U1855 ( .A(n3760), .B(n3759), .Z(n163) );
  NANDN U1856 ( .A(n3758), .B(n3757), .Z(n164) );
  AND U1857 ( .A(n163), .B(n164), .Z(n6395) );
  NANDN U1858 ( .A(n2273), .B(n2272), .Z(n165) );
  NANDN U1859 ( .A(n2271), .B(n2270), .Z(n166) );
  AND U1860 ( .A(n165), .B(n166), .Z(n6389) );
  NANDN U1861 ( .A(n999), .B(n998), .Z(n167) );
  NANDN U1862 ( .A(n1001), .B(n1000), .Z(n168) );
  NAND U1863 ( .A(n167), .B(n168), .Z(n5565) );
  NANDN U1864 ( .A(n1105), .B(n1104), .Z(n169) );
  NANDN U1865 ( .A(n1107), .B(n1106), .Z(n170) );
  NAND U1866 ( .A(n169), .B(n170), .Z(n5613) );
  NANDN U1867 ( .A(n907), .B(n906), .Z(n171) );
  NANDN U1868 ( .A(n909), .B(n908), .Z(n172) );
  NAND U1869 ( .A(n171), .B(n172), .Z(n5609) );
  NANDN U1870 ( .A(n1017), .B(n1016), .Z(n173) );
  NANDN U1871 ( .A(n1019), .B(n1018), .Z(n174) );
  NAND U1872 ( .A(n173), .B(n174), .Z(n5601) );
  NANDN U1873 ( .A(n911), .B(n910), .Z(n175) );
  NANDN U1874 ( .A(n913), .B(n912), .Z(n176) );
  NAND U1875 ( .A(n175), .B(n176), .Z(n5990) );
  XOR U1876 ( .A(n5977), .B(n5978), .Z(n5979) );
  NANDN U1877 ( .A(n3428), .B(n3427), .Z(n177) );
  NANDN U1878 ( .A(n3426), .B(n3425), .Z(n178) );
  AND U1879 ( .A(n177), .B(n178), .Z(n5959) );
  NANDN U1880 ( .A(n1397), .B(n1396), .Z(n179) );
  NANDN U1881 ( .A(n1395), .B(n1394), .Z(n180) );
  AND U1882 ( .A(n179), .B(n180), .Z(n7236) );
  NANDN U1883 ( .A(n1963), .B(n1962), .Z(n181) );
  NANDN U1884 ( .A(n1965), .B(n1964), .Z(n182) );
  NAND U1885 ( .A(n181), .B(n182), .Z(n7230) );
  NANDN U1886 ( .A(n4003), .B(n4002), .Z(n183) );
  NANDN U1887 ( .A(n4005), .B(n4004), .Z(n184) );
  NAND U1888 ( .A(n183), .B(n184), .Z(n7224) );
  NANDN U1889 ( .A(n2789), .B(n2788), .Z(n185) );
  NANDN U1890 ( .A(n2791), .B(n2790), .Z(n186) );
  NAND U1891 ( .A(n185), .B(n186), .Z(n6980) );
  NANDN U1892 ( .A(n3810), .B(n3809), .Z(n187) );
  NANDN U1893 ( .A(n3812), .B(n3811), .Z(n188) );
  NAND U1894 ( .A(n187), .B(n188), .Z(n6975) );
  XOR U1895 ( .A(n5328), .B(n5329), .Z(n5330) );
  NANDN U1896 ( .A(n1581), .B(n1580), .Z(n189) );
  NANDN U1897 ( .A(n1583), .B(n1582), .Z(n190) );
  NAND U1898 ( .A(n189), .B(n190), .Z(n5335) );
  NANDN U1899 ( .A(n3522), .B(n3521), .Z(n191) );
  NANDN U1900 ( .A(n3524), .B(n3523), .Z(n192) );
  NAND U1901 ( .A(n191), .B(n192), .Z(n6128) );
  NANDN U1902 ( .A(n2397), .B(n2396), .Z(n193) );
  NANDN U1903 ( .A(n2395), .B(n2394), .Z(n194) );
  AND U1904 ( .A(n193), .B(n194), .Z(n6131) );
  NANDN U1905 ( .A(n3917), .B(n3916), .Z(n195) );
  NANDN U1906 ( .A(n3915), .B(n3914), .Z(n196) );
  AND U1907 ( .A(n195), .B(n196), .Z(n6119) );
  NANDN U1908 ( .A(n2427), .B(n2426), .Z(n197) );
  NANDN U1909 ( .A(n2425), .B(n2424), .Z(n198) );
  AND U1910 ( .A(n197), .B(n198), .Z(n6644) );
  NANDN U1911 ( .A(n2487), .B(n2486), .Z(n199) );
  NANDN U1912 ( .A(n2489), .B(n2488), .Z(n200) );
  NAND U1913 ( .A(n199), .B(n200), .Z(n5541) );
  NANDN U1914 ( .A(n1829), .B(n1828), .Z(n201) );
  NANDN U1915 ( .A(n1827), .B(n1826), .Z(n202) );
  AND U1916 ( .A(n201), .B(n202), .Z(n6159) );
  NANDN U1917 ( .A(n4335), .B(n4334), .Z(n203) );
  NANDN U1918 ( .A(n4333), .B(n4332), .Z(n204) );
  AND U1919 ( .A(n203), .B(n204), .Z(n6461) );
  NANDN U1920 ( .A(n2355), .B(n2354), .Z(n205) );
  NANDN U1921 ( .A(n2353), .B(n2352), .Z(n206) );
  AND U1922 ( .A(n205), .B(n206), .Z(n6468) );
  NANDN U1923 ( .A(n4357), .B(n4356), .Z(n207) );
  NANDN U1924 ( .A(n4355), .B(n4354), .Z(n208) );
  AND U1925 ( .A(n207), .B(n208), .Z(n6426) );
  NANDN U1926 ( .A(n2305), .B(n2304), .Z(n209) );
  NANDN U1927 ( .A(n2303), .B(n2302), .Z(n210) );
  AND U1928 ( .A(n209), .B(n210), .Z(n6419) );
  NANDN U1929 ( .A(n2343), .B(n2342), .Z(n211) );
  NANDN U1930 ( .A(n2341), .B(n2340), .Z(n212) );
  AND U1931 ( .A(n211), .B(n212), .Z(n6432) );
  NANDN U1932 ( .A(n4675), .B(n4674), .Z(n213) );
  NANDN U1933 ( .A(n4673), .B(n4672), .Z(n214) );
  AND U1934 ( .A(n213), .B(n214), .Z(n6179) );
  NANDN U1935 ( .A(n2239), .B(n2238), .Z(n215) );
  NANDN U1936 ( .A(n2237), .B(n2236), .Z(n216) );
  AND U1937 ( .A(n215), .B(n216), .Z(n6089) );
  NANDN U1938 ( .A(n1853), .B(n1852), .Z(n217) );
  NANDN U1939 ( .A(n1851), .B(n1850), .Z(n218) );
  AND U1940 ( .A(n217), .B(n218), .Z(n6083) );
  XOR U1941 ( .A(n6077), .B(n6078), .Z(n6079) );
  NANDN U1942 ( .A(n2951), .B(n2950), .Z(n219) );
  NANDN U1943 ( .A(n2953), .B(n2952), .Z(n220) );
  NAND U1944 ( .A(n219), .B(n220), .Z(n6670) );
  NANDN U1945 ( .A(n4787), .B(n4786), .Z(n221) );
  NANDN U1946 ( .A(n4785), .B(n4784), .Z(n222) );
  AND U1947 ( .A(n221), .B(n222), .Z(n6269) );
  NANDN U1948 ( .A(n3548), .B(n3547), .Z(n223) );
  NANDN U1949 ( .A(n3550), .B(n3549), .Z(n224) );
  NAND U1950 ( .A(n223), .B(n224), .Z(n5888) );
  NANDN U1951 ( .A(n4815), .B(n4814), .Z(n225) );
  NANDN U1952 ( .A(n4817), .B(n4816), .Z(n226) );
  NAND U1953 ( .A(n225), .B(n226), .Z(n5936) );
  NANDN U1954 ( .A(n3372), .B(n3371), .Z(n227) );
  NANDN U1955 ( .A(n3374), .B(n3373), .Z(n228) );
  NAND U1956 ( .A(n227), .B(n228), .Z(n5929) );
  NANDN U1957 ( .A(n2291), .B(n2290), .Z(n229) );
  NANDN U1958 ( .A(n2289), .B(n2288), .Z(n230) );
  AND U1959 ( .A(n229), .B(n230), .Z(n7004) );
  NANDN U1960 ( .A(n2325), .B(n2324), .Z(n231) );
  NANDN U1961 ( .A(n2323), .B(n2322), .Z(n232) );
  AND U1962 ( .A(n231), .B(n232), .Z(n7010) );
  NANDN U1963 ( .A(n1981), .B(n1980), .Z(n233) );
  NANDN U1964 ( .A(n1979), .B(n1978), .Z(n234) );
  AND U1965 ( .A(n233), .B(n234), .Z(n6998) );
  NANDN U1966 ( .A(n4935), .B(n4934), .Z(n235) );
  NANDN U1967 ( .A(n4933), .B(n4932), .Z(n236) );
  AND U1968 ( .A(n235), .B(n236), .Z(n5244) );
  NANDN U1969 ( .A(n1779), .B(n1778), .Z(n237) );
  NANDN U1970 ( .A(n1781), .B(n1780), .Z(n238) );
  NAND U1971 ( .A(n237), .B(n238), .Z(n5235) );
  NANDN U1972 ( .A(n2737), .B(n2736), .Z(n239) );
  NANDN U1973 ( .A(n2735), .B(n2734), .Z(n240) );
  AND U1974 ( .A(n239), .B(n240), .Z(n5164) );
  NANDN U1975 ( .A(n2703), .B(n2702), .Z(n241) );
  NANDN U1976 ( .A(n2701), .B(n2700), .Z(n242) );
  AND U1977 ( .A(n241), .B(n242), .Z(n5158) );
  NANDN U1978 ( .A(n1913), .B(n1912), .Z(n243) );
  NANDN U1979 ( .A(n1911), .B(n1910), .Z(n244) );
  AND U1980 ( .A(n243), .B(n244), .Z(n5268) );
  NANDN U1981 ( .A(n1081), .B(n1080), .Z(n245) );
  NANDN U1982 ( .A(n1079), .B(n1078), .Z(n246) );
  AND U1983 ( .A(n245), .B(n246), .Z(n5256) );
  NANDN U1984 ( .A(n1901), .B(n1900), .Z(n247) );
  NANDN U1985 ( .A(n1899), .B(n1898), .Z(n248) );
  AND U1986 ( .A(n247), .B(n248), .Z(n5785) );
  NANDN U1987 ( .A(n867), .B(n866), .Z(n249) );
  NANDN U1988 ( .A(n865), .B(n864), .Z(n250) );
  AND U1989 ( .A(n249), .B(n250), .Z(n5779) );
  NANDN U1990 ( .A(n2011), .B(n2010), .Z(n251) );
  NANDN U1991 ( .A(n2013), .B(n2012), .Z(n252) );
  NAND U1992 ( .A(n251), .B(n252), .Z(n6335) );
  NANDN U1993 ( .A(n993), .B(n992), .Z(n253) );
  NANDN U1994 ( .A(n991), .B(n990), .Z(n254) );
  AND U1995 ( .A(n253), .B(n254), .Z(n5576) );
  NANDN U1996 ( .A(n4441), .B(n4440), .Z(n255) );
  NANDN U1997 ( .A(n4439), .B(n4438), .Z(n256) );
  AND U1998 ( .A(n255), .B(n256), .Z(n5869) );
  XOR U1999 ( .A(n6922), .B(n6923), .Z(n6924) );
  NAND U2000 ( .A(n2258), .B(n2259), .Z(n257) );
  NANDN U2001 ( .A(n2257), .B(n2256), .Z(n258) );
  NAND U2002 ( .A(n257), .B(n258), .Z(n6511) );
  NANDN U2003 ( .A(n4213), .B(n4212), .Z(n259) );
  NANDN U2004 ( .A(n4215), .B(n4214), .Z(n260) );
  NAND U2005 ( .A(n259), .B(n260), .Z(n6186) );
  NANDN U2006 ( .A(n4681), .B(n4680), .Z(n261) );
  NANDN U2007 ( .A(n4683), .B(n4682), .Z(n262) );
  NAND U2008 ( .A(n261), .B(n262), .Z(n6150) );
  NANDN U2009 ( .A(n4277), .B(n4276), .Z(n263) );
  NANDN U2010 ( .A(n4279), .B(n4278), .Z(n264) );
  NAND U2011 ( .A(n263), .B(n264), .Z(n6492) );
  NANDN U2012 ( .A(n4297), .B(n4296), .Z(n265) );
  NANDN U2013 ( .A(n4299), .B(n4298), .Z(n266) );
  NAND U2014 ( .A(n265), .B(n266), .Z(n6488) );
  NANDN U2015 ( .A(n4225), .B(n4224), .Z(n267) );
  NANDN U2016 ( .A(n4227), .B(n4226), .Z(n268) );
  NAND U2017 ( .A(n267), .B(n268), .Z(n6064) );
  NANDN U2018 ( .A(n2173), .B(n2172), .Z(n269) );
  NANDN U2019 ( .A(n2171), .B(n2170), .Z(n270) );
  AND U2020 ( .A(n269), .B(n270), .Z(n6055) );
  NANDN U2021 ( .A(n4017), .B(n4016), .Z(n271) );
  NANDN U2022 ( .A(n4019), .B(n4018), .Z(n272) );
  NAND U2023 ( .A(n271), .B(n272), .Z(n6049) );
  NANDN U2024 ( .A(n4627), .B(n4626), .Z(n273) );
  NANDN U2025 ( .A(n4625), .B(n4624), .Z(n274) );
  AND U2026 ( .A(n273), .B(n274), .Z(n6728) );
  NANDN U2027 ( .A(n2485), .B(n2484), .Z(n275) );
  NANDN U2028 ( .A(n2483), .B(n2482), .Z(n276) );
  AND U2029 ( .A(n275), .B(n276), .Z(n6723) );
  NAND U2030 ( .A(n5651), .B(n5650), .Z(n277) );
  NANDN U2031 ( .A(n5649), .B(n5648), .Z(n278) );
  AND U2032 ( .A(n277), .B(n278), .Z(n7618) );
  NANDN U2033 ( .A(n6158), .B(n6157), .Z(n279) );
  NANDN U2034 ( .A(n6156), .B(n6155), .Z(n280) );
  AND U2035 ( .A(n279), .B(n280), .Z(n7397) );
  NANDN U2036 ( .A(n6076), .B(n6075), .Z(n281) );
  NANDN U2037 ( .A(n6074), .B(n6073), .Z(n282) );
  AND U2038 ( .A(n281), .B(n282), .Z(n8127) );
  NANDN U2039 ( .A(n6062), .B(n6061), .Z(n283) );
  NANDN U2040 ( .A(n6060), .B(n6059), .Z(n284) );
  AND U2041 ( .A(n283), .B(n284), .Z(n8121) );
  NANDN U2042 ( .A(n5816), .B(n5815), .Z(n285) );
  NANDN U2043 ( .A(n5818), .B(n5817), .Z(n286) );
  NAND U2044 ( .A(n285), .B(n286), .Z(n8403) );
  NANDN U2045 ( .A(n5511), .B(n5510), .Z(n287) );
  NANDN U2046 ( .A(n5513), .B(n5512), .Z(n288) );
  NAND U2047 ( .A(n287), .B(n288), .Z(n8410) );
  NAND U2048 ( .A(n8270), .B(n8271), .Z(n289) );
  NANDN U2049 ( .A(n8269), .B(n8268), .Z(n290) );
  NAND U2050 ( .A(n289), .B(n290), .Z(n8943) );
  NAND U2051 ( .A(n7927), .B(n7925), .Z(n291) );
  XOR U2052 ( .A(n7925), .B(n7927), .Z(n292) );
  NANDN U2053 ( .A(n7926), .B(n292), .Z(n293) );
  NAND U2054 ( .A(n291), .B(n293), .Z(n8967) );
  XNOR U2055 ( .A(n9007), .B(n9006), .Z(n8683) );
  NAND U2056 ( .A(n7983), .B(n7982), .Z(n294) );
  NANDN U2057 ( .A(n7981), .B(n7980), .Z(n295) );
  AND U2058 ( .A(n294), .B(n295), .Z(n8549) );
  NANDN U2059 ( .A(n7985), .B(n7984), .Z(n296) );
  NANDN U2060 ( .A(n7987), .B(n7986), .Z(n297) );
  NAND U2061 ( .A(n296), .B(n297), .Z(n8715) );
  NAND U2062 ( .A(n7886), .B(n7887), .Z(n298) );
  NANDN U2063 ( .A(n7885), .B(n7884), .Z(n299) );
  NAND U2064 ( .A(n298), .B(n299), .Z(n8528) );
  XOR U2065 ( .A(n9250), .B(n9251), .Z(n9247) );
  NAND U2066 ( .A(n8541), .B(n8540), .Z(n300) );
  NAND U2067 ( .A(n8539), .B(n8538), .Z(n301) );
  NAND U2068 ( .A(n300), .B(n301), .Z(n9042) );
  NAND U2069 ( .A(n9149), .B(n9148), .Z(n302) );
  NANDN U2070 ( .A(n9147), .B(n9146), .Z(n303) );
  AND U2071 ( .A(n302), .B(n303), .Z(n9384) );
  NANDN U2072 ( .A(n9075), .B(n9074), .Z(n304) );
  NANDN U2073 ( .A(n9073), .B(n9072), .Z(n305) );
  AND U2074 ( .A(n304), .B(n305), .Z(n9412) );
  XNOR U2075 ( .A(n9508), .B(n9509), .Z(n9501) );
  NANDN U2076 ( .A(n9534), .B(n9533), .Z(n306) );
  NANDN U2077 ( .A(n9532), .B(n9531), .Z(n307) );
  AND U2078 ( .A(n306), .B(n307), .Z(n9561) );
  XNOR U2079 ( .A(n2260), .B(n2261), .Z(n2263) );
  XNOR U2080 ( .A(n1402), .B(n1403), .Z(n1405) );
  XOR U2081 ( .A(n4036), .B(n4037), .Z(n4038) );
  XOR U2082 ( .A(n2832), .B(n2833), .Z(n2834) );
  XOR U2083 ( .A(n1252), .B(n1253), .Z(n1254) );
  XNOR U2084 ( .A(n3677), .B(n3678), .Z(n3680) );
  XOR U2085 ( .A(n4482), .B(n4483), .Z(n4484) );
  XNOR U2086 ( .A(n2588), .B(n2589), .Z(n2591) );
  XOR U2087 ( .A(n4136), .B(n4137), .Z(n4138) );
  NANDN U2088 ( .A(n4915), .B(n4914), .Z(n308) );
  NANDN U2089 ( .A(n4917), .B(n4916), .Z(n309) );
  NAND U2090 ( .A(n308), .B(n309), .Z(n6252) );
  NANDN U2091 ( .A(n1521), .B(n1520), .Z(n310) );
  NANDN U2092 ( .A(n1523), .B(n1522), .Z(n311) );
  NAND U2093 ( .A(n310), .B(n311), .Z(n6246) );
  XOR U2094 ( .A(n6239), .B(n6240), .Z(n6241) );
  NANDN U2095 ( .A(n1729), .B(n1728), .Z(n312) );
  NANDN U2096 ( .A(n1731), .B(n1730), .Z(n313) );
  NAND U2097 ( .A(n312), .B(n313), .Z(n5313) );
  NANDN U2098 ( .A(n3696), .B(n3695), .Z(n314) );
  NANDN U2099 ( .A(n3694), .B(n3693), .Z(n315) );
  AND U2100 ( .A(n314), .B(n315), .Z(n6582) );
  NANDN U2101 ( .A(n2911), .B(n2910), .Z(n316) );
  NANDN U2102 ( .A(n2909), .B(n2908), .Z(n317) );
  AND U2103 ( .A(n316), .B(n317), .Z(n6576) );
  NANDN U2104 ( .A(n4719), .B(n4718), .Z(n318) );
  NANDN U2105 ( .A(n4721), .B(n4720), .Z(n319) );
  NAND U2106 ( .A(n318), .B(n319), .Z(n5447) );
  NANDN U2107 ( .A(n3027), .B(n3026), .Z(n320) );
  NANDN U2108 ( .A(n3029), .B(n3028), .Z(n321) );
  NAND U2109 ( .A(n320), .B(n321), .Z(n5453) );
  NANDN U2110 ( .A(n833), .B(n832), .Z(n322) );
  NANDN U2111 ( .A(n835), .B(n834), .Z(n323) );
  NAND U2112 ( .A(n322), .B(n323), .Z(n5439) );
  NANDN U2113 ( .A(n1871), .B(n1870), .Z(n324) );
  NANDN U2114 ( .A(n1873), .B(n1872), .Z(n325) );
  NAND U2115 ( .A(n324), .B(n325), .Z(n5397) );
  NANDN U2116 ( .A(n1153), .B(n1152), .Z(n326) );
  NANDN U2117 ( .A(n1155), .B(n1154), .Z(n327) );
  NAND U2118 ( .A(n326), .B(n327), .Z(n5390) );
  XOR U2119 ( .A(n5492), .B(n5493), .Z(n5494) );
  NANDN U2120 ( .A(n3211), .B(n3210), .Z(n328) );
  NANDN U2121 ( .A(n3213), .B(n3212), .Z(n329) );
  NAND U2122 ( .A(n328), .B(n329), .Z(n5487) );
  NANDN U2123 ( .A(n3716), .B(n3715), .Z(n330) );
  NANDN U2124 ( .A(n3718), .B(n3717), .Z(n331) );
  NAND U2125 ( .A(n330), .B(n331), .Z(n6110) );
  NANDN U2126 ( .A(n3656), .B(n3655), .Z(n332) );
  NANDN U2127 ( .A(n3654), .B(n3653), .Z(n333) );
  AND U2128 ( .A(n332), .B(n333), .Z(n6552) );
  NANDN U2129 ( .A(n3776), .B(n3775), .Z(n334) );
  NANDN U2130 ( .A(n3778), .B(n3777), .Z(n335) );
  NAND U2131 ( .A(n334), .B(n335), .Z(n6549) );
  NANDN U2132 ( .A(n1385), .B(n1384), .Z(n336) );
  NANDN U2133 ( .A(n1387), .B(n1386), .Z(n337) );
  NAND U2134 ( .A(n336), .B(n337), .Z(n6543) );
  NANDN U2135 ( .A(n1717), .B(n1716), .Z(n338) );
  NANDN U2136 ( .A(n1719), .B(n1718), .Z(n339) );
  NAND U2137 ( .A(n338), .B(n339), .Z(n6296) );
  NANDN U2138 ( .A(n4123), .B(n4122), .Z(n340) );
  NANDN U2139 ( .A(n4125), .B(n4124), .Z(n341) );
  NAND U2140 ( .A(n340), .B(n341), .Z(n6288) );
  NANDN U2141 ( .A(n3334), .B(n3333), .Z(n342) );
  NANDN U2142 ( .A(n3336), .B(n3335), .Z(n343) );
  NAND U2143 ( .A(n342), .B(n343), .Z(n5347) );
  NANDN U2144 ( .A(n3386), .B(n3385), .Z(n344) );
  NANDN U2145 ( .A(n3388), .B(n3387), .Z(n345) );
  NAND U2146 ( .A(n344), .B(n345), .Z(n5353) );
  NANDN U2147 ( .A(n4893), .B(n4892), .Z(n346) );
  NANDN U2148 ( .A(n4895), .B(n4894), .Z(n347) );
  NAND U2149 ( .A(n346), .B(n347), .Z(n5359) );
  XOR U2150 ( .A(n5748), .B(n5749), .Z(n5750) );
  XOR U2151 ( .A(n5754), .B(n5755), .Z(n5756) );
  XOR U2152 ( .A(n6019), .B(n6020), .Z(n6021) );
  NANDN U2153 ( .A(n3632), .B(n3631), .Z(n348) );
  NANDN U2154 ( .A(n3634), .B(n3633), .Z(n349) );
  NAND U2155 ( .A(n348), .B(n349), .Z(n7019) );
  NANDN U2156 ( .A(n3662), .B(n3661), .Z(n350) );
  NANDN U2157 ( .A(n3664), .B(n3663), .Z(n351) );
  NAND U2158 ( .A(n350), .B(n351), .Z(n7023) );
  XOR U2159 ( .A(n7028), .B(n7029), .Z(n7030) );
  NANDN U2160 ( .A(n3935), .B(n3934), .Z(n352) );
  NANDN U2161 ( .A(n3937), .B(n3936), .Z(n353) );
  NAND U2162 ( .A(n352), .B(n353), .Z(n7054) );
  NANDN U2163 ( .A(n1639), .B(n1638), .Z(n354) );
  NANDN U2164 ( .A(n1637), .B(n1636), .Z(n355) );
  AND U2165 ( .A(n354), .B(n355), .Z(n7041) );
  XOR U2166 ( .A(n5292), .B(n5293), .Z(n5294) );
  NANDN U2167 ( .A(n1567), .B(n1566), .Z(n356) );
  NANDN U2168 ( .A(n1569), .B(n1568), .Z(n357) );
  NAND U2169 ( .A(n356), .B(n357), .Z(n5299) );
  XOR U2170 ( .A(n6612), .B(n6613), .Z(n6614) );
  NANDN U2171 ( .A(n2895), .B(n2894), .Z(n358) );
  NANDN U2172 ( .A(n2897), .B(n2896), .Z(n359) );
  NAND U2173 ( .A(n358), .B(n359), .Z(n6573) );
  NANDN U2174 ( .A(n2019), .B(n2018), .Z(n360) );
  NANDN U2175 ( .A(n2021), .B(n2020), .Z(n361) );
  NAND U2176 ( .A(n360), .B(n361), .Z(n6378) );
  NANDN U2177 ( .A(n3780), .B(n3779), .Z(n362) );
  NANDN U2178 ( .A(n3782), .B(n3781), .Z(n363) );
  NAND U2179 ( .A(n362), .B(n363), .Z(n6366) );
  NANDN U2180 ( .A(n3754), .B(n3753), .Z(n364) );
  NANDN U2181 ( .A(n3756), .B(n3755), .Z(n365) );
  NAND U2182 ( .A(n364), .B(n365), .Z(n6396) );
  NANDN U2183 ( .A(n2267), .B(n2266), .Z(n366) );
  NANDN U2184 ( .A(n2269), .B(n2268), .Z(n367) );
  NAND U2185 ( .A(n366), .B(n367), .Z(n6390) );
  NANDN U2186 ( .A(n1007), .B(n1006), .Z(n368) );
  NANDN U2187 ( .A(n1009), .B(n1008), .Z(n369) );
  NAND U2188 ( .A(n368), .B(n369), .Z(n5567) );
  XOR U2189 ( .A(n5612), .B(n5613), .Z(n5614) );
  XOR U2190 ( .A(n5606), .B(n5607), .Z(n5608) );
  NANDN U2191 ( .A(n1027), .B(n1026), .Z(n370) );
  NANDN U2192 ( .A(n1029), .B(n1028), .Z(n371) );
  NAND U2193 ( .A(n370), .B(n371), .Z(n5603) );
  NANDN U2194 ( .A(n919), .B(n918), .Z(n372) );
  NANDN U2195 ( .A(n921), .B(n920), .Z(n373) );
  NAND U2196 ( .A(n372), .B(n373), .Z(n5992) );
  NANDN U2197 ( .A(n895), .B(n894), .Z(n374) );
  NANDN U2198 ( .A(n897), .B(n896), .Z(n375) );
  NAND U2199 ( .A(n374), .B(n375), .Z(n5980) );
  NANDN U2200 ( .A(n3460), .B(n3459), .Z(n376) );
  NANDN U2201 ( .A(n3462), .B(n3461), .Z(n377) );
  NAND U2202 ( .A(n376), .B(n377), .Z(n5956) );
  NANDN U2203 ( .A(n1687), .B(n1686), .Z(n378) );
  NANDN U2204 ( .A(n1689), .B(n1688), .Z(n379) );
  NAND U2205 ( .A(n378), .B(n379), .Z(n5209) );
  NANDN U2206 ( .A(n3294), .B(n3293), .Z(n380) );
  NANDN U2207 ( .A(n3296), .B(n3295), .Z(n381) );
  NAND U2208 ( .A(n380), .B(n381), .Z(n5197) );
  NANDN U2209 ( .A(n1495), .B(n1494), .Z(n382) );
  NANDN U2210 ( .A(n1497), .B(n1496), .Z(n383) );
  NAND U2211 ( .A(n382), .B(n383), .Z(n6210) );
  NANDN U2212 ( .A(n3195), .B(n3194), .Z(n384) );
  NANDN U2213 ( .A(n3197), .B(n3196), .Z(n385) );
  NAND U2214 ( .A(n384), .B(n385), .Z(n6204) );
  NANDN U2215 ( .A(n1399), .B(n1398), .Z(n386) );
  NANDN U2216 ( .A(n1401), .B(n1400), .Z(n387) );
  NAND U2217 ( .A(n386), .B(n387), .Z(n7239) );
  NANDN U2218 ( .A(n1959), .B(n1958), .Z(n388) );
  NANDN U2219 ( .A(n1961), .B(n1960), .Z(n389) );
  NAND U2220 ( .A(n388), .B(n389), .Z(n7231) );
  XOR U2221 ( .A(n7224), .B(n7225), .Z(n7226) );
  NANDN U2222 ( .A(n2793), .B(n2792), .Z(n390) );
  NANDN U2223 ( .A(n2795), .B(n2794), .Z(n391) );
  NAND U2224 ( .A(n390), .B(n391), .Z(n6983) );
  XOR U2225 ( .A(n6974), .B(n6975), .Z(n6976) );
  NANDN U2226 ( .A(n3149), .B(n3148), .Z(n392) );
  NANDN U2227 ( .A(n3151), .B(n3150), .Z(n393) );
  NAND U2228 ( .A(n392), .B(n393), .Z(n5331) );
  NANDN U2229 ( .A(n1589), .B(n1588), .Z(n394) );
  NANDN U2230 ( .A(n1591), .B(n1590), .Z(n395) );
  NAND U2231 ( .A(n394), .B(n395), .Z(n5337) );
  XOR U2232 ( .A(n6125), .B(n6126), .Z(n6127) );
  NANDN U2233 ( .A(n2399), .B(n2398), .Z(n396) );
  NANDN U2234 ( .A(n2401), .B(n2400), .Z(n397) );
  NAND U2235 ( .A(n396), .B(n397), .Z(n6134) );
  NANDN U2236 ( .A(n3911), .B(n3910), .Z(n398) );
  NANDN U2237 ( .A(n3913), .B(n3912), .Z(n399) );
  NAND U2238 ( .A(n398), .B(n399), .Z(n6120) );
  NANDN U2239 ( .A(n2421), .B(n2420), .Z(n400) );
  NANDN U2240 ( .A(n2423), .B(n2422), .Z(n401) );
  NAND U2241 ( .A(n400), .B(n401), .Z(n6643) );
  XOR U2242 ( .A(n6637), .B(n6638), .Z(n6639) );
  NANDN U2243 ( .A(n1225), .B(n1224), .Z(n402) );
  NANDN U2244 ( .A(n1227), .B(n1226), .Z(n403) );
  NAND U2245 ( .A(n402), .B(n403), .Z(n6631) );
  XOR U2246 ( .A(n6679), .B(n6680), .Z(n6681) );
  NANDN U2247 ( .A(n2961), .B(n2960), .Z(n404) );
  NANDN U2248 ( .A(n2963), .B(n2962), .Z(n405) );
  NAND U2249 ( .A(n404), .B(n405), .Z(n6673) );
  NANDN U2250 ( .A(n2473), .B(n2472), .Z(n406) );
  NANDN U2251 ( .A(n2471), .B(n2470), .Z(n407) );
  AND U2252 ( .A(n406), .B(n407), .Z(n6686) );
  XOR U2253 ( .A(n5534), .B(n5535), .Z(n5536) );
  NANDN U2254 ( .A(n2497), .B(n2496), .Z(n408) );
  NANDN U2255 ( .A(n2499), .B(n2498), .Z(n409) );
  NAND U2256 ( .A(n408), .B(n409), .Z(n5543) );
  NANDN U2257 ( .A(n4647), .B(n4646), .Z(n410) );
  NANDN U2258 ( .A(n4649), .B(n4648), .Z(n411) );
  NAND U2259 ( .A(n410), .B(n411), .Z(n6165) );
  NANDN U2260 ( .A(n1823), .B(n1822), .Z(n412) );
  NANDN U2261 ( .A(n1825), .B(n1824), .Z(n413) );
  NAND U2262 ( .A(n412), .B(n413), .Z(n6160) );
  NANDN U2263 ( .A(n4661), .B(n4660), .Z(n414) );
  NANDN U2264 ( .A(n4663), .B(n4662), .Z(n415) );
  NAND U2265 ( .A(n414), .B(n415), .Z(n6171) );
  NANDN U2266 ( .A(n4329), .B(n4328), .Z(n416) );
  NANDN U2267 ( .A(n4331), .B(n4330), .Z(n417) );
  NAND U2268 ( .A(n416), .B(n417), .Z(n6462) );
  NANDN U2269 ( .A(n2345), .B(n2344), .Z(n418) );
  NANDN U2270 ( .A(n2347), .B(n2346), .Z(n419) );
  NAND U2271 ( .A(n418), .B(n419), .Z(n6470) );
  NANDN U2272 ( .A(n4351), .B(n4350), .Z(n420) );
  NANDN U2273 ( .A(n4353), .B(n4352), .Z(n421) );
  NAND U2274 ( .A(n420), .B(n421), .Z(n6425) );
  NANDN U2275 ( .A(n2299), .B(n2298), .Z(n422) );
  NANDN U2276 ( .A(n2301), .B(n2300), .Z(n423) );
  NAND U2277 ( .A(n422), .B(n423), .Z(n6420) );
  NANDN U2278 ( .A(n2337), .B(n2336), .Z(n424) );
  NANDN U2279 ( .A(n2339), .B(n2338), .Z(n425) );
  NAND U2280 ( .A(n424), .B(n425), .Z(n6431) );
  NANDN U2281 ( .A(n4669), .B(n4668), .Z(n426) );
  NANDN U2282 ( .A(n4671), .B(n4670), .Z(n427) );
  NAND U2283 ( .A(n426), .B(n427), .Z(n6180) );
  NANDN U2284 ( .A(n4657), .B(n4656), .Z(n428) );
  NANDN U2285 ( .A(n4659), .B(n4658), .Z(n429) );
  NAND U2286 ( .A(n428), .B(n429), .Z(n6177) );
  NANDN U2287 ( .A(n2233), .B(n2232), .Z(n430) );
  NANDN U2288 ( .A(n2235), .B(n2234), .Z(n431) );
  NAND U2289 ( .A(n430), .B(n431), .Z(n6090) );
  NANDN U2290 ( .A(n1847), .B(n1846), .Z(n432) );
  NANDN U2291 ( .A(n1849), .B(n1848), .Z(n433) );
  NAND U2292 ( .A(n432), .B(n433), .Z(n6084) );
  NANDN U2293 ( .A(n1209), .B(n1208), .Z(n434) );
  NANDN U2294 ( .A(n1211), .B(n1210), .Z(n435) );
  NAND U2295 ( .A(n434), .B(n435), .Z(n6080) );
  XOR U2296 ( .A(n6667), .B(n6668), .Z(n6669) );
  XOR U2297 ( .A(n6655), .B(n6656), .Z(n6657) );
  NANDN U2298 ( .A(n4781), .B(n4780), .Z(n436) );
  NANDN U2299 ( .A(n4783), .B(n4782), .Z(n437) );
  NAND U2300 ( .A(n436), .B(n437), .Z(n6270) );
  NANDN U2301 ( .A(n4557), .B(n4556), .Z(n438) );
  NANDN U2302 ( .A(n4555), .B(n4554), .Z(n439) );
  AND U2303 ( .A(n438), .B(n439), .Z(n6263) );
  NANDN U2304 ( .A(n4805), .B(n4804), .Z(n440) );
  NANDN U2305 ( .A(n4807), .B(n4806), .Z(n441) );
  NAND U2306 ( .A(n440), .B(n441), .Z(n5893) );
  NANDN U2307 ( .A(n1031), .B(n1030), .Z(n442) );
  NANDN U2308 ( .A(n1033), .B(n1032), .Z(n443) );
  NAND U2309 ( .A(n442), .B(n443), .Z(n6698) );
  XOR U2310 ( .A(n6703), .B(n6704), .Z(n6705) );
  NANDN U2311 ( .A(n4825), .B(n4824), .Z(n444) );
  NANDN U2312 ( .A(n4827), .B(n4826), .Z(n445) );
  NAND U2313 ( .A(n444), .B(n445), .Z(n5938) );
  XOR U2314 ( .A(n5929), .B(n5930), .Z(n5931) );
  NANDN U2315 ( .A(n2285), .B(n2284), .Z(n446) );
  NANDN U2316 ( .A(n2287), .B(n2286), .Z(n447) );
  NAND U2317 ( .A(n446), .B(n447), .Z(n7005) );
  NANDN U2318 ( .A(n2327), .B(n2326), .Z(n448) );
  NANDN U2319 ( .A(n2329), .B(n2328), .Z(n449) );
  NAND U2320 ( .A(n448), .B(n449), .Z(n7013) );
  NANDN U2321 ( .A(n1983), .B(n1982), .Z(n450) );
  NANDN U2322 ( .A(n1985), .B(n1984), .Z(n451) );
  NAND U2323 ( .A(n450), .B(n451), .Z(n7001) );
  NANDN U2324 ( .A(n4929), .B(n4928), .Z(n452) );
  NANDN U2325 ( .A(n4931), .B(n4930), .Z(n453) );
  NAND U2326 ( .A(n452), .B(n453), .Z(n5245) );
  XOR U2327 ( .A(n5170), .B(n5171), .Z(n5172) );
  NANDN U2328 ( .A(n2731), .B(n2730), .Z(n454) );
  NANDN U2329 ( .A(n2733), .B(n2732), .Z(n455) );
  NAND U2330 ( .A(n454), .B(n455), .Z(n5165) );
  NANDN U2331 ( .A(n2705), .B(n2704), .Z(n456) );
  NANDN U2332 ( .A(n2707), .B(n2706), .Z(n457) );
  NAND U2333 ( .A(n456), .B(n457), .Z(n5161) );
  NANDN U2334 ( .A(n953), .B(n952), .Z(n458) );
  NANDN U2335 ( .A(n951), .B(n950), .Z(n459) );
  AND U2336 ( .A(n458), .B(n459), .Z(n5262) );
  NANDN U2337 ( .A(n1907), .B(n1906), .Z(n460) );
  NANDN U2338 ( .A(n1909), .B(n1908), .Z(n461) );
  NAND U2339 ( .A(n460), .B(n461), .Z(n5269) );
  NANDN U2340 ( .A(n1083), .B(n1082), .Z(n462) );
  NANDN U2341 ( .A(n1085), .B(n1084), .Z(n463) );
  NAND U2342 ( .A(n462), .B(n463), .Z(n5259) );
  NANDN U2343 ( .A(n1903), .B(n1902), .Z(n464) );
  NANDN U2344 ( .A(n1905), .B(n1904), .Z(n465) );
  NAND U2345 ( .A(n464), .B(n465), .Z(n5788) );
  NANDN U2346 ( .A(n869), .B(n868), .Z(n466) );
  NANDN U2347 ( .A(n871), .B(n870), .Z(n467) );
  NAND U2348 ( .A(n466), .B(n467), .Z(n5782) );
  XOR U2349 ( .A(n6335), .B(n6336), .Z(n6337) );
  NANDN U2350 ( .A(n3732), .B(n3731), .Z(n468) );
  NANDN U2351 ( .A(n3734), .B(n3733), .Z(n469) );
  NAND U2352 ( .A(n468), .B(n469), .Z(n6329) );
  NANDN U2353 ( .A(n995), .B(n994), .Z(n470) );
  NANDN U2354 ( .A(n997), .B(n996), .Z(n471) );
  NAND U2355 ( .A(n470), .B(n471), .Z(n5579) );
  NANDN U2356 ( .A(n4435), .B(n4434), .Z(n472) );
  NANDN U2357 ( .A(n4437), .B(n4436), .Z(n473) );
  NAND U2358 ( .A(n472), .B(n473), .Z(n5870) );
  NANDN U2359 ( .A(n1937), .B(n1936), .Z(n474) );
  NANDN U2360 ( .A(n1939), .B(n1938), .Z(n475) );
  NAND U2361 ( .A(n474), .B(n475), .Z(n5864) );
  NANDN U2362 ( .A(n3526), .B(n3525), .Z(n476) );
  NANDN U2363 ( .A(n3528), .B(n3527), .Z(n477) );
  NAND U2364 ( .A(n476), .B(n477), .Z(n5858) );
  XOR U2365 ( .A(n6710), .B(n6711), .Z(n6712) );
  XOR U2366 ( .A(n6437), .B(n6438), .Z(n6439) );
  NAND U2367 ( .A(n4262), .B(n4263), .Z(n478) );
  NANDN U2368 ( .A(n4261), .B(n4260), .Z(n479) );
  NAND U2369 ( .A(n478), .B(n479), .Z(n7152) );
  NAND U2370 ( .A(n1343), .B(n1342), .Z(n480) );
  NANDN U2371 ( .A(n1341), .B(n1340), .Z(n481) );
  AND U2372 ( .A(n480), .B(n481), .Z(n7085) );
  XOR U2373 ( .A(n5378), .B(n5379), .Z(n5380) );
  NANDN U2374 ( .A(n4285), .B(n4284), .Z(n482) );
  NANDN U2375 ( .A(n4287), .B(n4286), .Z(n483) );
  NAND U2376 ( .A(n482), .B(n483), .Z(n6494) );
  XOR U2377 ( .A(n6485), .B(n6486), .Z(n6487) );
  NANDN U2378 ( .A(n2435), .B(n2434), .Z(n484) );
  NANDN U2379 ( .A(n2437), .B(n2436), .Z(n485) );
  NAND U2380 ( .A(n484), .B(n485), .Z(n6479) );
  NANDN U2381 ( .A(n4637), .B(n4636), .Z(n486) );
  NANDN U2382 ( .A(n4639), .B(n4638), .Z(n487) );
  NAND U2383 ( .A(n486), .B(n487), .Z(n6074) );
  NANDN U2384 ( .A(n4233), .B(n4232), .Z(n488) );
  NANDN U2385 ( .A(n4235), .B(n4234), .Z(n489) );
  NAND U2386 ( .A(n488), .B(n489), .Z(n6066) );
  NANDN U2387 ( .A(n2249), .B(n2248), .Z(n490) );
  NANDN U2388 ( .A(n2251), .B(n2250), .Z(n491) );
  NAND U2389 ( .A(n490), .B(n491), .Z(n6060) );
  NANDN U2390 ( .A(n4021), .B(n4020), .Z(n492) );
  NANDN U2391 ( .A(n4023), .B(n4022), .Z(n493) );
  NAND U2392 ( .A(n492), .B(n493), .Z(n6052) );
  NANDN U2393 ( .A(n4621), .B(n4620), .Z(n494) );
  NANDN U2394 ( .A(n4623), .B(n4622), .Z(n495) );
  NAND U2395 ( .A(n494), .B(n495), .Z(n6729) );
  NANDN U2396 ( .A(n2479), .B(n2478), .Z(n496) );
  NANDN U2397 ( .A(n2481), .B(n2480), .Z(n497) );
  NAND U2398 ( .A(n496), .B(n497), .Z(n6722) );
  XOR U2399 ( .A(n7296), .B(n7297), .Z(n7298) );
  XOR U2400 ( .A(n1470), .B(n1471), .Z(n1472) );
  XNOR U2401 ( .A(n4512), .B(n4513), .Z(n4515) );
  NAND U2402 ( .A(n985), .B(n984), .Z(n498) );
  NANDN U2403 ( .A(n983), .B(n982), .Z(n499) );
  AND U2404 ( .A(n498), .B(n499), .Z(n5415) );
  XOR U2405 ( .A(n7544), .B(n7545), .Z(n7546) );
  XOR U2406 ( .A(n8162), .B(n8163), .Z(n8164) );
  NAND U2407 ( .A(n4977), .B(n4976), .Z(n500) );
  NANDN U2408 ( .A(n4979), .B(n4978), .Z(n501) );
  NAND U2409 ( .A(n500), .B(n501), .Z(n8015) );
  NAND U2410 ( .A(n5695), .B(n5694), .Z(n502) );
  NANDN U2411 ( .A(n5693), .B(n5692), .Z(n503) );
  AND U2412 ( .A(n502), .B(n503), .Z(n7988) );
  NAND U2413 ( .A(n5646), .B(n5647), .Z(n504) );
  NANDN U2414 ( .A(n5645), .B(n5644), .Z(n505) );
  NAND U2415 ( .A(n504), .B(n505), .Z(n7619) );
  NAND U2416 ( .A(n5729), .B(n5728), .Z(n506) );
  NAND U2417 ( .A(n5727), .B(n5726), .Z(n507) );
  NAND U2418 ( .A(n506), .B(n507), .Z(n7646) );
  XNOR U2419 ( .A(n8060), .B(n8061), .Z(n8063) );
  XNOR U2420 ( .A(n8054), .B(n8055), .Z(n8057) );
  XNOR U2421 ( .A(n7402), .B(n7403), .Z(n7405) );
  XOR U2422 ( .A(n7396), .B(n7397), .Z(n7398) );
  NANDN U2423 ( .A(n6070), .B(n6069), .Z(n508) );
  NANDN U2424 ( .A(n6072), .B(n6071), .Z(n509) );
  NAND U2425 ( .A(n508), .B(n509), .Z(n8126) );
  NANDN U2426 ( .A(n6056), .B(n6055), .Z(n510) );
  NANDN U2427 ( .A(n6058), .B(n6057), .Z(n511) );
  NAND U2428 ( .A(n510), .B(n511), .Z(n8120) );
  NANDN U2429 ( .A(n5822), .B(n5821), .Z(n512) );
  NANDN U2430 ( .A(n5820), .B(n5819), .Z(n513) );
  AND U2431 ( .A(n512), .B(n513), .Z(n8405) );
  XOR U2432 ( .A(n7830), .B(n7831), .Z(n7832) );
  NAND U2433 ( .A(n5109), .B(n5108), .Z(n514) );
  NAND U2434 ( .A(n5107), .B(n5106), .Z(n515) );
  NAND U2435 ( .A(n514), .B(n515), .Z(n7809) );
  NAND U2436 ( .A(n5179), .B(n5178), .Z(n516) );
  NANDN U2437 ( .A(n5177), .B(n5176), .Z(n517) );
  AND U2438 ( .A(n516), .B(n517), .Z(n7504) );
  NAND U2439 ( .A(n6860), .B(n6861), .Z(n518) );
  NANDN U2440 ( .A(n6859), .B(n6858), .Z(n519) );
  NAND U2441 ( .A(n518), .B(n519), .Z(n7427) );
  XOR U2442 ( .A(n8918), .B(n8919), .Z(n8920) );
  NAND U2443 ( .A(n7459), .B(n7458), .Z(n520) );
  XOR U2444 ( .A(n7458), .B(n7459), .Z(n521) );
  NAND U2445 ( .A(n521), .B(n7457), .Z(n522) );
  NAND U2446 ( .A(n520), .B(n522), .Z(n8609) );
  XOR U2447 ( .A(n8498), .B(n8499), .Z(n8500) );
  XOR U2448 ( .A(n8816), .B(n8817), .Z(n8818) );
  XOR U2449 ( .A(n8972), .B(n8973), .Z(n8974) );
  NAND U2450 ( .A(n7868), .B(n7869), .Z(n523) );
  NANDN U2451 ( .A(n7867), .B(n7866), .Z(n524) );
  NAND U2452 ( .A(n523), .B(n524), .Z(n8949) );
  XOR U2453 ( .A(n7924), .B(n7923), .Z(n525) );
  NANDN U2454 ( .A(n7922), .B(n525), .Z(n526) );
  NAND U2455 ( .A(n7924), .B(n7923), .Z(n527) );
  AND U2456 ( .A(n526), .B(n527), .Z(n8966) );
  XNOR U2457 ( .A(n8572), .B(n8573), .Z(n8575) );
  XOR U2458 ( .A(n8566), .B(n8567), .Z(n8568) );
  NAND U2459 ( .A(n7678), .B(n7679), .Z(n528) );
  NANDN U2460 ( .A(n7677), .B(n7676), .Z(n529) );
  NAND U2461 ( .A(n528), .B(n529), .Z(n8755) );
  NAND U2462 ( .A(n7603), .B(n7602), .Z(n530) );
  NANDN U2463 ( .A(n7605), .B(n7604), .Z(n531) );
  NAND U2464 ( .A(n530), .B(n531), .Z(n8674) );
  XOR U2465 ( .A(n7915), .B(n7914), .Z(n532) );
  NANDN U2466 ( .A(n7913), .B(n532), .Z(n533) );
  NAND U2467 ( .A(n7915), .B(n7914), .Z(n534) );
  AND U2468 ( .A(n533), .B(n534), .Z(n8931) );
  NAND U2469 ( .A(n8411), .B(n8410), .Z(n535) );
  NANDN U2470 ( .A(n8409), .B(n8408), .Z(n536) );
  AND U2471 ( .A(n535), .B(n536), .Z(n8835) );
  NAND U2472 ( .A(n8321), .B(n8320), .Z(n537) );
  NAND U2473 ( .A(n8318), .B(n8319), .Z(n538) );
  NAND U2474 ( .A(n537), .B(n538), .Z(n8658) );
  NAND U2475 ( .A(n1170), .B(n1171), .Z(n539) );
  NANDN U2476 ( .A(n1169), .B(n1168), .Z(n540) );
  NAND U2477 ( .A(n539), .B(n540), .Z(n6789) );
  NAND U2478 ( .A(n7416), .B(n7417), .Z(n541) );
  NANDN U2479 ( .A(n7415), .B(n7414), .Z(n542) );
  NAND U2480 ( .A(n541), .B(n542), .Z(n8711) );
  OR U2481 ( .A(n7880), .B(n7881), .Z(n543) );
  NAND U2482 ( .A(n7883), .B(n7882), .Z(n544) );
  NAND U2483 ( .A(n543), .B(n544), .Z(n8531) );
  NAND U2484 ( .A(n8683), .B(n8682), .Z(n545) );
  XOR U2485 ( .A(n8682), .B(n8683), .Z(n546) );
  NAND U2486 ( .A(n546), .B(n8681), .Z(n547) );
  NAND U2487 ( .A(n545), .B(n547), .Z(n9048) );
  NAND U2488 ( .A(n8536), .B(n8537), .Z(n548) );
  NANDN U2489 ( .A(n8535), .B(n8534), .Z(n549) );
  NAND U2490 ( .A(n548), .B(n549), .Z(n9045) );
  NAND U2491 ( .A(n9025), .B(n9024), .Z(n550) );
  NANDN U2492 ( .A(n9023), .B(n9022), .Z(n551) );
  AND U2493 ( .A(n550), .B(n551), .Z(n9118) );
  NAND U2494 ( .A(n8739), .B(n8738), .Z(n552) );
  NAND U2495 ( .A(n8736), .B(n8737), .Z(n553) );
  NAND U2496 ( .A(n552), .B(n553), .Z(n9057) );
  XOR U2497 ( .A(n9345), .B(n9346), .Z(n9355) );
  XOR U2498 ( .A(n9339), .B(n9340), .Z(n9341) );
  NAND U2499 ( .A(n9206), .B(n9207), .Z(n554) );
  NANDN U2500 ( .A(n9205), .B(n9204), .Z(n555) );
  NAND U2501 ( .A(n554), .B(n555), .Z(n9378) );
  NAND U2502 ( .A(n9278), .B(n9279), .Z(n556) );
  NANDN U2503 ( .A(n9277), .B(n9276), .Z(n557) );
  NAND U2504 ( .A(n556), .B(n557), .Z(n9443) );
  XOR U2505 ( .A(n9417), .B(n9418), .Z(n9419) );
  XOR U2506 ( .A(n9488), .B(n9489), .Z(n9490) );
  XOR U2507 ( .A(n9494), .B(n9495), .Z(n9496) );
  NAND U2508 ( .A(n9410), .B(n9409), .Z(n558) );
  NANDN U2509 ( .A(n9408), .B(n9407), .Z(n559) );
  AND U2510 ( .A(n558), .B(n559), .Z(n9512) );
  NAND U2511 ( .A(n9312), .B(n9313), .Z(n560) );
  NANDN U2512 ( .A(n9311), .B(n9310), .Z(n561) );
  NAND U2513 ( .A(n560), .B(n561), .Z(n9448) );
  NAND U2514 ( .A(n9486), .B(n9487), .Z(n562) );
  NANDN U2515 ( .A(n9485), .B(n9484), .Z(n563) );
  NAND U2516 ( .A(n562), .B(n563), .Z(n9548) );
  XOR U2517 ( .A(n9563), .B(n9562), .Z(n564) );
  NAND U2518 ( .A(n564), .B(n9561), .Z(n565) );
  NAND U2519 ( .A(n9563), .B(n9562), .Z(n566) );
  AND U2520 ( .A(n565), .B(n566), .Z(n9568) );
  XOR U2521 ( .A(n2310), .B(n2311), .Z(n2312) );
  XNOR U2522 ( .A(n4024), .B(n4025), .Z(n4027) );
  XNOR U2523 ( .A(n2064), .B(n2065), .Z(n2067) );
  XNOR U2524 ( .A(n2196), .B(n2197), .Z(n2199) );
  XOR U2525 ( .A(n2070), .B(n2071), .Z(n2072) );
  XNOR U2526 ( .A(n2100), .B(n2101), .Z(n2103) );
  XOR U2527 ( .A(n4394), .B(n4395), .Z(n4396) );
  XNOR U2528 ( .A(n2936), .B(n2937), .Z(n2939) );
  XOR U2529 ( .A(n1864), .B(n1865), .Z(n1866) );
  XNOR U2530 ( .A(n4908), .B(n4909), .Z(n4911) );
  XOR U2531 ( .A(n4446), .B(n4447), .Z(n4448) );
  XOR U2532 ( .A(n3505), .B(n3506), .Z(n3507) );
  XNOR U2533 ( .A(n3413), .B(n3414), .Z(n3416) );
  XOR U2534 ( .A(n1316), .B(n1317), .Z(n1318) );
  XOR U2535 ( .A(n3321), .B(n3322), .Z(n3323) );
  XOR U2536 ( .A(n2052), .B(n2053), .Z(n2054) );
  XNOR U2537 ( .A(n2094), .B(n2095), .Z(n2097) );
  XOR U2538 ( .A(n2278), .B(n2279), .Z(n2280) );
  XNOR U2539 ( .A(n4158), .B(n4159), .Z(n4161) );
  XNOR U2540 ( .A(n2148), .B(n2149), .Z(n2151) );
  XOR U2541 ( .A(n4428), .B(n4429), .Z(n4430) );
  XNOR U2542 ( .A(n4075), .B(n4074), .Z(n3791) );
  XOR U2543 ( .A(n6251), .B(n6252), .Z(n6253) );
  NANDN U2544 ( .A(n3318), .B(n3317), .Z(n567) );
  NANDN U2545 ( .A(n3320), .B(n3319), .Z(n568) );
  NAND U2546 ( .A(n567), .B(n568), .Z(n6242) );
  NANDN U2547 ( .A(n4107), .B(n4106), .Z(n569) );
  NANDN U2548 ( .A(n4109), .B(n4108), .Z(n570) );
  NAND U2549 ( .A(n569), .B(n570), .Z(n5317) );
  XOR U2550 ( .A(n5310), .B(n5311), .Z(n5312) );
  NANDN U2551 ( .A(n1419), .B(n1418), .Z(n571) );
  NANDN U2552 ( .A(n1421), .B(n1420), .Z(n572) );
  NAND U2553 ( .A(n571), .B(n572), .Z(n5305) );
  NANDN U2554 ( .A(n3690), .B(n3689), .Z(n573) );
  NANDN U2555 ( .A(n3692), .B(n3691), .Z(n574) );
  NAND U2556 ( .A(n573), .B(n574), .Z(n6583) );
  NANDN U2557 ( .A(n2905), .B(n2904), .Z(n575) );
  NANDN U2558 ( .A(n2907), .B(n2906), .Z(n576) );
  NAND U2559 ( .A(n575), .B(n576), .Z(n6577) );
  XOR U2560 ( .A(n5444), .B(n5445), .Z(n5446) );
  NANDN U2561 ( .A(n3019), .B(n3018), .Z(n577) );
  NANDN U2562 ( .A(n3021), .B(n3020), .Z(n578) );
  NAND U2563 ( .A(n577), .B(n578), .Z(n5451) );
  XOR U2564 ( .A(n5438), .B(n5439), .Z(n5440) );
  NANDN U2565 ( .A(n1879), .B(n1878), .Z(n579) );
  NANDN U2566 ( .A(n1881), .B(n1880), .Z(n580) );
  NAND U2567 ( .A(n579), .B(n580), .Z(n5399) );
  XOR U2568 ( .A(n5390), .B(n5391), .Z(n5392) );
  XOR U2569 ( .A(n5384), .B(n5385), .Z(n5386) );
  NANDN U2570 ( .A(n883), .B(n882), .Z(n581) );
  NANDN U2571 ( .A(n885), .B(n884), .Z(n582) );
  NAND U2572 ( .A(n581), .B(n582), .Z(n5495) );
  XOR U2573 ( .A(n5486), .B(n5487), .Z(n5488) );
  NANDN U2574 ( .A(n3658), .B(n3657), .Z(n583) );
  NANDN U2575 ( .A(n3660), .B(n3659), .Z(n584) );
  NAND U2576 ( .A(n583), .B(n584), .Z(n6555) );
  XOR U2577 ( .A(n6546), .B(n6547), .Z(n6548) );
  XOR U2578 ( .A(n6540), .B(n6541), .Z(n6542) );
  XOR U2579 ( .A(n5346), .B(n5347), .Z(n5348) );
  XOR U2580 ( .A(n5352), .B(n5353), .Z(n5354) );
  XOR U2581 ( .A(n5358), .B(n5359), .Z(n5360) );
  XOR U2582 ( .A(n6025), .B(n6026), .Z(n6027) );
  NANDN U2583 ( .A(n2859), .B(n2858), .Z(n585) );
  NANDN U2584 ( .A(n2861), .B(n2860), .Z(n586) );
  NAND U2585 ( .A(n585), .B(n586), .Z(n7062) );
  XOR U2586 ( .A(n7071), .B(n7072), .Z(n7073) );
  XOR U2587 ( .A(n7065), .B(n7066), .Z(n7067) );
  NANDN U2588 ( .A(n1641), .B(n1640), .Z(n587) );
  NANDN U2589 ( .A(n1643), .B(n1642), .Z(n588) );
  NAND U2590 ( .A(n587), .B(n588), .Z(n7044) );
  XOR U2591 ( .A(n6600), .B(n6601), .Z(n6602) );
  XOR U2592 ( .A(n6570), .B(n6571), .Z(n6572) );
  NANDN U2593 ( .A(n2385), .B(n2384), .Z(n589) );
  NANDN U2594 ( .A(n2387), .B(n2386), .Z(n590) );
  NAND U2595 ( .A(n589), .B(n590), .Z(n6567) );
  NANDN U2596 ( .A(n2027), .B(n2026), .Z(n591) );
  NANDN U2597 ( .A(n2029), .B(n2028), .Z(n592) );
  NAND U2598 ( .A(n591), .B(n592), .Z(n6380) );
  XOR U2599 ( .A(n6371), .B(n6372), .Z(n6373) );
  NANDN U2600 ( .A(n3788), .B(n3787), .Z(n593) );
  NANDN U2601 ( .A(n3790), .B(n3789), .Z(n594) );
  NAND U2602 ( .A(n593), .B(n594), .Z(n6368) );
  XOR U2603 ( .A(n6401), .B(n6402), .Z(n6403) );
  NANDN U2604 ( .A(n3762), .B(n3761), .Z(n595) );
  NANDN U2605 ( .A(n3764), .B(n3763), .Z(n596) );
  NAND U2606 ( .A(n595), .B(n596), .Z(n6398) );
  NANDN U2607 ( .A(n2275), .B(n2274), .Z(n597) );
  NANDN U2608 ( .A(n2277), .B(n2276), .Z(n598) );
  NAND U2609 ( .A(n597), .B(n598), .Z(n6392) );
  NANDN U2610 ( .A(n2743), .B(n2742), .Z(n599) );
  NANDN U2611 ( .A(n2745), .B(n2744), .Z(n600) );
  NAND U2612 ( .A(n599), .B(n600), .Z(n5559) );
  NANDN U2613 ( .A(n2715), .B(n2714), .Z(n601) );
  NANDN U2614 ( .A(n2717), .B(n2716), .Z(n602) );
  NAND U2615 ( .A(n601), .B(n602), .Z(n5553) );
  NANDN U2616 ( .A(n1113), .B(n1112), .Z(n603) );
  NANDN U2617 ( .A(n1115), .B(n1114), .Z(n604) );
  NAND U2618 ( .A(n603), .B(n604), .Z(n5615) );
  NANDN U2619 ( .A(n899), .B(n898), .Z(n605) );
  NANDN U2620 ( .A(n901), .B(n900), .Z(n606) );
  NAND U2621 ( .A(n605), .B(n606), .Z(n5607) );
  XOR U2622 ( .A(n5989), .B(n5990), .Z(n5991) );
  NANDN U2623 ( .A(n4877), .B(n4876), .Z(n607) );
  NANDN U2624 ( .A(n4879), .B(n4878), .Z(n608) );
  NAND U2625 ( .A(n607), .B(n608), .Z(n5966) );
  XOR U2626 ( .A(n5953), .B(n5954), .Z(n5955) );
  NANDN U2627 ( .A(n1697), .B(n1696), .Z(n609) );
  NANDN U2628 ( .A(n1699), .B(n1698), .Z(n610) );
  NAND U2629 ( .A(n609), .B(n610), .Z(n5211) );
  XOR U2630 ( .A(n5196), .B(n5197), .Z(n5198) );
  NANDN U2631 ( .A(n1505), .B(n1504), .Z(n611) );
  NANDN U2632 ( .A(n1507), .B(n1506), .Z(n612) );
  NAND U2633 ( .A(n611), .B(n612), .Z(n6212) );
  XOR U2634 ( .A(n6203), .B(n6204), .Z(n6205) );
  XOR U2635 ( .A(n6215), .B(n6216), .Z(n6217) );
  XOR U2636 ( .A(n7230), .B(n7231), .Z(n7232) );
  NANDN U2637 ( .A(n4007), .B(n4006), .Z(n613) );
  NANDN U2638 ( .A(n4009), .B(n4008), .Z(n614) );
  NAND U2639 ( .A(n613), .B(n614), .Z(n7227) );
  XOR U2640 ( .A(n6986), .B(n6987), .Z(n6988) );
  XOR U2641 ( .A(n6980), .B(n6981), .Z(n6982) );
  XOR U2642 ( .A(n5322), .B(n5323), .Z(n5324) );
  NANDN U2643 ( .A(n3919), .B(n3918), .Z(n615) );
  NANDN U2644 ( .A(n3921), .B(n3920), .Z(n616) );
  NAND U2645 ( .A(n615), .B(n616), .Z(n6122) );
  NANDN U2646 ( .A(n2417), .B(n2416), .Z(n617) );
  NANDN U2647 ( .A(n2419), .B(n2418), .Z(n618) );
  NAND U2648 ( .A(n617), .B(n618), .Z(n6646) );
  XOR U2649 ( .A(n6631), .B(n6632), .Z(n6633) );
  XOR U2650 ( .A(n6673), .B(n6674), .Z(n6675) );
  NANDN U2651 ( .A(n2467), .B(n2466), .Z(n619) );
  NANDN U2652 ( .A(n2469), .B(n2468), .Z(n620) );
  NAND U2653 ( .A(n619), .B(n620), .Z(n6685) );
  NANDN U2654 ( .A(n4653), .B(n4652), .Z(n621) );
  NANDN U2655 ( .A(n4651), .B(n4650), .Z(n622) );
  AND U2656 ( .A(n621), .B(n622), .Z(n6166) );
  NANDN U2657 ( .A(n1831), .B(n1830), .Z(n623) );
  NANDN U2658 ( .A(n1833), .B(n1832), .Z(n624) );
  NAND U2659 ( .A(n623), .B(n624), .Z(n6162) );
  NANDN U2660 ( .A(n4667), .B(n4666), .Z(n625) );
  NANDN U2661 ( .A(n4665), .B(n4664), .Z(n626) );
  AND U2662 ( .A(n625), .B(n626), .Z(n6172) );
  NANDN U2663 ( .A(n4337), .B(n4336), .Z(n627) );
  NANDN U2664 ( .A(n4339), .B(n4338), .Z(n628) );
  NAND U2665 ( .A(n627), .B(n628), .Z(n6464) );
  NANDN U2666 ( .A(n4419), .B(n4418), .Z(n629) );
  NANDN U2667 ( .A(n4421), .B(n4420), .Z(n630) );
  NAND U2668 ( .A(n629), .B(n630), .Z(n6458) );
  NANDN U2669 ( .A(n2349), .B(n2348), .Z(n631) );
  NANDN U2670 ( .A(n2351), .B(n2350), .Z(n632) );
  NAND U2671 ( .A(n631), .B(n632), .Z(n6467) );
  NANDN U2672 ( .A(n4347), .B(n4346), .Z(n633) );
  NANDN U2673 ( .A(n4349), .B(n4348), .Z(n634) );
  NAND U2674 ( .A(n633), .B(n634), .Z(n6428) );
  NANDN U2675 ( .A(n2307), .B(n2306), .Z(n635) );
  NANDN U2676 ( .A(n2309), .B(n2308), .Z(n636) );
  NAND U2677 ( .A(n635), .B(n636), .Z(n6422) );
  NANDN U2678 ( .A(n4679), .B(n4678), .Z(n637) );
  NANDN U2679 ( .A(n4677), .B(n4676), .Z(n638) );
  AND U2680 ( .A(n637), .B(n638), .Z(n6182) );
  NANDN U2681 ( .A(n4655), .B(n4654), .Z(n6178) );
  NANDN U2682 ( .A(n2241), .B(n2240), .Z(n639) );
  NANDN U2683 ( .A(n2243), .B(n2242), .Z(n640) );
  NAND U2684 ( .A(n639), .B(n640), .Z(n6092) );
  NANDN U2685 ( .A(n1855), .B(n1854), .Z(n641) );
  NANDN U2686 ( .A(n1857), .B(n1856), .Z(n642) );
  NAND U2687 ( .A(n641), .B(n642), .Z(n6086) );
  NANDN U2688 ( .A(n2357), .B(n2356), .Z(n643) );
  NANDN U2689 ( .A(n2359), .B(n2358), .Z(n644) );
  NAND U2690 ( .A(n643), .B(n644), .Z(n6662) );
  NANDN U2691 ( .A(n2943), .B(n2942), .Z(n645) );
  NANDN U2692 ( .A(n2945), .B(n2944), .Z(n646) );
  NAND U2693 ( .A(n645), .B(n646), .Z(n6668) );
  NANDN U2694 ( .A(n2875), .B(n2874), .Z(n647) );
  NANDN U2695 ( .A(n2877), .B(n2876), .Z(n648) );
  NAND U2696 ( .A(n647), .B(n648), .Z(n6656) );
  NANDN U2697 ( .A(n4789), .B(n4788), .Z(n649) );
  NANDN U2698 ( .A(n4791), .B(n4790), .Z(n650) );
  NAND U2699 ( .A(n649), .B(n650), .Z(n6272) );
  NANDN U2700 ( .A(n4559), .B(n4558), .Z(n651) );
  NANDN U2701 ( .A(n4561), .B(n4560), .Z(n652) );
  NAND U2702 ( .A(n651), .B(n652), .Z(n6266) );
  XOR U2703 ( .A(n5899), .B(n5900), .Z(n5901) );
  XOR U2704 ( .A(n5893), .B(n5894), .Z(n5895) );
  XOR U2705 ( .A(n5887), .B(n5888), .Z(n5889) );
  NANDN U2706 ( .A(n1037), .B(n1036), .Z(n653) );
  NANDN U2707 ( .A(n1035), .B(n1034), .Z(n654) );
  AND U2708 ( .A(n653), .B(n654), .Z(n6697) );
  XOR U2709 ( .A(n5935), .B(n5936), .Z(n5937) );
  NANDN U2710 ( .A(n3376), .B(n3375), .Z(n655) );
  NANDN U2711 ( .A(n3378), .B(n3377), .Z(n656) );
  NAND U2712 ( .A(n655), .B(n656), .Z(n5932) );
  XOR U2713 ( .A(n5923), .B(n5924), .Z(n5925) );
  NANDN U2714 ( .A(n1611), .B(n1610), .Z(n657) );
  NANDN U2715 ( .A(n1613), .B(n1612), .Z(n658) );
  NAND U2716 ( .A(n657), .B(n658), .Z(n6531) );
  NANDN U2717 ( .A(n1623), .B(n1622), .Z(n659) );
  NANDN U2718 ( .A(n1621), .B(n1620), .Z(n660) );
  AND U2719 ( .A(n659), .B(n660), .Z(n6522) );
  NANDN U2720 ( .A(n4937), .B(n4936), .Z(n661) );
  NANDN U2721 ( .A(n4939), .B(n4938), .Z(n662) );
  NAND U2722 ( .A(n661), .B(n662), .Z(n5247) );
  NANDN U2723 ( .A(n1771), .B(n1770), .Z(n663) );
  NANDN U2724 ( .A(n1773), .B(n1772), .Z(n664) );
  NAND U2725 ( .A(n663), .B(n664), .Z(n5233) );
  NANDN U2726 ( .A(n4735), .B(n4734), .Z(n665) );
  NANDN U2727 ( .A(n4737), .B(n4736), .Z(n666) );
  NAND U2728 ( .A(n665), .B(n666), .Z(n5173) );
  NANDN U2729 ( .A(n2739), .B(n2738), .Z(n667) );
  NANDN U2730 ( .A(n2741), .B(n2740), .Z(n668) );
  NAND U2731 ( .A(n667), .B(n668), .Z(n5167) );
  NANDN U2732 ( .A(n2697), .B(n2696), .Z(n669) );
  NANDN U2733 ( .A(n2699), .B(n2698), .Z(n670) );
  NAND U2734 ( .A(n669), .B(n670), .Z(n5159) );
  NANDN U2735 ( .A(n947), .B(n946), .Z(n671) );
  NANDN U2736 ( .A(n949), .B(n948), .Z(n672) );
  NAND U2737 ( .A(n671), .B(n672), .Z(n5263) );
  NANDN U2738 ( .A(n1915), .B(n1914), .Z(n673) );
  NANDN U2739 ( .A(n1917), .B(n1916), .Z(n674) );
  NAND U2740 ( .A(n673), .B(n674), .Z(n5271) );
  NANDN U2741 ( .A(n1075), .B(n1074), .Z(n675) );
  NANDN U2742 ( .A(n1077), .B(n1076), .Z(n676) );
  NAND U2743 ( .A(n675), .B(n676), .Z(n5257) );
  NANDN U2744 ( .A(n1895), .B(n1894), .Z(n677) );
  NANDN U2745 ( .A(n1897), .B(n1896), .Z(n678) );
  NAND U2746 ( .A(n677), .B(n678), .Z(n5786) );
  NANDN U2747 ( .A(n861), .B(n860), .Z(n679) );
  NANDN U2748 ( .A(n863), .B(n862), .Z(n680) );
  NAND U2749 ( .A(n679), .B(n680), .Z(n5780) );
  NANDN U2750 ( .A(n961), .B(n960), .Z(n681) );
  NANDN U2751 ( .A(n963), .B(n962), .Z(n682) );
  NAND U2752 ( .A(n681), .B(n682), .Z(n5774) );
  NANDN U2753 ( .A(n2015), .B(n2014), .Z(n683) );
  NANDN U2754 ( .A(n2017), .B(n2016), .Z(n684) );
  NAND U2755 ( .A(n683), .B(n684), .Z(n6338) );
  XOR U2756 ( .A(n6329), .B(n6330), .Z(n6331) );
  NANDN U2757 ( .A(n987), .B(n986), .Z(n685) );
  NANDN U2758 ( .A(n989), .B(n988), .Z(n686) );
  NAND U2759 ( .A(n685), .B(n686), .Z(n5577) );
  NANDN U2760 ( .A(n4443), .B(n4442), .Z(n687) );
  NANDN U2761 ( .A(n4445), .B(n4444), .Z(n688) );
  NAND U2762 ( .A(n687), .B(n688), .Z(n5872) );
  XOR U2763 ( .A(n5863), .B(n5864), .Z(n5865) );
  XOR U2764 ( .A(n5857), .B(n5858), .Z(n5859) );
  XNOR U2765 ( .A(n6649), .B(n6650), .Z(n6652) );
  NAND U2766 ( .A(n1740), .B(n1741), .Z(n689) );
  NANDN U2767 ( .A(n1739), .B(n1738), .Z(n690) );
  NAND U2768 ( .A(n689), .B(n690), .Z(n5619) );
  XNOR U2769 ( .A(n5594), .B(n5595), .Z(n5597) );
  XOR U2770 ( .A(n6383), .B(n6384), .Z(n6385) );
  XOR U2771 ( .A(n6359), .B(n6360), .Z(n6361) );
  XOR U2772 ( .A(n6353), .B(n6354), .Z(n6355) );
  XOR U2773 ( .A(n7152), .B(n7153), .Z(n7154) );
  XOR U2774 ( .A(n6892), .B(n6893), .Z(n6894) );
  XOR U2775 ( .A(n6962), .B(n6963), .Z(n6964) );
  XOR U2776 ( .A(n5468), .B(n5469), .Z(n5470) );
  XOR U2777 ( .A(n7102), .B(n7103), .Z(n7104) );
  XOR U2778 ( .A(n6618), .B(n6619), .Z(n6620) );
  XOR U2779 ( .A(n6594), .B(n6595), .Z(n6596) );
  XOR U2780 ( .A(n7124), .B(n7125), .Z(n7126) );
  NAND U2781 ( .A(n3908), .B(n3909), .Z(n691) );
  NANDN U2782 ( .A(n3907), .B(n3906), .Z(n692) );
  NAND U2783 ( .A(n691), .B(n692), .Z(n5013) );
  NAND U2784 ( .A(n3601), .B(n3602), .Z(n693) );
  NANDN U2785 ( .A(n3600), .B(n3599), .Z(n694) );
  NAND U2786 ( .A(n693), .B(n694), .Z(n5686) );
  NAND U2787 ( .A(n1416), .B(n1417), .Z(n695) );
  NANDN U2788 ( .A(n1415), .B(n1414), .Z(n696) );
  NAND U2789 ( .A(n695), .B(n696), .Z(n5140) );
  NAND U2790 ( .A(n4144), .B(n4145), .Z(n697) );
  NANDN U2791 ( .A(n4143), .B(n4142), .Z(n698) );
  NAND U2792 ( .A(n697), .B(n698), .Z(n5671) );
  NAND U2793 ( .A(n4315), .B(n4314), .Z(n699) );
  NANDN U2794 ( .A(n4313), .B(n4312), .Z(n700) );
  AND U2795 ( .A(n699), .B(n700), .Z(n5017) );
  NANDN U2796 ( .A(n1193), .B(n1192), .Z(n701) );
  NANDN U2797 ( .A(n1191), .B(n1190), .Z(n702) );
  NAND U2798 ( .A(n701), .B(n702), .Z(n5058) );
  NAND U2799 ( .A(n4582), .B(n4583), .Z(n703) );
  NANDN U2800 ( .A(n4581), .B(n4580), .Z(n704) );
  NAND U2801 ( .A(n703), .B(n704), .Z(n6305) );
  NANDN U2802 ( .A(n2043), .B(n2042), .Z(n705) );
  NANDN U2803 ( .A(n2045), .B(n2044), .Z(n706) );
  NAND U2804 ( .A(n705), .B(n706), .Z(n6095) );
  XNOR U2805 ( .A(n7206), .B(n7207), .Z(n7209) );
  NANDN U2806 ( .A(n4221), .B(n4220), .Z(n707) );
  NANDN U2807 ( .A(n4223), .B(n4222), .Z(n708) );
  NAND U2808 ( .A(n707), .B(n708), .Z(n6188) );
  NANDN U2809 ( .A(n1819), .B(n1818), .Z(n709) );
  NANDN U2810 ( .A(n1821), .B(n1820), .Z(n710) );
  NAND U2811 ( .A(n709), .B(n710), .Z(n6194) );
  NANDN U2812 ( .A(n4691), .B(n4690), .Z(n711) );
  NANDN U2813 ( .A(n4689), .B(n4688), .Z(n712) );
  AND U2814 ( .A(n711), .B(n712), .Z(n6152) );
  NANDN U2815 ( .A(n4867), .B(n4866), .Z(n713) );
  NANDN U2816 ( .A(n4869), .B(n4868), .Z(n714) );
  NAND U2817 ( .A(n713), .B(n714), .Z(n6158) );
  XOR U2818 ( .A(n6491), .B(n6492), .Z(n6493) );
  NANDN U2819 ( .A(n2441), .B(n2440), .Z(n715) );
  NANDN U2820 ( .A(n2439), .B(n2438), .Z(n716) );
  AND U2821 ( .A(n715), .B(n716), .Z(n6480) );
  NANDN U2822 ( .A(n4633), .B(n4632), .Z(n717) );
  NANDN U2823 ( .A(n4635), .B(n4634), .Z(n718) );
  NAND U2824 ( .A(n717), .B(n718), .Z(n6076) );
  NANDN U2825 ( .A(n4849), .B(n4848), .Z(n719) );
  NANDN U2826 ( .A(n4847), .B(n4846), .Z(n720) );
  AND U2827 ( .A(n719), .B(n720), .Z(n6069) );
  NANDN U2828 ( .A(n2245), .B(n2244), .Z(n721) );
  NANDN U2829 ( .A(n2247), .B(n2246), .Z(n722) );
  NAND U2830 ( .A(n721), .B(n722), .Z(n6062) );
  NANDN U2831 ( .A(n2175), .B(n2174), .Z(n723) );
  NANDN U2832 ( .A(n2177), .B(n2176), .Z(n724) );
  NAND U2833 ( .A(n723), .B(n724), .Z(n6058) );
  NANDN U2834 ( .A(n4629), .B(n4628), .Z(n725) );
  NANDN U2835 ( .A(n4631), .B(n4630), .Z(n726) );
  NAND U2836 ( .A(n725), .B(n726), .Z(n6731) );
  NANDN U2837 ( .A(n2475), .B(n2474), .Z(n727) );
  NANDN U2838 ( .A(n2477), .B(n2476), .Z(n728) );
  NAND U2839 ( .A(n727), .B(n728), .Z(n6725) );
  NANDN U2840 ( .A(n2537), .B(n2536), .Z(n729) );
  NANDN U2841 ( .A(n2539), .B(n2538), .Z(n730) );
  NAND U2842 ( .A(n729), .B(n730), .Z(n5815) );
  XOR U2843 ( .A(n5809), .B(n5810), .Z(n5811) );
  NANDN U2844 ( .A(n1745), .B(n1744), .Z(n731) );
  NANDN U2845 ( .A(n1743), .B(n1742), .Z(n732) );
  AND U2846 ( .A(n731), .B(n732), .Z(n5521) );
  NANDN U2847 ( .A(n3073), .B(n3072), .Z(n733) );
  NANDN U2848 ( .A(n3075), .B(n3074), .Z(n734) );
  NAND U2849 ( .A(n733), .B(n734), .Z(n5515) );
  NANDN U2850 ( .A(n2403), .B(n2402), .Z(n735) );
  NANDN U2851 ( .A(n2405), .B(n2404), .Z(n736) );
  NAND U2852 ( .A(n735), .B(n736), .Z(n5513) );
  XNOR U2853 ( .A(n5803), .B(n5804), .Z(n5806) );
  XNOR U2854 ( .A(n5797), .B(n5798), .Z(n5800) );
  XNOR U2855 ( .A(n5917), .B(n5918), .Z(n5920) );
  XNOR U2856 ( .A(n4518), .B(n4519), .Z(n4521) );
  XOR U2857 ( .A(n4422), .B(n4423), .Z(n4424) );
  XOR U2858 ( .A(n4744), .B(n4745), .Z(n4746) );
  XOR U2859 ( .A(n4506), .B(n4507), .Z(n4508) );
  XNOR U2860 ( .A(n4045), .B(n4044), .Z(n4695) );
  XNOR U2861 ( .A(n1310), .B(n1311), .Z(n1313) );
  XOR U2862 ( .A(n1304), .B(n1305), .Z(n1306) );
  XOR U2863 ( .A(n4164), .B(n4165), .Z(n4166) );
  XOR U2864 ( .A(n3435), .B(n3436), .Z(n3437) );
  XOR U2865 ( .A(n7572), .B(n7573), .Z(n7574) );
  XNOR U2866 ( .A(n7566), .B(n7567), .Z(n7569) );
  XNOR U2867 ( .A(n7448), .B(n7449), .Z(n7451) );
  XNOR U2868 ( .A(n7442), .B(n7443), .Z(n7445) );
  XOR U2869 ( .A(n7526), .B(n7527), .Z(n7528) );
  XNOR U2870 ( .A(n7520), .B(n7521), .Z(n7523) );
  XOR U2871 ( .A(n7484), .B(n7485), .Z(n7486) );
  XNOR U2872 ( .A(n8138), .B(n8139), .Z(n8141) );
  XNOR U2873 ( .A(n8000), .B(n8001), .Z(n8003) );
  XOR U2874 ( .A(n7956), .B(n7957), .Z(n7958) );
  XOR U2875 ( .A(n7944), .B(n7945), .Z(n7946) );
  XOR U2876 ( .A(n8084), .B(n8085), .Z(n8086) );
  NAND U2877 ( .A(n5639), .B(n5638), .Z(n737) );
  NANDN U2878 ( .A(n5637), .B(n5636), .Z(n738) );
  AND U2879 ( .A(n737), .B(n738), .Z(n7671) );
  NAND U2880 ( .A(n5642), .B(n5643), .Z(n739) );
  NANDN U2881 ( .A(n5641), .B(n5640), .Z(n740) );
  NAND U2882 ( .A(n739), .B(n740), .Z(n7621) );
  NAND U2883 ( .A(n6943), .B(n6942), .Z(n741) );
  NAND U2884 ( .A(n6941), .B(n6940), .Z(n742) );
  NAND U2885 ( .A(n741), .B(n742), .Z(n7971) );
  NAND U2886 ( .A(n7116), .B(n7117), .Z(n743) );
  NANDN U2887 ( .A(n7115), .B(n7114), .Z(n744) );
  NAND U2888 ( .A(n743), .B(n744), .Z(n7965) );
  NAND U2889 ( .A(n5655), .B(n5654), .Z(n745) );
  NAND U2890 ( .A(n5653), .B(n5652), .Z(n746) );
  NAND U2891 ( .A(n745), .B(n746), .Z(n7466) );
  XNOR U2892 ( .A(n8050), .B(n8051), .Z(n8021) );
  XOR U2893 ( .A(n7514), .B(n7515), .Z(n7516) );
  XNOR U2894 ( .A(n7508), .B(n7509), .Z(n7511) );
  XOR U2895 ( .A(n8202), .B(n8203), .Z(n8204) );
  XOR U2896 ( .A(n7824), .B(n7825), .Z(n7826) );
  XNOR U2897 ( .A(n2533), .B(n2532), .Z(n3990) );
  XOR U2898 ( .A(n1554), .B(n1555), .Z(n1556) );
  XNOR U2899 ( .A(n4152), .B(n4153), .Z(n4155) );
  XOR U2900 ( .A(n976), .B(n977), .Z(n978) );
  XNOR U2901 ( .A(n1782), .B(n1783), .Z(n1785) );
  XOR U2902 ( .A(n1536), .B(n1537), .Z(n1538) );
  XOR U2903 ( .A(n1668), .B(n1669), .Z(n1670) );
  XOR U2904 ( .A(n4452), .B(n4453), .Z(n4454) );
  OR U2905 ( .A(n4090), .B(n4091), .Z(n747) );
  NANDN U2906 ( .A(n4093), .B(n4092), .Z(n748) );
  NAND U2907 ( .A(n747), .B(n748), .Z(n6937) );
  NAND U2908 ( .A(n7144), .B(n7145), .Z(n749) );
  NANDN U2909 ( .A(n7143), .B(n7142), .Z(n750) );
  NAND U2910 ( .A(n749), .B(n750), .Z(n7851) );
  NAND U2911 ( .A(n1260), .B(n1261), .Z(n751) );
  NANDN U2912 ( .A(n1259), .B(n1258), .Z(n752) );
  NAND U2913 ( .A(n751), .B(n752), .Z(n6824) );
  NAND U2914 ( .A(n5831), .B(n5832), .Z(n753) );
  NANDN U2915 ( .A(n5830), .B(n5829), .Z(n754) );
  NAND U2916 ( .A(n753), .B(n754), .Z(n7843) );
  XNOR U2917 ( .A(n8912), .B(n8913), .Z(n8915) );
  NAND U2918 ( .A(n7551), .B(n7550), .Z(n755) );
  XOR U2919 ( .A(n7550), .B(n7551), .Z(n756) );
  NANDN U2920 ( .A(n7552), .B(n756), .Z(n757) );
  NAND U2921 ( .A(n755), .B(n757), .Z(n8615) );
  NAND U2922 ( .A(n7456), .B(n7455), .Z(n758) );
  XOR U2923 ( .A(n7455), .B(n7456), .Z(n759) );
  NAND U2924 ( .A(n759), .B(n7454), .Z(n760) );
  NAND U2925 ( .A(n758), .B(n760), .Z(n8610) );
  XOR U2926 ( .A(n8627), .B(n8628), .Z(n8629) );
  XOR U2927 ( .A(n8621), .B(n8622), .Z(n8623) );
  XOR U2928 ( .A(n8828), .B(n8829), .Z(n8830) );
  XOR U2929 ( .A(n8822), .B(n8823), .Z(n8824) );
  XOR U2930 ( .A(n8978), .B(n8979), .Z(n8980) );
  XOR U2931 ( .A(n8948), .B(n8949), .Z(n8950) );
  XNOR U2932 ( .A(n8942), .B(n8943), .Z(n8945) );
  XOR U2933 ( .A(n8804), .B(n8805), .Z(n8806) );
  XNOR U2934 ( .A(n8960), .B(n8961), .Z(n8963) );
  XNOR U2935 ( .A(n8998), .B(n8999), .Z(n9001) );
  NAND U2936 ( .A(n8176), .B(n8177), .Z(n761) );
  NANDN U2937 ( .A(n8175), .B(n8174), .Z(n762) );
  NAND U2938 ( .A(n761), .B(n762), .Z(n9016) );
  NAND U2939 ( .A(n7930), .B(n7931), .Z(n763) );
  NANDN U2940 ( .A(n7929), .B(n7928), .Z(n764) );
  NAND U2941 ( .A(n763), .B(n764), .Z(n8932) );
  NAND U2942 ( .A(n7388), .B(n7389), .Z(n765) );
  NANDN U2943 ( .A(n7387), .B(n7386), .Z(n766) );
  NAND U2944 ( .A(n765), .B(n766), .Z(n8482) );
  XOR U2945 ( .A(n8516), .B(n8517), .Z(n8518) );
  XOR U2946 ( .A(n8522), .B(n8523), .Z(n8524) );
  XNOR U2947 ( .A(n8510), .B(n8511), .Z(n8513) );
  XNOR U2948 ( .A(n8846), .B(n8847), .Z(n8849) );
  XOR U2949 ( .A(n8840), .B(n8841), .Z(n8842) );
  XOR U2950 ( .A(n8834), .B(n8835), .Z(n8836) );
  XOR U2951 ( .A(n8578), .B(n8579), .Z(n8580) );
  XNOR U2952 ( .A(n8989), .B(n8988), .Z(n8596) );
  XOR U2953 ( .A(n8590), .B(n8591), .Z(n8592) );
  XOR U2954 ( .A(n8852), .B(n8853), .Z(n8854) );
  NAND U2955 ( .A(n7911), .B(n7910), .Z(n767) );
  XOR U2956 ( .A(n7910), .B(n7911), .Z(n768) );
  NANDN U2957 ( .A(n7912), .B(n768), .Z(n769) );
  NAND U2958 ( .A(n767), .B(n769), .Z(n8554) );
  XNOR U2959 ( .A(n3722), .B(n3721), .Z(n2868) );
  NANDN U2960 ( .A(n5183), .B(n5182), .Z(n770) );
  NANDN U2961 ( .A(n5181), .B(n5180), .Z(n771) );
  AND U2962 ( .A(n770), .B(n771), .Z(n7694) );
  NANDN U2963 ( .A(n7877), .B(n7876), .Z(n772) );
  NANDN U2964 ( .A(n7879), .B(n7878), .Z(n773) );
  NAND U2965 ( .A(n772), .B(n773), .Z(n8638) );
  NAND U2966 ( .A(n7639), .B(n7638), .Z(n774) );
  NANDN U2967 ( .A(n7637), .B(n7636), .Z(n775) );
  AND U2968 ( .A(n774), .B(n775), .Z(n8781) );
  XNOR U2969 ( .A(n9168), .B(n9169), .Z(n9171) );
  XNOR U2970 ( .A(n9180), .B(n9181), .Z(n9183) );
  NAND U2971 ( .A(n8636), .B(n8635), .Z(n776) );
  NANDN U2972 ( .A(n8634), .B(n8633), .Z(n777) );
  AND U2973 ( .A(n776), .B(n777), .Z(n9193) );
  NAND U2974 ( .A(n8679), .B(n8680), .Z(n778) );
  NANDN U2975 ( .A(n8678), .B(n8677), .Z(n779) );
  NAND U2976 ( .A(n778), .B(n779), .Z(n9125) );
  NAND U2977 ( .A(n8657), .B(n8658), .Z(n780) );
  NANDN U2978 ( .A(n8656), .B(n8655), .Z(n781) );
  NAND U2979 ( .A(n780), .B(n781), .Z(n9098) );
  NAND U2980 ( .A(n8761), .B(n8760), .Z(n782) );
  NANDN U2981 ( .A(n8759), .B(n8758), .Z(n783) );
  AND U2982 ( .A(n782), .B(n783), .Z(n9055) );
  OR U2983 ( .A(n6788), .B(n6789), .Z(n784) );
  NAND U2984 ( .A(n6790), .B(n6791), .Z(n785) );
  AND U2985 ( .A(n784), .B(n785), .Z(n8306) );
  NAND U2986 ( .A(n8717), .B(n8716), .Z(n786) );
  NANDN U2987 ( .A(n8715), .B(n8714), .Z(n787) );
  AND U2988 ( .A(n786), .B(n787), .Z(n9265) );
  XOR U2989 ( .A(n9347), .B(n9348), .Z(n9349) );
  XOR U2990 ( .A(n9383), .B(n9384), .Z(n9385) );
  XNOR U2991 ( .A(n9356), .B(n9355), .Z(n9390) );
  XOR U2992 ( .A(n9377), .B(n9378), .Z(n9379) );
  NAND U2993 ( .A(n9034), .B(n9035), .Z(n788) );
  NANDN U2994 ( .A(n9033), .B(n9032), .Z(n789) );
  NAND U2995 ( .A(n788), .B(n789), .Z(n9404) );
  NAND U2996 ( .A(n8292), .B(n8293), .Z(n790) );
  NANDN U2997 ( .A(n8291), .B(n8290), .Z(n791) );
  NAND U2998 ( .A(n790), .B(n791), .Z(n8469) );
  NAND U2999 ( .A(n9097), .B(n9096), .Z(n792) );
  NANDN U3000 ( .A(n9095), .B(n9094), .Z(n793) );
  AND U3001 ( .A(n792), .B(n793), .Z(n9436) );
  XOR U3002 ( .A(n9502), .B(n9503), .Z(n9486) );
  XOR U3003 ( .A(n9512), .B(n9513), .Z(n9514) );
  OR U3004 ( .A(n9432), .B(n9433), .Z(n794) );
  NAND U3005 ( .A(n9435), .B(n9434), .Z(n795) );
  NAND U3006 ( .A(n794), .B(n795), .Z(n9475) );
  XOR U3007 ( .A(n9542), .B(n9541), .Z(n9551) );
  XOR U3008 ( .A(n9425), .B(n9424), .Z(n796) );
  NANDN U3009 ( .A(n9423), .B(n796), .Z(n797) );
  NAND U3010 ( .A(n9425), .B(n9424), .Z(n798) );
  AND U3011 ( .A(n797), .B(n798), .Z(n9454) );
  XOR U3012 ( .A(n9567), .B(n9568), .Z(n799) );
  NANDN U3013 ( .A(n9569), .B(n799), .Z(n800) );
  NAND U3014 ( .A(n9567), .B(n9568), .Z(n801) );
  AND U3015 ( .A(n800), .B(n801), .Z(o[10]) );
  XNOR U3016 ( .A(x[1159]), .B(y[1159]), .Z(n929) );
  XNOR U3017 ( .A(x[91]), .B(y[91]), .Z(n927) );
  XOR U3018 ( .A(x[1161]), .B(y[1161]), .Z(n926) );
  XNOR U3019 ( .A(n927), .B(n926), .Z(n928) );
  XOR U3020 ( .A(n929), .B(n928), .Z(n4485) );
  XNOR U3021 ( .A(x[1151]), .B(y[1151]), .Z(n3320) );
  XNOR U3022 ( .A(x[85]), .B(y[85]), .Z(n3318) );
  XOR U3023 ( .A(x[1153]), .B(y[1153]), .Z(n3317) );
  XNOR U3024 ( .A(n3318), .B(n3317), .Z(n3319) );
  XNOR U3025 ( .A(n3320), .B(n3319), .Z(n4482) );
  XNOR U3026 ( .A(x[1155]), .B(y[1155]), .Z(n3316) );
  XNOR U3027 ( .A(x[280]), .B(y[280]), .Z(n3314) );
  XOR U3028 ( .A(x[1157]), .B(y[1157]), .Z(n3313) );
  XNOR U3029 ( .A(n3314), .B(n3313), .Z(n3315) );
  XNOR U3030 ( .A(n3316), .B(n3315), .Z(n4483) );
  XNOR U3031 ( .A(n4485), .B(n4484), .Z(n2839) );
  XNOR U3032 ( .A(x[1171]), .B(y[1171]), .Z(n839) );
  XNOR U3033 ( .A(x[101]), .B(y[101]), .Z(n836) );
  XNOR U3034 ( .A(x[1173]), .B(y[1173]), .Z(n837) );
  XOR U3035 ( .A(n836), .B(n837), .Z(n838) );
  XOR U3036 ( .A(n839), .B(n838), .Z(n4303) );
  XNOR U3037 ( .A(x[1167]), .B(y[1167]), .Z(n845) );
  XNOR U3038 ( .A(x[1169]), .B(y[1169]), .Z(n842) );
  XNOR U3039 ( .A(x[1548]), .B(y[1548]), .Z(n843) );
  XOR U3040 ( .A(n842), .B(n843), .Z(n844) );
  XOR U3041 ( .A(n845), .B(n844), .Z(n4300) );
  XNOR U3042 ( .A(x[1163]), .B(y[1163]), .Z(n1159) );
  XNOR U3043 ( .A(x[95]), .B(y[95]), .Z(n1156) );
  XNOR U3044 ( .A(x[1165]), .B(y[1165]), .Z(n1157) );
  XOR U3045 ( .A(n1156), .B(n1157), .Z(n1158) );
  XNOR U3046 ( .A(n1159), .B(n1158), .Z(n4301) );
  XNOR U3047 ( .A(n4300), .B(n4301), .Z(n4302) );
  XOR U3048 ( .A(n4303), .B(n4302), .Z(n2838) );
  XOR U3049 ( .A(n2839), .B(n2838), .Z(n2841) );
  XNOR U3050 ( .A(x[1147]), .B(y[1147]), .Z(n3280) );
  XNOR U3051 ( .A(x[286]), .B(y[286]), .Z(n3278) );
  XOR U3052 ( .A(x[1149]), .B(y[1149]), .Z(n3276) );
  XNOR U3053 ( .A(n3278), .B(n3276), .Z(n3279) );
  XOR U3054 ( .A(n3280), .B(n3279), .Z(n4051) );
  XNOR U3055 ( .A(x[1139]), .B(y[1139]), .Z(n3378) );
  XNOR U3056 ( .A(x[79]), .B(y[79]), .Z(n3376) );
  XOR U3057 ( .A(x[1141]), .B(y[1141]), .Z(n3375) );
  XNOR U3058 ( .A(n3376), .B(n3375), .Z(n3377) );
  XOR U3059 ( .A(n3378), .B(n3377), .Z(n4048) );
  XNOR U3060 ( .A(x[1143]), .B(y[1143]), .Z(n3340) );
  XNOR U3061 ( .A(x[1145]), .B(y[1145]), .Z(n3338) );
  XOR U3062 ( .A(x[1546]), .B(y[1546]), .Z(n3337) );
  XNOR U3063 ( .A(n3338), .B(n3337), .Z(n3339) );
  XNOR U3064 ( .A(n3340), .B(n3339), .Z(n4049) );
  XNOR U3065 ( .A(n4048), .B(n4049), .Z(n4050) );
  XNOR U3066 ( .A(n4051), .B(n4050), .Z(n2840) );
  XNOR U3067 ( .A(n2841), .B(n2840), .Z(n823) );
  XNOR U3068 ( .A(x[1107]), .B(y[1107]), .Z(n2493) );
  XNOR U3069 ( .A(x[57]), .B(y[57]), .Z(n2490) );
  XNOR U3070 ( .A(x[1109]), .B(y[1109]), .Z(n2491) );
  XOR U3071 ( .A(n2490), .B(n2491), .Z(n2492) );
  XOR U3072 ( .A(n2493), .B(n2492), .Z(n4073) );
  XNOR U3073 ( .A(x[1103]), .B(y[1103]), .Z(n3612) );
  XNOR U3074 ( .A(x[1105]), .B(y[1105]), .Z(n3609) );
  XNOR U3075 ( .A(x[1540]), .B(y[1540]), .Z(n3610) );
  XOR U3076 ( .A(n3609), .B(n3610), .Z(n3611) );
  XNOR U3077 ( .A(n3612), .B(n3611), .Z(n4072) );
  XOR U3078 ( .A(n4073), .B(n4072), .Z(n4075) );
  XNOR U3079 ( .A(x[1111]), .B(y[1111]), .Z(n1577) );
  XNOR U3080 ( .A(x[1113]), .B(y[1113]), .Z(n1574) );
  XNOR U3081 ( .A(x[1542]), .B(y[1542]), .Z(n1575) );
  XOR U3082 ( .A(n1574), .B(n1575), .Z(n1576) );
  XNOR U3083 ( .A(n1577), .B(n1576), .Z(n4074) );
  XNOR U3084 ( .A(x[1123]), .B(y[1123]), .Z(n3450) );
  XNOR U3085 ( .A(x[300]), .B(y[300]), .Z(n3447) );
  XNOR U3086 ( .A(x[1125]), .B(y[1125]), .Z(n3448) );
  XOR U3087 ( .A(n3447), .B(n3448), .Z(n3449) );
  XOR U3088 ( .A(n3450), .B(n3449), .Z(n1319) );
  XNOR U3089 ( .A(x[1115]), .B(y[1115]), .Z(n1949) );
  XNOR U3090 ( .A(x[306]), .B(y[306]), .Z(n1946) );
  XNOR U3091 ( .A(x[1117]), .B(y[1117]), .Z(n1947) );
  XOR U3092 ( .A(n1946), .B(n1947), .Z(n1948) );
  XNOR U3093 ( .A(n1949), .B(n1948), .Z(n1316) );
  XNOR U3094 ( .A(x[1119]), .B(y[1119]), .Z(n1943) );
  XNOR U3095 ( .A(x[63]), .B(y[63]), .Z(n1940) );
  XNOR U3096 ( .A(x[1121]), .B(y[1121]), .Z(n1941) );
  XOR U3097 ( .A(n1940), .B(n1941), .Z(n1942) );
  XNOR U3098 ( .A(n1943), .B(n1942), .Z(n1317) );
  XNOR U3099 ( .A(n1319), .B(n1318), .Z(n3792) );
  XOR U3100 ( .A(n3791), .B(n3792), .Z(n3793) );
  XNOR U3101 ( .A(x[1135]), .B(y[1135]), .Z(n3392) );
  XNOR U3102 ( .A(x[1137]), .B(y[1137]), .Z(n3389) );
  XNOR U3103 ( .A(x[1544]), .B(y[1544]), .Z(n3390) );
  XOR U3104 ( .A(n3389), .B(n3390), .Z(n3391) );
  XOR U3105 ( .A(n3392), .B(n3391), .Z(n4431) );
  XNOR U3106 ( .A(x[1127]), .B(y[1127]), .Z(n3554) );
  XNOR U3107 ( .A(x[69]), .B(y[69]), .Z(n3551) );
  XNOR U3108 ( .A(x[1129]), .B(y[1129]), .Z(n3552) );
  XOR U3109 ( .A(n3551), .B(n3552), .Z(n3553) );
  XNOR U3110 ( .A(n3554), .B(n3553), .Z(n4428) );
  XNOR U3111 ( .A(x[1131]), .B(y[1131]), .Z(n3432) );
  XNOR U3112 ( .A(x[73]), .B(y[73]), .Z(n3429) );
  XNOR U3113 ( .A(x[1133]), .B(y[1133]), .Z(n3430) );
  XOR U3114 ( .A(n3429), .B(n3430), .Z(n3431) );
  XNOR U3115 ( .A(n3432), .B(n3431), .Z(n4429) );
  XNOR U3116 ( .A(n4431), .B(n4430), .Z(n3794) );
  XOR U3117 ( .A(n3793), .B(n3794), .Z(n820) );
  XNOR U3118 ( .A(x[1419]), .B(y[1419]), .Z(n1719) );
  XNOR U3119 ( .A(x[271]), .B(y[271]), .Z(n1717) );
  XOR U3120 ( .A(x[1421]), .B(y[1421]), .Z(n1716) );
  XNOR U3121 ( .A(n1717), .B(n1716), .Z(n1718) );
  XOR U3122 ( .A(n1719), .B(n1718), .Z(n1511) );
  XNOR U3123 ( .A(x[1323]), .B(y[1323]), .Z(n1809) );
  XNOR U3124 ( .A(x[205]), .B(y[205]), .Z(n1807) );
  XNOR U3125 ( .A(x[1325]), .B(y[1325]), .Z(n1806) );
  XNOR U3126 ( .A(n1807), .B(n1806), .Z(n1808) );
  XNOR U3127 ( .A(n1809), .B(n1808), .Z(n1508) );
  XNOR U3128 ( .A(x[1423]), .B(y[1423]), .Z(n1587) );
  XNOR U3129 ( .A(x[1425]), .B(y[1425]), .Z(n1585) );
  XOR U3130 ( .A(x[1580]), .B(y[1580]), .Z(n1584) );
  XNOR U3131 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U3132 ( .A(n1587), .B(n1586), .Z(n1509) );
  XNOR U3133 ( .A(n1508), .B(n1509), .Z(n1510) );
  XNOR U3134 ( .A(n1511), .B(n1510), .Z(n1269) );
  XNOR U3135 ( .A(x[1331]), .B(y[1331]), .Z(n2255) );
  XNOR U3136 ( .A(x[211]), .B(y[211]), .Z(n2253) );
  XOR U3137 ( .A(x[1333]), .B(y[1333]), .Z(n2252) );
  XNOR U3138 ( .A(n2253), .B(n2252), .Z(n2254) );
  XOR U3139 ( .A(n2255), .B(n2254), .Z(n2503) );
  XNOR U3140 ( .A(x[1363]), .B(y[1363]), .Z(n4679) );
  XNOR U3141 ( .A(x[233]), .B(y[233]), .Z(n4677) );
  XOR U3142 ( .A(x[1365]), .B(y[1365]), .Z(n4676) );
  XNOR U3143 ( .A(n4677), .B(n4676), .Z(n4678) );
  XOR U3144 ( .A(n4679), .B(n4678), .Z(n2500) );
  XNOR U3145 ( .A(x[1327]), .B(y[1327]), .Z(n2235) );
  XNOR U3146 ( .A(x[1329]), .B(y[1329]), .Z(n2233) );
  XOR U3147 ( .A(x[1568]), .B(y[1568]), .Z(n2232) );
  XNOR U3148 ( .A(n2233), .B(n2232), .Z(n2234) );
  XNOR U3149 ( .A(n2235), .B(n2234), .Z(n2501) );
  XNOR U3150 ( .A(n2500), .B(n2501), .Z(n2502) );
  XOR U3151 ( .A(n2503), .B(n2502), .Z(n1268) );
  XOR U3152 ( .A(n1269), .B(n1268), .Z(n1271) );
  XNOR U3153 ( .A(x[1319]), .B(y[1319]), .Z(n4849) );
  XNOR U3154 ( .A(x[201]), .B(y[201]), .Z(n4847) );
  XOR U3155 ( .A(x[1321]), .B(y[1321]), .Z(n4846) );
  XNOR U3156 ( .A(n4847), .B(n4846), .Z(n4848) );
  XOR U3157 ( .A(n4849), .B(n4848), .Z(n1047) );
  XNOR U3158 ( .A(x[1315]), .B(y[1315]), .Z(n1833) );
  XNOR U3159 ( .A(x[180]), .B(y[180]), .Z(n1831) );
  XOR U3160 ( .A(x[1317]), .B(y[1317]), .Z(n1830) );
  XNOR U3161 ( .A(n1831), .B(n1830), .Z(n1832) );
  XOR U3162 ( .A(n1833), .B(n1832), .Z(n1044) );
  XNOR U3163 ( .A(x[1427]), .B(y[1427]), .Z(n1573) );
  XNOR U3164 ( .A(x[277]), .B(y[277]), .Z(n1571) );
  XOR U3165 ( .A(x[1429]), .B(y[1429]), .Z(n1570) );
  XNOR U3166 ( .A(n1571), .B(n1570), .Z(n1572) );
  XNOR U3167 ( .A(n1573), .B(n1572), .Z(n1045) );
  XNOR U3168 ( .A(n1044), .B(n1045), .Z(n1046) );
  XNOR U3169 ( .A(n1047), .B(n1046), .Z(n1270) );
  XOR U3170 ( .A(n1271), .B(n1270), .Z(n821) );
  XNOR U3171 ( .A(n820), .B(n821), .Z(n822) );
  XNOR U3172 ( .A(n823), .B(n822), .Z(n1181) );
  XNOR U3173 ( .A(x[1287]), .B(y[1287]), .Z(n4787) );
  XNOR U3174 ( .A(x[179]), .B(y[179]), .Z(n4785) );
  XOR U3175 ( .A(x[1289]), .B(y[1289]), .Z(n4784) );
  XNOR U3176 ( .A(n4785), .B(n4784), .Z(n4786) );
  XOR U3177 ( .A(n4787), .B(n4786), .Z(n1791) );
  XNOR U3178 ( .A(x[1283]), .B(y[1283]), .Z(n4935) );
  XNOR U3179 ( .A(x[200]), .B(y[200]), .Z(n4933) );
  XOR U3180 ( .A(x[1285]), .B(y[1285]), .Z(n4932) );
  XNOR U3181 ( .A(n4933), .B(n4932), .Z(n4934) );
  XOR U3182 ( .A(n4935), .B(n4934), .Z(n1788) );
  XNOR U3183 ( .A(x[1443]), .B(y[1443]), .Z(n989) );
  XNOR U3184 ( .A(x[100]), .B(y[100]), .Z(n987) );
  XOR U3185 ( .A(x[1445]), .B(y[1445]), .Z(n986) );
  XNOR U3186 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U3187 ( .A(n989), .B(n988), .Z(n1789) );
  XNOR U3188 ( .A(n1788), .B(n1789), .Z(n1790) );
  XNOR U3189 ( .A(n1791), .B(n1790), .Z(n2209) );
  XNOR U3190 ( .A(x[1279]), .B(y[1279]), .Z(n4921) );
  XNOR U3191 ( .A(x[173]), .B(y[173]), .Z(n4918) );
  XNOR U3192 ( .A(x[1281]), .B(y[1281]), .Z(n4919) );
  XOR U3193 ( .A(n4918), .B(n4919), .Z(n4920) );
  XOR U3194 ( .A(n4921), .B(n4920), .Z(n4741) );
  XNOR U3195 ( .A(x[1275]), .B(y[1275]), .Z(n1709) );
  XNOR U3196 ( .A(x[206]), .B(y[206]), .Z(n1706) );
  XNOR U3197 ( .A(x[1277]), .B(y[1277]), .Z(n1707) );
  XOR U3198 ( .A(n1706), .B(n1707), .Z(n1708) );
  XOR U3199 ( .A(n1709), .B(n1708), .Z(n4738) );
  XNOR U3200 ( .A(x[1447]), .B(y[1447]), .Z(n1041) );
  XNOR U3201 ( .A(x[289]), .B(y[289]), .Z(n1038) );
  XNOR U3202 ( .A(x[1449]), .B(y[1449]), .Z(n1039) );
  XOR U3203 ( .A(n1038), .B(n1039), .Z(n1040) );
  XNOR U3204 ( .A(n1041), .B(n1040), .Z(n4739) );
  XNOR U3205 ( .A(n4738), .B(n4739), .Z(n4740) );
  XOR U3206 ( .A(n4741), .B(n4740), .Z(n2208) );
  XOR U3207 ( .A(n2209), .B(n2208), .Z(n2211) );
  XNOR U3208 ( .A(x[1271]), .B(y[1271]), .Z(n1497) );
  XNOR U3209 ( .A(x[1273]), .B(y[1273]), .Z(n1495) );
  XOR U3210 ( .A(x[1562]), .B(y[1562]), .Z(n1494) );
  XNOR U3211 ( .A(n1495), .B(n1494), .Z(n1496) );
  XOR U3212 ( .A(n1497), .B(n1496), .Z(n1803) );
  XNOR U3213 ( .A(x[1267]), .B(y[1267]), .Z(n1689) );
  XNOR U3214 ( .A(x[167]), .B(y[167]), .Z(n1687) );
  XOR U3215 ( .A(x[1269]), .B(y[1269]), .Z(n1686) );
  XNOR U3216 ( .A(n1687), .B(n1686), .Z(n1688) );
  XOR U3217 ( .A(n1689), .B(n1688), .Z(n1800) );
  XNOR U3218 ( .A(x[1451]), .B(y[1451]), .Z(n3514) );
  XNOR U3219 ( .A(x[293]), .B(y[293]), .Z(n3512) );
  XOR U3220 ( .A(x[1453]), .B(y[1453]), .Z(n3511) );
  XNOR U3221 ( .A(n3512), .B(n3511), .Z(n3513) );
  XNOR U3222 ( .A(n3514), .B(n3513), .Z(n1801) );
  XNOR U3223 ( .A(n1800), .B(n1801), .Z(n1802) );
  XNOR U3224 ( .A(n1803), .B(n1802), .Z(n2210) );
  XNOR U3225 ( .A(n2211), .B(n2210), .Z(n1178) );
  XNOR U3226 ( .A(x[1263]), .B(y[1263]), .Z(n1001) );
  XNOR U3227 ( .A(x[1265]), .B(y[1265]), .Z(n999) );
  XOR U3228 ( .A(x[1560]), .B(y[1560]), .Z(n998) );
  XNOR U3229 ( .A(n999), .B(n998), .Z(n1000) );
  XOR U3230 ( .A(n1001), .B(n1000), .Z(n1797) );
  XNOR U3231 ( .A(x[1259]), .B(y[1259]), .Z(n2489) );
  XNOR U3232 ( .A(x[161]), .B(y[161]), .Z(n2487) );
  XOR U3233 ( .A(x[1261]), .B(y[1261]), .Z(n2486) );
  XNOR U3234 ( .A(n2487), .B(n2486), .Z(n2488) );
  XOR U3235 ( .A(n2489), .B(n2488), .Z(n1794) );
  XNOR U3236 ( .A(x[1455]), .B(y[1455]), .Z(n3867) );
  XNOR U3237 ( .A(x[1457]), .B(y[1457]), .Z(n3865) );
  XOR U3238 ( .A(x[1584]), .B(y[1584]), .Z(n3864) );
  XNOR U3239 ( .A(n3865), .B(n3864), .Z(n3866) );
  XNOR U3240 ( .A(n3867), .B(n3866), .Z(n1795) );
  XNOR U3241 ( .A(n1794), .B(n1795), .Z(n1796) );
  XNOR U3242 ( .A(n1797), .B(n1796), .Z(n1925) );
  XNOR U3243 ( .A(x[1255]), .B(y[1255]), .Z(n1569) );
  XNOR U3244 ( .A(x[157]), .B(y[157]), .Z(n1567) );
  XOR U3245 ( .A(x[1257]), .B(y[1257]), .Z(n1566) );
  XNOR U3246 ( .A(n1567), .B(n1566), .Z(n1568) );
  XOR U3247 ( .A(n1569), .B(n1568), .Z(n4611) );
  XNOR U3248 ( .A(x[1251]), .B(y[1251]), .Z(n1583) );
  XNOR U3249 ( .A(x[220]), .B(y[220]), .Z(n1581) );
  XOR U3250 ( .A(x[1253]), .B(y[1253]), .Z(n1580) );
  XNOR U3251 ( .A(n1581), .B(n1580), .Z(n1582) );
  XOR U3252 ( .A(n1583), .B(n1582), .Z(n4608) );
  XNOR U3253 ( .A(x[1459]), .B(y[1459]), .Z(n1961) );
  XNOR U3254 ( .A(x[299]), .B(y[299]), .Z(n1959) );
  XOR U3255 ( .A(x[1461]), .B(y[1461]), .Z(n1958) );
  XNOR U3256 ( .A(n1959), .B(n1958), .Z(n1960) );
  XNOR U3257 ( .A(n1961), .B(n1960), .Z(n4609) );
  XNOR U3258 ( .A(n4608), .B(n4609), .Z(n4610) );
  XOR U3259 ( .A(n4611), .B(n4610), .Z(n1924) );
  XOR U3260 ( .A(n1925), .B(n1924), .Z(n1927) );
  XNOR U3261 ( .A(x[1247]), .B(y[1247]), .Z(n1715) );
  XNOR U3262 ( .A(x[151]), .B(y[151]), .Z(n1713) );
  XOR U3263 ( .A(x[1249]), .B(y[1249]), .Z(n1712) );
  XNOR U3264 ( .A(n1713), .B(n1712), .Z(n1714) );
  XOR U3265 ( .A(n1715), .B(n1714), .Z(n1761) );
  XNOR U3266 ( .A(x[1243]), .B(y[1243]), .Z(n1507) );
  XNOR U3267 ( .A(x[226]), .B(y[226]), .Z(n1505) );
  XOR U3268 ( .A(x[1245]), .B(y[1245]), .Z(n1504) );
  XNOR U3269 ( .A(n1505), .B(n1504), .Z(n1506) );
  XOR U3270 ( .A(n1507), .B(n1506), .Z(n1758) );
  XNOR U3271 ( .A(x[1463]), .B(y[1463]), .Z(n2045) );
  XNOR U3272 ( .A(x[1465]), .B(y[1465]), .Z(n2043) );
  XOR U3273 ( .A(x[1586]), .B(y[1586]), .Z(n2042) );
  XNOR U3274 ( .A(n2043), .B(n2042), .Z(n2044) );
  XNOR U3275 ( .A(n2045), .B(n2044), .Z(n1759) );
  XNOR U3276 ( .A(n1758), .B(n1759), .Z(n1760) );
  XNOR U3277 ( .A(n1761), .B(n1760), .Z(n1926) );
  XOR U3278 ( .A(n1927), .B(n1926), .Z(n1179) );
  XNOR U3279 ( .A(n1178), .B(n1179), .Z(n1180) );
  XNOR U3280 ( .A(n1181), .B(n1180), .Z(n1170) );
  XNOR U3281 ( .A(x[701]), .B(y[701]), .Z(n3398) );
  XNOR U3282 ( .A(x[274]), .B(y[274]), .Z(n3395) );
  XNOR U3283 ( .A(x[703]), .B(y[703]), .Z(n3396) );
  XOR U3284 ( .A(n3395), .B(n3396), .Z(n3397) );
  XOR U3285 ( .A(n3398), .B(n3397), .Z(n3855) );
  XNOR U3286 ( .A(x[693]), .B(y[693]), .Z(n3422) );
  XNOR U3287 ( .A(x[695]), .B(y[695]), .Z(n3419) );
  XNOR U3288 ( .A(x[1490]), .B(y[1490]), .Z(n3420) );
  XOR U3289 ( .A(n3419), .B(n3420), .Z(n3421) );
  XOR U3290 ( .A(n3422), .B(n3421), .Z(n3852) );
  XNOR U3291 ( .A(x[697]), .B(y[697]), .Z(n1089) );
  XNOR U3292 ( .A(x[566]), .B(y[566]), .Z(n1086) );
  XNOR U3293 ( .A(x[699]), .B(y[699]), .Z(n1087) );
  XOR U3294 ( .A(n1086), .B(n1087), .Z(n1088) );
  XNOR U3295 ( .A(n1089), .B(n1088), .Z(n3853) );
  XNOR U3296 ( .A(n3852), .B(n3853), .Z(n3854) );
  XNOR U3297 ( .A(n3855), .B(n3854), .Z(n4313) );
  XNOR U3298 ( .A(x[713]), .B(y[713]), .Z(n3344) );
  XNOR U3299 ( .A(x[262]), .B(y[262]), .Z(n3341) );
  XNOR U3300 ( .A(x[715]), .B(y[715]), .Z(n3342) );
  XOR U3301 ( .A(n3341), .B(n3342), .Z(n3343) );
  XOR U3302 ( .A(n3344), .B(n3343), .Z(n3849) );
  XNOR U3303 ( .A(x[705]), .B(y[705]), .Z(n3368) );
  XNOR U3304 ( .A(x[560]), .B(y[560]), .Z(n3365) );
  XNOR U3305 ( .A(x[707]), .B(y[707]), .Z(n3366) );
  XOR U3306 ( .A(n3365), .B(n3366), .Z(n3367) );
  XOR U3307 ( .A(n3368), .B(n3367), .Z(n3846) );
  XNOR U3308 ( .A(x[709]), .B(y[709]), .Z(n3578) );
  XNOR U3309 ( .A(x[268]), .B(y[268]), .Z(n3575) );
  XNOR U3310 ( .A(x[711]), .B(y[711]), .Z(n3576) );
  XOR U3311 ( .A(n3575), .B(n3576), .Z(n3577) );
  XNOR U3312 ( .A(n3578), .B(n3577), .Z(n3847) );
  XNOR U3313 ( .A(n3846), .B(n3847), .Z(n3848) );
  XOR U3314 ( .A(n3849), .B(n3848), .Z(n4312) );
  XNOR U3315 ( .A(n4313), .B(n4312), .Z(n4314) );
  XNOR U3316 ( .A(x[689]), .B(y[689]), .Z(n3456) );
  XNOR U3317 ( .A(x[282]), .B(y[282]), .Z(n3453) );
  XNOR U3318 ( .A(x[691]), .B(y[691]), .Z(n3454) );
  XOR U3319 ( .A(n3453), .B(n3454), .Z(n3455) );
  XOR U3320 ( .A(n3456), .B(n3455), .Z(n3879) );
  XNOR U3321 ( .A(x[681]), .B(y[681]), .Z(n1101) );
  XNOR U3322 ( .A(x[290]), .B(y[290]), .Z(n1098) );
  XNOR U3323 ( .A(x[683]), .B(y[683]), .Z(n1099) );
  XOR U3324 ( .A(n1098), .B(n1099), .Z(n1100) );
  XOR U3325 ( .A(n1101), .B(n1100), .Z(n3876) );
  XNOR U3326 ( .A(x[685]), .B(y[685]), .Z(n1095) );
  XNOR U3327 ( .A(x[687]), .B(y[687]), .Z(n1092) );
  XNOR U3328 ( .A(x[1488]), .B(y[1488]), .Z(n1093) );
  XOR U3329 ( .A(n1092), .B(n1093), .Z(n1094) );
  XNOR U3330 ( .A(n1095), .B(n1094), .Z(n3877) );
  XNOR U3331 ( .A(n3876), .B(n3877), .Z(n3878) );
  XOR U3332 ( .A(n3879), .B(n3878), .Z(n4315) );
  XOR U3333 ( .A(n4314), .B(n4315), .Z(n1164) );
  XNOR U3334 ( .A(x[629]), .B(y[629]), .Z(n4391) );
  XNOR U3335 ( .A(x[631]), .B(y[631]), .Z(n4388) );
  XNOR U3336 ( .A(x[1482]), .B(y[1482]), .Z(n4389) );
  XOR U3337 ( .A(n4388), .B(n4389), .Z(n4390) );
  XOR U3338 ( .A(n4391), .B(n4390), .Z(n3897) );
  XNOR U3339 ( .A(x[621]), .B(y[621]), .Z(n4367) );
  XNOR U3340 ( .A(x[623]), .B(y[623]), .Z(n4364) );
  XNOR U3341 ( .A(x[1480]), .B(y[1480]), .Z(n4365) );
  XOR U3342 ( .A(n4364), .B(n4365), .Z(n4366) );
  XOR U3343 ( .A(n4367), .B(n4366), .Z(n3894) );
  XNOR U3344 ( .A(x[625]), .B(y[625]), .Z(n4379) );
  XNOR U3345 ( .A(x[336]), .B(y[336]), .Z(n4376) );
  XNOR U3346 ( .A(x[627]), .B(y[627]), .Z(n4377) );
  XOR U3347 ( .A(n4376), .B(n4377), .Z(n4378) );
  XNOR U3348 ( .A(n4379), .B(n4378), .Z(n3895) );
  XNOR U3349 ( .A(n3894), .B(n3895), .Z(n3896) );
  XNOR U3350 ( .A(n3897), .B(n3896), .Z(n1191) );
  XNOR U3351 ( .A(x[641]), .B(y[641]), .Z(n1377) );
  XNOR U3352 ( .A(x[600]), .B(y[600]), .Z(n1374) );
  XNOR U3353 ( .A(x[643]), .B(y[643]), .Z(n1375) );
  XOR U3354 ( .A(n1374), .B(n1375), .Z(n1376) );
  XOR U3355 ( .A(n1377), .B(n1376), .Z(n3903) );
  XNOR U3356 ( .A(x[637]), .B(y[637]), .Z(n4491) );
  XNOR U3357 ( .A(x[330]), .B(y[330]), .Z(n4488) );
  XNOR U3358 ( .A(x[639]), .B(y[639]), .Z(n4489) );
  XOR U3359 ( .A(n4488), .B(n4489), .Z(n4490) );
  XOR U3360 ( .A(n4491), .B(n4490), .Z(n3900) );
  XNOR U3361 ( .A(x[633]), .B(y[633]), .Z(n4385) );
  XNOR U3362 ( .A(x[606]), .B(y[606]), .Z(n4382) );
  XNOR U3363 ( .A(x[635]), .B(y[635]), .Z(n4383) );
  XOR U3364 ( .A(n4382), .B(n4383), .Z(n4384) );
  XNOR U3365 ( .A(n4385), .B(n4384), .Z(n3901) );
  XNOR U3366 ( .A(n3900), .B(n3901), .Z(n3902) );
  XOR U3367 ( .A(n3903), .B(n3902), .Z(n1190) );
  XNOR U3368 ( .A(n1191), .B(n1190), .Z(n1192) );
  XNOR U3369 ( .A(x[617]), .B(y[617]), .Z(n4373) );
  XNOR U3370 ( .A(x[344]), .B(y[344]), .Z(n4370) );
  XNOR U3371 ( .A(x[619]), .B(y[619]), .Z(n4371) );
  XOR U3372 ( .A(n4370), .B(n4371), .Z(n4372) );
  XOR U3373 ( .A(n4373), .B(n4372), .Z(n3924) );
  XNOR U3374 ( .A(x[609]), .B(y[609]), .Z(n4353) );
  XNOR U3375 ( .A(x[611]), .B(y[611]), .Z(n4351) );
  XOR U3376 ( .A(x[620]), .B(y[620]), .Z(n4350) );
  XNOR U3377 ( .A(n4351), .B(n4350), .Z(n4352) );
  XNOR U3378 ( .A(n4353), .B(n4352), .Z(n3922) );
  XNOR U3379 ( .A(x[613]), .B(y[613]), .Z(n4361) );
  XNOR U3380 ( .A(x[350]), .B(y[350]), .Z(n4358) );
  XNOR U3381 ( .A(x[615]), .B(y[615]), .Z(n4359) );
  XOR U3382 ( .A(n4358), .B(n4359), .Z(n4360) );
  XNOR U3383 ( .A(n4361), .B(n4360), .Z(n3923) );
  XOR U3384 ( .A(n3924), .B(n3925), .Z(n1193) );
  XNOR U3385 ( .A(n1192), .B(n1193), .Z(n1162) );
  XNOR U3386 ( .A(x[665]), .B(y[665]), .Z(n3528) );
  XNOR U3387 ( .A(x[586]), .B(y[586]), .Z(n3526) );
  XOR U3388 ( .A(x[667]), .B(y[667]), .Z(n3525) );
  XNOR U3389 ( .A(n3526), .B(n3525), .Z(n3527) );
  XOR U3390 ( .A(n3528), .B(n3527), .Z(n1989) );
  XNOR U3391 ( .A(x[657]), .B(y[657]), .Z(n1939) );
  XNOR U3392 ( .A(x[310]), .B(y[310]), .Z(n1937) );
  XOR U3393 ( .A(x[659]), .B(y[659]), .Z(n1936) );
  XNOR U3394 ( .A(n1937), .B(n1936), .Z(n1938) );
  XOR U3395 ( .A(n1939), .B(n1938), .Z(n1986) );
  XNOR U3396 ( .A(x[661]), .B(y[661]), .Z(n3734) );
  XNOR U3397 ( .A(x[663]), .B(y[663]), .Z(n3732) );
  XOR U3398 ( .A(x[1486]), .B(y[1486]), .Z(n3731) );
  XNOR U3399 ( .A(n3732), .B(n3731), .Z(n3733) );
  XNOR U3400 ( .A(n3734), .B(n3733), .Z(n1987) );
  XNOR U3401 ( .A(n1986), .B(n1987), .Z(n1988) );
  XNOR U3402 ( .A(n1989), .B(n1988), .Z(n4581) );
  XNOR U3403 ( .A(x[677]), .B(y[677]), .Z(n3572) );
  XNOR U3404 ( .A(x[294]), .B(y[294]), .Z(n3569) );
  XNOR U3405 ( .A(x[679]), .B(y[679]), .Z(n3570) );
  XOR U3406 ( .A(n3569), .B(n3570), .Z(n3571) );
  XOR U3407 ( .A(n3572), .B(n3571), .Z(n3806) );
  XNOR U3408 ( .A(x[669]), .B(y[669]), .Z(n3560) );
  XNOR U3409 ( .A(x[302]), .B(y[302]), .Z(n3557) );
  XNOR U3410 ( .A(x[671]), .B(y[671]), .Z(n3558) );
  XOR U3411 ( .A(n3557), .B(n3558), .Z(n3559) );
  XOR U3412 ( .A(n3560), .B(n3559), .Z(n3803) );
  XNOR U3413 ( .A(x[673]), .B(y[673]), .Z(n3532) );
  XNOR U3414 ( .A(x[580]), .B(y[580]), .Z(n3529) );
  XNOR U3415 ( .A(x[675]), .B(y[675]), .Z(n3530) );
  XOR U3416 ( .A(n3529), .B(n3530), .Z(n3531) );
  XNOR U3417 ( .A(n3532), .B(n3531), .Z(n3804) );
  XNOR U3418 ( .A(n3803), .B(n3804), .Z(n3805) );
  XOR U3419 ( .A(n3806), .B(n3805), .Z(n4580) );
  XNOR U3420 ( .A(n4581), .B(n4580), .Z(n4582) );
  XNOR U3421 ( .A(x[653]), .B(y[653]), .Z(n3728) );
  XNOR U3422 ( .A(x[655]), .B(y[655]), .Z(n3725) );
  XNOR U3423 ( .A(x[1484]), .B(y[1484]), .Z(n3726) );
  XOR U3424 ( .A(n3725), .B(n3726), .Z(n3727) );
  XOR U3425 ( .A(n3728), .B(n3727), .Z(n3828) );
  XNOR U3426 ( .A(x[645]), .B(y[645]), .Z(n2007) );
  XNOR U3427 ( .A(x[322]), .B(y[322]), .Z(n2004) );
  XNOR U3428 ( .A(x[647]), .B(y[647]), .Z(n2005) );
  XOR U3429 ( .A(n2004), .B(n2005), .Z(n2006) );
  XOR U3430 ( .A(n2007), .B(n2006), .Z(n3825) );
  XNOR U3431 ( .A(x[649]), .B(y[649]), .Z(n4503) );
  XNOR U3432 ( .A(x[316]), .B(y[316]), .Z(n4500) );
  XNOR U3433 ( .A(x[651]), .B(y[651]), .Z(n4501) );
  XOR U3434 ( .A(n4500), .B(n4501), .Z(n4502) );
  XNOR U3435 ( .A(n4503), .B(n4502), .Z(n3826) );
  XNOR U3436 ( .A(n3825), .B(n3826), .Z(n3827) );
  XOR U3437 ( .A(n3828), .B(n3827), .Z(n4583) );
  XOR U3438 ( .A(n4582), .B(n4583), .Z(n1163) );
  XOR U3439 ( .A(n1162), .B(n1163), .Z(n1165) );
  XNOR U3440 ( .A(n1164), .B(n1165), .Z(n1168) );
  XNOR U3441 ( .A(x[983]), .B(y[983]), .Z(n2543) );
  XNOR U3442 ( .A(x[985]), .B(y[985]), .Z(n2541) );
  XNOR U3443 ( .A(x[1526]), .B(y[1526]), .Z(n2540) );
  XNOR U3444 ( .A(n2541), .B(n2540), .Z(n2542) );
  XNOR U3445 ( .A(n2543), .B(n2542), .Z(n4197) );
  XNOR U3446 ( .A(x[975]), .B(y[975]), .Z(n4725) );
  XNOR U3447 ( .A(x[977]), .B(y[977]), .Z(n4722) );
  XNOR U3448 ( .A(x[1524]), .B(y[1524]), .Z(n4723) );
  XOR U3449 ( .A(n4722), .B(n4723), .Z(n4724) );
  XOR U3450 ( .A(n4725), .B(n4724), .Z(n4194) );
  XNOR U3451 ( .A(x[967]), .B(y[967]), .Z(n4731) );
  XNOR U3452 ( .A(x[48]), .B(y[48]), .Z(n4728) );
  XNOR U3453 ( .A(x[969]), .B(y[969]), .Z(n4729) );
  XOR U3454 ( .A(n4728), .B(n4729), .Z(n4730) );
  XNOR U3455 ( .A(n4731), .B(n4730), .Z(n4195) );
  XNOR U3456 ( .A(n4194), .B(n4195), .Z(n4196) );
  XOR U3457 ( .A(n4197), .B(n4196), .Z(n1992) );
  XNOR U3458 ( .A(x[959]), .B(y[959]), .Z(n4721) );
  XNOR U3459 ( .A(x[54]), .B(y[54]), .Z(n4719) );
  XOR U3460 ( .A(x[961]), .B(y[961]), .Z(n4718) );
  XNOR U3461 ( .A(n4719), .B(n4718), .Z(n4720) );
  XOR U3462 ( .A(n4721), .B(n4720), .Z(n4160) );
  XNOR U3463 ( .A(x[943]), .B(y[943]), .Z(n1873) );
  XNOR U3464 ( .A(x[945]), .B(y[945]), .Z(n1871) );
  XOR U3465 ( .A(x[1520]), .B(y[1520]), .Z(n1870) );
  XNOR U3466 ( .A(n1871), .B(n1870), .Z(n1872) );
  XNOR U3467 ( .A(n1873), .B(n1872), .Z(n4158) );
  XNOR U3468 ( .A(x[951]), .B(y[951]), .Z(n1877) );
  XNOR U3469 ( .A(x[953]), .B(y[953]), .Z(n1875) );
  XOR U3470 ( .A(x[1522]), .B(y[1522]), .Z(n1874) );
  XNOR U3471 ( .A(n1875), .B(n1874), .Z(n1876) );
  XNOR U3472 ( .A(n1877), .B(n1876), .Z(n4159) );
  XOR U3473 ( .A(n4160), .B(n4161), .Z(n1993) );
  XNOR U3474 ( .A(n1992), .B(n1993), .Z(n1994) );
  XNOR U3475 ( .A(x[935]), .B(y[935]), .Z(n4593) );
  XNOR U3476 ( .A(x[74]), .B(y[74]), .Z(n4590) );
  XNOR U3477 ( .A(x[937]), .B(y[937]), .Z(n4591) );
  XOR U3478 ( .A(n4590), .B(n4591), .Z(n4592) );
  XOR U3479 ( .A(n4593), .B(n4592), .Z(n4167) );
  XNOR U3480 ( .A(x[919]), .B(y[919]), .Z(n3885) );
  XNOR U3481 ( .A(x[921]), .B(y[921]), .Z(n3883) );
  XOR U3482 ( .A(x[1518]), .B(y[1518]), .Z(n3882) );
  XNOR U3483 ( .A(n3883), .B(n3882), .Z(n3884) );
  XNOR U3484 ( .A(n3885), .B(n3884), .Z(n4164) );
  XNOR U3485 ( .A(x[927]), .B(y[927]), .Z(n4905) );
  XNOR U3486 ( .A(x[82]), .B(y[82]), .Z(n4902) );
  XNOR U3487 ( .A(x[929]), .B(y[929]), .Z(n4903) );
  XOR U3488 ( .A(n4902), .B(n4903), .Z(n4904) );
  XNOR U3489 ( .A(n4905), .B(n4904), .Z(n4165) );
  XNOR U3490 ( .A(n4167), .B(n4166), .Z(n1995) );
  XOR U3491 ( .A(n1994), .B(n1995), .Z(n2669) );
  XNOR U3492 ( .A(x[1395]), .B(y[1395]), .Z(n4939) );
  XNOR U3493 ( .A(x[255]), .B(y[255]), .Z(n4937) );
  XOR U3494 ( .A(x[1397]), .B(y[1397]), .Z(n4936) );
  XNOR U3495 ( .A(n4937), .B(n4936), .Z(n4938) );
  XOR U3496 ( .A(n4939), .B(n4938), .Z(n4873) );
  XNOR U3497 ( .A(x[1379]), .B(y[1379]), .Z(n4843) );
  XNOR U3498 ( .A(x[140]), .B(y[140]), .Z(n4841) );
  XNOR U3499 ( .A(x[1381]), .B(y[1381]), .Z(n4840) );
  XNOR U3500 ( .A(n4841), .B(n4840), .Z(n4842) );
  XNOR U3501 ( .A(n4843), .B(n4842), .Z(n4870) );
  XNOR U3502 ( .A(x[1399]), .B(y[1399]), .Z(n4931) );
  XNOR U3503 ( .A(x[1401]), .B(y[1401]), .Z(n4929) );
  XOR U3504 ( .A(x[1578]), .B(y[1578]), .Z(n4928) );
  XNOR U3505 ( .A(n4929), .B(n4928), .Z(n4930) );
  XNOR U3506 ( .A(n4931), .B(n4930), .Z(n4871) );
  XNOR U3507 ( .A(n4870), .B(n4871), .Z(n4872) );
  XNOR U3508 ( .A(n4873), .B(n4872), .Z(n941) );
  XNOR U3509 ( .A(x[1407]), .B(y[1407]), .Z(n4927) );
  XNOR U3510 ( .A(x[261]), .B(y[261]), .Z(n4925) );
  XOR U3511 ( .A(x[1409]), .B(y[1409]), .Z(n4924) );
  XNOR U3512 ( .A(n4925), .B(n4924), .Z(n4926) );
  XOR U3513 ( .A(n4927), .B(n4926), .Z(n4795) );
  XNOR U3514 ( .A(x[1355]), .B(y[1355]), .Z(n1731) );
  XNOR U3515 ( .A(x[227]), .B(y[227]), .Z(n1729) );
  XOR U3516 ( .A(x[1357]), .B(y[1357]), .Z(n1728) );
  XNOR U3517 ( .A(n1729), .B(n1728), .Z(n1730) );
  XOR U3518 ( .A(n1731), .B(n1730), .Z(n4792) );
  XNOR U3519 ( .A(x[1371]), .B(y[1371]), .Z(n1821) );
  XNOR U3520 ( .A(x[146]), .B(y[146]), .Z(n1819) );
  XOR U3521 ( .A(x[1373]), .B(y[1373]), .Z(n1818) );
  XNOR U3522 ( .A(n1819), .B(n1818), .Z(n1820) );
  XNOR U3523 ( .A(n1821), .B(n1820), .Z(n4793) );
  XNOR U3524 ( .A(n4792), .B(n4793), .Z(n4794) );
  XOR U3525 ( .A(n4795), .B(n4794), .Z(n940) );
  XOR U3526 ( .A(n941), .B(n940), .Z(n943) );
  XNOR U3527 ( .A(x[1339]), .B(y[1339]), .Z(n1829) );
  XNOR U3528 ( .A(x[166]), .B(y[166]), .Z(n1827) );
  XOR U3529 ( .A(x[1341]), .B(y[1341]), .Z(n1826) );
  XNOR U3530 ( .A(n1827), .B(n1826), .Z(n1828) );
  XOR U3531 ( .A(n1829), .B(n1828), .Z(n1703) );
  XNOR U3532 ( .A(x[1411]), .B(y[1411]), .Z(n1727) );
  XNOR U3533 ( .A(x[120]), .B(y[120]), .Z(n1725) );
  XOR U3534 ( .A(x[1413]), .B(y[1413]), .Z(n1724) );
  XNOR U3535 ( .A(n1725), .B(n1724), .Z(n1726) );
  XOR U3536 ( .A(n1727), .B(n1726), .Z(n1700) );
  XNOR U3537 ( .A(x[1359]), .B(y[1359]), .Z(n4663) );
  XNOR U3538 ( .A(x[1361]), .B(y[1361]), .Z(n4661) );
  XOR U3539 ( .A(x[1572]), .B(y[1572]), .Z(n4660) );
  XNOR U3540 ( .A(n4661), .B(n4660), .Z(n4662) );
  XNOR U3541 ( .A(n4663), .B(n4662), .Z(n1701) );
  XNOR U3542 ( .A(n1700), .B(n1701), .Z(n1702) );
  XNOR U3543 ( .A(n1703), .B(n1702), .Z(n942) );
  XNOR U3544 ( .A(n943), .B(n942), .Z(n2666) );
  XNOR U3545 ( .A(x[863]), .B(y[863]), .Z(n2445) );
  XNOR U3546 ( .A(x[136]), .B(y[136]), .Z(n2442) );
  XNOR U3547 ( .A(x[865]), .B(y[865]), .Z(n2443) );
  XOR U3548 ( .A(n2442), .B(n2443), .Z(n2444) );
  XOR U3549 ( .A(n2445), .B(n2444), .Z(n2281) );
  XNOR U3550 ( .A(x[847]), .B(y[847]), .Z(n3674) );
  XNOR U3551 ( .A(x[849]), .B(y[849]), .Z(n3671) );
  XNOR U3552 ( .A(x[1508]), .B(y[1508]), .Z(n3672) );
  XOR U3553 ( .A(n3671), .B(n3672), .Z(n3673) );
  XNOR U3554 ( .A(n3674), .B(n3673), .Z(n2278) );
  XNOR U3555 ( .A(x[855]), .B(y[855]), .Z(n1633) );
  XNOR U3556 ( .A(x[857]), .B(y[857]), .Z(n1630) );
  XNOR U3557 ( .A(x[1510]), .B(y[1510]), .Z(n1631) );
  XOR U3558 ( .A(n1630), .B(n1631), .Z(n1632) );
  XNOR U3559 ( .A(n1633), .B(n1632), .Z(n2279) );
  XNOR U3560 ( .A(n2281), .B(n2280), .Z(n3800) );
  XNOR U3561 ( .A(x[911]), .B(y[911]), .Z(n3812) );
  XNOR U3562 ( .A(x[913]), .B(y[913]), .Z(n3810) );
  XOR U3563 ( .A(x[1516]), .B(y[1516]), .Z(n3809) );
  XNOR U3564 ( .A(n3810), .B(n3809), .Z(n3811) );
  XOR U3565 ( .A(n3812), .B(n3811), .Z(n2313) );
  XNOR U3566 ( .A(x[903]), .B(y[903]), .Z(n3834) );
  XNOR U3567 ( .A(x[102]), .B(y[102]), .Z(n3832) );
  XOR U3568 ( .A(x[905]), .B(y[905]), .Z(n3831) );
  XNOR U3569 ( .A(n3832), .B(n3831), .Z(n3833) );
  XNOR U3570 ( .A(n3834), .B(n3833), .Z(n2310) );
  XNOR U3571 ( .A(x[895]), .B(y[895]), .Z(n1975) );
  XNOR U3572 ( .A(x[110]), .B(y[110]), .Z(n1972) );
  XNOR U3573 ( .A(x[897]), .B(y[897]), .Z(n1973) );
  XOR U3574 ( .A(n1972), .B(n1973), .Z(n1974) );
  XNOR U3575 ( .A(n1975), .B(n1974), .Z(n2311) );
  XNOR U3576 ( .A(n2313), .B(n2312), .Z(n3797) );
  XNOR U3577 ( .A(x[887]), .B(y[887]), .Z(n3768) );
  XNOR U3578 ( .A(x[889]), .B(y[889]), .Z(n3765) );
  XNOR U3579 ( .A(x[1514]), .B(y[1514]), .Z(n3766) );
  XOR U3580 ( .A(n3765), .B(n3766), .Z(n3767) );
  XOR U3581 ( .A(n3768), .B(n3767), .Z(n2262) );
  XNOR U3582 ( .A(x[879]), .B(y[879]), .Z(n3706) );
  XNOR U3583 ( .A(x[881]), .B(y[881]), .Z(n3703) );
  XNOR U3584 ( .A(x[1512]), .B(y[1512]), .Z(n3704) );
  XOR U3585 ( .A(n3703), .B(n3704), .Z(n3705) );
  XNOR U3586 ( .A(n3706), .B(n3705), .Z(n2260) );
  XNOR U3587 ( .A(x[871]), .B(y[871]), .Z(n2319) );
  XNOR U3588 ( .A(x[130]), .B(y[130]), .Z(n2316) );
  XNOR U3589 ( .A(x[873]), .B(y[873]), .Z(n2317) );
  XOR U3590 ( .A(n2316), .B(n2317), .Z(n2318) );
  XNOR U3591 ( .A(n2319), .B(n2318), .Z(n2261) );
  XOR U3592 ( .A(n2262), .B(n2263), .Z(n3798) );
  XOR U3593 ( .A(n3797), .B(n3798), .Z(n3799) );
  XNOR U3594 ( .A(n3800), .B(n3799), .Z(n2667) );
  XNOR U3595 ( .A(n2666), .B(n2667), .Z(n2668) );
  XNOR U3596 ( .A(n2669), .B(n2668), .Z(n1169) );
  XNOR U3597 ( .A(n1168), .B(n1169), .Z(n1171) );
  XOR U3598 ( .A(n1170), .B(n1171), .Z(n811) );
  XNOR U3599 ( .A(x[497]), .B(y[497]), .Z(n4577) );
  XNOR U3600 ( .A(x[499]), .B(y[499]), .Z(n4574) );
  XNOR U3601 ( .A(x[501]), .B(y[501]), .Z(n4575) );
  XOR U3602 ( .A(n4574), .B(n4575), .Z(n4576) );
  XOR U3603 ( .A(n4577), .B(n4576), .Z(n2799) );
  XNOR U3604 ( .A(x[493]), .B(y[493]), .Z(n4565) );
  XNOR U3605 ( .A(x[76]), .B(y[76]), .Z(n4562) );
  XNOR U3606 ( .A(x[495]), .B(y[495]), .Z(n4563) );
  XOR U3607 ( .A(n4562), .B(n4563), .Z(n4564) );
  XOR U3608 ( .A(n4565), .B(n4564), .Z(n2796) );
  XNOR U3609 ( .A(x[1051]), .B(y[1051]), .Z(n2561) );
  XNOR U3610 ( .A(x[346]), .B(y[346]), .Z(n2558) );
  XNOR U3611 ( .A(x[1053]), .B(y[1053]), .Z(n2559) );
  XOR U3612 ( .A(n2558), .B(n2559), .Z(n2560) );
  XNOR U3613 ( .A(n2561), .B(n2560), .Z(n2797) );
  XNOR U3614 ( .A(n2796), .B(n2797), .Z(n2798) );
  XNOR U3615 ( .A(n2799), .B(n2798), .Z(n1363) );
  XNOR U3616 ( .A(x[489]), .B(y[489]), .Z(n4571) );
  XNOR U3617 ( .A(x[84]), .B(y[84]), .Z(n4568) );
  XNOR U3618 ( .A(x[491]), .B(y[491]), .Z(n4569) );
  XOR U3619 ( .A(n4568), .B(n4569), .Z(n4570) );
  XOR U3620 ( .A(n4571), .B(n4570), .Z(n2805) );
  XNOR U3621 ( .A(x[483]), .B(y[483]), .Z(n4539) );
  XNOR U3622 ( .A(x[485]), .B(y[485]), .Z(n4536) );
  XNOR U3623 ( .A(x[487]), .B(y[487]), .Z(n4537) );
  XOR U3624 ( .A(n4536), .B(n4537), .Z(n4538) );
  XOR U3625 ( .A(n4539), .B(n4538), .Z(n2802) );
  XNOR U3626 ( .A(x[1479]), .B(y[1479]), .Z(n2391) );
  XNOR U3627 ( .A(x[311]), .B(y[311]), .Z(n2388) );
  XNOR U3628 ( .A(x[1481]), .B(y[1481]), .Z(n2389) );
  XOR U3629 ( .A(n2388), .B(n2389), .Z(n2390) );
  XNOR U3630 ( .A(n2391), .B(n2390), .Z(n2803) );
  XNOR U3631 ( .A(n2802), .B(n2803), .Z(n2804) );
  XOR U3632 ( .A(n2805), .B(n2804), .Z(n1362) );
  XOR U3633 ( .A(n1363), .B(n1362), .Z(n1365) );
  XNOR U3634 ( .A(x[477]), .B(y[477]), .Z(n4533) );
  XNOR U3635 ( .A(x[479]), .B(y[479]), .Z(n4530) );
  XNOR U3636 ( .A(x[481]), .B(y[481]), .Z(n4531) );
  XOR U3637 ( .A(n4530), .B(n4531), .Z(n4532) );
  XOR U3638 ( .A(n4533), .B(n4532), .Z(n2973) );
  XNOR U3639 ( .A(x[473]), .B(y[473]), .Z(n4545) );
  XNOR U3640 ( .A(x[112]), .B(y[112]), .Z(n4542) );
  XNOR U3641 ( .A(x[475]), .B(y[475]), .Z(n4543) );
  XOR U3642 ( .A(n4542), .B(n4543), .Z(n4544) );
  XOR U3643 ( .A(n4545), .B(n4544), .Z(n2970) );
  XNOR U3644 ( .A(x[1043]), .B(y[1043]), .Z(n963) );
  XNOR U3645 ( .A(x[13]), .B(y[13]), .Z(n961) );
  XOR U3646 ( .A(x[1045]), .B(y[1045]), .Z(n960) );
  XNOR U3647 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U3648 ( .A(n963), .B(n962), .Z(n2971) );
  XNOR U3649 ( .A(n2970), .B(n2971), .Z(n2972) );
  XNOR U3650 ( .A(n2973), .B(n2972), .Z(n1364) );
  XNOR U3651 ( .A(n1365), .B(n1364), .Z(n4473) );
  XNOR U3652 ( .A(x[449]), .B(y[449]), .Z(n2945) );
  XNOR U3653 ( .A(x[154]), .B(y[154]), .Z(n2943) );
  XOR U3654 ( .A(x[451]), .B(y[451]), .Z(n2942) );
  XNOR U3655 ( .A(n2943), .B(n2942), .Z(n2944) );
  XOR U3656 ( .A(n2945), .B(n2944), .Z(n3508) );
  XNOR U3657 ( .A(x[443]), .B(y[443]), .Z(n2949) );
  XNOR U3658 ( .A(x[445]), .B(y[445]), .Z(n2947) );
  XOR U3659 ( .A(x[447]), .B(y[447]), .Z(n2946) );
  XNOR U3660 ( .A(n2947), .B(n2946), .Z(n2948) );
  XNOR U3661 ( .A(n2949), .B(n2948), .Z(n3505) );
  XNOR U3662 ( .A(x[1487]), .B(y[1487]), .Z(n2181) );
  XNOR U3663 ( .A(x[1489]), .B(y[1489]), .Z(n2178) );
  XNOR U3664 ( .A(x[1588]), .B(y[1588]), .Z(n2179) );
  XOR U3665 ( .A(n2178), .B(n2179), .Z(n2180) );
  XNOR U3666 ( .A(n2181), .B(n2180), .Z(n3506) );
  XNOR U3667 ( .A(n3508), .B(n3507), .Z(n1371) );
  XNOR U3668 ( .A(x[469]), .B(y[469]), .Z(n2967) );
  XNOR U3669 ( .A(x[118]), .B(y[118]), .Z(n2964) );
  XNOR U3670 ( .A(x[471]), .B(y[471]), .Z(n2965) );
  XOR U3671 ( .A(n2964), .B(n2965), .Z(n2966) );
  XOR U3672 ( .A(n2967), .B(n2966), .Z(n2901) );
  XNOR U3673 ( .A(x[463]), .B(y[463]), .Z(n2957) );
  XNOR U3674 ( .A(x[465]), .B(y[465]), .Z(n2954) );
  XNOR U3675 ( .A(x[467]), .B(y[467]), .Z(n2955) );
  XOR U3676 ( .A(n2954), .B(n2955), .Z(n2956) );
  XOR U3677 ( .A(n2957), .B(n2956), .Z(n2898) );
  XNOR U3678 ( .A(x[1483]), .B(y[1483]), .Z(n3624) );
  XNOR U3679 ( .A(x[315]), .B(y[315]), .Z(n3622) );
  XOR U3680 ( .A(x[1485]), .B(y[1485]), .Z(n3621) );
  XNOR U3681 ( .A(n3622), .B(n3621), .Z(n3623) );
  XNOR U3682 ( .A(n3624), .B(n3623), .Z(n2899) );
  XNOR U3683 ( .A(n2898), .B(n2899), .Z(n2900) );
  XNOR U3684 ( .A(n2901), .B(n2900), .Z(n1368) );
  XNOR U3685 ( .A(x[457]), .B(y[457]), .Z(n2963) );
  XNOR U3686 ( .A(x[459]), .B(y[459]), .Z(n2961) );
  XOR U3687 ( .A(x[461]), .B(y[461]), .Z(n2960) );
  XNOR U3688 ( .A(n2961), .B(n2960), .Z(n2962) );
  XOR U3689 ( .A(n2963), .B(n2962), .Z(n2938) );
  XNOR U3690 ( .A(x[453]), .B(y[453]), .Z(n2953) );
  XNOR U3691 ( .A(x[148]), .B(y[148]), .Z(n2951) );
  XOR U3692 ( .A(x[455]), .B(y[455]), .Z(n2950) );
  XNOR U3693 ( .A(n2951), .B(n2950), .Z(n2952) );
  XNOR U3694 ( .A(n2953), .B(n2952), .Z(n2936) );
  XNOR U3695 ( .A(x[1035]), .B(y[1035]), .Z(n953) );
  XNOR U3696 ( .A(x[7]), .B(y[7]), .Z(n951) );
  XOR U3697 ( .A(x[1037]), .B(y[1037]), .Z(n950) );
  XNOR U3698 ( .A(n951), .B(n950), .Z(n952) );
  XNOR U3699 ( .A(n953), .B(n952), .Z(n2937) );
  XOR U3700 ( .A(n2938), .B(n2939), .Z(n1369) );
  XOR U3701 ( .A(n1368), .B(n1369), .Z(n1370) );
  XOR U3702 ( .A(n1371), .B(n1370), .Z(n4470) );
  XNOR U3703 ( .A(x[417]), .B(y[417]), .Z(n2889) );
  XNOR U3704 ( .A(x[419]), .B(y[419]), .Z(n2887) );
  XOR U3705 ( .A(x[421]), .B(y[421]), .Z(n2886) );
  XNOR U3706 ( .A(n2887), .B(n2886), .Z(n2888) );
  XOR U3707 ( .A(n2889), .B(n2888), .Z(n3584) );
  XNOR U3708 ( .A(x[413]), .B(y[413]), .Z(n2893) );
  XNOR U3709 ( .A(x[216]), .B(y[216]), .Z(n2891) );
  XOR U3710 ( .A(x[415]), .B(y[415]), .Z(n2890) );
  XNOR U3711 ( .A(n2891), .B(n2890), .Z(n2892) );
  XOR U3712 ( .A(n2893), .B(n2892), .Z(n3581) );
  XNOR U3713 ( .A(x[1019]), .B(y[1019]), .Z(n1745) );
  XNOR U3714 ( .A(x[366]), .B(y[366]), .Z(n1743) );
  XOR U3715 ( .A(x[1021]), .B(y[1021]), .Z(n1742) );
  XNOR U3716 ( .A(n1743), .B(n1742), .Z(n1744) );
  XNOR U3717 ( .A(n1745), .B(n1744), .Z(n3582) );
  XNOR U3718 ( .A(n3581), .B(n3582), .Z(n3583) );
  XNOR U3719 ( .A(n3584), .B(n3583), .Z(n4033) );
  XNOR U3720 ( .A(x[437]), .B(y[437]), .Z(n2885) );
  XNOR U3721 ( .A(x[439]), .B(y[439]), .Z(n2883) );
  XOR U3722 ( .A(x[441]), .B(y[441]), .Z(n2882) );
  XNOR U3723 ( .A(n2883), .B(n2882), .Z(n2884) );
  XOR U3724 ( .A(n2885), .B(n2884), .Z(n3544) );
  XNOR U3725 ( .A(x[433]), .B(y[433]), .Z(n2877) );
  XNOR U3726 ( .A(x[182]), .B(y[182]), .Z(n2875) );
  XOR U3727 ( .A(x[435]), .B(y[435]), .Z(n2874) );
  XNOR U3728 ( .A(n2875), .B(n2874), .Z(n2876) );
  XOR U3729 ( .A(n2877), .B(n2876), .Z(n3541) );
  XNOR U3730 ( .A(x[1027]), .B(y[1027]), .Z(n949) );
  XNOR U3731 ( .A(x[360]), .B(y[360]), .Z(n947) );
  XOR U3732 ( .A(x[1029]), .B(y[1029]), .Z(n946) );
  XNOR U3733 ( .A(n947), .B(n946), .Z(n948) );
  XNOR U3734 ( .A(n949), .B(n948), .Z(n3542) );
  XNOR U3735 ( .A(n3541), .B(n3542), .Z(n3543) );
  XNOR U3736 ( .A(n3544), .B(n3543), .Z(n4030) );
  XNOR U3737 ( .A(x[429]), .B(y[429]), .Z(n2881) );
  XNOR U3738 ( .A(x[190]), .B(y[190]), .Z(n2879) );
  XOR U3739 ( .A(x[431]), .B(y[431]), .Z(n2878) );
  XNOR U3740 ( .A(n2879), .B(n2878), .Z(n2880) );
  XOR U3741 ( .A(n2881), .B(n2880), .Z(n3415) );
  XNOR U3742 ( .A(x[423]), .B(y[423]), .Z(n2897) );
  XNOR U3743 ( .A(x[425]), .B(y[425]), .Z(n2895) );
  XOR U3744 ( .A(x[427]), .B(y[427]), .Z(n2894) );
  XNOR U3745 ( .A(n2895), .B(n2894), .Z(n2896) );
  XNOR U3746 ( .A(n2897), .B(n2896), .Z(n3413) );
  XNOR U3747 ( .A(x[1491]), .B(y[1491]), .Z(n4125) );
  XNOR U3748 ( .A(x[321]), .B(y[321]), .Z(n4123) );
  XOR U3749 ( .A(x[1493]), .B(y[1493]), .Z(n4122) );
  XNOR U3750 ( .A(n4123), .B(n4122), .Z(n4124) );
  XNOR U3751 ( .A(n4125), .B(n4124), .Z(n3414) );
  XOR U3752 ( .A(n3415), .B(n3416), .Z(n4031) );
  XOR U3753 ( .A(n4030), .B(n4031), .Z(n4032) );
  XNOR U3754 ( .A(n4033), .B(n4032), .Z(n4471) );
  XNOR U3755 ( .A(n4470), .B(n4471), .Z(n4472) );
  XNOR U3756 ( .A(n4473), .B(n4472), .Z(n3587) );
  XNOR U3757 ( .A(x[569]), .B(y[569]), .Z(n4409) );
  XNOR U3758 ( .A(x[376]), .B(y[376]), .Z(n4406) );
  XNOR U3759 ( .A(x[571]), .B(y[571]), .Z(n4407) );
  XOR U3760 ( .A(n4406), .B(n4407), .Z(n4408) );
  XOR U3761 ( .A(n4409), .B(n4408), .Z(n2865) );
  XNOR U3762 ( .A(x[561]), .B(y[561]), .Z(n4295) );
  XNOR U3763 ( .A(x[384]), .B(y[384]), .Z(n4293) );
  XOR U3764 ( .A(x[563]), .B(y[563]), .Z(n4292) );
  XNOR U3765 ( .A(n4293), .B(n4292), .Z(n4294) );
  XOR U3766 ( .A(n4295), .B(n4294), .Z(n2862) );
  XNOR U3767 ( .A(x[565]), .B(y[565]), .Z(n4415) );
  XNOR U3768 ( .A(x[567]), .B(y[567]), .Z(n4412) );
  XNOR U3769 ( .A(x[640]), .B(y[640]), .Z(n4413) );
  XOR U3770 ( .A(n4412), .B(n4413), .Z(n4414) );
  XNOR U3771 ( .A(n4415), .B(n4414), .Z(n2863) );
  XNOR U3772 ( .A(n2862), .B(n2863), .Z(n2864) );
  XNOR U3773 ( .A(n2865), .B(n2864), .Z(n4459) );
  XNOR U3774 ( .A(x[581]), .B(y[581]), .Z(n4331) );
  XNOR U3775 ( .A(x[364]), .B(y[364]), .Z(n4329) );
  XOR U3776 ( .A(x[583]), .B(y[583]), .Z(n4328) );
  XNOR U3777 ( .A(n4329), .B(n4328), .Z(n4330) );
  XOR U3778 ( .A(n4331), .B(n4330), .Z(n3931) );
  XNOR U3779 ( .A(x[573]), .B(y[573]), .Z(n4421) );
  XNOR U3780 ( .A(x[372]), .B(y[372]), .Z(n4419) );
  XOR U3781 ( .A(x[575]), .B(y[575]), .Z(n4418) );
  XNOR U3782 ( .A(n4419), .B(n4418), .Z(n4420) );
  XOR U3783 ( .A(n4421), .B(n4420), .Z(n3928) );
  XNOR U3784 ( .A(x[577]), .B(y[577]), .Z(n4335) );
  XNOR U3785 ( .A(x[579]), .B(y[579]), .Z(n4333) );
  XOR U3786 ( .A(x[1476]), .B(y[1476]), .Z(n4332) );
  XNOR U3787 ( .A(n4333), .B(n4332), .Z(n4334) );
  XNOR U3788 ( .A(n4335), .B(n4334), .Z(n3929) );
  XNOR U3789 ( .A(n3928), .B(n3929), .Z(n3930) );
  XOR U3790 ( .A(n3931), .B(n3930), .Z(n4458) );
  XOR U3791 ( .A(n4459), .B(n4458), .Z(n4461) );
  XNOR U3792 ( .A(x[605]), .B(y[605]), .Z(n4349) );
  XNOR U3793 ( .A(x[356]), .B(y[356]), .Z(n4347) );
  XOR U3794 ( .A(x[607]), .B(y[607]), .Z(n4346) );
  XNOR U3795 ( .A(n4347), .B(n4346), .Z(n4348) );
  XOR U3796 ( .A(n4349), .B(n4348), .Z(n3951) );
  XNOR U3797 ( .A(x[585]), .B(y[585]), .Z(n4339) );
  XNOR U3798 ( .A(x[593]), .B(y[593]), .Z(n4337) );
  XOR U3799 ( .A(x[1478]), .B(y[1478]), .Z(n4336) );
  XNOR U3800 ( .A(n4337), .B(n4336), .Z(n4338) );
  XOR U3801 ( .A(n4339), .B(n4338), .Z(n3948) );
  XNOR U3802 ( .A(x[601]), .B(y[601]), .Z(n4357) );
  XNOR U3803 ( .A(x[603]), .B(y[603]), .Z(n4355) );
  XOR U3804 ( .A(x[626]), .B(y[626]), .Z(n4354) );
  XNOR U3805 ( .A(n4355), .B(n4354), .Z(n4356) );
  XNOR U3806 ( .A(n4357), .B(n4356), .Z(n3949) );
  XNOR U3807 ( .A(n3948), .B(n3949), .Z(n3950) );
  XNOR U3808 ( .A(n3951), .B(n3950), .Z(n4460) );
  XOR U3809 ( .A(n4461), .B(n4460), .Z(n4093) );
  XNOR U3810 ( .A(x[533]), .B(y[533]), .Z(n1237) );
  XNOR U3811 ( .A(x[535]), .B(y[535]), .Z(n1234) );
  XNOR U3812 ( .A(x[660]), .B(y[660]), .Z(n1235) );
  XOR U3813 ( .A(n1234), .B(n1235), .Z(n1236) );
  XOR U3814 ( .A(n1237), .B(n1236), .Z(n2779) );
  XNOR U3815 ( .A(x[529]), .B(y[529]), .Z(n1249) );
  XNOR U3816 ( .A(x[412]), .B(y[412]), .Z(n1246) );
  XNOR U3817 ( .A(x[531]), .B(y[531]), .Z(n1247) );
  XOR U3818 ( .A(n1246), .B(n1247), .Z(n1248) );
  XOR U3819 ( .A(n1249), .B(n1248), .Z(n2776) );
  XNOR U3820 ( .A(x[1067]), .B(y[1067]), .Z(n2573) );
  XNOR U3821 ( .A(x[29]), .B(y[29]), .Z(n2570) );
  XNOR U3822 ( .A(x[1069]), .B(y[1069]), .Z(n2571) );
  XOR U3823 ( .A(n2570), .B(n2571), .Z(n2572) );
  XNOR U3824 ( .A(n2573), .B(n2572), .Z(n2777) );
  XNOR U3825 ( .A(n2776), .B(n2777), .Z(n2778) );
  XNOR U3826 ( .A(n2779), .B(n2778), .Z(n1410) );
  XNOR U3827 ( .A(x[557]), .B(y[557]), .Z(n4299) );
  XNOR U3828 ( .A(x[559]), .B(y[559]), .Z(n4297) );
  XOR U3829 ( .A(x[646]), .B(y[646]), .Z(n4296) );
  XNOR U3830 ( .A(n4297), .B(n4296), .Z(n4298) );
  XOR U3831 ( .A(n4299), .B(n4298), .Z(n3981) );
  XNOR U3832 ( .A(x[549]), .B(y[549]), .Z(n4283) );
  XNOR U3833 ( .A(x[392]), .B(y[392]), .Z(n4281) );
  XOR U3834 ( .A(x[551]), .B(y[551]), .Z(n4280) );
  XNOR U3835 ( .A(n4281), .B(n4280), .Z(n4282) );
  XOR U3836 ( .A(n4283), .B(n4282), .Z(n3978) );
  XNOR U3837 ( .A(x[553]), .B(y[553]), .Z(n4291) );
  XNOR U3838 ( .A(x[555]), .B(y[555]), .Z(n4289) );
  XOR U3839 ( .A(x[1474]), .B(y[1474]), .Z(n4288) );
  XNOR U3840 ( .A(n4289), .B(n4288), .Z(n4290) );
  XNOR U3841 ( .A(n4291), .B(n4290), .Z(n3979) );
  XNOR U3842 ( .A(n3978), .B(n3979), .Z(n3980) );
  XNOR U3843 ( .A(n3981), .B(n3980), .Z(n1409) );
  XNOR U3844 ( .A(x[545]), .B(y[545]), .Z(n4287) );
  XNOR U3845 ( .A(x[547]), .B(y[547]), .Z(n4285) );
  XOR U3846 ( .A(x[1472]), .B(y[1472]), .Z(n4284) );
  XNOR U3847 ( .A(n4285), .B(n4284), .Z(n4286) );
  XOR U3848 ( .A(n4287), .B(n4286), .Z(n3957) );
  XNOR U3849 ( .A(x[537]), .B(y[537]), .Z(n1243) );
  XNOR U3850 ( .A(x[404]), .B(y[404]), .Z(n1240) );
  XNOR U3851 ( .A(x[539]), .B(y[539]), .Z(n1241) );
  XOR U3852 ( .A(n1240), .B(n1241), .Z(n1242) );
  XOR U3853 ( .A(n1243), .B(n1242), .Z(n3954) );
  XNOR U3854 ( .A(x[541]), .B(y[541]), .Z(n4279) );
  XNOR U3855 ( .A(x[398]), .B(y[398]), .Z(n4277) );
  XOR U3856 ( .A(x[543]), .B(y[543]), .Z(n4276) );
  XNOR U3857 ( .A(n4277), .B(n4276), .Z(n4278) );
  XNOR U3858 ( .A(n4279), .B(n4278), .Z(n3955) );
  XNOR U3859 ( .A(n3954), .B(n3955), .Z(n3956) );
  XOR U3860 ( .A(n3957), .B(n3956), .Z(n1408) );
  XOR U3861 ( .A(n1409), .B(n1408), .Z(n1411) );
  XOR U3862 ( .A(n1410), .B(n1411), .Z(n4090) );
  XNOR U3863 ( .A(x[509]), .B(y[509]), .Z(n4623) );
  XNOR U3864 ( .A(x[50]), .B(y[50]), .Z(n4621) );
  XOR U3865 ( .A(x[511]), .B(y[511]), .Z(n4620) );
  XNOR U3866 ( .A(n4621), .B(n4620), .Z(n4622) );
  XOR U3867 ( .A(n4623), .B(n4622), .Z(n2835) );
  XNOR U3868 ( .A(x[503]), .B(y[503]), .Z(n4627) );
  XNOR U3869 ( .A(x[505]), .B(y[505]), .Z(n4625) );
  XOR U3870 ( .A(x[507]), .B(y[507]), .Z(n4624) );
  XNOR U3871 ( .A(n4625), .B(n4624), .Z(n4626) );
  XNOR U3872 ( .A(n4627), .B(n4626), .Z(n2832) );
  XNOR U3873 ( .A(x[1475]), .B(y[1475]), .Z(n2405) );
  XNOR U3874 ( .A(x[80]), .B(y[80]), .Z(n2403) );
  XOR U3875 ( .A(x[1477]), .B(y[1477]), .Z(n2402) );
  XNOR U3876 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3877 ( .A(n2405), .B(n2404), .Z(n2833) );
  XNOR U3878 ( .A(n2835), .B(n2834), .Z(n1485) );
  XNOR U3879 ( .A(x[1059]), .B(y[1059]), .Z(n2567) );
  XNOR U3880 ( .A(x[340]), .B(y[340]), .Z(n2564) );
  XNOR U3881 ( .A(x[1061]), .B(y[1061]), .Z(n2565) );
  XOR U3882 ( .A(n2564), .B(n2565), .Z(n2566) );
  XOR U3883 ( .A(n2567), .B(n2566), .Z(n2827) );
  XNOR U3884 ( .A(x[513]), .B(y[513]), .Z(n4631) );
  XNOR U3885 ( .A(x[515]), .B(y[515]), .Z(n4629) );
  XOR U3886 ( .A(x[1468]), .B(y[1468]), .Z(n4628) );
  XNOR U3887 ( .A(n4629), .B(n4628), .Z(n4630) );
  XNOR U3888 ( .A(n4631), .B(n4630), .Z(n2826) );
  XOR U3889 ( .A(n2827), .B(n2826), .Z(n2829) );
  XNOR U3890 ( .A(x[517]), .B(y[517]), .Z(n1227) );
  XNOR U3891 ( .A(x[418]), .B(y[418]), .Z(n1225) );
  XOR U3892 ( .A(x[519]), .B(y[519]), .Z(n1224) );
  XNOR U3893 ( .A(n1225), .B(n1224), .Z(n1226) );
  XNOR U3894 ( .A(n1227), .B(n1226), .Z(n2828) );
  XNOR U3895 ( .A(x[525]), .B(y[525]), .Z(n1231) );
  XNOR U3896 ( .A(x[527]), .B(y[527]), .Z(n1228) );
  XNOR U3897 ( .A(x[666]), .B(y[666]), .Z(n1229) );
  XOR U3898 ( .A(n1228), .B(n1229), .Z(n1230) );
  XOR U3899 ( .A(n1231), .B(n1230), .Z(n2761) );
  XNOR U3900 ( .A(x[521]), .B(y[521]), .Z(n1221) );
  XNOR U3901 ( .A(x[523]), .B(y[523]), .Z(n1218) );
  XNOR U3902 ( .A(x[1470]), .B(y[1470]), .Z(n1219) );
  XOR U3903 ( .A(n1218), .B(n1219), .Z(n1220) );
  XOR U3904 ( .A(n1221), .B(n1220), .Z(n2758) );
  XNOR U3905 ( .A(x[1471]), .B(y[1471]), .Z(n2287) );
  XNOR U3906 ( .A(x[305]), .B(y[305]), .Z(n2285) );
  XOR U3907 ( .A(x[1473]), .B(y[1473]), .Z(n2284) );
  XNOR U3908 ( .A(n2285), .B(n2284), .Z(n2286) );
  XNOR U3909 ( .A(n2287), .B(n2286), .Z(n2759) );
  XNOR U3910 ( .A(n2758), .B(n2759), .Z(n2760) );
  XNOR U3911 ( .A(n2761), .B(n2760), .Z(n1483) );
  XOR U3912 ( .A(n1482), .B(n1483), .Z(n1484) );
  XNOR U3913 ( .A(n1485), .B(n1484), .Z(n4091) );
  XOR U3914 ( .A(n4090), .B(n4091), .Z(n4092) );
  XNOR U3915 ( .A(n4093), .B(n4092), .Z(n3588) );
  XNOR U3916 ( .A(n3587), .B(n3588), .Z(n3589) );
  XNOR U3917 ( .A(x[389]), .B(y[389]), .Z(n2907) );
  XNOR U3918 ( .A(x[258]), .B(y[258]), .Z(n2905) );
  XOR U3919 ( .A(x[391]), .B(y[391]), .Z(n2904) );
  XNOR U3920 ( .A(n2905), .B(n2904), .Z(n2906) );
  XOR U3921 ( .A(n2907), .B(n2906), .Z(n3438) );
  XNOR U3922 ( .A(x[383]), .B(y[383]), .Z(n2911) );
  XNOR U3923 ( .A(x[385]), .B(y[385]), .Z(n2909) );
  XOR U3924 ( .A(x[387]), .B(y[387]), .Z(n2908) );
  XNOR U3925 ( .A(n2909), .B(n2908), .Z(n2910) );
  XNOR U3926 ( .A(n2911), .B(n2910), .Z(n3435) );
  XNOR U3927 ( .A(x[1499]), .B(y[1499]), .Z(n4219) );
  XNOR U3928 ( .A(x[66]), .B(y[66]), .Z(n4217) );
  XOR U3929 ( .A(x[1501]), .B(y[1501]), .Z(n4216) );
  XNOR U3930 ( .A(n4217), .B(n4216), .Z(n4218) );
  XNOR U3931 ( .A(n4219), .B(n4218), .Z(n3436) );
  XNOR U3932 ( .A(n3438), .B(n3437), .Z(n1448) );
  XNOR U3933 ( .A(x[409]), .B(y[409]), .Z(n2933) );
  XNOR U3934 ( .A(x[224]), .B(y[224]), .Z(n2930) );
  XNOR U3935 ( .A(x[411]), .B(y[411]), .Z(n2931) );
  XOR U3936 ( .A(n2930), .B(n2931), .Z(n2932) );
  XOR U3937 ( .A(n2933), .B(n2932), .Z(n3466) );
  XNOR U3938 ( .A(x[403]), .B(y[403]), .Z(n2921) );
  XNOR U3939 ( .A(x[405]), .B(y[405]), .Z(n2918) );
  XNOR U3940 ( .A(x[407]), .B(y[407]), .Z(n2919) );
  XOR U3941 ( .A(n2918), .B(n2919), .Z(n2920) );
  XOR U3942 ( .A(n2921), .B(n2920), .Z(n3463) );
  XNOR U3943 ( .A(x[1495]), .B(y[1495]), .Z(n2115) );
  XNOR U3944 ( .A(x[1497]), .B(y[1497]), .Z(n2112) );
  XNOR U3945 ( .A(x[1590]), .B(y[1590]), .Z(n2113) );
  XOR U3946 ( .A(n2112), .B(n2113), .Z(n2114) );
  XNOR U3947 ( .A(n2115), .B(n2114), .Z(n3464) );
  XNOR U3948 ( .A(n3463), .B(n3464), .Z(n3465) );
  XNOR U3949 ( .A(n3466), .B(n3465), .Z(n1447) );
  XNOR U3950 ( .A(x[397]), .B(y[397]), .Z(n2927) );
  XNOR U3951 ( .A(x[399]), .B(y[399]), .Z(n2924) );
  XNOR U3952 ( .A(x[401]), .B(y[401]), .Z(n2925) );
  XOR U3953 ( .A(n2924), .B(n2925), .Z(n2926) );
  XOR U3954 ( .A(n2927), .B(n2926), .Z(n3444) );
  XNOR U3955 ( .A(x[393]), .B(y[393]), .Z(n2915) );
  XNOR U3956 ( .A(x[252]), .B(y[252]), .Z(n2912) );
  XNOR U3957 ( .A(x[395]), .B(y[395]), .Z(n2913) );
  XOR U3958 ( .A(n2912), .B(n2913), .Z(n2914) );
  XOR U3959 ( .A(n2915), .B(n2914), .Z(n3441) );
  XNOR U3960 ( .A(x[1011]), .B(y[1011]), .Z(n2521) );
  XNOR U3961 ( .A(x[8]), .B(y[8]), .Z(n2518) );
  XNOR U3962 ( .A(x[1013]), .B(y[1013]), .Z(n2519) );
  XOR U3963 ( .A(n2518), .B(n2519), .Z(n2520) );
  XNOR U3964 ( .A(n2521), .B(n2520), .Z(n3442) );
  XNOR U3965 ( .A(n3441), .B(n3442), .Z(n3443) );
  XOR U3966 ( .A(n3444), .B(n3443), .Z(n1446) );
  XOR U3967 ( .A(n1447), .B(n1446), .Z(n1449) );
  XOR U3968 ( .A(n1448), .B(n1449), .Z(n1346) );
  XNOR U3969 ( .A(x[319]), .B(y[319]), .Z(n2785) );
  XNOR U3970 ( .A(x[323]), .B(y[323]), .Z(n2782) );
  XNOR U3971 ( .A(x[325]), .B(y[325]), .Z(n2783) );
  XOR U3972 ( .A(n2782), .B(n2783), .Z(n2784) );
  XOR U3973 ( .A(n2785), .B(n2784), .Z(n3362) );
  XNOR U3974 ( .A(x[303]), .B(y[303]), .Z(n2823) );
  XNOR U3975 ( .A(x[307]), .B(y[307]), .Z(n2820) );
  XNOR U3976 ( .A(x[358]), .B(y[358]), .Z(n2821) );
  XOR U3977 ( .A(n2820), .B(n2821), .Z(n2822) );
  XOR U3978 ( .A(n2823), .B(n2822), .Z(n3359) );
  XNOR U3979 ( .A(x[1507]), .B(y[1507]), .Z(n1391) );
  XNOR U3980 ( .A(x[60]), .B(y[60]), .Z(n1388) );
  XNOR U3981 ( .A(x[1509]), .B(y[1509]), .Z(n1389) );
  XOR U3982 ( .A(n1388), .B(n1389), .Z(n1390) );
  XNOR U3983 ( .A(n1391), .B(n1390), .Z(n3360) );
  XNOR U3984 ( .A(n3359), .B(n3360), .Z(n3361) );
  XNOR U3985 ( .A(n3362), .B(n3361), .Z(n3600) );
  XNOR U3986 ( .A(x[297]), .B(y[297]), .Z(n2811) );
  XNOR U3987 ( .A(x[301]), .B(y[301]), .Z(n2808) );
  XNOR U3988 ( .A(x[368]), .B(y[368]), .Z(n2809) );
  XOR U3989 ( .A(n2808), .B(n2809), .Z(n2810) );
  XOR U3990 ( .A(n2811), .B(n2810), .Z(n3263) );
  XNOR U3991 ( .A(x[287]), .B(y[287]), .Z(n2817) );
  XNOR U3992 ( .A(x[291]), .B(y[291]), .Z(n2814) );
  XNOR U3993 ( .A(x[295]), .B(y[295]), .Z(n2815) );
  XOR U3994 ( .A(n2814), .B(n2815), .Z(n2816) );
  XOR U3995 ( .A(n2817), .B(n2816), .Z(n3260) );
  XNOR U3996 ( .A(x[987]), .B(y[987]), .Z(n2549) );
  XNOR U3997 ( .A(x[386]), .B(y[386]), .Z(n2546) );
  XNOR U3998 ( .A(x[989]), .B(y[989]), .Z(n2547) );
  XOR U3999 ( .A(n2546), .B(n2547), .Z(n2548) );
  XNOR U4000 ( .A(n2549), .B(n2548), .Z(n3261) );
  XNOR U4001 ( .A(n3260), .B(n3261), .Z(n3262) );
  XOR U4002 ( .A(n3263), .B(n3262), .Z(n3599) );
  XNOR U4003 ( .A(n3600), .B(n3599), .Z(n3601) );
  XNOR U4004 ( .A(x[279]), .B(y[279]), .Z(n2775) );
  XNOR U4005 ( .A(x[281]), .B(y[281]), .Z(n2773) );
  XOR U4006 ( .A(x[285]), .B(y[285]), .Z(n2772) );
  XNOR U4007 ( .A(n2773), .B(n2772), .Z(n2774) );
  XOR U4008 ( .A(n2775), .B(n2774), .Z(n3356) );
  XNOR U4009 ( .A(x[273]), .B(y[273]), .Z(n2767) );
  XNOR U4010 ( .A(x[275]), .B(y[275]), .Z(n2765) );
  XOR U4011 ( .A(x[394]), .B(y[394]), .Z(n2764) );
  XNOR U4012 ( .A(n2765), .B(n2764), .Z(n2766) );
  XOR U4013 ( .A(n2767), .B(n2766), .Z(n3353) );
  XNOR U4014 ( .A(x[1511]), .B(y[1511]), .Z(n3650) );
  XNOR U4015 ( .A(x[333]), .B(y[333]), .Z(n3647) );
  XNOR U4016 ( .A(x[1513]), .B(y[1513]), .Z(n3648) );
  XOR U4017 ( .A(n3647), .B(n3648), .Z(n3649) );
  XNOR U4018 ( .A(n3650), .B(n3649), .Z(n3354) );
  XNOR U4019 ( .A(n3353), .B(n3354), .Z(n3355) );
  XOR U4020 ( .A(n3356), .B(n3355), .Z(n3602) );
  XOR U4021 ( .A(n3601), .B(n3602), .Z(n1344) );
  XNOR U4022 ( .A(x[373]), .B(y[373]), .Z(n3484) );
  XNOR U4023 ( .A(x[375]), .B(y[375]), .Z(n3481) );
  XNOR U4024 ( .A(x[379]), .B(y[379]), .Z(n3482) );
  XOR U4025 ( .A(n3481), .B(n3482), .Z(n3483) );
  XOR U4026 ( .A(n3484), .B(n3483), .Z(n3382) );
  XNOR U4027 ( .A(x[367]), .B(y[367]), .Z(n3472) );
  XNOR U4028 ( .A(x[288]), .B(y[288]), .Z(n3469) );
  XNOR U4029 ( .A(x[369]), .B(y[369]), .Z(n3470) );
  XOR U4030 ( .A(n3469), .B(n3470), .Z(n3471) );
  XOR U4031 ( .A(n3472), .B(n3471), .Z(n3379) );
  XNOR U4032 ( .A(x[1003]), .B(y[1003]), .Z(n2369) );
  XNOR U4033 ( .A(x[14]), .B(y[14]), .Z(n2366) );
  XNOR U4034 ( .A(x[1005]), .B(y[1005]), .Z(n2367) );
  XOR U4035 ( .A(n2366), .B(n2367), .Z(n2368) );
  XNOR U4036 ( .A(n2369), .B(n2368), .Z(n3380) );
  XNOR U4037 ( .A(n3379), .B(n3380), .Z(n3381) );
  XNOR U4038 ( .A(n3382), .B(n3381), .Z(n1415) );
  XNOR U4039 ( .A(x[361]), .B(y[361]), .Z(n3478) );
  XNOR U4040 ( .A(x[296]), .B(y[296]), .Z(n3475) );
  XNOR U4041 ( .A(x[363]), .B(y[363]), .Z(n3476) );
  XOR U4042 ( .A(n3475), .B(n3476), .Z(n3477) );
  XOR U4043 ( .A(n3478), .B(n3477), .Z(n3404) );
  XNOR U4044 ( .A(x[351]), .B(y[351]), .Z(n3502) );
  XNOR U4045 ( .A(x[353]), .B(y[353]), .Z(n3499) );
  XNOR U4046 ( .A(x[357]), .B(y[357]), .Z(n3500) );
  XOR U4047 ( .A(n3499), .B(n3500), .Z(n3501) );
  XOR U4048 ( .A(n3502), .B(n3501), .Z(n3401) );
  XNOR U4049 ( .A(x[1503]), .B(y[1503]), .Z(n4013) );
  XNOR U4050 ( .A(x[327]), .B(y[327]), .Z(n4010) );
  XNOR U4051 ( .A(x[1505]), .B(y[1505]), .Z(n4011) );
  XOR U4052 ( .A(n4010), .B(n4011), .Z(n4012) );
  XNOR U4053 ( .A(n4013), .B(n4012), .Z(n3402) );
  XNOR U4054 ( .A(n3401), .B(n3402), .Z(n3403) );
  XOR U4055 ( .A(n3404), .B(n3403), .Z(n1414) );
  XNOR U4056 ( .A(n1415), .B(n1414), .Z(n1416) );
  XNOR U4057 ( .A(x[341]), .B(y[341]), .Z(n3490) );
  XNOR U4058 ( .A(x[345]), .B(y[345]), .Z(n3487) );
  XNOR U4059 ( .A(x[347]), .B(y[347]), .Z(n3488) );
  XOR U4060 ( .A(n3487), .B(n3488), .Z(n3489) );
  XOR U4061 ( .A(n3490), .B(n3489), .Z(n3410) );
  XNOR U4062 ( .A(x[335]), .B(y[335]), .Z(n3496) );
  XNOR U4063 ( .A(x[324]), .B(y[324]), .Z(n3493) );
  XNOR U4064 ( .A(x[339]), .B(y[339]), .Z(n3494) );
  XOR U4065 ( .A(n3493), .B(n3494), .Z(n3495) );
  XOR U4066 ( .A(n3496), .B(n3495), .Z(n3407) );
  XNOR U4067 ( .A(x[995]), .B(y[995]), .Z(n2539) );
  XNOR U4068 ( .A(x[380]), .B(y[380]), .Z(n2537) );
  XOR U4069 ( .A(x[997]), .B(y[997]), .Z(n2536) );
  XNOR U4070 ( .A(n2537), .B(n2536), .Z(n2538) );
  XNOR U4071 ( .A(n2539), .B(n2538), .Z(n3408) );
  XNOR U4072 ( .A(n3407), .B(n3408), .Z(n3409) );
  XOR U4073 ( .A(n3410), .B(n3409), .Z(n1417) );
  XOR U4074 ( .A(n1416), .B(n1417), .Z(n1345) );
  XOR U4075 ( .A(n1344), .B(n1345), .Z(n1347) );
  XOR U4076 ( .A(n1346), .B(n1347), .Z(n3590) );
  XOR U4077 ( .A(n3589), .B(n3590), .Z(n808) );
  XNOR U4078 ( .A(x[816]), .B(y[816]), .Z(n1917) );
  XNOR U4079 ( .A(x[814]), .B(y[814]), .Z(n1915) );
  XOR U4080 ( .A(x[1146]), .B(y[1146]), .Z(n1914) );
  XNOR U4081 ( .A(n1915), .B(n1914), .Z(n1916) );
  XOR U4082 ( .A(n1917), .B(n1916), .Z(n1071) );
  XNOR U4083 ( .A(x[828]), .B(y[828]), .Z(n1913) );
  XNOR U4084 ( .A(x[826]), .B(y[826]), .Z(n1911) );
  XOR U4085 ( .A(x[1150]), .B(y[1150]), .Z(n1910) );
  XNOR U4086 ( .A(n1911), .B(n1910), .Z(n1912) );
  XOR U4087 ( .A(n1913), .B(n1912), .Z(n1068) );
  XNOR U4088 ( .A(x[824]), .B(y[824]), .Z(n1909) );
  XNOR U4089 ( .A(x[820]), .B(y[820]), .Z(n1907) );
  XOR U4090 ( .A(x[1428]), .B(y[1428]), .Z(n1906) );
  XNOR U4091 ( .A(n1907), .B(n1906), .Z(n1908) );
  XNOR U4092 ( .A(n1909), .B(n1908), .Z(n1069) );
  XNOR U4093 ( .A(n1068), .B(n1069), .Z(n1070) );
  XNOR U4094 ( .A(n1071), .B(n1070), .Z(n2155) );
  XNOR U4095 ( .A(x[1314]), .B(y[1314]), .Z(n1295) );
  XNOR U4096 ( .A(x[1322]), .B(y[1322]), .Z(n1293) );
  XNOR U4097 ( .A(x[1358]), .B(y[1358]), .Z(n1292) );
  XNOR U4098 ( .A(n1293), .B(n1292), .Z(n1294) );
  XNOR U4099 ( .A(n1295), .B(n1294), .Z(n2259) );
  XNOR U4100 ( .A(x[1354]), .B(y[1354]), .Z(n1289) );
  XNOR U4101 ( .A(x[1342]), .B(y[1342]), .Z(n1287) );
  XNOR U4102 ( .A(x[1356]), .B(y[1356]), .Z(n1286) );
  XNOR U4103 ( .A(n1287), .B(n1286), .Z(n1288) );
  XNOR U4104 ( .A(n1289), .B(n1288), .Z(n2256) );
  XNOR U4105 ( .A(x[548]), .B(y[548]), .Z(n4223) );
  XNOR U4106 ( .A(x[542]), .B(y[542]), .Z(n4221) );
  XOR U4107 ( .A(x[840]), .B(y[840]), .Z(n4220) );
  XNOR U4108 ( .A(n4221), .B(n4220), .Z(n4222) );
  XNOR U4109 ( .A(n4223), .B(n4222), .Z(n2257) );
  XNOR U4110 ( .A(n2256), .B(n2257), .Z(n2258) );
  XOR U4111 ( .A(n2259), .B(n2258), .Z(n2154) );
  XOR U4112 ( .A(n2155), .B(n2154), .Z(n2157) );
  XNOR U4113 ( .A(x[832]), .B(y[832]), .Z(n1085) );
  XNOR U4114 ( .A(x[830]), .B(y[830]), .Z(n1083) );
  XOR U4115 ( .A(x[1426]), .B(y[1426]), .Z(n1082) );
  XNOR U4116 ( .A(n1083), .B(n1082), .Z(n1084) );
  XOR U4117 ( .A(n1085), .B(n1084), .Z(n2217) );
  XNOR U4118 ( .A(x[844]), .B(y[844]), .Z(n1081) );
  XNOR U4119 ( .A(x[842]), .B(y[842]), .Z(n1079) );
  XOR U4120 ( .A(x[1424]), .B(y[1424]), .Z(n1078) );
  XNOR U4121 ( .A(n1079), .B(n1078), .Z(n1080) );
  XOR U4122 ( .A(n1081), .B(n1080), .Z(n2214) );
  XNOR U4123 ( .A(x[838]), .B(y[838]), .Z(n1077) );
  XNOR U4124 ( .A(x[834]), .B(y[834]), .Z(n1075) );
  XOR U4125 ( .A(x[1154]), .B(y[1154]), .Z(n1074) );
  XNOR U4126 ( .A(n1075), .B(n1074), .Z(n1076) );
  XNOR U4127 ( .A(n1077), .B(n1076), .Z(n2215) );
  XNOR U4128 ( .A(n2214), .B(n2215), .Z(n2216) );
  XNOR U4129 ( .A(n2217), .B(n2216), .Z(n2156) );
  XNOR U4130 ( .A(n2157), .B(n2156), .Z(n1491) );
  XNOR U4131 ( .A(x[868]), .B(y[868]), .Z(n859) );
  XNOR U4132 ( .A(x[866]), .B(y[866]), .Z(n857) );
  XOR U4133 ( .A(x[1166]), .B(y[1166]), .Z(n856) );
  XNOR U4134 ( .A(n857), .B(n856), .Z(n858) );
  XOR U4135 ( .A(n859), .B(n858), .Z(n3033) );
  XNOR U4136 ( .A(x[878]), .B(y[878]), .Z(n855) );
  XNOR U4137 ( .A(x[876]), .B(y[876]), .Z(n853) );
  XOR U4138 ( .A(x[1170]), .B(y[1170]), .Z(n852) );
  XNOR U4139 ( .A(n853), .B(n852), .Z(n854) );
  XOR U4140 ( .A(n855), .B(n854), .Z(n3030) );
  XNOR U4141 ( .A(x[874]), .B(y[874]), .Z(n851) );
  XNOR U4142 ( .A(x[870]), .B(y[870]), .Z(n849) );
  XOR U4143 ( .A(x[1418]), .B(y[1418]), .Z(n848) );
  XNOR U4144 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U4145 ( .A(n851), .B(n850), .Z(n3031) );
  XNOR U4146 ( .A(n3030), .B(n3031), .Z(n3032) );
  XNOR U4147 ( .A(n3033), .B(n3032), .Z(n4147) );
  XNOR U4148 ( .A(x[1366]), .B(y[1366]), .Z(n1857) );
  XNOR U4149 ( .A(x[1282]), .B(y[1282]), .Z(n1855) );
  XOR U4150 ( .A(x[1326]), .B(y[1326]), .Z(n1854) );
  XNOR U4151 ( .A(n1855), .B(n1854), .Z(n1856) );
  XOR U4152 ( .A(n1857), .B(n1856), .Z(n1517) );
  XNOR U4153 ( .A(x[1286]), .B(y[1286]), .Z(n1853) );
  XNOR U4154 ( .A(x[1284]), .B(y[1284]), .Z(n1851) );
  XOR U4155 ( .A(x[1320]), .B(y[1320]), .Z(n1850) );
  XNOR U4156 ( .A(n1851), .B(n1850), .Z(n1852) );
  XOR U4157 ( .A(n1853), .B(n1852), .Z(n1514) );
  XNOR U4158 ( .A(x[1362]), .B(y[1362]), .Z(n1849) );
  XNOR U4159 ( .A(x[1324]), .B(y[1324]), .Z(n1847) );
  XOR U4160 ( .A(x[1364]), .B(y[1364]), .Z(n1846) );
  XNOR U4161 ( .A(n1847), .B(n1846), .Z(n1848) );
  XNOR U4162 ( .A(n1849), .B(n1848), .Z(n1515) );
  XNOR U4163 ( .A(n1514), .B(n1515), .Z(n1516) );
  XOR U4164 ( .A(n1517), .B(n1516), .Z(n4146) );
  XOR U4165 ( .A(n4147), .B(n4146), .Z(n4149) );
  XNOR U4166 ( .A(x[882]), .B(y[882]), .Z(n1145) );
  XNOR U4167 ( .A(x[880]), .B(y[880]), .Z(n1143) );
  XOR U4168 ( .A(x[1416]), .B(y[1416]), .Z(n1142) );
  XNOR U4169 ( .A(n1143), .B(n1142), .Z(n1144) );
  XOR U4170 ( .A(n1145), .B(n1144), .Z(n2979) );
  XNOR U4171 ( .A(x[890]), .B(y[890]), .Z(n1141) );
  XNOR U4172 ( .A(x[888]), .B(y[888]), .Z(n1139) );
  XOR U4173 ( .A(x[1414]), .B(y[1414]), .Z(n1138) );
  XNOR U4174 ( .A(n1139), .B(n1138), .Z(n1140) );
  XOR U4175 ( .A(n1141), .B(n1140), .Z(n2976) );
  XNOR U4176 ( .A(x[886]), .B(y[886]), .Z(n1137) );
  XNOR U4177 ( .A(x[884]), .B(y[884]), .Z(n1135) );
  XOR U4178 ( .A(x[1174]), .B(y[1174]), .Z(n1134) );
  XNOR U4179 ( .A(n1135), .B(n1134), .Z(n1136) );
  XNOR U4180 ( .A(n1137), .B(n1136), .Z(n2977) );
  XNOR U4181 ( .A(n2976), .B(n2977), .Z(n2978) );
  XNOR U4182 ( .A(n2979), .B(n2978), .Z(n4148) );
  XNOR U4183 ( .A(n4149), .B(n4148), .Z(n1488) );
  XNOR U4184 ( .A(x[1294]), .B(y[1294]), .Z(n4639) );
  XNOR U4185 ( .A(x[1318]), .B(y[1318]), .Z(n4637) );
  XOR U4186 ( .A(x[1360]), .B(y[1360]), .Z(n4636) );
  XNOR U4187 ( .A(n4637), .B(n4636), .Z(n4638) );
  XOR U4188 ( .A(n4639), .B(n4638), .Z(n4943) );
  XNOR U4189 ( .A(x[1312]), .B(y[1312]), .Z(n4635) );
  XNOR U4190 ( .A(x[1298]), .B(y[1298]), .Z(n4633) );
  XOR U4191 ( .A(x[1316]), .B(y[1316]), .Z(n4632) );
  XNOR U4192 ( .A(n4633), .B(n4632), .Z(n4634) );
  XOR U4193 ( .A(n4635), .B(n4634), .Z(n4940) );
  XNOR U4194 ( .A(x[532]), .B(y[532]), .Z(n4227) );
  XNOR U4195 ( .A(x[528]), .B(y[528]), .Z(n4225) );
  XOR U4196 ( .A(x[530]), .B(y[530]), .Z(n4224) );
  XNOR U4197 ( .A(n4225), .B(n4224), .Z(n4226) );
  XNOR U4198 ( .A(n4227), .B(n4226), .Z(n4941) );
  XNOR U4199 ( .A(n4940), .B(n4941), .Z(n4942) );
  XNOR U4200 ( .A(n4943), .B(n4942), .Z(n4095) );
  XNOR U4201 ( .A(x[848]), .B(y[848]), .Z(n1905) );
  XNOR U4202 ( .A(x[846]), .B(y[846]), .Z(n1903) );
  XOR U4203 ( .A(x[1158]), .B(y[1158]), .Z(n1902) );
  XNOR U4204 ( .A(n1903), .B(n1902), .Z(n1904) );
  XOR U4205 ( .A(n1905), .B(n1904), .Z(n829) );
  XNOR U4206 ( .A(x[852]), .B(y[852]), .Z(n1901) );
  XNOR U4207 ( .A(x[850]), .B(y[850]), .Z(n1899) );
  XOR U4208 ( .A(x[1422]), .B(y[1422]), .Z(n1898) );
  XNOR U4209 ( .A(n1899), .B(n1898), .Z(n1900) );
  XOR U4210 ( .A(n1901), .B(n1900), .Z(n826) );
  XNOR U4211 ( .A(x[185]), .B(y[185]), .Z(n2857) );
  XNOR U4212 ( .A(x[187]), .B(y[187]), .Z(n2855) );
  XOR U4213 ( .A(x[191]), .B(y[191]), .Z(n2854) );
  XNOR U4214 ( .A(n2855), .B(n2854), .Z(n2856) );
  XNOR U4215 ( .A(n2857), .B(n2856), .Z(n827) );
  XNOR U4216 ( .A(n826), .B(n827), .Z(n828) );
  XOR U4217 ( .A(n829), .B(n828), .Z(n4094) );
  XOR U4218 ( .A(n4095), .B(n4094), .Z(n4097) );
  XNOR U4219 ( .A(x[860]), .B(y[860]), .Z(n871) );
  XNOR U4220 ( .A(x[856]), .B(y[856]), .Z(n869) );
  XOR U4221 ( .A(x[1162]), .B(y[1162]), .Z(n868) );
  XNOR U4222 ( .A(n869), .B(n868), .Z(n870) );
  XOR U4223 ( .A(n871), .B(n870), .Z(n2711) );
  XNOR U4224 ( .A(x[864]), .B(y[864]), .Z(n867) );
  XNOR U4225 ( .A(x[862]), .B(y[862]), .Z(n865) );
  XOR U4226 ( .A(x[1420]), .B(y[1420]), .Z(n864) );
  XNOR U4227 ( .A(n865), .B(n864), .Z(n866) );
  XOR U4228 ( .A(n867), .B(n866), .Z(n2708) );
  XNOR U4229 ( .A(x[171]), .B(y[171]), .Z(n3945) );
  XNOR U4230 ( .A(x[175]), .B(y[175]), .Z(n3942) );
  XNOR U4231 ( .A(x[476]), .B(y[476]), .Z(n3943) );
  XOR U4232 ( .A(n3942), .B(n3943), .Z(n3944) );
  XNOR U4233 ( .A(n3945), .B(n3944), .Z(n2709) );
  XNOR U4234 ( .A(n2708), .B(n2709), .Z(n2710) );
  XNOR U4235 ( .A(n2711), .B(n2710), .Z(n4096) );
  XOR U4236 ( .A(n4097), .B(n4096), .Z(n1489) );
  XNOR U4237 ( .A(n1488), .B(n1489), .Z(n1490) );
  XNOR U4238 ( .A(n1491), .B(n1490), .Z(n1353) );
  XNOR U4239 ( .A(x[1250]), .B(y[1250]), .Z(n1533) );
  XNOR U4240 ( .A(x[1246]), .B(y[1246]), .Z(n1530) );
  XNOR U4241 ( .A(x[1248]), .B(y[1248]), .Z(n1531) );
  XOR U4242 ( .A(n1530), .B(n1531), .Z(n1532) );
  XOR U4243 ( .A(n1533), .B(n1532), .Z(n1867) );
  XNOR U4244 ( .A(x[1256]), .B(y[1256]), .Z(n1527) );
  XNOR U4245 ( .A(x[1252]), .B(y[1252]), .Z(n1524) );
  XNOR U4246 ( .A(x[1254]), .B(y[1254]), .Z(n1525) );
  XOR U4247 ( .A(n1524), .B(n1525), .Z(n1526) );
  XNOR U4248 ( .A(n1527), .B(n1526), .Z(n1864) );
  XNOR U4249 ( .A(x[390]), .B(y[390]), .Z(n3668) );
  XNOR U4250 ( .A(x[382]), .B(y[382]), .Z(n3665) );
  XNOR U4251 ( .A(x[388]), .B(y[388]), .Z(n3666) );
  XOR U4252 ( .A(n3665), .B(n3666), .Z(n3667) );
  XNOR U4253 ( .A(n3668), .B(n3667), .Z(n1865) );
  XNOR U4254 ( .A(n1867), .B(n1866), .Z(n4242) );
  XNOR U4255 ( .A(x[1034]), .B(y[1034]), .Z(n3167) );
  XNOR U4256 ( .A(x[1030]), .B(y[1030]), .Z(n3164) );
  XNOR U4257 ( .A(x[1032]), .B(y[1032]), .Z(n3165) );
  XOR U4258 ( .A(n3164), .B(n3165), .Z(n3166) );
  XOR U4259 ( .A(n3167), .B(n3166), .Z(n4026) );
  XNOR U4260 ( .A(x[1046]), .B(y[1046]), .Z(n3161) );
  XNOR U4261 ( .A(x[1042]), .B(y[1042]), .Z(n3158) );
  XNOR U4262 ( .A(x[1044]), .B(y[1044]), .Z(n3159) );
  XOR U4263 ( .A(n3158), .B(n3159), .Z(n3160) );
  XNOR U4264 ( .A(n3161), .B(n3160), .Z(n4024) );
  XNOR U4265 ( .A(x[1040]), .B(y[1040]), .Z(n3155) );
  XNOR U4266 ( .A(x[1036]), .B(y[1036]), .Z(n3152) );
  XNOR U4267 ( .A(x[1038]), .B(y[1038]), .Z(n3153) );
  XOR U4268 ( .A(n3152), .B(n3153), .Z(n3154) );
  XNOR U4269 ( .A(n3155), .B(n3154), .Z(n4025) );
  XOR U4270 ( .A(n4026), .B(n4027), .Z(n4243) );
  XOR U4271 ( .A(n4242), .B(n4243), .Z(n4244) );
  XNOR U4272 ( .A(x[1016]), .B(y[1016]), .Z(n3045) );
  XNOR U4273 ( .A(x[1012]), .B(y[1012]), .Z(n3042) );
  XNOR U4274 ( .A(x[1014]), .B(y[1014]), .Z(n3043) );
  XOR U4275 ( .A(n3042), .B(n3043), .Z(n3044) );
  XOR U4276 ( .A(n3045), .B(n3044), .Z(n4069) );
  XNOR U4277 ( .A(x[1022]), .B(y[1022]), .Z(n3039) );
  XNOR U4278 ( .A(x[1018]), .B(y[1018]), .Z(n3036) );
  XNOR U4279 ( .A(x[1020]), .B(y[1020]), .Z(n3037) );
  XOR U4280 ( .A(n3036), .B(n3037), .Z(n3038) );
  XOR U4281 ( .A(n3039), .B(n3038), .Z(n4066) );
  XNOR U4282 ( .A(x[1028]), .B(y[1028]), .Z(n3051) );
  XNOR U4283 ( .A(x[1024]), .B(y[1024]), .Z(n3048) );
  XNOR U4284 ( .A(x[1026]), .B(y[1026]), .Z(n3049) );
  XOR U4285 ( .A(n3048), .B(n3049), .Z(n3050) );
  XNOR U4286 ( .A(n3051), .B(n3050), .Z(n4067) );
  XNOR U4287 ( .A(n4066), .B(n4067), .Z(n4068) );
  XNOR U4288 ( .A(n4069), .B(n4068), .Z(n4245) );
  XOR U4289 ( .A(n4244), .B(n4245), .Z(n2597) );
  XNOR U4290 ( .A(x[1220]), .B(y[1220]), .Z(n1467) );
  XNOR U4291 ( .A(x[1216]), .B(y[1216]), .Z(n1464) );
  XNOR U4292 ( .A(x[1218]), .B(y[1218]), .Z(n1465) );
  XOR U4293 ( .A(n1464), .B(n1465), .Z(n1466) );
  XOR U4294 ( .A(n1467), .B(n1466), .Z(n4449) );
  XNOR U4295 ( .A(x[1232]), .B(y[1232]), .Z(n1461) );
  XNOR U4296 ( .A(x[1228]), .B(y[1228]), .Z(n1458) );
  XNOR U4297 ( .A(x[1230]), .B(y[1230]), .Z(n1459) );
  XOR U4298 ( .A(n1458), .B(n1459), .Z(n1460) );
  XNOR U4299 ( .A(n1461), .B(n1460), .Z(n4446) );
  XNOR U4300 ( .A(x[1226]), .B(y[1226]), .Z(n1455) );
  XNOR U4301 ( .A(x[1222]), .B(y[1222]), .Z(n1452) );
  XNOR U4302 ( .A(x[1224]), .B(y[1224]), .Z(n1453) );
  XOR U4303 ( .A(n1452), .B(n1453), .Z(n1454) );
  XNOR U4304 ( .A(n1455), .B(n1454), .Z(n4447) );
  XNOR U4305 ( .A(n4449), .B(n4448), .Z(n4209) );
  XNOR U4306 ( .A(x[1052]), .B(y[1052]), .Z(n2997) );
  XNOR U4307 ( .A(x[1048]), .B(y[1048]), .Z(n2994) );
  XNOR U4308 ( .A(x[1050]), .B(y[1050]), .Z(n2995) );
  XOR U4309 ( .A(n2994), .B(n2995), .Z(n2996) );
  XOR U4310 ( .A(n2997), .B(n2996), .Z(n4039) );
  XNOR U4311 ( .A(x[1058]), .B(y[1058]), .Z(n2991) );
  XNOR U4312 ( .A(x[1054]), .B(y[1054]), .Z(n2988) );
  XNOR U4313 ( .A(x[1056]), .B(y[1056]), .Z(n2989) );
  XOR U4314 ( .A(n2988), .B(n2989), .Z(n2990) );
  XNOR U4315 ( .A(n2991), .B(n2990), .Z(n4036) );
  XNOR U4316 ( .A(x[138]), .B(y[138]), .Z(n3712) );
  XNOR U4317 ( .A(x[132]), .B(y[132]), .Z(n3709) );
  XNOR U4318 ( .A(x[134]), .B(y[134]), .Z(n3710) );
  XOR U4319 ( .A(n3709), .B(n3710), .Z(n3711) );
  XNOR U4320 ( .A(n3712), .B(n3711), .Z(n4037) );
  XNOR U4321 ( .A(n4039), .B(n4038), .Z(n4206) );
  XNOR U4322 ( .A(x[1238]), .B(y[1238]), .Z(n1431) );
  XNOR U4323 ( .A(x[1234]), .B(y[1234]), .Z(n1428) );
  XNOR U4324 ( .A(x[1236]), .B(y[1236]), .Z(n1429) );
  XOR U4325 ( .A(n1428), .B(n1429), .Z(n1430) );
  XOR U4326 ( .A(n1431), .B(n1430), .Z(n4910) );
  XNOR U4327 ( .A(x[362]), .B(y[362]), .Z(n3628) );
  XNOR U4328 ( .A(x[354]), .B(y[354]), .Z(n3625) );
  XNOR U4329 ( .A(x[750]), .B(y[750]), .Z(n3626) );
  XOR U4330 ( .A(n3625), .B(n3626), .Z(n3627) );
  XNOR U4331 ( .A(n3628), .B(n3627), .Z(n4908) );
  XNOR U4332 ( .A(x[1244]), .B(y[1244]), .Z(n1425) );
  XNOR U4333 ( .A(x[1240]), .B(y[1240]), .Z(n1422) );
  XNOR U4334 ( .A(x[1242]), .B(y[1242]), .Z(n1423) );
  XOR U4335 ( .A(n1422), .B(n1423), .Z(n1424) );
  XNOR U4336 ( .A(n1425), .B(n1424), .Z(n4909) );
  XOR U4337 ( .A(n4910), .B(n4911), .Z(n4207) );
  XOR U4338 ( .A(n4206), .B(n4207), .Z(n4208) );
  XOR U4339 ( .A(n4209), .B(n4208), .Z(n2594) );
  XNOR U4340 ( .A(x[1156]), .B(y[1156]), .Z(n3306) );
  XNOR U4341 ( .A(x[1148]), .B(y[1148]), .Z(n3303) );
  XNOR U4342 ( .A(x[1152]), .B(y[1152]), .Z(n3304) );
  XOR U4343 ( .A(n3303), .B(n3304), .Z(n3305) );
  XOR U4344 ( .A(n3306), .B(n3305), .Z(n1255) );
  XNOR U4345 ( .A(x[1168]), .B(y[1168]), .Z(n3300) );
  XNOR U4346 ( .A(x[1160]), .B(y[1160]), .Z(n3297) );
  XNOR U4347 ( .A(x[1164]), .B(y[1164]), .Z(n3298) );
  XOR U4348 ( .A(n3297), .B(n3298), .Z(n3299) );
  XNOR U4349 ( .A(n3300), .B(n3299), .Z(n1252) );
  XNOR U4350 ( .A(x[250]), .B(y[250]), .Z(n2457) );
  XNOR U4351 ( .A(x[244]), .B(y[244]), .Z(n2454) );
  XNOR U4352 ( .A(x[710]), .B(y[710]), .Z(n2455) );
  XOR U4353 ( .A(n2454), .B(n2455), .Z(n2456) );
  XNOR U4354 ( .A(n2457), .B(n2456), .Z(n1253) );
  XNOR U4355 ( .A(n1255), .B(n1254), .Z(n4200) );
  XNOR U4356 ( .A(x[1064]), .B(y[1064]), .Z(n3119) );
  XNOR U4357 ( .A(x[1060]), .B(y[1060]), .Z(n3116) );
  XNOR U4358 ( .A(x[1062]), .B(y[1062]), .Z(n3117) );
  XOR U4359 ( .A(n3116), .B(n3117), .Z(n3118) );
  XOR U4360 ( .A(n3119), .B(n3118), .Z(n1404) );
  XNOR U4361 ( .A(x[1072]), .B(y[1072]), .Z(n3113) );
  XNOR U4362 ( .A(x[1066]), .B(y[1066]), .Z(n3110) );
  XNOR U4363 ( .A(x[1068]), .B(y[1068]), .Z(n3111) );
  XOR U4364 ( .A(n3110), .B(n3111), .Z(n3112) );
  XNOR U4365 ( .A(n3113), .B(n3112), .Z(n1402) );
  XNOR U4366 ( .A(x[162]), .B(y[162]), .Z(n2295) );
  XNOR U4367 ( .A(x[158]), .B(y[158]), .Z(n2292) );
  XNOR U4368 ( .A(x[678]), .B(y[678]), .Z(n2293) );
  XOR U4369 ( .A(n2292), .B(n2293), .Z(n2294) );
  XNOR U4370 ( .A(n2295), .B(n2294), .Z(n1403) );
  XOR U4371 ( .A(n1404), .B(n1405), .Z(n4201) );
  XOR U4372 ( .A(n4200), .B(n4201), .Z(n4202) );
  XNOR U4373 ( .A(x[1202]), .B(y[1202]), .Z(n3185) );
  XNOR U4374 ( .A(x[1196]), .B(y[1196]), .Z(n3182) );
  XNOR U4375 ( .A(x[1200]), .B(y[1200]), .Z(n3183) );
  XOR U4376 ( .A(n3182), .B(n3183), .Z(n3184) );
  XOR U4377 ( .A(n3185), .B(n3184), .Z(n4397) );
  XNOR U4378 ( .A(x[1208]), .B(y[1208]), .Z(n3179) );
  XNOR U4379 ( .A(x[1204]), .B(y[1204]), .Z(n3176) );
  XNOR U4380 ( .A(x[1206]), .B(y[1206]), .Z(n3177) );
  XOR U4381 ( .A(n3176), .B(n3177), .Z(n3178) );
  XNOR U4382 ( .A(n3179), .B(n3178), .Z(n4394) );
  XNOR U4383 ( .A(x[1214]), .B(y[1214]), .Z(n3191) );
  XNOR U4384 ( .A(x[1210]), .B(y[1210]), .Z(n3188) );
  XNOR U4385 ( .A(x[1212]), .B(y[1212]), .Z(n3189) );
  XOR U4386 ( .A(n3188), .B(n3189), .Z(n3190) );
  XNOR U4387 ( .A(n3191), .B(n3190), .Z(n4395) );
  XNOR U4388 ( .A(n4397), .B(n4396), .Z(n4203) );
  XNOR U4389 ( .A(n4202), .B(n4203), .Z(n2595) );
  XNOR U4390 ( .A(n2594), .B(n2595), .Z(n2596) );
  XNOR U4391 ( .A(n2597), .B(n2596), .Z(n1351) );
  XNOR U4392 ( .A(x[894]), .B(y[894]), .Z(n897) );
  XNOR U4393 ( .A(x[892]), .B(y[892]), .Z(n895) );
  XOR U4394 ( .A(x[1178]), .B(y[1178]), .Z(n894) );
  XNOR U4395 ( .A(n895), .B(n894), .Z(n896) );
  XOR U4396 ( .A(n897), .B(n896), .Z(n3173) );
  XNOR U4397 ( .A(x[898]), .B(y[898]), .Z(n893) );
  XNOR U4398 ( .A(x[896]), .B(y[896]), .Z(n891) );
  XOR U4399 ( .A(x[1412]), .B(y[1412]), .Z(n890) );
  XNOR U4400 ( .A(n891), .B(n890), .Z(n892) );
  XOR U4401 ( .A(n893), .B(n892), .Z(n3170) );
  XNOR U4402 ( .A(x[115]), .B(y[115]), .Z(n3893) );
  XNOR U4403 ( .A(x[119]), .B(y[119]), .Z(n3891) );
  XOR U4404 ( .A(x[516]), .B(y[516]), .Z(n3890) );
  XNOR U4405 ( .A(n3891), .B(n3890), .Z(n3892) );
  XNOR U4406 ( .A(n3893), .B(n3892), .Z(n3171) );
  XNOR U4407 ( .A(n3170), .B(n3171), .Z(n3172) );
  XNOR U4408 ( .A(n3173), .B(n3172), .Z(n4143) );
  XNOR U4409 ( .A(x[1370]), .B(y[1370]), .Z(n1211) );
  XNOR U4410 ( .A(x[1292]), .B(y[1292]), .Z(n1209) );
  XOR U4411 ( .A(x[1372]), .B(y[1372]), .Z(n1208) );
  XNOR U4412 ( .A(n1209), .B(n1208), .Z(n1210) );
  XOR U4413 ( .A(n1211), .B(n1210), .Z(n1595) );
  XNOR U4414 ( .A(x[1280]), .B(y[1280]), .Z(n1207) );
  XNOR U4415 ( .A(x[1278]), .B(y[1278]), .Z(n1205) );
  XOR U4416 ( .A(x[1290]), .B(y[1290]), .Z(n1204) );
  XNOR U4417 ( .A(n1205), .B(n1204), .Z(n1206) );
  XOR U4418 ( .A(n1207), .B(n1206), .Z(n1592) );
  XNOR U4419 ( .A(x[1276]), .B(y[1276]), .Z(n1203) );
  XNOR U4420 ( .A(x[1288]), .B(y[1288]), .Z(n1201) );
  XOR U4421 ( .A(x[1368]), .B(y[1368]), .Z(n1200) );
  XNOR U4422 ( .A(n1201), .B(n1200), .Z(n1202) );
  XNOR U4423 ( .A(n1203), .B(n1202), .Z(n1593) );
  XNOR U4424 ( .A(n1592), .B(n1593), .Z(n1594) );
  XOR U4425 ( .A(n1595), .B(n1594), .Z(n4142) );
  XNOR U4426 ( .A(n4143), .B(n4142), .Z(n4144) );
  XNOR U4427 ( .A(x[902]), .B(y[902]), .Z(n921) );
  XNOR U4428 ( .A(x[900]), .B(y[900]), .Z(n919) );
  XOR U4429 ( .A(x[1182]), .B(y[1182]), .Z(n918) );
  XNOR U4430 ( .A(n919), .B(n918), .Z(n920) );
  XOR U4431 ( .A(n921), .B(n920), .Z(n3638) );
  XNOR U4432 ( .A(x[906]), .B(y[906]), .Z(n917) );
  XNOR U4433 ( .A(x[904]), .B(y[904]), .Z(n915) );
  XOR U4434 ( .A(x[1410]), .B(y[1410]), .Z(n914) );
  XNOR U4435 ( .A(n915), .B(n914), .Z(n916) );
  XOR U4436 ( .A(n917), .B(n916), .Z(n3635) );
  XNOR U4437 ( .A(x[99]), .B(y[99]), .Z(n3889) );
  XNOR U4438 ( .A(x[103]), .B(y[103]), .Z(n3887) );
  XOR U4439 ( .A(x[105]), .B(y[105]), .Z(n3886) );
  XNOR U4440 ( .A(n3887), .B(n3886), .Z(n3888) );
  XNOR U4441 ( .A(n3889), .B(n3888), .Z(n3636) );
  XNOR U4442 ( .A(n3635), .B(n3636), .Z(n3637) );
  XOR U4443 ( .A(n3638), .B(n3637), .Z(n4145) );
  XOR U4444 ( .A(n4144), .B(n4145), .Z(n4478) );
  XNOR U4445 ( .A(x[1378]), .B(y[1378]), .Z(n4561) );
  XNOR U4446 ( .A(x[1308]), .B(y[1308]), .Z(n4559) );
  XOR U4447 ( .A(x[1380]), .B(y[1380]), .Z(n4558) );
  XNOR U4448 ( .A(n4559), .B(n4558), .Z(n4560) );
  XOR U4449 ( .A(n4561), .B(n4560), .Z(n1013) );
  XNOR U4450 ( .A(x[1374]), .B(y[1374]), .Z(n4557) );
  XNOR U4451 ( .A(x[1296]), .B(y[1296]), .Z(n4555) );
  XOR U4452 ( .A(x[1376]), .B(y[1376]), .Z(n4554) );
  XNOR U4453 ( .A(n4555), .B(n4554), .Z(n4556) );
  XNOR U4454 ( .A(n4557), .B(n4556), .Z(n1010) );
  XNOR U4455 ( .A(x[474]), .B(y[474]), .Z(n4129) );
  XNOR U4456 ( .A(x[470]), .B(y[470]), .Z(n4127) );
  XOR U4457 ( .A(x[800]), .B(y[800]), .Z(n4126) );
  XNOR U4458 ( .A(n4127), .B(n4126), .Z(n4128) );
  XNOR U4459 ( .A(n4129), .B(n4128), .Z(n1011) );
  XNOR U4460 ( .A(n1013), .B(n1012), .Z(n4054) );
  XNOR U4461 ( .A(x[910]), .B(y[910]), .Z(n909) );
  XNOR U4462 ( .A(x[908]), .B(y[908]), .Z(n907) );
  XOR U4463 ( .A(x[1186]), .B(y[1186]), .Z(n906) );
  XNOR U4464 ( .A(n907), .B(n906), .Z(n908) );
  XOR U4465 ( .A(n909), .B(n908), .Z(n3679) );
  XNOR U4466 ( .A(x[914]), .B(y[914]), .Z(n901) );
  XNOR U4467 ( .A(x[912]), .B(y[912]), .Z(n899) );
  XOR U4468 ( .A(x[1408]), .B(y[1408]), .Z(n898) );
  XNOR U4469 ( .A(n899), .B(n898), .Z(n900) );
  XNOR U4470 ( .A(n901), .B(n900), .Z(n3677) );
  XNOR U4471 ( .A(x[918]), .B(y[918]), .Z(n905) );
  XNOR U4472 ( .A(x[916]), .B(y[916]), .Z(n903) );
  XOR U4473 ( .A(x[1190]), .B(y[1190]), .Z(n902) );
  XNOR U4474 ( .A(n903), .B(n902), .Z(n904) );
  XNOR U4475 ( .A(n905), .B(n904), .Z(n3678) );
  XOR U4476 ( .A(n3679), .B(n3680), .Z(n4055) );
  XOR U4477 ( .A(n4054), .B(n4055), .Z(n4056) );
  XNOR U4478 ( .A(x[922]), .B(y[922]), .Z(n1115) );
  XNOR U4479 ( .A(x[920]), .B(y[920]), .Z(n1113) );
  XOR U4480 ( .A(x[1406]), .B(y[1406]), .Z(n1112) );
  XNOR U4481 ( .A(n1113), .B(n1112), .Z(n1114) );
  XOR U4482 ( .A(n1115), .B(n1114), .Z(n2198) );
  XNOR U4483 ( .A(x[930]), .B(y[930]), .Z(n1111) );
  XNOR U4484 ( .A(x[928]), .B(y[928]), .Z(n1109) );
  XOR U4485 ( .A(x[1404]), .B(y[1404]), .Z(n1108) );
  XNOR U4486 ( .A(n1109), .B(n1108), .Z(n1110) );
  XNOR U4487 ( .A(n1111), .B(n1110), .Z(n2196) );
  XNOR U4488 ( .A(x[926]), .B(y[926]), .Z(n1107) );
  XNOR U4489 ( .A(x[924]), .B(y[924]), .Z(n1105) );
  XOR U4490 ( .A(x[1194]), .B(y[1194]), .Z(n1104) );
  XNOR U4491 ( .A(n1105), .B(n1104), .Z(n1106) );
  XNOR U4492 ( .A(n1107), .B(n1106), .Z(n2197) );
  XOR U4493 ( .A(n2198), .B(n2199), .Z(n4057) );
  XNOR U4494 ( .A(n4056), .B(n4057), .Z(n4476) );
  XNOR U4495 ( .A(x[944]), .B(y[944]), .Z(n3103) );
  XNOR U4496 ( .A(x[940]), .B(y[940]), .Z(n3100) );
  XNOR U4497 ( .A(x[942]), .B(y[942]), .Z(n3101) );
  XOR U4498 ( .A(n3100), .B(n3101), .Z(n3102) );
  XOR U4499 ( .A(n3103), .B(n3102), .Z(n4139) );
  XNOR U4500 ( .A(x[950]), .B(y[950]), .Z(n3097) );
  XNOR U4501 ( .A(x[946]), .B(y[946]), .Z(n3094) );
  XNOR U4502 ( .A(x[948]), .B(y[948]), .Z(n3095) );
  XOR U4503 ( .A(n3094), .B(n3095), .Z(n3096) );
  XNOR U4504 ( .A(n3097), .B(n3096), .Z(n4136) );
  XNOR U4505 ( .A(x[27]), .B(y[27]), .Z(n3845) );
  XNOR U4506 ( .A(x[31]), .B(y[31]), .Z(n3843) );
  XOR U4507 ( .A(x[33]), .B(y[33]), .Z(n3842) );
  XNOR U4508 ( .A(n3843), .B(n3842), .Z(n3844) );
  XNOR U4509 ( .A(n3845), .B(n3844), .Z(n4137) );
  XNOR U4510 ( .A(n4139), .B(n4138), .Z(n4060) );
  XNOR U4511 ( .A(x[1384]), .B(y[1384]), .Z(n4765) );
  XNOR U4512 ( .A(x[1310]), .B(y[1310]), .Z(n4762) );
  XNOR U4513 ( .A(x[1386]), .B(y[1386]), .Z(n4763) );
  XOR U4514 ( .A(n4762), .B(n4763), .Z(n4764) );
  XOR U4515 ( .A(n4765), .B(n4764), .Z(n2590) );
  XNOR U4516 ( .A(x[458]), .B(y[458]), .Z(n4133) );
  XNOR U4517 ( .A(x[452]), .B(y[452]), .Z(n4130) );
  XNOR U4518 ( .A(x[456]), .B(y[456]), .Z(n4131) );
  XOR U4519 ( .A(n4130), .B(n4131), .Z(n4132) );
  XNOR U4520 ( .A(n4133), .B(n4132), .Z(n2588) );
  XNOR U4521 ( .A(x[1274]), .B(y[1274]), .Z(n4759) );
  XNOR U4522 ( .A(x[1300]), .B(y[1300]), .Z(n4756) );
  XNOR U4523 ( .A(x[1382]), .B(y[1382]), .Z(n4757) );
  XOR U4524 ( .A(n4756), .B(n4757), .Z(n4758) );
  XNOR U4525 ( .A(n4759), .B(n4758), .Z(n2589) );
  XOR U4526 ( .A(n2590), .B(n2591), .Z(n4061) );
  XOR U4527 ( .A(n4060), .B(n4061), .Z(n4062) );
  XNOR U4528 ( .A(x[934]), .B(y[934]), .Z(n3069) );
  XNOR U4529 ( .A(x[932]), .B(y[932]), .Z(n3066) );
  XNOR U4530 ( .A(x[1198]), .B(y[1198]), .Z(n3067) );
  XOR U4531 ( .A(n3066), .B(n3067), .Z(n3068) );
  XOR U4532 ( .A(n3069), .B(n3068), .Z(n2150) );
  XNOR U4533 ( .A(x[938]), .B(y[938]), .Z(n3063) );
  XNOR U4534 ( .A(x[936]), .B(y[936]), .Z(n3060) );
  XNOR U4535 ( .A(x[1402]), .B(y[1402]), .Z(n3061) );
  XOR U4536 ( .A(n3060), .B(n3061), .Z(n3062) );
  XNOR U4537 ( .A(n3063), .B(n3062), .Z(n2148) );
  XNOR U4538 ( .A(x[45]), .B(y[45]), .Z(n3871) );
  XNOR U4539 ( .A(x[49]), .B(y[49]), .Z(n3869) );
  XOR U4540 ( .A(x[568]), .B(y[568]), .Z(n3868) );
  XNOR U4541 ( .A(n3869), .B(n3868), .Z(n3870) );
  XNOR U4542 ( .A(n3871), .B(n3870), .Z(n2149) );
  XOR U4543 ( .A(n2150), .B(n2151), .Z(n4063) );
  XNOR U4544 ( .A(n4062), .B(n4063), .Z(n4477) );
  XOR U4545 ( .A(n4476), .B(n4477), .Z(n4479) );
  XOR U4546 ( .A(n4478), .B(n4479), .Z(n1350) );
  XOR U4547 ( .A(n1351), .B(n1350), .Z(n1352) );
  XOR U4548 ( .A(n1353), .B(n1352), .Z(n809) );
  XOR U4549 ( .A(n808), .B(n809), .Z(n810) );
  XOR U4550 ( .A(n811), .B(n810), .Z(n802) );
  XNOR U4551 ( .A(x[807]), .B(y[807]), .Z(n2477) );
  XNOR U4552 ( .A(x[184]), .B(y[184]), .Z(n2475) );
  XOR U4553 ( .A(x[809]), .B(y[809]), .Z(n2474) );
  XNOR U4554 ( .A(n2475), .B(n2474), .Z(n2476) );
  XOR U4555 ( .A(n2477), .B(n2476), .Z(n3720) );
  XNOR U4556 ( .A(x[803]), .B(y[803]), .Z(n2375) );
  XNOR U4557 ( .A(x[500]), .B(y[500]), .Z(n2372) );
  XNOR U4558 ( .A(x[805]), .B(y[805]), .Z(n2373) );
  XOR U4559 ( .A(n2372), .B(n2373), .Z(n2374) );
  XNOR U4560 ( .A(n2375), .B(n2374), .Z(n3719) );
  XOR U4561 ( .A(n3720), .B(n3719), .Z(n3722) );
  XNOR U4562 ( .A(x[815]), .B(y[815]), .Z(n4649) );
  XNOR U4563 ( .A(x[817]), .B(y[817]), .Z(n4647) );
  XOR U4564 ( .A(x[1504]), .B(y[1504]), .Z(n4646) );
  XNOR U4565 ( .A(n4647), .B(n4646), .Z(n4648) );
  XNOR U4566 ( .A(n4649), .B(n4648), .Z(n3721) );
  XNOR U4567 ( .A(x[839]), .B(y[839]), .Z(n2133) );
  XNOR U4568 ( .A(x[156]), .B(y[156]), .Z(n2130) );
  XNOR U4569 ( .A(x[841]), .B(y[841]), .Z(n2131) );
  XOR U4570 ( .A(n2130), .B(n2131), .Z(n2132) );
  XOR U4571 ( .A(n2133), .B(n2132), .Z(n4701) );
  XNOR U4572 ( .A(x[831]), .B(y[831]), .Z(n4109) );
  XNOR U4573 ( .A(x[164]), .B(y[164]), .Z(n4107) );
  XOR U4574 ( .A(x[833]), .B(y[833]), .Z(n4106) );
  XNOR U4575 ( .A(n4107), .B(n4106), .Z(n4108) );
  XOR U4576 ( .A(n4109), .B(n4108), .Z(n4698) );
  XNOR U4577 ( .A(x[823]), .B(y[823]), .Z(n4235) );
  XNOR U4578 ( .A(x[825]), .B(y[825]), .Z(n4233) );
  XOR U4579 ( .A(x[1506]), .B(y[1506]), .Z(n4232) );
  XNOR U4580 ( .A(n4233), .B(n4232), .Z(n4234) );
  XNOR U4581 ( .A(n4235), .B(n4234), .Z(n4699) );
  XNOR U4582 ( .A(n4698), .B(n4699), .Z(n4700) );
  XNOR U4583 ( .A(n4701), .B(n4700), .Z(n2869) );
  XOR U4584 ( .A(n2868), .B(n2869), .Z(n2870) );
  XNOR U4585 ( .A(x[799]), .B(y[799]), .Z(n2431) );
  XNOR U4586 ( .A(x[192]), .B(y[192]), .Z(n2428) );
  XNOR U4587 ( .A(x[801]), .B(y[801]), .Z(n2429) );
  XOR U4588 ( .A(n2428), .B(n2429), .Z(n2430) );
  XOR U4589 ( .A(n2431), .B(n2430), .Z(n2847) );
  XNOR U4590 ( .A(x[791]), .B(y[791]), .Z(n2333) );
  XNOR U4591 ( .A(x[793]), .B(y[793]), .Z(n2330) );
  XNOR U4592 ( .A(x[1502]), .B(y[1502]), .Z(n2331) );
  XOR U4593 ( .A(n2330), .B(n2331), .Z(n2332) );
  XOR U4594 ( .A(n2333), .B(n2332), .Z(n2844) );
  XNOR U4595 ( .A(x[795]), .B(y[795]), .Z(n4497) );
  XNOR U4596 ( .A(x[506]), .B(y[506]), .Z(n4494) );
  XNOR U4597 ( .A(x[797]), .B(y[797]), .Z(n4495) );
  XOR U4598 ( .A(n4494), .B(n4495), .Z(n4496) );
  XNOR U4599 ( .A(n4497), .B(n4496), .Z(n2845) );
  XNOR U4600 ( .A(n2844), .B(n2845), .Z(n2846) );
  XNOR U4601 ( .A(n2847), .B(n2846), .Z(n2871) );
  XOR U4602 ( .A(n2870), .B(n2871), .Z(n985) );
  XNOR U4603 ( .A(x[773]), .B(y[773]), .Z(n3221) );
  XNOR U4604 ( .A(x[212]), .B(y[212]), .Z(n3218) );
  XNOR U4605 ( .A(x[775]), .B(y[775]), .Z(n3219) );
  XOR U4606 ( .A(n3218), .B(n3219), .Z(n3220) );
  XOR U4607 ( .A(n3221), .B(n3220), .Z(n3861) );
  XNOR U4608 ( .A(x[765]), .B(y[765]), .Z(n3085) );
  XNOR U4609 ( .A(x[218]), .B(y[218]), .Z(n3082) );
  XNOR U4610 ( .A(x[767]), .B(y[767]), .Z(n3083) );
  XOR U4611 ( .A(n3082), .B(n3083), .Z(n3084) );
  XOR U4612 ( .A(n3085), .B(n3084), .Z(n3858) );
  XNOR U4613 ( .A(x[769]), .B(y[769]), .Z(n3079) );
  XNOR U4614 ( .A(x[520]), .B(y[520]), .Z(n3076) );
  XNOR U4615 ( .A(x[771]), .B(y[771]), .Z(n3077) );
  XOR U4616 ( .A(n3076), .B(n3077), .Z(n3078) );
  XNOR U4617 ( .A(n3079), .B(n3078), .Z(n3859) );
  XNOR U4618 ( .A(n3858), .B(n3859), .Z(n3860) );
  XNOR U4619 ( .A(n3861), .B(n3860), .Z(n1334) );
  XNOR U4620 ( .A(x[785]), .B(y[785]), .Z(n3029) );
  XNOR U4621 ( .A(x[198]), .B(y[198]), .Z(n3027) );
  XOR U4622 ( .A(x[787]), .B(y[787]), .Z(n3026) );
  XNOR U4623 ( .A(n3027), .B(n3026), .Z(n3028) );
  XOR U4624 ( .A(n3029), .B(n3028), .Z(n3909) );
  XNOR U4625 ( .A(x[777]), .B(y[777]), .Z(n3131) );
  XNOR U4626 ( .A(x[208]), .B(y[208]), .Z(n3129) );
  XNOR U4627 ( .A(x[779]), .B(y[779]), .Z(n3128) );
  XNOR U4628 ( .A(n3129), .B(n3128), .Z(n3130) );
  XNOR U4629 ( .A(n3131), .B(n3130), .Z(n3906) );
  XNOR U4630 ( .A(x[781]), .B(y[781]), .Z(n3025) );
  XNOR U4631 ( .A(x[783]), .B(y[783]), .Z(n3023) );
  XOR U4632 ( .A(x[1500]), .B(y[1500]), .Z(n3022) );
  XNOR U4633 ( .A(n3023), .B(n3022), .Z(n3024) );
  XNOR U4634 ( .A(n3025), .B(n3024), .Z(n3907) );
  XNOR U4635 ( .A(n3906), .B(n3907), .Z(n3908) );
  XNOR U4636 ( .A(n3909), .B(n3908), .Z(n1335) );
  XOR U4637 ( .A(n1334), .B(n1335), .Z(n1336) );
  XNOR U4638 ( .A(x[761]), .B(y[761]), .Z(n3137) );
  XNOR U4639 ( .A(x[526]), .B(y[526]), .Z(n3135) );
  XNOR U4640 ( .A(x[763]), .B(y[763]), .Z(n3134) );
  XNOR U4641 ( .A(n3135), .B(n3134), .Z(n3136) );
  XNOR U4642 ( .A(n3137), .B(n3136), .Z(n1933) );
  XNOR U4643 ( .A(x[753]), .B(y[753]), .Z(n2277) );
  XNOR U4644 ( .A(x[228]), .B(y[228]), .Z(n2275) );
  XOR U4645 ( .A(x[755]), .B(y[755]), .Z(n2274) );
  XNOR U4646 ( .A(n2275), .B(n2274), .Z(n2276) );
  XOR U4647 ( .A(n2277), .B(n2276), .Z(n1930) );
  XNOR U4648 ( .A(x[757]), .B(y[757]), .Z(n3999) );
  XNOR U4649 ( .A(x[759]), .B(y[759]), .Z(n3996) );
  XNOR U4650 ( .A(x[1498]), .B(y[1498]), .Z(n3997) );
  XOR U4651 ( .A(n3996), .B(n3997), .Z(n3998) );
  XNOR U4652 ( .A(n3999), .B(n3998), .Z(n1931) );
  XNOR U4653 ( .A(n1930), .B(n1931), .Z(n1932) );
  XOR U4654 ( .A(n1933), .B(n1932), .Z(n1337) );
  XNOR U4655 ( .A(n1336), .B(n1337), .Z(n982) );
  XNOR U4656 ( .A(x[737]), .B(y[737]), .Z(n933) );
  XNOR U4657 ( .A(x[540]), .B(y[540]), .Z(n931) );
  XOR U4658 ( .A(x[739]), .B(y[739]), .Z(n930) );
  XNOR U4659 ( .A(n931), .B(n930), .Z(n932) );
  XOR U4660 ( .A(n933), .B(n932), .Z(n3744) );
  XNOR U4661 ( .A(x[729]), .B(y[729]), .Z(n3312) );
  XNOR U4662 ( .A(x[546]), .B(y[546]), .Z(n3310) );
  XOR U4663 ( .A(x[731]), .B(y[731]), .Z(n3309) );
  XNOR U4664 ( .A(n3310), .B(n3309), .Z(n3311) );
  XOR U4665 ( .A(n3312), .B(n3311), .Z(n3741) );
  XNOR U4666 ( .A(x[733]), .B(y[733]), .Z(n3255) );
  XNOR U4667 ( .A(x[248]), .B(y[248]), .Z(n3253) );
  XOR U4668 ( .A(x[735]), .B(y[735]), .Z(n3252) );
  XNOR U4669 ( .A(n3253), .B(n3252), .Z(n3254) );
  XNOR U4670 ( .A(n3255), .B(n3254), .Z(n3742) );
  XNOR U4671 ( .A(n3741), .B(n3742), .Z(n3743) );
  XNOR U4672 ( .A(n3744), .B(n3743), .Z(n1329) );
  XNOR U4673 ( .A(x[749]), .B(y[749]), .Z(n1617) );
  XNOR U4674 ( .A(x[751]), .B(y[751]), .Z(n1614) );
  XNOR U4675 ( .A(x[1496]), .B(y[1496]), .Z(n1615) );
  XOR U4676 ( .A(n1614), .B(n1615), .Z(n1616) );
  XOR U4677 ( .A(n1617), .B(n1616), .Z(n1955) );
  XNOR U4678 ( .A(x[745]), .B(y[745]), .Z(n3756) );
  XNOR U4679 ( .A(x[234]), .B(y[234]), .Z(n3754) );
  XOR U4680 ( .A(x[747]), .B(y[747]), .Z(n3753) );
  XNOR U4681 ( .A(n3754), .B(n3753), .Z(n3755) );
  XOR U4682 ( .A(n3756), .B(n3755), .Z(n1952) );
  XNOR U4683 ( .A(x[741]), .B(y[741]), .Z(n1149) );
  XNOR U4684 ( .A(x[238]), .B(y[238]), .Z(n1146) );
  XNOR U4685 ( .A(x[743]), .B(y[743]), .Z(n1147) );
  XOR U4686 ( .A(n1146), .B(n1147), .Z(n1148) );
  XNOR U4687 ( .A(n1149), .B(n1148), .Z(n1953) );
  XNOR U4688 ( .A(n1952), .B(n1953), .Z(n1954) );
  XOR U4689 ( .A(n1955), .B(n1954), .Z(n1328) );
  XOR U4690 ( .A(n1329), .B(n1328), .Z(n1331) );
  XNOR U4691 ( .A(x[725]), .B(y[725]), .Z(n3286) );
  XNOR U4692 ( .A(x[727]), .B(y[727]), .Z(n3284) );
  XOR U4693 ( .A(x[1494]), .B(y[1494]), .Z(n3283) );
  XNOR U4694 ( .A(n3284), .B(n3283), .Z(n3285) );
  XOR U4695 ( .A(n3286), .B(n3285), .Z(n3750) );
  XNOR U4696 ( .A(x[717]), .B(y[717]), .Z(n3251) );
  XNOR U4697 ( .A(x[719]), .B(y[719]), .Z(n3249) );
  XOR U4698 ( .A(x[1492]), .B(y[1492]), .Z(n3248) );
  XNOR U4699 ( .A(n3249), .B(n3248), .Z(n3250) );
  XOR U4700 ( .A(n3251), .B(n3250), .Z(n3747) );
  XNOR U4701 ( .A(x[721]), .B(y[721]), .Z(n3259) );
  XNOR U4702 ( .A(x[254]), .B(y[254]), .Z(n3257) );
  XOR U4703 ( .A(x[723]), .B(y[723]), .Z(n3256) );
  XNOR U4704 ( .A(n3257), .B(n3256), .Z(n3258) );
  XNOR U4705 ( .A(n3259), .B(n3258), .Z(n3748) );
  XNOR U4706 ( .A(n3747), .B(n3748), .Z(n3749) );
  XNOR U4707 ( .A(n3750), .B(n3749), .Z(n1330) );
  XOR U4708 ( .A(n1331), .B(n1330), .Z(n983) );
  XNOR U4709 ( .A(n982), .B(n983), .Z(n984) );
  XNOR U4710 ( .A(n985), .B(n984), .Z(n4325) );
  XNOR U4711 ( .A(x[1075]), .B(y[1075]), .Z(n1023) );
  XNOR U4712 ( .A(x[35]), .B(y[35]), .Z(n1020) );
  XNOR U4713 ( .A(x[1077]), .B(y[1077]), .Z(n1021) );
  XOR U4714 ( .A(n1020), .B(n1021), .Z(n1022) );
  XOR U4715 ( .A(n1023), .B(n1022), .Z(n4081) );
  XNOR U4716 ( .A(x[1063]), .B(y[1063]), .Z(n2579) );
  XNOR U4717 ( .A(x[25]), .B(y[25]), .Z(n2576) );
  XNOR U4718 ( .A(x[1065]), .B(y[1065]), .Z(n2577) );
  XOR U4719 ( .A(n2576), .B(n2577), .Z(n2578) );
  XOR U4720 ( .A(n2579), .B(n2578), .Z(n4078) );
  XNOR U4721 ( .A(x[1071]), .B(y[1071]), .Z(n2585) );
  XNOR U4722 ( .A(x[1073]), .B(y[1073]), .Z(n2582) );
  XNOR U4723 ( .A(x[1536]), .B(y[1536]), .Z(n2583) );
  XOR U4724 ( .A(n2582), .B(n2583), .Z(n2584) );
  XNOR U4725 ( .A(n2585), .B(n2584), .Z(n4079) );
  XNOR U4726 ( .A(n4078), .B(n4079), .Z(n4080) );
  XNOR U4727 ( .A(n4081), .B(n4080), .Z(n2001) );
  XNOR U4728 ( .A(x[1099]), .B(y[1099]), .Z(n993) );
  XNOR U4729 ( .A(x[51]), .B(y[51]), .Z(n991) );
  XOR U4730 ( .A(x[1101]), .B(y[1101]), .Z(n990) );
  XNOR U4731 ( .A(n991), .B(n990), .Z(n992) );
  XOR U4732 ( .A(n993), .B(n992), .Z(n1307) );
  XNOR U4733 ( .A(x[1091]), .B(y[1091]), .Z(n1033) );
  XNOR U4734 ( .A(x[320]), .B(y[320]), .Z(n1031) );
  XOR U4735 ( .A(x[1093]), .B(y[1093]), .Z(n1030) );
  XNOR U4736 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4737 ( .A(n1033), .B(n1032), .Z(n1304) );
  XNOR U4738 ( .A(x[1095]), .B(y[1095]), .Z(n997) );
  XNOR U4739 ( .A(x[47]), .B(y[47]), .Z(n995) );
  XOR U4740 ( .A(x[1097]), .B(y[1097]), .Z(n994) );
  XNOR U4741 ( .A(n995), .B(n994), .Z(n996) );
  XNOR U4742 ( .A(n997), .B(n996), .Z(n1305) );
  XNOR U4743 ( .A(n1307), .B(n1306), .Z(n1998) );
  XNOR U4744 ( .A(x[1087]), .B(y[1087]), .Z(n1037) );
  XNOR U4745 ( .A(x[41]), .B(y[41]), .Z(n1035) );
  XOR U4746 ( .A(x[1089]), .B(y[1089]), .Z(n1034) );
  XNOR U4747 ( .A(n1035), .B(n1034), .Z(n1036) );
  XOR U4748 ( .A(n1037), .B(n1036), .Z(n1312) );
  XNOR U4749 ( .A(x[1079]), .B(y[1079]), .Z(n1019) );
  XNOR U4750 ( .A(x[1081]), .B(y[1081]), .Z(n1017) );
  XOR U4751 ( .A(x[1538]), .B(y[1538]), .Z(n1016) );
  XNOR U4752 ( .A(n1017), .B(n1016), .Z(n1018) );
  XNOR U4753 ( .A(n1019), .B(n1018), .Z(n1310) );
  XNOR U4754 ( .A(x[1083]), .B(y[1083]), .Z(n1029) );
  XNOR U4755 ( .A(x[326]), .B(y[326]), .Z(n1027) );
  XOR U4756 ( .A(x[1085]), .B(y[1085]), .Z(n1026) );
  XNOR U4757 ( .A(n1027), .B(n1026), .Z(n1028) );
  XNOR U4758 ( .A(n1029), .B(n1028), .Z(n1311) );
  XOR U4759 ( .A(n1312), .B(n1313), .Z(n1999) );
  XOR U4760 ( .A(n1998), .B(n1999), .Z(n2000) );
  XOR U4761 ( .A(n2001), .B(n2000), .Z(n817) );
  XNOR U4762 ( .A(x[1007]), .B(y[1007]), .Z(n2527) );
  XNOR U4763 ( .A(x[1009]), .B(y[1009]), .Z(n2524) );
  XNOR U4764 ( .A(x[1528]), .B(y[1528]), .Z(n2525) );
  XOR U4765 ( .A(n2524), .B(n2525), .Z(n2526) );
  XOR U4766 ( .A(n2527), .B(n2526), .Z(n4191) );
  XNOR U4767 ( .A(x[991]), .B(y[991]), .Z(n1601) );
  XNOR U4768 ( .A(x[28]), .B(y[28]), .Z(n1598) );
  XNOR U4769 ( .A(x[993]), .B(y[993]), .Z(n1599) );
  XOR U4770 ( .A(n1598), .B(n1599), .Z(n1600) );
  XOR U4771 ( .A(n1601), .B(n1600), .Z(n4188) );
  XNOR U4772 ( .A(x[999]), .B(y[999]), .Z(n2515) );
  XNOR U4773 ( .A(x[18]), .B(y[18]), .Z(n2512) );
  XNOR U4774 ( .A(x[1001]), .B(y[1001]), .Z(n2513) );
  XOR U4775 ( .A(n2512), .B(n2513), .Z(n2514) );
  XNOR U4776 ( .A(n2515), .B(n2514), .Z(n4189) );
  XNOR U4777 ( .A(n4188), .B(n4189), .Z(n4190) );
  XNOR U4778 ( .A(n4191), .B(n4190), .Z(n2049) );
  XNOR U4779 ( .A(x[1055]), .B(y[1055]), .Z(n2555) );
  XNOR U4780 ( .A(x[19]), .B(y[19]), .Z(n2552) );
  XNOR U4781 ( .A(x[1057]), .B(y[1057]), .Z(n2553) );
  XOR U4782 ( .A(n2552), .B(n2553), .Z(n2554) );
  XOR U4783 ( .A(n2555), .B(n2554), .Z(n4257) );
  XNOR U4784 ( .A(x[1039]), .B(y[1039]), .Z(n967) );
  XNOR U4785 ( .A(x[1041]), .B(y[1041]), .Z(n964) );
  XNOR U4786 ( .A(x[1532]), .B(y[1532]), .Z(n965) );
  XOR U4787 ( .A(n964), .B(n965), .Z(n966) );
  XOR U4788 ( .A(n967), .B(n966), .Z(n4254) );
  XNOR U4789 ( .A(x[1047]), .B(y[1047]), .Z(n973) );
  XNOR U4790 ( .A(x[1049]), .B(y[1049]), .Z(n970) );
  XNOR U4791 ( .A(x[1534]), .B(y[1534]), .Z(n971) );
  XOR U4792 ( .A(n970), .B(n971), .Z(n972) );
  XNOR U4793 ( .A(n973), .B(n972), .Z(n4255) );
  XNOR U4794 ( .A(n4254), .B(n4255), .Z(n4256) );
  XNOR U4795 ( .A(n4257), .B(n4256), .Z(n2046) );
  XNOR U4796 ( .A(x[1031]), .B(y[1031]), .Z(n957) );
  XNOR U4797 ( .A(x[3]), .B(y[3]), .Z(n954) );
  XNOR U4798 ( .A(x[1033]), .B(y[1033]), .Z(n955) );
  XOR U4799 ( .A(n954), .B(n955), .Z(n956) );
  XOR U4800 ( .A(n957), .B(n956), .Z(n4263) );
  XNOR U4801 ( .A(x[1015]), .B(y[1015]), .Z(n1755) );
  XNOR U4802 ( .A(x[1017]), .B(y[1017]), .Z(n1753) );
  XNOR U4803 ( .A(x[1530]), .B(y[1530]), .Z(n1752) );
  XNOR U4804 ( .A(n1753), .B(n1752), .Z(n1754) );
  XNOR U4805 ( .A(n1755), .B(n1754), .Z(n4260) );
  XNOR U4806 ( .A(x[1023]), .B(y[1023]), .Z(n1749) );
  XNOR U4807 ( .A(x[2]), .B(y[2]), .Z(n1747) );
  XNOR U4808 ( .A(x[1025]), .B(y[1025]), .Z(n1746) );
  XNOR U4809 ( .A(n1747), .B(n1746), .Z(n1748) );
  XOR U4810 ( .A(n1749), .B(n1748), .Z(n4261) );
  XNOR U4811 ( .A(n4260), .B(n4261), .Z(n4262) );
  XNOR U4812 ( .A(n4263), .B(n4262), .Z(n2047) );
  XOR U4813 ( .A(n2046), .B(n2047), .Z(n2048) );
  XOR U4814 ( .A(n2049), .B(n2048), .Z(n814) );
  XNOR U4815 ( .A(x[1387]), .B(y[1387]), .Z(n2247) );
  XNOR U4816 ( .A(x[249]), .B(y[249]), .Z(n2245) );
  XOR U4817 ( .A(x[1389]), .B(y[1389]), .Z(n2244) );
  XNOR U4818 ( .A(n2245), .B(n2244), .Z(n2246) );
  XOR U4819 ( .A(n2247), .B(n2246), .Z(n4692) );
  XNOR U4820 ( .A(x[1383]), .B(y[1383]), .Z(n2251) );
  XNOR U4821 ( .A(x[245]), .B(y[245]), .Z(n2249) );
  XOR U4822 ( .A(x[1385]), .B(y[1385]), .Z(n2248) );
  XNOR U4823 ( .A(n2249), .B(n2248), .Z(n2250) );
  XNOR U4824 ( .A(n2251), .B(n2250), .Z(n4693) );
  XNOR U4825 ( .A(n4692), .B(n4693), .Z(n4694) );
  XNOR U4826 ( .A(x[1375]), .B(y[1375]), .Z(n1815) );
  XNOR U4827 ( .A(x[239]), .B(y[239]), .Z(n1813) );
  XNOR U4828 ( .A(x[1377]), .B(y[1377]), .Z(n1812) );
  XNOR U4829 ( .A(n1813), .B(n1812), .Z(n1814) );
  XNOR U4830 ( .A(n1815), .B(n1814), .Z(n4044) );
  XNOR U4831 ( .A(x[1391]), .B(y[1391]), .Z(n4791) );
  XNOR U4832 ( .A(x[1393]), .B(y[1393]), .Z(n4789) );
  XOR U4833 ( .A(x[1576]), .B(y[1576]), .Z(n4788) );
  XNOR U4834 ( .A(n4789), .B(n4788), .Z(n4790) );
  XNOR U4835 ( .A(n4791), .B(n4790), .Z(n4042) );
  XNOR U4836 ( .A(x[1403]), .B(y[1403]), .Z(n4917) );
  XNOR U4837 ( .A(x[126]), .B(y[126]), .Z(n4915) );
  XOR U4838 ( .A(x[1405]), .B(y[1405]), .Z(n4914) );
  XNOR U4839 ( .A(n4915), .B(n4914), .Z(n4916) );
  XNOR U4840 ( .A(n4917), .B(n4916), .Z(n4043) );
  XNOR U4841 ( .A(n4694), .B(n4695), .Z(n1053) );
  XNOR U4842 ( .A(x[1347]), .B(y[1347]), .Z(n4671) );
  XNOR U4843 ( .A(x[160]), .B(y[160]), .Z(n4669) );
  XOR U4844 ( .A(x[1349]), .B(y[1349]), .Z(n4668) );
  XNOR U4845 ( .A(n4669), .B(n4668), .Z(n4670) );
  XOR U4846 ( .A(n4671), .B(n4670), .Z(n1735) );
  XNOR U4847 ( .A(x[1351]), .B(y[1351]), .Z(n1825) );
  XNOR U4848 ( .A(x[223]), .B(y[223]), .Z(n1823) );
  XOR U4849 ( .A(x[1353]), .B(y[1353]), .Z(n1822) );
  XNOR U4850 ( .A(n1823), .B(n1822), .Z(n1824) );
  XOR U4851 ( .A(n1825), .B(n1824), .Z(n1732) );
  XNOR U4852 ( .A(x[1343]), .B(y[1343]), .Z(n4667) );
  XNOR U4853 ( .A(x[217]), .B(y[217]), .Z(n4665) );
  XOR U4854 ( .A(x[1345]), .B(y[1345]), .Z(n4664) );
  XNOR U4855 ( .A(n4665), .B(n4664), .Z(n4666) );
  XNOR U4856 ( .A(n4667), .B(n4666), .Z(n1733) );
  XNOR U4857 ( .A(n1732), .B(n1733), .Z(n1734) );
  XNOR U4858 ( .A(n1735), .B(n1734), .Z(n1050) );
  XNOR U4859 ( .A(x[1415]), .B(y[1415]), .Z(n1723) );
  XNOR U4860 ( .A(x[267]), .B(y[267]), .Z(n1721) );
  XOR U4861 ( .A(x[1417]), .B(y[1417]), .Z(n1720) );
  XNOR U4862 ( .A(n1721), .B(n1720), .Z(n1722) );
  XOR U4863 ( .A(n1723), .B(n1722), .Z(n4777) );
  XNOR U4864 ( .A(x[1335]), .B(y[1335]), .Z(n4783) );
  XNOR U4865 ( .A(x[1337]), .B(y[1337]), .Z(n4781) );
  XOR U4866 ( .A(x[1570]), .B(y[1570]), .Z(n4780) );
  XNOR U4867 ( .A(n4781), .B(n4780), .Z(n4782) );
  XOR U4868 ( .A(n4783), .B(n4782), .Z(n4774) );
  XNOR U4869 ( .A(x[1367]), .B(y[1367]), .Z(n4675) );
  XNOR U4870 ( .A(x[1369]), .B(y[1369]), .Z(n4673) );
  XOR U4871 ( .A(x[1574]), .B(y[1574]), .Z(n4672) );
  XNOR U4872 ( .A(n4673), .B(n4672), .Z(n4674) );
  XNOR U4873 ( .A(n4675), .B(n4674), .Z(n4775) );
  XNOR U4874 ( .A(n4774), .B(n4775), .Z(n4776) );
  XOR U4875 ( .A(n4777), .B(n4776), .Z(n1051) );
  XNOR U4876 ( .A(n1050), .B(n1051), .Z(n1052) );
  XNOR U4877 ( .A(n1053), .B(n1052), .Z(n815) );
  XNOR U4878 ( .A(n814), .B(n815), .Z(n816) );
  XNOR U4879 ( .A(n817), .B(n816), .Z(n4322) );
  XNOR U4880 ( .A(x[1195]), .B(y[1195]), .Z(n3015) );
  XNOR U4881 ( .A(x[117]), .B(y[117]), .Z(n3013) );
  XNOR U4882 ( .A(x[1197]), .B(y[1197]), .Z(n3012) );
  XNOR U4883 ( .A(n3013), .B(n3012), .Z(n3014) );
  XNOR U4884 ( .A(n3015), .B(n3014), .Z(n4343) );
  XNOR U4885 ( .A(x[1187]), .B(y[1187]), .Z(n2737) );
  XNOR U4886 ( .A(x[260]), .B(y[260]), .Z(n2735) );
  XOR U4887 ( .A(x[1189]), .B(y[1189]), .Z(n2734) );
  XNOR U4888 ( .A(n2735), .B(n2734), .Z(n2736) );
  XOR U4889 ( .A(n2737), .B(n2736), .Z(n4340) );
  XNOR U4890 ( .A(x[1191]), .B(y[1191]), .Z(n3009) );
  XNOR U4891 ( .A(x[113]), .B(y[113]), .Z(n3007) );
  XNOR U4892 ( .A(x[1193]), .B(y[1193]), .Z(n3006) );
  XNOR U4893 ( .A(n3007), .B(n3006), .Z(n3008) );
  XOR U4894 ( .A(n3009), .B(n3008), .Z(n4341) );
  XNOR U4895 ( .A(n4340), .B(n4341), .Z(n4342) );
  XOR U4896 ( .A(n4343), .B(n4342), .Z(n3327) );
  XNOR U4897 ( .A(x[1207]), .B(y[1207]), .Z(n3374) );
  XNOR U4898 ( .A(x[1209]), .B(y[1209]), .Z(n3372) );
  XOR U4899 ( .A(x[1554]), .B(y[1554]), .Z(n3371) );
  XNOR U4900 ( .A(n3372), .B(n3371), .Z(n3373) );
  XOR U4901 ( .A(n3374), .B(n3373), .Z(n4587) );
  XNOR U4902 ( .A(x[1203]), .B(y[1203]), .Z(n1155) );
  XNOR U4903 ( .A(x[123]), .B(y[123]), .Z(n1153) );
  XOR U4904 ( .A(x[1205]), .B(y[1205]), .Z(n1152) );
  XNOR U4905 ( .A(n1153), .B(n1152), .Z(n1154) );
  XOR U4906 ( .A(n1155), .B(n1154), .Z(n4584) );
  XNOR U4907 ( .A(x[1199]), .B(y[1199]), .Z(n2741) );
  XNOR U4908 ( .A(x[1201]), .B(y[1201]), .Z(n2739) );
  XOR U4909 ( .A(x[1552]), .B(y[1552]), .Z(n2738) );
  XNOR U4910 ( .A(n2739), .B(n2738), .Z(n2740) );
  XNOR U4911 ( .A(n2741), .B(n2740), .Z(n4585) );
  XNOR U4912 ( .A(n4584), .B(n4585), .Z(n4586) );
  XOR U4913 ( .A(n4587), .B(n4586), .Z(n3328) );
  XOR U4914 ( .A(n3327), .B(n3328), .Z(n3329) );
  XNOR U4915 ( .A(x[1183]), .B(y[1183]), .Z(n3217) );
  XNOR U4916 ( .A(x[107]), .B(y[107]), .Z(n3215) );
  XOR U4917 ( .A(x[1185]), .B(y[1185]), .Z(n3214) );
  XNOR U4918 ( .A(n3215), .B(n3214), .Z(n3216) );
  XOR U4919 ( .A(n3217), .B(n3216), .Z(n4455) );
  XNOR U4920 ( .A(x[1175]), .B(y[1175]), .Z(n2707) );
  XNOR U4921 ( .A(x[1177]), .B(y[1177]), .Z(n2705) );
  XOR U4922 ( .A(x[1550]), .B(y[1550]), .Z(n2704) );
  XNOR U4923 ( .A(n2705), .B(n2704), .Z(n2706) );
  XNOR U4924 ( .A(n2707), .B(n2706), .Z(n4452) );
  XNOR U4925 ( .A(x[1179]), .B(y[1179]), .Z(n2703) );
  XNOR U4926 ( .A(x[266]), .B(y[266]), .Z(n2701) );
  XOR U4927 ( .A(x[1181]), .B(y[1181]), .Z(n2700) );
  XNOR U4928 ( .A(n2701), .B(n2700), .Z(n2702) );
  XNOR U4929 ( .A(n2703), .B(n2702), .Z(n4453) );
  XNOR U4930 ( .A(n4455), .B(n4454), .Z(n3330) );
  XOR U4931 ( .A(n3329), .B(n3330), .Z(n2663) );
  XNOR U4932 ( .A(x[1219]), .B(y[1219]), .Z(n2387) );
  XNOR U4933 ( .A(x[240]), .B(y[240]), .Z(n2385) );
  XOR U4934 ( .A(x[1221]), .B(y[1221]), .Z(n2384) );
  XNOR U4935 ( .A(n2385), .B(n2384), .Z(n2386) );
  XOR U4936 ( .A(n2387), .B(n2386), .Z(n4509) );
  XNOR U4937 ( .A(x[1211]), .B(y[1211]), .Z(n3428) );
  XNOR U4938 ( .A(x[246]), .B(y[246]), .Z(n3426) );
  XOR U4939 ( .A(x[1213]), .B(y[1213]), .Z(n3425) );
  XNOR U4940 ( .A(n3426), .B(n3425), .Z(n3427) );
  XNOR U4941 ( .A(n3428), .B(n3427), .Z(n4506) );
  XNOR U4942 ( .A(x[1215]), .B(y[1215]), .Z(n3550) );
  XNOR U4943 ( .A(x[129]), .B(y[129]), .Z(n3548) );
  XOR U4944 ( .A(x[1217]), .B(y[1217]), .Z(n3547) );
  XNOR U4945 ( .A(n3548), .B(n3547), .Z(n3549) );
  XNOR U4946 ( .A(n3550), .B(n3549), .Z(n4507) );
  XNOR U4947 ( .A(n4509), .B(n4508), .Z(n2674) );
  XNOR U4948 ( .A(x[1239]), .B(y[1239]), .Z(n1501) );
  XNOR U4949 ( .A(x[1241]), .B(y[1241]), .Z(n1498) );
  XNOR U4950 ( .A(x[1558]), .B(y[1558]), .Z(n1499) );
  XOR U4951 ( .A(n1498), .B(n1499), .Z(n1500) );
  XOR U4952 ( .A(n1501), .B(n1500), .Z(n4831) );
  XNOR U4953 ( .A(x[1235]), .B(y[1235]), .Z(n1693) );
  XNOR U4954 ( .A(x[145]), .B(y[145]), .Z(n1690) );
  XNOR U4955 ( .A(x[1237]), .B(y[1237]), .Z(n1691) );
  XOR U4956 ( .A(n1690), .B(n1691), .Z(n1692) );
  XOR U4957 ( .A(n1693), .B(n1692), .Z(n4828) );
  XNOR U4958 ( .A(x[1467]), .B(y[1467]), .Z(n3700) );
  XNOR U4959 ( .A(x[86]), .B(y[86]), .Z(n3697) );
  XNOR U4960 ( .A(x[1469]), .B(y[1469]), .Z(n3698) );
  XOR U4961 ( .A(n3697), .B(n3698), .Z(n3699) );
  XNOR U4962 ( .A(n3700), .B(n3699), .Z(n4829) );
  XNOR U4963 ( .A(n4828), .B(n4829), .Z(n4830) );
  XNOR U4964 ( .A(n4831), .B(n4830), .Z(n2673) );
  XNOR U4965 ( .A(x[1231]), .B(y[1231]), .Z(n1699) );
  XNOR U4966 ( .A(x[1233]), .B(y[1233]), .Z(n1697) );
  XOR U4967 ( .A(x[1556]), .B(y[1556]), .Z(n1696) );
  XNOR U4968 ( .A(n1697), .B(n1696), .Z(n1698) );
  XOR U4969 ( .A(n1699), .B(n1698), .Z(n1885) );
  XNOR U4970 ( .A(x[1223]), .B(y[1223]), .Z(n2381) );
  XNOR U4971 ( .A(x[135]), .B(y[135]), .Z(n2378) );
  XNOR U4972 ( .A(x[1225]), .B(y[1225]), .Z(n2379) );
  XOR U4973 ( .A(n2378), .B(n2379), .Z(n2380) );
  XOR U4974 ( .A(n2381), .B(n2380), .Z(n1882) );
  XNOR U4975 ( .A(x[1227]), .B(y[1227]), .Z(n1591) );
  XNOR U4976 ( .A(x[139]), .B(y[139]), .Z(n1589) );
  XOR U4977 ( .A(x[1229]), .B(y[1229]), .Z(n1588) );
  XNOR U4978 ( .A(n1589), .B(n1588), .Z(n1590) );
  XNOR U4979 ( .A(n1591), .B(n1590), .Z(n1883) );
  XNOR U4980 ( .A(n1882), .B(n1883), .Z(n1884) );
  XOR U4981 ( .A(n1885), .B(n1884), .Z(n2672) );
  XOR U4982 ( .A(n2673), .B(n2672), .Z(n2675) );
  XNOR U4983 ( .A(n2674), .B(n2675), .Z(n2660) );
  XNOR U4984 ( .A(x[1311]), .B(y[1311]), .Z(n4865) );
  XNOR U4985 ( .A(x[195]), .B(y[195]), .Z(n4863) );
  XOR U4986 ( .A(x[1313]), .B(y[1313]), .Z(n4862) );
  XNOR U4987 ( .A(n4863), .B(n4862), .Z(n4864) );
  XOR U4988 ( .A(n4865), .B(n4864), .Z(n1683) );
  XNOR U4989 ( .A(x[1307]), .B(y[1307]), .Z(n4869) );
  XNOR U4990 ( .A(x[186]), .B(y[186]), .Z(n4867) );
  XOR U4991 ( .A(x[1309]), .B(y[1309]), .Z(n4866) );
  XNOR U4992 ( .A(n4867), .B(n4866), .Z(n4868) );
  XOR U4993 ( .A(n4869), .B(n4868), .Z(n1680) );
  XNOR U4994 ( .A(x[1431]), .B(y[1431]), .Z(n2499) );
  XNOR U4995 ( .A(x[1433]), .B(y[1433]), .Z(n2497) );
  XOR U4996 ( .A(x[1582]), .B(y[1582]), .Z(n2496) );
  XNOR U4997 ( .A(n2497), .B(n2496), .Z(n2498) );
  XNOR U4998 ( .A(n2499), .B(n2498), .Z(n1681) );
  XNOR U4999 ( .A(n1680), .B(n1681), .Z(n1682) );
  XNOR U5000 ( .A(n1683), .B(n1682), .Z(n1889) );
  XNOR U5001 ( .A(x[1303]), .B(y[1303]), .Z(n4859) );
  XNOR U5002 ( .A(x[1305]), .B(y[1305]), .Z(n4857) );
  XNOR U5003 ( .A(x[1566]), .B(y[1566]), .Z(n4856) );
  XNOR U5004 ( .A(n4857), .B(n4856), .Z(n4858) );
  XNOR U5005 ( .A(n4859), .B(n4858), .Z(n1741) );
  XNOR U5006 ( .A(x[1299]), .B(y[1299]), .Z(n4853) );
  XNOR U5007 ( .A(x[189]), .B(y[189]), .Z(n4851) );
  XNOR U5008 ( .A(x[1301]), .B(y[1301]), .Z(n4850) );
  XNOR U5009 ( .A(n4851), .B(n4850), .Z(n4852) );
  XNOR U5010 ( .A(n4853), .B(n4852), .Z(n1738) );
  XNOR U5011 ( .A(x[1435]), .B(y[1435]), .Z(n1009) );
  XNOR U5012 ( .A(x[106]), .B(y[106]), .Z(n1007) );
  XOR U5013 ( .A(x[1437]), .B(y[1437]), .Z(n1006) );
  XNOR U5014 ( .A(n1007), .B(n1006), .Z(n1008) );
  XNOR U5015 ( .A(n1009), .B(n1008), .Z(n1739) );
  XNOR U5016 ( .A(n1738), .B(n1739), .Z(n1740) );
  XOR U5017 ( .A(n1741), .B(n1740), .Z(n1888) );
  XOR U5018 ( .A(n1889), .B(n1888), .Z(n1891) );
  XNOR U5019 ( .A(x[1295]), .B(y[1295]), .Z(n2243) );
  XNOR U5020 ( .A(x[1297]), .B(y[1297]), .Z(n2241) );
  XOR U5021 ( .A(x[1564]), .B(y[1564]), .Z(n2240) );
  XNOR U5022 ( .A(n2241), .B(n2240), .Z(n2242) );
  XOR U5023 ( .A(n2243), .B(n2242), .Z(n2509) );
  XNOR U5024 ( .A(x[1291]), .B(y[1291]), .Z(n2239) );
  XNOR U5025 ( .A(x[183]), .B(y[183]), .Z(n2237) );
  XOR U5026 ( .A(x[1293]), .B(y[1293]), .Z(n2236) );
  XNOR U5027 ( .A(n2237), .B(n2236), .Z(n2238) );
  XOR U5028 ( .A(n2239), .B(n2238), .Z(n2506) );
  XNOR U5029 ( .A(x[1439]), .B(y[1439]), .Z(n1005) );
  XNOR U5030 ( .A(x[283]), .B(y[283]), .Z(n1003) );
  XOR U5031 ( .A(x[1441]), .B(y[1441]), .Z(n1002) );
  XNOR U5032 ( .A(n1003), .B(n1002), .Z(n1004) );
  XNOR U5033 ( .A(n1005), .B(n1004), .Z(n2507) );
  XNOR U5034 ( .A(n2506), .B(n2507), .Z(n2508) );
  XNOR U5035 ( .A(n2509), .B(n2508), .Z(n1890) );
  XOR U5036 ( .A(n1891), .B(n1890), .Z(n2661) );
  XNOR U5037 ( .A(n2660), .B(n2661), .Z(n2662) );
  XOR U5038 ( .A(n2663), .B(n2662), .Z(n4323) );
  XNOR U5039 ( .A(n4322), .B(n4323), .Z(n4324) );
  XOR U5040 ( .A(n4325), .B(n4324), .Z(n803) );
  XOR U5041 ( .A(n802), .B(n803), .Z(n805) );
  XNOR U5042 ( .A(x[378]), .B(y[378]), .Z(n1421) );
  XNOR U5043 ( .A(x[370]), .B(y[370]), .Z(n1419) );
  XOR U5044 ( .A(x[374]), .B(y[374]), .Z(n1418) );
  XNOR U5045 ( .A(n1419), .B(n1418), .Z(n1420) );
  XOR U5046 ( .A(n1421), .B(n1420), .Z(n1539) );
  XNOR U5047 ( .A(x[408]), .B(y[408]), .Z(n1523) );
  XNOR U5048 ( .A(x[396]), .B(y[396]), .Z(n1521) );
  XOR U5049 ( .A(x[764]), .B(y[764]), .Z(n1520) );
  XNOR U5050 ( .A(n1521), .B(n1520), .Z(n1522) );
  XNOR U5051 ( .A(n1523), .B(n1522), .Z(n1536) );
  XNOR U5052 ( .A(x[1563]), .B(y[1563]), .Z(n2021) );
  XNOR U5053 ( .A(x[26]), .B(y[26]), .Z(n2019) );
  XOR U5054 ( .A(x[1565]), .B(y[1565]), .Z(n2018) );
  XNOR U5055 ( .A(n2019), .B(n2018), .Z(n2020) );
  XNOR U5056 ( .A(n2021), .B(n2020), .Z(n1537) );
  XNOR U5057 ( .A(n1539), .B(n1538), .Z(n3984) );
  XNOR U5058 ( .A(x[342]), .B(y[342]), .Z(n1639) );
  XNOR U5059 ( .A(x[334]), .B(y[334]), .Z(n1637) );
  XOR U5060 ( .A(x[338]), .B(y[338]), .Z(n1636) );
  XNOR U5061 ( .A(n1637), .B(n1636), .Z(n1638) );
  XOR U5062 ( .A(n1639), .B(n1638), .Z(n1784) );
  XNOR U5063 ( .A(x[352]), .B(y[352]), .Z(n3634) );
  XNOR U5064 ( .A(x[348]), .B(y[348]), .Z(n3632) );
  XOR U5065 ( .A(x[746]), .B(y[746]), .Z(n3631) );
  XNOR U5066 ( .A(n3632), .B(n3631), .Z(n3633) );
  XNOR U5067 ( .A(n3634), .B(n3633), .Z(n1782) );
  XNOR U5068 ( .A(x[883]), .B(y[883]), .Z(n4827) );
  XNOR U5069 ( .A(x[116]), .B(y[116]), .Z(n4825) );
  XOR U5070 ( .A(x[885]), .B(y[885]), .Z(n4824) );
  XNOR U5071 ( .A(n4825), .B(n4824), .Z(n4826) );
  XNOR U5072 ( .A(n4827), .B(n4826), .Z(n1783) );
  XOR U5073 ( .A(n1784), .B(n1785), .Z(n3985) );
  XOR U5074 ( .A(n3984), .B(n3985), .Z(n3986) );
  XNOR U5075 ( .A(x[414]), .B(y[414]), .Z(n3664) );
  XNOR U5076 ( .A(x[410]), .B(y[410]), .Z(n3662) );
  XOR U5077 ( .A(x[768]), .B(y[768]), .Z(n3661) );
  XNOR U5078 ( .A(n3662), .B(n3661), .Z(n3663) );
  XOR U5079 ( .A(n3664), .B(n3663), .Z(n1437) );
  XNOR U5080 ( .A(x[424]), .B(y[424]), .Z(n2193) );
  XNOR U5081 ( .A(x[416]), .B(y[416]), .Z(n2190) );
  XNOR U5082 ( .A(x[422]), .B(y[422]), .Z(n2191) );
  XOR U5083 ( .A(n2190), .B(n2191), .Z(n2192) );
  XOR U5084 ( .A(n2193), .B(n2192), .Z(n1434) );
  XNOR U5085 ( .A(x[875]), .B(y[875]), .Z(n4817) );
  XNOR U5086 ( .A(x[124]), .B(y[124]), .Z(n4815) );
  XOR U5087 ( .A(x[877]), .B(y[877]), .Z(n4814) );
  XNOR U5088 ( .A(n4815), .B(n4814), .Z(n4816) );
  XNOR U5089 ( .A(n4817), .B(n4816), .Z(n1435) );
  XNOR U5090 ( .A(n1434), .B(n1435), .Z(n1436) );
  XNOR U5091 ( .A(n1437), .B(n1436), .Z(n3987) );
  XOR U5092 ( .A(n3986), .B(n3987), .Z(n4273) );
  XNOR U5093 ( .A(x[292]), .B(y[292]), .Z(n3197) );
  XNOR U5094 ( .A(x[278]), .B(y[278]), .Z(n3195) );
  XOR U5095 ( .A(x[284]), .B(y[284]), .Z(n3194) );
  XNOR U5096 ( .A(n3195), .B(n3194), .Z(n3196) );
  XOR U5097 ( .A(n3197), .B(n3196), .Z(n4771) );
  XNOR U5098 ( .A(x[304]), .B(y[304]), .Z(n2401) );
  XNOR U5099 ( .A(x[298]), .B(y[298]), .Z(n2399) );
  XOR U5100 ( .A(x[728]), .B(y[728]), .Z(n2398) );
  XNOR U5101 ( .A(n2399), .B(n2398), .Z(n2400) );
  XOR U5102 ( .A(n2401), .B(n2400), .Z(n4768) );
  XNOR U5103 ( .A(x[891]), .B(y[891]), .Z(n4879) );
  XNOR U5104 ( .A(x[446]), .B(y[446]), .Z(n4877) );
  XOR U5105 ( .A(x[893]), .B(y[893]), .Z(n4876) );
  XNOR U5106 ( .A(n4877), .B(n4876), .Z(n4878) );
  XNOR U5107 ( .A(n4879), .B(n4878), .Z(n4769) );
  XNOR U5108 ( .A(n4768), .B(n4769), .Z(n4770) );
  XNOR U5109 ( .A(n4771), .B(n4770), .Z(n1341) );
  XNOR U5110 ( .A(x[312]), .B(y[312]), .Z(n2397) );
  XNOR U5111 ( .A(x[308]), .B(y[308]), .Z(n2395) );
  XOR U5112 ( .A(x[732]), .B(y[732]), .Z(n2394) );
  XNOR U5113 ( .A(n2395), .B(n2394), .Z(n2396) );
  XOR U5114 ( .A(n2397), .B(n2396), .Z(n1677) );
  XNOR U5115 ( .A(x[328]), .B(y[328]), .Z(n1643) );
  XNOR U5116 ( .A(x[314]), .B(y[314]), .Z(n1641) );
  XOR U5117 ( .A(x[318]), .B(y[318]), .Z(n1640) );
  XNOR U5118 ( .A(n1641), .B(n1640), .Z(n1642) );
  XOR U5119 ( .A(n1643), .B(n1642), .Z(n1674) );
  XNOR U5120 ( .A(x[1559]), .B(y[1559]), .Z(n3790) );
  XNOR U5121 ( .A(x[1561]), .B(y[1561]), .Z(n3788) );
  XOR U5122 ( .A(x[1598]), .B(y[1598]), .Z(n3787) );
  XNOR U5123 ( .A(n3788), .B(n3787), .Z(n3789) );
  XNOR U5124 ( .A(n3790), .B(n3789), .Z(n1675) );
  XNOR U5125 ( .A(n1674), .B(n1675), .Z(n1676) );
  XOR U5126 ( .A(n1677), .B(n1676), .Z(n1340) );
  XNOR U5127 ( .A(n1341), .B(n1340), .Z(n1342) );
  XNOR U5128 ( .A(x[242]), .B(y[242]), .Z(n2409) );
  XNOR U5129 ( .A(x[232]), .B(y[232]), .Z(n2407) );
  XNOR U5130 ( .A(x[236]), .B(y[236]), .Z(n2406) );
  XNOR U5131 ( .A(n2407), .B(n2406), .Z(n2408) );
  XNOR U5132 ( .A(n2409), .B(n2408), .Z(n4527) );
  XNOR U5133 ( .A(x[1555]), .B(y[1555]), .Z(n2301) );
  XNOR U5134 ( .A(x[365]), .B(y[365]), .Z(n2299) );
  XOR U5135 ( .A(x[1557]), .B(y[1557]), .Z(n2298) );
  XNOR U5136 ( .A(n2299), .B(n2298), .Z(n2300) );
  XOR U5137 ( .A(n2301), .B(n2300), .Z(n4524) );
  XNOR U5138 ( .A(x[264]), .B(y[264]), .Z(n3296) );
  XNOR U5139 ( .A(x[256]), .B(y[256]), .Z(n3294) );
  XOR U5140 ( .A(x[714]), .B(y[714]), .Z(n3293) );
  XNOR U5141 ( .A(n3294), .B(n3293), .Z(n3295) );
  XNOR U5142 ( .A(n3296), .B(n3295), .Z(n4525) );
  XNOR U5143 ( .A(n4524), .B(n4525), .Z(n4526) );
  XOR U5144 ( .A(n4527), .B(n4526), .Z(n1343) );
  XOR U5145 ( .A(n1342), .B(n1343), .Z(n4270) );
  XNOR U5146 ( .A(x[150]), .B(y[150]), .Z(n2985) );
  XNOR U5147 ( .A(x[142]), .B(y[142]), .Z(n2982) );
  XNOR U5148 ( .A(x[674]), .B(y[674]), .Z(n2983) );
  XOR U5149 ( .A(n2982), .B(n2983), .Z(n2984) );
  XOR U5150 ( .A(n2985), .B(n2984), .Z(n4617) );
  XNOR U5151 ( .A(x[174]), .B(y[174]), .Z(n3109) );
  XNOR U5152 ( .A(x[168]), .B(y[168]), .Z(n3107) );
  XOR U5153 ( .A(x[170]), .B(y[170]), .Z(n3106) );
  XNOR U5154 ( .A(n3107), .B(n3106), .Z(n3108) );
  XOR U5155 ( .A(n3109), .B(n3108), .Z(n4614) );
  XNOR U5156 ( .A(x[907]), .B(y[907]), .Z(n4883) );
  XNOR U5157 ( .A(x[96]), .B(y[96]), .Z(n4880) );
  XNOR U5158 ( .A(x[909]), .B(y[909]), .Z(n4881) );
  XOR U5159 ( .A(n4880), .B(n4881), .Z(n4882) );
  XNOR U5160 ( .A(n4883), .B(n4882), .Z(n4615) );
  XNOR U5161 ( .A(n4614), .B(n4615), .Z(n4616) );
  XNOR U5162 ( .A(n4617), .B(n4616), .Z(n4465) );
  XNOR U5163 ( .A(x[194]), .B(y[194]), .Z(n2291) );
  XNOR U5164 ( .A(x[176]), .B(y[176]), .Z(n2289) );
  XOR U5165 ( .A(x[188]), .B(y[188]), .Z(n2288) );
  XNOR U5166 ( .A(n2289), .B(n2288), .Z(n2290) );
  XOR U5167 ( .A(n2291), .B(n2290), .Z(n1861) );
  XNOR U5168 ( .A(x[1551]), .B(y[1551]), .Z(n2347) );
  XNOR U5169 ( .A(x[1553]), .B(y[1553]), .Z(n2345) );
  XOR U5170 ( .A(x[1596]), .B(y[1596]), .Z(n2344) );
  XNOR U5171 ( .A(n2345), .B(n2344), .Z(n2346) );
  XOR U5172 ( .A(n2347), .B(n2346), .Z(n1858) );
  XNOR U5173 ( .A(x[202]), .B(y[202]), .Z(n2329) );
  XNOR U5174 ( .A(x[196]), .B(y[196]), .Z(n2327) );
  XOR U5175 ( .A(x[692]), .B(y[692]), .Z(n2326) );
  XNOR U5176 ( .A(n2327), .B(n2326), .Z(n2328) );
  XNOR U5177 ( .A(n2329), .B(n2328), .Z(n1859) );
  XNOR U5178 ( .A(n1858), .B(n1859), .Z(n1860) );
  XNOR U5179 ( .A(n1861), .B(n1860), .Z(n4464) );
  XNOR U5180 ( .A(n4465), .B(n4464), .Z(n4467) );
  XNOR U5181 ( .A(x[210]), .B(y[210]), .Z(n2325) );
  XNOR U5182 ( .A(x[204]), .B(y[204]), .Z(n2323) );
  XOR U5183 ( .A(x[696]), .B(y[696]), .Z(n2322) );
  XNOR U5184 ( .A(n2323), .B(n2322), .Z(n2324) );
  XOR U5185 ( .A(n2325), .B(n2324), .Z(n1215) );
  XNOR U5186 ( .A(x[230]), .B(y[230]), .Z(n2415) );
  XNOR U5187 ( .A(x[214]), .B(y[214]), .Z(n2413) );
  XOR U5188 ( .A(x[222]), .B(y[222]), .Z(n2412) );
  XNOR U5189 ( .A(n2413), .B(n2412), .Z(n2414) );
  XOR U5190 ( .A(n2415), .B(n2414), .Z(n1212) );
  XNOR U5191 ( .A(x[899]), .B(y[899]), .Z(n4889) );
  XNOR U5192 ( .A(x[440]), .B(y[440]), .Z(n4886) );
  XNOR U5193 ( .A(x[901]), .B(y[901]), .Z(n4887) );
  XOR U5194 ( .A(n4886), .B(n4887), .Z(n4888) );
  XNOR U5195 ( .A(n4889), .B(n4888), .Z(n1213) );
  XNOR U5196 ( .A(n1212), .B(n1213), .Z(n1214) );
  XNOR U5197 ( .A(n1215), .B(n1214), .Z(n4466) );
  XOR U5198 ( .A(n4467), .B(n4466), .Z(n4271) );
  XOR U5199 ( .A(n4270), .B(n4271), .Z(n4272) );
  XNOR U5200 ( .A(n4273), .B(n4272), .Z(n2656) );
  XNOR U5201 ( .A(x[265]), .B(y[265]), .Z(n2771) );
  XNOR U5202 ( .A(x[269]), .B(y[269]), .Z(n2769) );
  XOR U5203 ( .A(x[402]), .B(y[402]), .Z(n2768) );
  XNOR U5204 ( .A(n2769), .B(n2768), .Z(n2770) );
  XOR U5205 ( .A(n2771), .B(n2770), .Z(n3350) );
  XNOR U5206 ( .A(x[247]), .B(y[247]), .Z(n3075) );
  XNOR U5207 ( .A(x[251]), .B(y[251]), .Z(n3073) );
  XOR U5208 ( .A(x[253]), .B(y[253]), .Z(n3072) );
  XNOR U5209 ( .A(n3073), .B(n3072), .Z(n3074) );
  XOR U5210 ( .A(n3075), .B(n3074), .Z(n3347) );
  XNOR U5211 ( .A(x[979]), .B(y[979]), .Z(n4737) );
  XNOR U5212 ( .A(x[34]), .B(y[34]), .Z(n4735) );
  XOR U5213 ( .A(x[981]), .B(y[981]), .Z(n4734) );
  XNOR U5214 ( .A(n4735), .B(n4734), .Z(n4736) );
  XNOR U5215 ( .A(n4737), .B(n4736), .Z(n3348) );
  XNOR U5216 ( .A(n3347), .B(n3348), .Z(n3349) );
  XNOR U5217 ( .A(n3350), .B(n3349), .Z(n1645) );
  XNOR U5218 ( .A(x[235]), .B(y[235]), .Z(n875) );
  XNOR U5219 ( .A(x[237]), .B(y[237]), .Z(n872) );
  XNOR U5220 ( .A(x[432]), .B(y[432]), .Z(n873) );
  XOR U5221 ( .A(n872), .B(n873), .Z(n874) );
  XOR U5222 ( .A(n875), .B(n874), .Z(n3245) );
  XNOR U5223 ( .A(x[225]), .B(y[225]), .Z(n3975) );
  XNOR U5224 ( .A(x[229]), .B(y[229]), .Z(n3972) );
  XNOR U5225 ( .A(x[231]), .B(y[231]), .Z(n3973) );
  XOR U5226 ( .A(n3972), .B(n3973), .Z(n3974) );
  XOR U5227 ( .A(n3975), .B(n3974), .Z(n3242) );
  XNOR U5228 ( .A(x[1515]), .B(y[1515]), .Z(n3618) );
  XNOR U5229 ( .A(x[337]), .B(y[337]), .Z(n3615) );
  XNOR U5230 ( .A(x[1517]), .B(y[1517]), .Z(n3616) );
  XOR U5231 ( .A(n3615), .B(n3616), .Z(n3617) );
  XNOR U5232 ( .A(n3618), .B(n3617), .Z(n3243) );
  XNOR U5233 ( .A(n3242), .B(n3243), .Z(n3244) );
  XOR U5234 ( .A(n3245), .B(n3244), .Z(n1644) );
  XOR U5235 ( .A(n1645), .B(n1644), .Z(n1647) );
  XNOR U5236 ( .A(x[215]), .B(y[215]), .Z(n3963) );
  XNOR U5237 ( .A(x[219]), .B(y[219]), .Z(n3960) );
  XNOR U5238 ( .A(x[221]), .B(y[221]), .Z(n3961) );
  XOR U5239 ( .A(n3960), .B(n3961), .Z(n3962) );
  XOR U5240 ( .A(n3963), .B(n3962), .Z(n3290) );
  XNOR U5241 ( .A(x[209]), .B(y[209]), .Z(n3969) );
  XNOR U5242 ( .A(x[213]), .B(y[213]), .Z(n3966) );
  XNOR U5243 ( .A(x[450]), .B(y[450]), .Z(n3967) );
  XOR U5244 ( .A(n3966), .B(n3967), .Z(n3968) );
  XOR U5245 ( .A(n3969), .B(n3968), .Z(n3287) );
  XNOR U5246 ( .A(x[971]), .B(y[971]), .Z(n3606) );
  XNOR U5247 ( .A(x[42]), .B(y[42]), .Z(n3603) );
  XNOR U5248 ( .A(x[973]), .B(y[973]), .Z(n3604) );
  XOR U5249 ( .A(n3603), .B(n3604), .Z(n3605) );
  XNOR U5250 ( .A(n3606), .B(n3605), .Z(n3288) );
  XNOR U5251 ( .A(n3287), .B(n3288), .Z(n3289) );
  XNOR U5252 ( .A(n3290), .B(n3289), .Z(n1646) );
  XNOR U5253 ( .A(n1647), .B(n1646), .Z(n1187) );
  XNOR U5254 ( .A(x[141]), .B(y[141]), .Z(n3921) );
  XNOR U5255 ( .A(x[143]), .B(y[143]), .Z(n3919) );
  XOR U5256 ( .A(x[498]), .B(y[498]), .Z(n3918) );
  XNOR U5257 ( .A(n3919), .B(n3918), .Z(n3920) );
  XOR U5258 ( .A(n3921), .B(n3920), .Z(n1443) );
  XNOR U5259 ( .A(x[131]), .B(y[131]), .Z(n3913) );
  XNOR U5260 ( .A(x[133]), .B(y[133]), .Z(n3911) );
  XOR U5261 ( .A(x[137]), .B(y[137]), .Z(n3910) );
  XNOR U5262 ( .A(n3911), .B(n3910), .Z(n3912) );
  XOR U5263 ( .A(n3913), .B(n3912), .Z(n1440) );
  XNOR U5264 ( .A(x[955]), .B(y[955]), .Z(n4713) );
  XNOR U5265 ( .A(x[406]), .B(y[406]), .Z(n4711) );
  XOR U5266 ( .A(x[957]), .B(y[957]), .Z(n4710) );
  XNOR U5267 ( .A(n4711), .B(n4710), .Z(n4712) );
  XNOR U5268 ( .A(n4713), .B(n4712), .Z(n1441) );
  XNOR U5269 ( .A(n1440), .B(n1441), .Z(n1442) );
  XNOR U5270 ( .A(n1443), .B(n1442), .Z(n4959) );
  XNOR U5271 ( .A(x[121]), .B(y[121]), .Z(n3917) );
  XNOR U5272 ( .A(x[125]), .B(y[125]), .Z(n3915) );
  XOR U5273 ( .A(x[127]), .B(y[127]), .Z(n3914) );
  XNOR U5274 ( .A(n3915), .B(n3914), .Z(n3916) );
  XOR U5275 ( .A(n3917), .B(n3916), .Z(n1545) );
  XNOR U5276 ( .A(x[109]), .B(y[109]), .Z(n889) );
  XNOR U5277 ( .A(x[111]), .B(y[111]), .Z(n887) );
  XOR U5278 ( .A(x[522]), .B(y[522]), .Z(n886) );
  XNOR U5279 ( .A(n887), .B(n886), .Z(n888) );
  XOR U5280 ( .A(n889), .B(n888), .Z(n1542) );
  XNOR U5281 ( .A(x[1527]), .B(y[1527]), .Z(n1613) );
  XNOR U5282 ( .A(x[1529]), .B(y[1529]), .Z(n1611) );
  XOR U5283 ( .A(x[1594]), .B(y[1594]), .Z(n1610) );
  XNOR U5284 ( .A(n1611), .B(n1610), .Z(n1612) );
  XNOR U5285 ( .A(n1613), .B(n1612), .Z(n1543) );
  XNOR U5286 ( .A(n1542), .B(n1543), .Z(n1544) );
  XOR U5287 ( .A(n1545), .B(n1544), .Z(n4958) );
  XOR U5288 ( .A(n4959), .B(n4958), .Z(n4961) );
  XNOR U5289 ( .A(x[89]), .B(y[89]), .Z(n913) );
  XNOR U5290 ( .A(x[93]), .B(y[93]), .Z(n911) );
  XOR U5291 ( .A(x[97]), .B(y[97]), .Z(n910) );
  XNOR U5292 ( .A(n911), .B(n910), .Z(n912) );
  XOR U5293 ( .A(n913), .B(n912), .Z(n1767) );
  XNOR U5294 ( .A(x[83]), .B(y[83]), .Z(n3524) );
  XNOR U5295 ( .A(x[87]), .B(y[87]), .Z(n3522) );
  XOR U5296 ( .A(x[538]), .B(y[538]), .Z(n3521) );
  XNOR U5297 ( .A(n3522), .B(n3521), .Z(n3523) );
  XOR U5298 ( .A(n3524), .B(n3523), .Z(n1764) );
  XNOR U5299 ( .A(x[947]), .B(y[947]), .Z(n1881) );
  XNOR U5300 ( .A(x[62]), .B(y[62]), .Z(n1879) );
  XOR U5301 ( .A(x[949]), .B(y[949]), .Z(n1878) );
  XNOR U5302 ( .A(n1879), .B(n1878), .Z(n1880) );
  XNOR U5303 ( .A(n1881), .B(n1880), .Z(n1765) );
  XNOR U5304 ( .A(n1764), .B(n1765), .Z(n1766) );
  XNOR U5305 ( .A(n1767), .B(n1766), .Z(n4960) );
  XNOR U5306 ( .A(n4961), .B(n4960), .Z(n1184) );
  XNOR U5307 ( .A(x[203]), .B(y[203]), .Z(n2861) );
  XNOR U5308 ( .A(x[207]), .B(y[207]), .Z(n2859) );
  XOR U5309 ( .A(x[454]), .B(y[454]), .Z(n2858) );
  XNOR U5310 ( .A(n2859), .B(n2858), .Z(n2860) );
  XOR U5311 ( .A(n2861), .B(n2860), .Z(n3269) );
  XNOR U5312 ( .A(x[193]), .B(y[193]), .Z(n2853) );
  XNOR U5313 ( .A(x[197]), .B(y[197]), .Z(n2851) );
  XOR U5314 ( .A(x[199]), .B(y[199]), .Z(n2850) );
  XNOR U5315 ( .A(n2851), .B(n2850), .Z(n2852) );
  XOR U5316 ( .A(n2853), .B(n2852), .Z(n3266) );
  XNOR U5317 ( .A(x[1519]), .B(y[1519]), .Z(n1627) );
  XNOR U5318 ( .A(x[1521]), .B(y[1521]), .Z(n1624) );
  XNOR U5319 ( .A(x[1592]), .B(y[1592]), .Z(n1625) );
  XOR U5320 ( .A(n1624), .B(n1625), .Z(n1626) );
  XNOR U5321 ( .A(n1627), .B(n1626), .Z(n3267) );
  XNOR U5322 ( .A(n3266), .B(n3267), .Z(n3268) );
  XNOR U5323 ( .A(n3269), .B(n3268), .Z(n4953) );
  XNOR U5324 ( .A(x[177]), .B(y[177]), .Z(n1897) );
  XNOR U5325 ( .A(x[181]), .B(y[181]), .Z(n1895) );
  XOR U5326 ( .A(x[472]), .B(y[472]), .Z(n1894) );
  XNOR U5327 ( .A(n1895), .B(n1894), .Z(n1896) );
  XOR U5328 ( .A(n1897), .B(n1896), .Z(n2229) );
  XNOR U5329 ( .A(x[163]), .B(y[163]), .Z(n863) );
  XNOR U5330 ( .A(x[165]), .B(y[165]), .Z(n861) );
  XOR U5331 ( .A(x[169]), .B(y[169]), .Z(n860) );
  XNOR U5332 ( .A(n861), .B(n860), .Z(n862) );
  XOR U5333 ( .A(n863), .B(n862), .Z(n2226) );
  XNOR U5334 ( .A(x[963]), .B(y[963]), .Z(n4717) );
  XNOR U5335 ( .A(x[400]), .B(y[400]), .Z(n4715) );
  XOR U5336 ( .A(x[965]), .B(y[965]), .Z(n4714) );
  XNOR U5337 ( .A(n4715), .B(n4714), .Z(n4716) );
  XNOR U5338 ( .A(n4717), .B(n4716), .Z(n2227) );
  XNOR U5339 ( .A(n2226), .B(n2227), .Z(n2228) );
  XOR U5340 ( .A(n2229), .B(n2228), .Z(n4952) );
  XOR U5341 ( .A(n4953), .B(n4952), .Z(n4955) );
  XNOR U5342 ( .A(x[153]), .B(y[153]), .Z(n3937) );
  XNOR U5343 ( .A(x[155]), .B(y[155]), .Z(n3935) );
  XOR U5344 ( .A(x[159]), .B(y[159]), .Z(n3934) );
  XNOR U5345 ( .A(n3935), .B(n3934), .Z(n3936) );
  XOR U5346 ( .A(n3937), .B(n3936), .Z(n1479) );
  XNOR U5347 ( .A(x[147]), .B(y[147]), .Z(n3941) );
  XNOR U5348 ( .A(x[149]), .B(y[149]), .Z(n3939) );
  XOR U5349 ( .A(x[494]), .B(y[494]), .Z(n3938) );
  XNOR U5350 ( .A(n3939), .B(n3938), .Z(n3940) );
  XOR U5351 ( .A(n3941), .B(n3940), .Z(n1476) );
  XNOR U5352 ( .A(x[1523]), .B(y[1523]), .Z(n1623) );
  XNOR U5353 ( .A(x[343]), .B(y[343]), .Z(n1621) );
  XOR U5354 ( .A(x[1525]), .B(y[1525]), .Z(n1620) );
  XNOR U5355 ( .A(n1621), .B(n1620), .Z(n1622) );
  XNOR U5356 ( .A(n1623), .B(n1622), .Z(n1477) );
  XNOR U5357 ( .A(n1476), .B(n1477), .Z(n1478) );
  XNOR U5358 ( .A(n1479), .B(n1478), .Z(n4954) );
  XOR U5359 ( .A(n4955), .B(n4954), .Z(n1185) );
  XNOR U5360 ( .A(n1184), .B(n1185), .Z(n1186) );
  XNOR U5361 ( .A(n1187), .B(n1186), .Z(n2655) );
  XNOR U5362 ( .A(x[59]), .B(y[59]), .Z(n3816) );
  XNOR U5363 ( .A(x[61]), .B(y[61]), .Z(n3813) );
  XNOR U5364 ( .A(x[65]), .B(y[65]), .Z(n3814) );
  XOR U5365 ( .A(n3813), .B(n3814), .Z(n3815) );
  XOR U5366 ( .A(n3816), .B(n3815), .Z(n4747) );
  XNOR U5367 ( .A(x[53]), .B(y[53]), .Z(n3875) );
  XNOR U5368 ( .A(x[55]), .B(y[55]), .Z(n3873) );
  XOR U5369 ( .A(x[562]), .B(y[562]), .Z(n3872) );
  XNOR U5370 ( .A(n3873), .B(n3872), .Z(n3874) );
  XNOR U5371 ( .A(n3875), .B(n3874), .Z(n4744) );
  XNOR U5372 ( .A(x[939]), .B(y[939]), .Z(n4605) );
  XNOR U5373 ( .A(x[70]), .B(y[70]), .Z(n4602) );
  XNOR U5374 ( .A(x[941]), .B(y[941]), .Z(n4603) );
  XOR U5375 ( .A(n4602), .B(n4603), .Z(n4604) );
  XNOR U5376 ( .A(n4605), .B(n4604), .Z(n4745) );
  XNOR U5377 ( .A(n4747), .B(n4746), .Z(n4306) );
  XNOR U5378 ( .A(x[37]), .B(y[37]), .Z(n3057) );
  XNOR U5379 ( .A(x[39]), .B(y[39]), .Z(n3054) );
  XNOR U5380 ( .A(x[43]), .B(y[43]), .Z(n3055) );
  XOR U5381 ( .A(n3054), .B(n3055), .Z(n3056) );
  XOR U5382 ( .A(n3057), .B(n3056), .Z(n4514) );
  XNOR U5383 ( .A(x[21]), .B(y[21]), .Z(n3091) );
  XNOR U5384 ( .A(x[23]), .B(y[23]), .Z(n3088) );
  XNOR U5385 ( .A(x[584]), .B(y[584]), .Z(n3089) );
  XOR U5386 ( .A(n3088), .B(n3089), .Z(n3090) );
  XNOR U5387 ( .A(n3091), .B(n3090), .Z(n4512) );
  XNOR U5388 ( .A(x[1535]), .B(y[1535]), .Z(n2363) );
  XNOR U5389 ( .A(x[349]), .B(y[349]), .Z(n2360) );
  XNOR U5390 ( .A(x[1537]), .B(y[1537]), .Z(n2361) );
  XOR U5391 ( .A(n2360), .B(n2361), .Z(n2362) );
  XNOR U5392 ( .A(n2363), .B(n2362), .Z(n4513) );
  XOR U5393 ( .A(n4514), .B(n4515), .Z(n4307) );
  XOR U5394 ( .A(n4306), .B(n4307), .Z(n4308) );
  XNOR U5395 ( .A(x[77]), .B(y[77]), .Z(n3518) );
  XNOR U5396 ( .A(x[81]), .B(y[81]), .Z(n3515) );
  XNOR U5397 ( .A(x[544]), .B(y[544]), .Z(n3516) );
  XOR U5398 ( .A(n3515), .B(n3516), .Z(n3517) );
  XOR U5399 ( .A(n3518), .B(n3517), .Z(n1671) );
  XNOR U5400 ( .A(x[67]), .B(y[67]), .Z(n3822) );
  XNOR U5401 ( .A(x[71]), .B(y[71]), .Z(n3819) );
  XNOR U5402 ( .A(x[75]), .B(y[75]), .Z(n3820) );
  XOR U5403 ( .A(n3819), .B(n3820), .Z(n3821) );
  XNOR U5404 ( .A(n3822), .B(n3821), .Z(n1668) );
  XNOR U5405 ( .A(x[1531]), .B(y[1531]), .Z(n1607) );
  XNOR U5406 ( .A(x[46]), .B(y[46]), .Z(n1604) );
  XNOR U5407 ( .A(x[1533]), .B(y[1533]), .Z(n1605) );
  XOR U5408 ( .A(n1604), .B(n1605), .Z(n1606) );
  XNOR U5409 ( .A(n1607), .B(n1606), .Z(n1669) );
  XNOR U5410 ( .A(n1671), .B(n1670), .Z(n4309) );
  XOR U5411 ( .A(n4308), .B(n4309), .Z(n4319) );
  XNOR U5412 ( .A(x[15]), .B(y[15]), .Z(n3839) );
  XNOR U5413 ( .A(x[17]), .B(y[17]), .Z(n3837) );
  XOR U5414 ( .A(x[590]), .B(y[590]), .Z(n3835) );
  XNOR U5415 ( .A(n3837), .B(n3835), .Z(n3838) );
  XOR U5416 ( .A(n3839), .B(n3838), .Z(n1197) );
  XNOR U5417 ( .A(x[5]), .B(y[5]), .Z(n1969) );
  XNOR U5418 ( .A(x[9]), .B(y[9]), .Z(n1966) );
  XNOR U5419 ( .A(x[11]), .B(y[11]), .Z(n1967) );
  XOR U5420 ( .A(n1966), .B(n1967), .Z(n1968) );
  XOR U5421 ( .A(n1969), .B(n1968), .Z(n1194) );
  XNOR U5422 ( .A(x[931]), .B(y[931]), .Z(n4599) );
  XNOR U5423 ( .A(x[420]), .B(y[420]), .Z(n4596) );
  XNOR U5424 ( .A(x[933]), .B(y[933]), .Z(n4597) );
  XOR U5425 ( .A(n4596), .B(n4597), .Z(n4598) );
  XNOR U5426 ( .A(n4599), .B(n4598), .Z(n1195) );
  XNOR U5427 ( .A(n1194), .B(n1195), .Z(n1196) );
  XNOR U5428 ( .A(n1197), .B(n1196), .Z(n4947) );
  XNOR U5429 ( .A(x[4]), .B(y[4]), .Z(n1965) );
  XNOR U5430 ( .A(x[0]), .B(y[0]), .Z(n1963) );
  XOR U5431 ( .A(x[1]), .B(y[1]), .Z(n1962) );
  XNOR U5432 ( .A(n1963), .B(n1962), .Z(n1964) );
  XOR U5433 ( .A(n1965), .B(n1964), .Z(n1843) );
  XNOR U5434 ( .A(x[10]), .B(y[10]), .Z(n1985) );
  XNOR U5435 ( .A(x[6]), .B(y[6]), .Z(n1983) );
  XOR U5436 ( .A(x[608]), .B(y[608]), .Z(n1982) );
  XNOR U5437 ( .A(n1983), .B(n1982), .Z(n1984) );
  XOR U5438 ( .A(n1985), .B(n1984), .Z(n1840) );
  XNOR U5439 ( .A(x[1539]), .B(y[1539]), .Z(n2359) );
  XNOR U5440 ( .A(x[40]), .B(y[40]), .Z(n2357) );
  XOR U5441 ( .A(x[1541]), .B(y[1541]), .Z(n2356) );
  XNOR U5442 ( .A(n2357), .B(n2356), .Z(n2358) );
  XNOR U5443 ( .A(n2359), .B(n2358), .Z(n1841) );
  XNOR U5444 ( .A(n1840), .B(n1841), .Z(n1842) );
  XOR U5445 ( .A(n1843), .B(n1842), .Z(n4946) );
  XOR U5446 ( .A(n4947), .B(n4946), .Z(n4949) );
  XNOR U5447 ( .A(x[16]), .B(y[16]), .Z(n1981) );
  XNOR U5448 ( .A(x[12]), .B(y[12]), .Z(n1979) );
  XOR U5449 ( .A(x[612]), .B(y[612]), .Z(n1978) );
  XNOR U5450 ( .A(n1979), .B(n1978), .Z(n1980) );
  XOR U5451 ( .A(n1981), .B(n1980), .Z(n1277) );
  XNOR U5452 ( .A(x[38]), .B(y[38]), .Z(n2745) );
  XNOR U5453 ( .A(x[32]), .B(y[32]), .Z(n2743) );
  XOR U5454 ( .A(x[36]), .B(y[36]), .Z(n2742) );
  XNOR U5455 ( .A(n2743), .B(n2742), .Z(n2744) );
  XOR U5456 ( .A(n2745), .B(n2744), .Z(n1274) );
  XNOR U5457 ( .A(x[923]), .B(y[923]), .Z(n4895) );
  XNOR U5458 ( .A(x[426]), .B(y[426]), .Z(n4893) );
  XOR U5459 ( .A(x[925]), .B(y[925]), .Z(n4892) );
  XNOR U5460 ( .A(n4893), .B(n4892), .Z(n4894) );
  XNOR U5461 ( .A(n4895), .B(n4894), .Z(n1275) );
  XNOR U5462 ( .A(n1274), .B(n1275), .Z(n1276) );
  XNOR U5463 ( .A(n1277), .B(n1276), .Z(n4948) );
  XNOR U5464 ( .A(n4949), .B(n4948), .Z(n4316) );
  XNOR U5465 ( .A(x[58]), .B(y[58]), .Z(n2717) );
  XNOR U5466 ( .A(x[56]), .B(y[56]), .Z(n2715) );
  XOR U5467 ( .A(x[634]), .B(y[634]), .Z(n2714) );
  XNOR U5468 ( .A(n2715), .B(n2714), .Z(n2716) );
  XOR U5469 ( .A(n2717), .B(n2716), .Z(n1563) );
  XNOR U5470 ( .A(x[72]), .B(y[72]), .Z(n3778) );
  XNOR U5471 ( .A(x[64]), .B(y[64]), .Z(n3776) );
  XOR U5472 ( .A(x[68]), .B(y[68]), .Z(n3775) );
  XNOR U5473 ( .A(n3776), .B(n3775), .Z(n3777) );
  XOR U5474 ( .A(n3778), .B(n3777), .Z(n1560) );
  XNOR U5475 ( .A(x[1543]), .B(y[1543]), .Z(n2463) );
  XNOR U5476 ( .A(x[355]), .B(y[355]), .Z(n2460) );
  XNOR U5477 ( .A(x[1545]), .B(y[1545]), .Z(n2461) );
  XOR U5478 ( .A(n2460), .B(n2461), .Z(n2462) );
  XNOR U5479 ( .A(n2463), .B(n2462), .Z(n1561) );
  XNOR U5480 ( .A(n1560), .B(n1561), .Z(n1562) );
  XNOR U5481 ( .A(n1563), .B(n1562), .Z(n4401) );
  XNOR U5482 ( .A(x[92]), .B(y[92]), .Z(n3774) );
  XNOR U5483 ( .A(x[78]), .B(y[78]), .Z(n3772) );
  XOR U5484 ( .A(x[88]), .B(y[88]), .Z(n3771) );
  XNOR U5485 ( .A(n3772), .B(n3771), .Z(n3773) );
  XOR U5486 ( .A(n3774), .B(n3773), .Z(n1551) );
  XNOR U5487 ( .A(x[98]), .B(y[98]), .Z(n3696) );
  XNOR U5488 ( .A(x[94]), .B(y[94]), .Z(n3694) );
  XOR U5489 ( .A(x[652]), .B(y[652]), .Z(n3693) );
  XNOR U5490 ( .A(n3694), .B(n3693), .Z(n3695) );
  XOR U5491 ( .A(n3696), .B(n3695), .Z(n1548) );
  XNOR U5492 ( .A(x[915]), .B(y[915]), .Z(n4899) );
  XNOR U5493 ( .A(x[90]), .B(y[90]), .Z(n4896) );
  XNOR U5494 ( .A(x[917]), .B(y[917]), .Z(n4897) );
  XOR U5495 ( .A(n4896), .B(n4897), .Z(n4898) );
  XNOR U5496 ( .A(n4899), .B(n4898), .Z(n1549) );
  XNOR U5497 ( .A(n1548), .B(n1549), .Z(n1550) );
  XOR U5498 ( .A(n1551), .B(n1550), .Z(n4400) );
  XOR U5499 ( .A(n4401), .B(n4400), .Z(n4403) );
  XNOR U5500 ( .A(x[108]), .B(y[108]), .Z(n3692) );
  XNOR U5501 ( .A(x[104]), .B(y[104]), .Z(n3690) );
  XOR U5502 ( .A(x[656]), .B(y[656]), .Z(n3689) );
  XNOR U5503 ( .A(n3690), .B(n3689), .Z(n3691) );
  XOR U5504 ( .A(n3692), .B(n3691), .Z(n1301) );
  XNOR U5505 ( .A(x[128]), .B(y[128]), .Z(n3718) );
  XNOR U5506 ( .A(x[114]), .B(y[114]), .Z(n3716) );
  XOR U5507 ( .A(x[122]), .B(y[122]), .Z(n3715) );
  XNOR U5508 ( .A(n3716), .B(n3715), .Z(n3717) );
  XOR U5509 ( .A(n3718), .B(n3717), .Z(n1298) );
  XNOR U5510 ( .A(x[1547]), .B(y[1547]), .Z(n2419) );
  XNOR U5511 ( .A(x[359]), .B(y[359]), .Z(n2417) );
  XOR U5512 ( .A(x[1549]), .B(y[1549]), .Z(n2416) );
  XNOR U5513 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U5514 ( .A(n2419), .B(n2418), .Z(n1299) );
  XNOR U5515 ( .A(n1298), .B(n1299), .Z(n1300) );
  XNOR U5516 ( .A(n1301), .B(n1300), .Z(n4402) );
  XOR U5517 ( .A(n4403), .B(n4402), .Z(n4317) );
  XNOR U5518 ( .A(n4316), .B(n4317), .Z(n4318) );
  XOR U5519 ( .A(n4319), .B(n4318), .Z(n2654) );
  XOR U5520 ( .A(n2655), .B(n2654), .Z(n2657) );
  XNOR U5521 ( .A(n2656), .B(n2657), .Z(n1175) );
  XNOR U5522 ( .A(x[974]), .B(y[974]), .Z(n2693) );
  XNOR U5523 ( .A(x[970]), .B(y[970]), .Z(n2690) );
  XNOR U5524 ( .A(x[972]), .B(y[972]), .Z(n2691) );
  XOR U5525 ( .A(n2690), .B(n2691), .Z(n2692) );
  XOR U5526 ( .A(n2693), .B(n2692), .Z(n4185) );
  XNOR U5527 ( .A(x[986]), .B(y[986]), .Z(n2687) );
  XNOR U5528 ( .A(x[982]), .B(y[982]), .Z(n2684) );
  XNOR U5529 ( .A(x[984]), .B(y[984]), .Z(n2685) );
  XOR U5530 ( .A(n2684), .B(n2685), .Z(n2686) );
  XOR U5531 ( .A(n2687), .B(n2686), .Z(n4182) );
  XNOR U5532 ( .A(x[980]), .B(y[980]), .Z(n2681) );
  XNOR U5533 ( .A(x[976]), .B(y[976]), .Z(n2678) );
  XNOR U5534 ( .A(x[978]), .B(y[978]), .Z(n2679) );
  XOR U5535 ( .A(n2678), .B(n2679), .Z(n2680) );
  XNOR U5536 ( .A(n2681), .B(n2680), .Z(n4183) );
  XNOR U5537 ( .A(n4182), .B(n4183), .Z(n4184) );
  XNOR U5538 ( .A(n4185), .B(n4184), .Z(n4087) );
  XNOR U5539 ( .A(x[1266]), .B(y[1266]), .Z(n1665) );
  XNOR U5540 ( .A(x[1306]), .B(y[1306]), .Z(n1662) );
  XNOR U5541 ( .A(x[1392]), .B(y[1392]), .Z(n1663) );
  XOR U5542 ( .A(n1662), .B(n1663), .Z(n1664) );
  XOR U5543 ( .A(n1665), .B(n1664), .Z(n979) );
  XNOR U5544 ( .A(x[1272]), .B(y[1272]), .Z(n1659) );
  XNOR U5545 ( .A(x[1270]), .B(y[1270]), .Z(n1656) );
  XNOR U5546 ( .A(x[1302]), .B(y[1302]), .Z(n1657) );
  XOR U5547 ( .A(n1656), .B(n1657), .Z(n1658) );
  XNOR U5548 ( .A(n1659), .B(n1658), .Z(n976) );
  XNOR U5549 ( .A(x[1268]), .B(y[1268]), .Z(n1653) );
  XNOR U5550 ( .A(x[1304]), .B(y[1304]), .Z(n1650) );
  XNOR U5551 ( .A(x[1388]), .B(y[1388]), .Z(n1651) );
  XOR U5552 ( .A(n1650), .B(n1651), .Z(n1652) );
  XNOR U5553 ( .A(n1653), .B(n1652), .Z(n977) );
  XNOR U5554 ( .A(n979), .B(n978), .Z(n4084) );
  XNOR U5555 ( .A(x[956]), .B(y[956]), .Z(n1131) );
  XNOR U5556 ( .A(x[952]), .B(y[952]), .Z(n1128) );
  XNOR U5557 ( .A(x[954]), .B(y[954]), .Z(n1129) );
  XOR U5558 ( .A(n1128), .B(n1129), .Z(n1130) );
  XOR U5559 ( .A(n1131), .B(n1130), .Z(n4154) );
  XNOR U5560 ( .A(x[968]), .B(y[968]), .Z(n1125) );
  XNOR U5561 ( .A(x[964]), .B(y[964]), .Z(n1122) );
  XNOR U5562 ( .A(x[966]), .B(y[966]), .Z(n1123) );
  XOR U5563 ( .A(n1122), .B(n1123), .Z(n1124) );
  XNOR U5564 ( .A(n1125), .B(n1124), .Z(n4152) );
  XNOR U5565 ( .A(x[962]), .B(y[962]), .Z(n1119) );
  XNOR U5566 ( .A(x[958]), .B(y[958]), .Z(n1116) );
  XNOR U5567 ( .A(x[960]), .B(y[960]), .Z(n1117) );
  XOR U5568 ( .A(n1116), .B(n1117), .Z(n1118) );
  XNOR U5569 ( .A(n1119), .B(n1118), .Z(n4153) );
  XOR U5570 ( .A(n4154), .B(n4155), .Z(n4085) );
  XOR U5571 ( .A(n4084), .B(n4085), .Z(n4086) );
  XOR U5572 ( .A(n4087), .B(n4086), .Z(n4837) );
  XNOR U5573 ( .A(x[1120]), .B(y[1120]), .Z(n3239) );
  XNOR U5574 ( .A(x[1112]), .B(y[1112]), .Z(n3236) );
  XNOR U5575 ( .A(x[1116]), .B(y[1116]), .Z(n3237) );
  XOR U5576 ( .A(n3236), .B(n3237), .Z(n3238) );
  XOR U5577 ( .A(n3239), .B(n3238), .Z(n1557) );
  XNOR U5578 ( .A(x[1144]), .B(y[1144]), .Z(n3233) );
  XNOR U5579 ( .A(x[1136]), .B(y[1136]), .Z(n3230) );
  XNOR U5580 ( .A(x[1140]), .B(y[1140]), .Z(n3231) );
  XOR U5581 ( .A(n3230), .B(n3231), .Z(n3232) );
  XNOR U5582 ( .A(n3233), .B(n3232), .Z(n1554) );
  XNOR U5583 ( .A(x[1132]), .B(y[1132]), .Z(n3227) );
  XNOR U5584 ( .A(x[1124]), .B(y[1124]), .Z(n3224) );
  XNOR U5585 ( .A(x[1128]), .B(y[1128]), .Z(n3225) );
  XOR U5586 ( .A(n3224), .B(n3225), .Z(n3226) );
  XNOR U5587 ( .A(n3227), .B(n3226), .Z(n1555) );
  XNOR U5588 ( .A(n1557), .B(n1556), .Z(n4267) );
  XNOR U5589 ( .A(x[1180]), .B(y[1180]), .Z(n3207) );
  XNOR U5590 ( .A(x[1172]), .B(y[1172]), .Z(n3204) );
  XNOR U5591 ( .A(x[1176]), .B(y[1176]), .Z(n3205) );
  XOR U5592 ( .A(n3204), .B(n3205), .Z(n3206) );
  XOR U5593 ( .A(n3207), .B(n3206), .Z(n4425) );
  XNOR U5594 ( .A(x[1192]), .B(y[1192]), .Z(n3201) );
  XNOR U5595 ( .A(x[1184]), .B(y[1184]), .Z(n3198) );
  XNOR U5596 ( .A(x[1188]), .B(y[1188]), .Z(n3199) );
  XOR U5597 ( .A(n3198), .B(n3199), .Z(n3200) );
  XNOR U5598 ( .A(n3201), .B(n3200), .Z(n4422) );
  XNOR U5599 ( .A(x[276]), .B(y[276]), .Z(n2451) );
  XNOR U5600 ( .A(x[270]), .B(y[270]), .Z(n2448) );
  XNOR U5601 ( .A(x[272]), .B(y[272]), .Z(n2449) );
  XOR U5602 ( .A(n2448), .B(n2449), .Z(n2450) );
  XNOR U5603 ( .A(n2451), .B(n2450), .Z(n4423) );
  XNOR U5604 ( .A(n4425), .B(n4424), .Z(n4264) );
  XNOR U5605 ( .A(x[1084]), .B(y[1084]), .Z(n3147) );
  XNOR U5606 ( .A(x[1076]), .B(y[1076]), .Z(n3145) );
  XOR U5607 ( .A(x[1080]), .B(y[1080]), .Z(n3144) );
  XNOR U5608 ( .A(n3145), .B(n3144), .Z(n3146) );
  XOR U5609 ( .A(n3147), .B(n3146), .Z(n4520) );
  XNOR U5610 ( .A(x[1096]), .B(y[1096]), .Z(n3143) );
  XNOR U5611 ( .A(x[1088]), .B(y[1088]), .Z(n3141) );
  XOR U5612 ( .A(x[1092]), .B(y[1092]), .Z(n3140) );
  XNOR U5613 ( .A(n3141), .B(n3140), .Z(n3142) );
  XNOR U5614 ( .A(n3143), .B(n3142), .Z(n4518) );
  XNOR U5615 ( .A(x[1108]), .B(y[1108]), .Z(n3151) );
  XNOR U5616 ( .A(x[1100]), .B(y[1100]), .Z(n3149) );
  XOR U5617 ( .A(x[1104]), .B(y[1104]), .Z(n3148) );
  XNOR U5618 ( .A(n3149), .B(n3148), .Z(n3150) );
  XNOR U5619 ( .A(n3151), .B(n3150), .Z(n4519) );
  XOR U5620 ( .A(n4520), .B(n4521), .Z(n4265) );
  XOR U5621 ( .A(n4264), .B(n4265), .Z(n4266) );
  XOR U5622 ( .A(n4267), .B(n4266), .Z(n4834) );
  XNOR U5623 ( .A(x[1004]), .B(y[1004]), .Z(n2727) );
  XNOR U5624 ( .A(x[1000]), .B(y[1000]), .Z(n2724) );
  XNOR U5625 ( .A(x[1002]), .B(y[1002]), .Z(n2725) );
  XOR U5626 ( .A(n2724), .B(n2725), .Z(n2726) );
  XOR U5627 ( .A(n2727), .B(n2726), .Z(n4251) );
  XNOR U5628 ( .A(x[1010]), .B(y[1010]), .Z(n2721) );
  XNOR U5629 ( .A(x[1006]), .B(y[1006]), .Z(n2718) );
  XNOR U5630 ( .A(x[1008]), .B(y[1008]), .Z(n2719) );
  XOR U5631 ( .A(n2718), .B(n2719), .Z(n2720) );
  XOR U5632 ( .A(n2721), .B(n2720), .Z(n4248) );
  XNOR U5633 ( .A(x[52]), .B(y[52]), .Z(n2039) );
  XNOR U5634 ( .A(x[44]), .B(y[44]), .Z(n2036) );
  XNOR U5635 ( .A(x[630]), .B(y[630]), .Z(n2037) );
  XOR U5636 ( .A(n2036), .B(n2037), .Z(n2038) );
  XNOR U5637 ( .A(n2039), .B(n2038), .Z(n4249) );
  XNOR U5638 ( .A(n4248), .B(n4249), .Z(n4250) );
  XNOR U5639 ( .A(n4251), .B(n4250), .Z(n3993) );
  XNOR U5640 ( .A(x[1396]), .B(y[1396]), .Z(n1773) );
  XNOR U5641 ( .A(x[1260]), .B(y[1260]), .Z(n1771) );
  XOR U5642 ( .A(x[1394]), .B(y[1394]), .Z(n1770) );
  XNOR U5643 ( .A(n1771), .B(n1770), .Z(n1772) );
  XOR U5644 ( .A(n1773), .B(n1772), .Z(n2531) );
  XNOR U5645 ( .A(x[1264]), .B(y[1264]), .Z(n1777) );
  XNOR U5646 ( .A(x[1262]), .B(y[1262]), .Z(n1775) );
  XOR U5647 ( .A(x[1390]), .B(y[1390]), .Z(n1774) );
  XNOR U5648 ( .A(n1775), .B(n1774), .Z(n1776) );
  XNOR U5649 ( .A(n1777), .B(n1776), .Z(n2530) );
  XOR U5650 ( .A(n2531), .B(n2530), .Z(n2533) );
  XNOR U5651 ( .A(x[1400]), .B(y[1400]), .Z(n1781) );
  XNOR U5652 ( .A(x[1258]), .B(y[1258]), .Z(n1779) );
  XOR U5653 ( .A(x[1398]), .B(y[1398]), .Z(n1778) );
  XNOR U5654 ( .A(n1779), .B(n1778), .Z(n1780) );
  XNOR U5655 ( .A(n1781), .B(n1780), .Z(n2532) );
  XNOR U5656 ( .A(x[992]), .B(y[992]), .Z(n2755) );
  XNOR U5657 ( .A(x[988]), .B(y[988]), .Z(n2752) );
  XNOR U5658 ( .A(x[990]), .B(y[990]), .Z(n2753) );
  XOR U5659 ( .A(n2752), .B(n2753), .Z(n2754) );
  XOR U5660 ( .A(n2755), .B(n2754), .Z(n4239) );
  XNOR U5661 ( .A(x[998]), .B(y[998]), .Z(n2749) );
  XNOR U5662 ( .A(x[994]), .B(y[994]), .Z(n2746) );
  XNOR U5663 ( .A(x[996]), .B(y[996]), .Z(n2747) );
  XOR U5664 ( .A(n2746), .B(n2747), .Z(n2748) );
  XOR U5665 ( .A(n2749), .B(n2748), .Z(n4236) );
  XNOR U5666 ( .A(x[30]), .B(y[30]), .Z(n2033) );
  XNOR U5667 ( .A(x[22]), .B(y[22]), .Z(n2030) );
  XNOR U5668 ( .A(x[24]), .B(y[24]), .Z(n2031) );
  XOR U5669 ( .A(n2030), .B(n2031), .Z(n2032) );
  XNOR U5670 ( .A(n2033), .B(n2032), .Z(n4237) );
  XNOR U5671 ( .A(n4236), .B(n4237), .Z(n4238) );
  XNOR U5672 ( .A(n4239), .B(n4238), .Z(n3991) );
  XOR U5673 ( .A(n3990), .B(n3991), .Z(n3992) );
  XNOR U5674 ( .A(n3993), .B(n3992), .Z(n4835) );
  XNOR U5675 ( .A(n4834), .B(n4835), .Z(n4836) );
  XNOR U5676 ( .A(n4837), .B(n4836), .Z(n1172) );
  XNOR U5677 ( .A(x[448]), .B(y[448]), .Z(n2145) );
  XNOR U5678 ( .A(x[444]), .B(y[444]), .Z(n2142) );
  XNOR U5679 ( .A(x[786]), .B(y[786]), .Z(n2143) );
  XOR U5680 ( .A(n2142), .B(n2143), .Z(n2144) );
  XOR U5681 ( .A(n2145), .B(n2144), .Z(n2055) );
  XNOR U5682 ( .A(x[468]), .B(y[468]), .Z(n4753) );
  XNOR U5683 ( .A(x[462]), .B(y[462]), .Z(n4750) );
  XNOR U5684 ( .A(x[464]), .B(y[464]), .Z(n4751) );
  XOR U5685 ( .A(n4750), .B(n4751), .Z(n4752) );
  XNOR U5686 ( .A(n4753), .B(n4752), .Z(n2052) );
  XNOR U5687 ( .A(x[867]), .B(y[867]), .Z(n4821) );
  XNOR U5688 ( .A(x[460]), .B(y[460]), .Z(n4818) );
  XNOR U5689 ( .A(x[869]), .B(y[869]), .Z(n4819) );
  XOR U5690 ( .A(n4818), .B(n4819), .Z(n4820) );
  XNOR U5691 ( .A(n4821), .B(n4820), .Z(n2053) );
  XNOR U5692 ( .A(n2055), .B(n2054), .Z(n4170) );
  XNOR U5693 ( .A(x[482]), .B(y[482]), .Z(n4551) );
  XNOR U5694 ( .A(x[478]), .B(y[478]), .Z(n4548) );
  XNOR U5695 ( .A(x[804]), .B(y[804]), .Z(n4549) );
  XOR U5696 ( .A(n4548), .B(n4549), .Z(n4550) );
  XOR U5697 ( .A(n4551), .B(n4550), .Z(n2096) );
  XNOR U5698 ( .A(x[490]), .B(y[490]), .Z(n4119) );
  XNOR U5699 ( .A(x[484]), .B(y[484]), .Z(n4116) );
  XNOR U5700 ( .A(x[488]), .B(y[488]), .Z(n4117) );
  XOR U5701 ( .A(n4116), .B(n4117), .Z(n4118) );
  XNOR U5702 ( .A(n4119), .B(n4118), .Z(n2094) );
  XNOR U5703 ( .A(x[1571]), .B(y[1571]), .Z(n3538) );
  XNOR U5704 ( .A(x[20]), .B(y[20]), .Z(n3535) );
  XNOR U5705 ( .A(x[1573]), .B(y[1573]), .Z(n3536) );
  XOR U5706 ( .A(n3535), .B(n3536), .Z(n3537) );
  XNOR U5707 ( .A(n3538), .B(n3537), .Z(n2095) );
  XOR U5708 ( .A(n2096), .B(n2097), .Z(n4171) );
  XOR U5709 ( .A(n4170), .B(n4171), .Z(n4172) );
  XNOR U5710 ( .A(x[436]), .B(y[436]), .Z(n2187) );
  XNOR U5711 ( .A(x[430]), .B(y[430]), .Z(n2184) );
  XNOR U5712 ( .A(x[434]), .B(y[434]), .Z(n2185) );
  XOR U5713 ( .A(n2184), .B(n2185), .Z(n2186) );
  XOR U5714 ( .A(n2187), .B(n2186), .Z(n1473) );
  XNOR U5715 ( .A(x[1567]), .B(y[1567]), .Z(n3738) );
  XNOR U5716 ( .A(x[371]), .B(y[371]), .Z(n3735) );
  XNOR U5717 ( .A(x[1569]), .B(y[1569]), .Z(n3736) );
  XOR U5718 ( .A(n3735), .B(n3736), .Z(n3737) );
  XNOR U5719 ( .A(n3738), .B(n3737), .Z(n1470) );
  XNOR U5720 ( .A(x[442]), .B(y[442]), .Z(n2139) );
  XNOR U5721 ( .A(x[438]), .B(y[438]), .Z(n2136) );
  XNOR U5722 ( .A(x[782]), .B(y[782]), .Z(n2137) );
  XOR U5723 ( .A(n2136), .B(n2137), .Z(n2138) );
  XNOR U5724 ( .A(n2139), .B(n2138), .Z(n1471) );
  XNOR U5725 ( .A(n1473), .B(n1472), .Z(n4173) );
  XOR U5726 ( .A(n4172), .B(n4173), .Z(n1261) );
  XNOR U5727 ( .A(x[536]), .B(y[536]), .Z(n4643) );
  XNOR U5728 ( .A(x[534]), .B(y[534]), .Z(n4641) );
  XNOR U5729 ( .A(x[836]), .B(y[836]), .Z(n4640) );
  XNOR U5730 ( .A(n4641), .B(n4640), .Z(n4642) );
  XNOR U5731 ( .A(n4643), .B(n4642), .Z(n2090) );
  XNOR U5732 ( .A(x[554]), .B(y[554]), .Z(n1283) );
  XNOR U5733 ( .A(x[550]), .B(y[550]), .Z(n1281) );
  XNOR U5734 ( .A(x[552]), .B(y[552]), .Z(n1280) );
  XNOR U5735 ( .A(n1281), .B(n1280), .Z(n1282) );
  XNOR U5736 ( .A(n1283), .B(n1282), .Z(n2088) );
  XNOR U5737 ( .A(x[851]), .B(y[851]), .Z(n4801) );
  XNOR U5738 ( .A(x[144]), .B(y[144]), .Z(n4798) );
  XNOR U5739 ( .A(x[853]), .B(y[853]), .Z(n4799) );
  XOR U5740 ( .A(n4798), .B(n4799), .Z(n4800) );
  XNOR U5741 ( .A(n4801), .B(n4800), .Z(n2089) );
  XOR U5742 ( .A(n2088), .B(n2089), .Z(n2091) );
  XNOR U5743 ( .A(n2090), .B(n2091), .Z(n4178) );
  XNOR U5744 ( .A(x[502]), .B(y[502]), .Z(n4113) );
  XNOR U5745 ( .A(x[492]), .B(y[492]), .Z(n4110) );
  XNOR U5746 ( .A(x[496]), .B(y[496]), .Z(n4111) );
  XOR U5747 ( .A(n4110), .B(n4111), .Z(n4112) );
  XOR U5748 ( .A(n4113), .B(n4112), .Z(n3324) );
  XNOR U5749 ( .A(x[508]), .B(y[508]), .Z(n2127) );
  XNOR U5750 ( .A(x[504]), .B(y[504]), .Z(n2124) );
  XNOR U5751 ( .A(x[818]), .B(y[818]), .Z(n2125) );
  XOR U5752 ( .A(n2124), .B(n2125), .Z(n2126) );
  XNOR U5753 ( .A(n2127), .B(n2126), .Z(n3321) );
  XNOR U5754 ( .A(x[859]), .B(y[859]), .Z(n4811) );
  XNOR U5755 ( .A(x[466]), .B(y[466]), .Z(n4808) );
  XNOR U5756 ( .A(x[861]), .B(y[861]), .Z(n4809) );
  XOR U5757 ( .A(n4808), .B(n4809), .Z(n4810) );
  XNOR U5758 ( .A(n4811), .B(n4810), .Z(n3322) );
  XNOR U5759 ( .A(n3324), .B(n3323), .Z(n4176) );
  XNOR U5760 ( .A(x[512]), .B(y[512]), .Z(n2121) );
  XNOR U5761 ( .A(x[510]), .B(y[510]), .Z(n2118) );
  XNOR U5762 ( .A(x[822]), .B(y[822]), .Z(n2119) );
  XOR U5763 ( .A(n2118), .B(n2119), .Z(n2120) );
  XOR U5764 ( .A(n2121), .B(n2120), .Z(n2102) );
  XNOR U5765 ( .A(x[524]), .B(y[524]), .Z(n4231) );
  XNOR U5766 ( .A(x[514]), .B(y[514]), .Z(n4229) );
  XOR U5767 ( .A(x[518]), .B(y[518]), .Z(n4228) );
  XNOR U5768 ( .A(n4229), .B(n4228), .Z(n4230) );
  XNOR U5769 ( .A(n4231), .B(n4230), .Z(n2100) );
  XNOR U5770 ( .A(x[1575]), .B(y[1575]), .Z(n3566) );
  XNOR U5771 ( .A(x[377]), .B(y[377]), .Z(n3563) );
  XNOR U5772 ( .A(x[1577]), .B(y[1577]), .Z(n3564) );
  XOR U5773 ( .A(n3563), .B(n3564), .Z(n3565) );
  XNOR U5774 ( .A(n3566), .B(n3565), .Z(n2101) );
  XOR U5775 ( .A(n2102), .B(n2103), .Z(n4177) );
  XOR U5776 ( .A(n4176), .B(n4177), .Z(n4179) );
  XNOR U5777 ( .A(n4178), .B(n4179), .Z(n1258) );
  XNOR U5778 ( .A(x[610]), .B(y[610]), .Z(n4009) );
  XNOR U5779 ( .A(x[604]), .B(y[604]), .Z(n4007) );
  XOR U5780 ( .A(x[1070]), .B(y[1070]), .Z(n4006) );
  XNOR U5781 ( .A(n4007), .B(n4006), .Z(n4008) );
  XOR U5782 ( .A(n4009), .B(n4008), .Z(n2079) );
  XNOR U5783 ( .A(x[616]), .B(y[616]), .Z(n4005) );
  XNOR U5784 ( .A(x[614]), .B(y[614]), .Z(n4003) );
  XOR U5785 ( .A(x[1466]), .B(y[1466]), .Z(n4002) );
  XNOR U5786 ( .A(n4003), .B(n4002), .Z(n4004) );
  XNOR U5787 ( .A(n4005), .B(n4004), .Z(n2076) );
  XNOR U5788 ( .A(x[1583]), .B(y[1583]), .Z(n3388) );
  XNOR U5789 ( .A(x[789]), .B(y[789]), .Z(n3386) );
  XOR U5790 ( .A(x[1585]), .B(y[1585]), .Z(n3385) );
  XNOR U5791 ( .A(n3386), .B(n3385), .Z(n3387) );
  XNOR U5792 ( .A(n3388), .B(n3387), .Z(n2077) );
  XNOR U5793 ( .A(n2079), .B(n2078), .Z(n4103) );
  XNOR U5794 ( .A(x[564]), .B(y[564]), .Z(n4215) );
  XNOR U5795 ( .A(x[556]), .B(y[556]), .Z(n4213) );
  XOR U5796 ( .A(x[558]), .B(y[558]), .Z(n4212) );
  XNOR U5797 ( .A(n4213), .B(n4212), .Z(n4214) );
  XOR U5798 ( .A(n4215), .B(n4214), .Z(n2073) );
  XNOR U5799 ( .A(x[588]), .B(y[588]), .Z(n2169) );
  XNOR U5800 ( .A(x[578]), .B(y[578]), .Z(n2167) );
  XOR U5801 ( .A(x[582]), .B(y[582]), .Z(n2166) );
  XNOR U5802 ( .A(n2167), .B(n2166), .Z(n2168) );
  XNOR U5803 ( .A(n2169), .B(n2168), .Z(n2070) );
  XNOR U5804 ( .A(x[1579]), .B(y[1579]), .Z(n3462) );
  XNOR U5805 ( .A(x[381]), .B(y[381]), .Z(n3460) );
  XOR U5806 ( .A(x[1581]), .B(y[1581]), .Z(n3459) );
  XNOR U5807 ( .A(n3460), .B(n3459), .Z(n3461) );
  XNOR U5808 ( .A(n3462), .B(n3461), .Z(n2071) );
  XNOR U5809 ( .A(n2073), .B(n2072), .Z(n4100) );
  XNOR U5810 ( .A(x[596]), .B(y[596]), .Z(n4019) );
  XNOR U5811 ( .A(x[592]), .B(y[592]), .Z(n4017) );
  XOR U5812 ( .A(x[594]), .B(y[594]), .Z(n4016) );
  XNOR U5813 ( .A(n4017), .B(n4016), .Z(n4018) );
  XOR U5814 ( .A(n4019), .B(n4018), .Z(n2066) );
  XNOR U5815 ( .A(x[843]), .B(y[843]), .Z(n4807) );
  XNOR U5816 ( .A(x[152]), .B(y[152]), .Z(n4805) );
  XOR U5817 ( .A(x[845]), .B(y[845]), .Z(n4804) );
  XNOR U5818 ( .A(n4805), .B(n4804), .Z(n4806) );
  XNOR U5819 ( .A(n4807), .B(n4806), .Z(n2064) );
  XNOR U5820 ( .A(x[602]), .B(y[602]), .Z(n4023) );
  XNOR U5821 ( .A(x[598]), .B(y[598]), .Z(n4021) );
  XOR U5822 ( .A(x[872]), .B(y[872]), .Z(n4020) );
  XNOR U5823 ( .A(n4021), .B(n4020), .Z(n4022) );
  XNOR U5824 ( .A(n4023), .B(n4022), .Z(n2065) );
  XOR U5825 ( .A(n2066), .B(n2067), .Z(n4101) );
  XOR U5826 ( .A(n4100), .B(n4101), .Z(n4102) );
  XNOR U5827 ( .A(n4103), .B(n4102), .Z(n1259) );
  XNOR U5828 ( .A(n1258), .B(n1259), .Z(n1260) );
  XNOR U5829 ( .A(n1261), .B(n1260), .Z(n1357) );
  XNOR U5830 ( .A(x[622]), .B(y[622]), .Z(n1397) );
  XNOR U5831 ( .A(x[618]), .B(y[618]), .Z(n1395) );
  XOR U5832 ( .A(x[1074]), .B(y[1074]), .Z(n1394) );
  XNOR U5833 ( .A(n1395), .B(n1394), .Z(n1396) );
  XOR U5834 ( .A(n1397), .B(n1396), .Z(n1065) );
  XNOR U5835 ( .A(x[628]), .B(y[628]), .Z(n1401) );
  XNOR U5836 ( .A(x[624]), .B(y[624]), .Z(n1399) );
  XOR U5837 ( .A(x[1464]), .B(y[1464]), .Z(n1398) );
  XNOR U5838 ( .A(n1399), .B(n1398), .Z(n1400) );
  XOR U5839 ( .A(n1401), .B(n1400), .Z(n1062) );
  XNOR U5840 ( .A(x[835]), .B(y[835]), .Z(n4441) );
  XNOR U5841 ( .A(x[480]), .B(y[480]), .Z(n4439) );
  XOR U5842 ( .A(x[837]), .B(y[837]), .Z(n4438) );
  XNOR U5843 ( .A(n4439), .B(n4438), .Z(n4440) );
  XNOR U5844 ( .A(n4441), .B(n4440), .Z(n1063) );
  XNOR U5845 ( .A(n1062), .B(n1063), .Z(n1064) );
  XNOR U5846 ( .A(n1065), .B(n1064), .Z(n2203) );
  XNOR U5847 ( .A(x[636]), .B(y[636]), .Z(n1387) );
  XNOR U5848 ( .A(x[632]), .B(y[632]), .Z(n1385) );
  XOR U5849 ( .A(x[1078]), .B(y[1078]), .Z(n1384) );
  XNOR U5850 ( .A(n1385), .B(n1384), .Z(n1386) );
  XOR U5851 ( .A(n1387), .B(n1386), .Z(n2223) );
  XNOR U5852 ( .A(x[642]), .B(y[642]), .Z(n1383) );
  XNOR U5853 ( .A(x[638]), .B(y[638]), .Z(n1381) );
  XOR U5854 ( .A(x[1462]), .B(y[1462]), .Z(n1380) );
  XNOR U5855 ( .A(n1381), .B(n1380), .Z(n1382) );
  XOR U5856 ( .A(n1383), .B(n1382), .Z(n2220) );
  XNOR U5857 ( .A(x[1587]), .B(y[1587]), .Z(n3336) );
  XNOR U5858 ( .A(x[1589]), .B(y[1589]), .Z(n3334) );
  XOR U5859 ( .A(x[1591]), .B(y[1591]), .Z(n3333) );
  XNOR U5860 ( .A(n3334), .B(n3333), .Z(n3335) );
  XNOR U5861 ( .A(n3336), .B(n3335), .Z(n2221) );
  XNOR U5862 ( .A(n2220), .B(n2221), .Z(n2222) );
  XOR U5863 ( .A(n2223), .B(n2222), .Z(n2202) );
  XOR U5864 ( .A(n2203), .B(n2202), .Z(n2205) );
  XNOR U5865 ( .A(x[648]), .B(y[648]), .Z(n3660) );
  XNOR U5866 ( .A(x[644]), .B(y[644]), .Z(n3658) );
  XOR U5867 ( .A(x[1082]), .B(y[1082]), .Z(n3657) );
  XNOR U5868 ( .A(n3658), .B(n3657), .Z(n3659) );
  XOR U5869 ( .A(n3660), .B(n3659), .Z(n1921) );
  XNOR U5870 ( .A(x[654]), .B(y[654]), .Z(n3656) );
  XNOR U5871 ( .A(x[650]), .B(y[650]), .Z(n3654) );
  XOR U5872 ( .A(x[1460]), .B(y[1460]), .Z(n3653) );
  XNOR U5873 ( .A(n3654), .B(n3653), .Z(n3655) );
  XOR U5874 ( .A(n3656), .B(n3655), .Z(n1918) );
  XNOR U5875 ( .A(x[827]), .B(y[827]), .Z(n4445) );
  XNOR U5876 ( .A(x[486]), .B(y[486]), .Z(n4443) );
  XOR U5877 ( .A(x[829]), .B(y[829]), .Z(n4442) );
  XNOR U5878 ( .A(n4443), .B(n4442), .Z(n4444) );
  XNOR U5879 ( .A(n4445), .B(n4444), .Z(n1919) );
  XNOR U5880 ( .A(n1918), .B(n1919), .Z(n1920) );
  XNOR U5881 ( .A(n1921), .B(n1920), .Z(n2204) );
  XNOR U5882 ( .A(n2205), .B(n2204), .Z(n1325) );
  XNOR U5883 ( .A(x[694]), .B(y[694]), .Z(n2437) );
  XNOR U5884 ( .A(x[690]), .B(y[690]), .Z(n2435) );
  XOR U5885 ( .A(x[1098]), .B(y[1098]), .Z(n2434) );
  XNOR U5886 ( .A(n2435), .B(n2434), .Z(n2436) );
  XOR U5887 ( .A(n2437), .B(n2436), .Z(n2627) );
  XNOR U5888 ( .A(x[700]), .B(y[700]), .Z(n2441) );
  XNOR U5889 ( .A(x[698]), .B(y[698]), .Z(n2439) );
  XOR U5890 ( .A(x[1452]), .B(y[1452]), .Z(n2438) );
  XNOR U5891 ( .A(n2439), .B(n2438), .Z(n2440) );
  XOR U5892 ( .A(n2441), .B(n2440), .Z(n2624) );
  XNOR U5893 ( .A(x[811]), .B(y[811]), .Z(n2177) );
  XNOR U5894 ( .A(x[178]), .B(y[178]), .Z(n2175) );
  XOR U5895 ( .A(x[813]), .B(y[813]), .Z(n2174) );
  XNOR U5896 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U5897 ( .A(n2177), .B(n2176), .Z(n2625) );
  XNOR U5898 ( .A(n2624), .B(n2625), .Z(n2626) );
  XNOR U5899 ( .A(n2627), .B(n2626), .Z(n3594) );
  XNOR U5900 ( .A(x[704]), .B(y[704]), .Z(n2351) );
  XNOR U5901 ( .A(x[702]), .B(y[702]), .Z(n2349) );
  XOR U5902 ( .A(x[1102]), .B(y[1102]), .Z(n2348) );
  XNOR U5903 ( .A(n2349), .B(n2348), .Z(n2350) );
  XOR U5904 ( .A(n2351), .B(n2350), .Z(n2639) );
  XNOR U5905 ( .A(x[708]), .B(y[708]), .Z(n2355) );
  XNOR U5906 ( .A(x[706]), .B(y[706]), .Z(n2353) );
  XOR U5907 ( .A(x[1450]), .B(y[1450]), .Z(n2352) );
  XNOR U5908 ( .A(n2353), .B(n2352), .Z(n2354) );
  XOR U5909 ( .A(n2355), .B(n2354), .Z(n2636) );
  XNOR U5910 ( .A(x[591]), .B(y[591]), .Z(n835) );
  XNOR U5911 ( .A(x[599]), .B(y[599]), .Z(n833) );
  XOR U5912 ( .A(x[1599]), .B(y[1599]), .Z(n832) );
  XNOR U5913 ( .A(n833), .B(n832), .Z(n834) );
  XNOR U5914 ( .A(n835), .B(n834), .Z(n2637) );
  XNOR U5915 ( .A(n2636), .B(n2637), .Z(n2638) );
  XOR U5916 ( .A(n2639), .B(n2638), .Z(n3593) );
  XOR U5917 ( .A(n3594), .B(n3593), .Z(n3596) );
  XNOR U5918 ( .A(x[716]), .B(y[716]), .Z(n2339) );
  XNOR U5919 ( .A(x[712]), .B(y[712]), .Z(n2337) );
  XOR U5920 ( .A(x[1106]), .B(y[1106]), .Z(n2336) );
  XNOR U5921 ( .A(n2337), .B(n2336), .Z(n2338) );
  XOR U5922 ( .A(n2339), .B(n2338), .Z(n2603) );
  XNOR U5923 ( .A(x[724]), .B(y[724]), .Z(n2309) );
  XNOR U5924 ( .A(x[722]), .B(y[722]), .Z(n2307) );
  XOR U5925 ( .A(x[1110]), .B(y[1110]), .Z(n2306) );
  XNOR U5926 ( .A(n2307), .B(n2306), .Z(n2308) );
  XOR U5927 ( .A(n2309), .B(n2308), .Z(n2600) );
  XNOR U5928 ( .A(x[720]), .B(y[720]), .Z(n2343) );
  XNOR U5929 ( .A(x[718]), .B(y[718]), .Z(n2341) );
  XOR U5930 ( .A(x[1448]), .B(y[1448]), .Z(n2340) );
  XNOR U5931 ( .A(n2341), .B(n2340), .Z(n2342) );
  XNOR U5932 ( .A(n2343), .B(n2342), .Z(n2601) );
  XNOR U5933 ( .A(n2600), .B(n2601), .Z(n2602) );
  XNOR U5934 ( .A(n2603), .B(n2602), .Z(n3595) );
  XNOR U5935 ( .A(n3596), .B(n3595), .Z(n1322) );
  XNOR U5936 ( .A(x[662]), .B(y[662]), .Z(n2469) );
  XNOR U5937 ( .A(x[658]), .B(y[658]), .Z(n2467) );
  XOR U5938 ( .A(x[1086]), .B(y[1086]), .Z(n2466) );
  XNOR U5939 ( .A(n2467), .B(n2466), .Z(n2468) );
  XOR U5940 ( .A(n2469), .B(n2468), .Z(n2645) );
  XNOR U5941 ( .A(x[668]), .B(y[668]), .Z(n2473) );
  XNOR U5942 ( .A(x[664]), .B(y[664]), .Z(n2471) );
  XOR U5943 ( .A(x[1458]), .B(y[1458]), .Z(n2470) );
  XNOR U5944 ( .A(n2471), .B(n2470), .Z(n2472) );
  XOR U5945 ( .A(n2473), .B(n2472), .Z(n2642) );
  XNOR U5946 ( .A(x[1593]), .B(y[1593]), .Z(n3275) );
  XNOR U5947 ( .A(x[587]), .B(y[587]), .Z(n3273) );
  XOR U5948 ( .A(x[1595]), .B(y[1595]), .Z(n3272) );
  XNOR U5949 ( .A(n3273), .B(n3272), .Z(n3274) );
  XNOR U5950 ( .A(n3275), .B(n3274), .Z(n2643) );
  XNOR U5951 ( .A(n2642), .B(n2643), .Z(n2644) );
  XNOR U5952 ( .A(n2645), .B(n2644), .Z(n3684) );
  XNOR U5953 ( .A(x[672]), .B(y[672]), .Z(n2481) );
  XNOR U5954 ( .A(x[670]), .B(y[670]), .Z(n2479) );
  XOR U5955 ( .A(x[1090]), .B(y[1090]), .Z(n2478) );
  XNOR U5956 ( .A(n2479), .B(n2478), .Z(n2480) );
  XOR U5957 ( .A(n2481), .B(n2480), .Z(n2651) );
  XNOR U5958 ( .A(x[680]), .B(y[680]), .Z(n2485) );
  XNOR U5959 ( .A(x[676]), .B(y[676]), .Z(n2483) );
  XOR U5960 ( .A(x[1456]), .B(y[1456]), .Z(n2482) );
  XNOR U5961 ( .A(n2483), .B(n2482), .Z(n2484) );
  XOR U5962 ( .A(n2485), .B(n2484), .Z(n2648) );
  XNOR U5963 ( .A(x[819]), .B(y[819]), .Z(n4437) );
  XNOR U5964 ( .A(x[172]), .B(y[172]), .Z(n4435) );
  XOR U5965 ( .A(x[821]), .B(y[821]), .Z(n4434) );
  XNOR U5966 ( .A(n4435), .B(n4434), .Z(n4436) );
  XNOR U5967 ( .A(n4437), .B(n4436), .Z(n2649) );
  XNOR U5968 ( .A(n2648), .B(n2649), .Z(n2650) );
  XOR U5969 ( .A(n2651), .B(n2650), .Z(n3683) );
  XOR U5970 ( .A(n3684), .B(n3683), .Z(n3686) );
  XNOR U5971 ( .A(x[684]), .B(y[684]), .Z(n2423) );
  XNOR U5972 ( .A(x[682]), .B(y[682]), .Z(n2421) );
  XOR U5973 ( .A(x[1094]), .B(y[1094]), .Z(n2420) );
  XNOR U5974 ( .A(n2421), .B(n2420), .Z(n2422) );
  XOR U5975 ( .A(n2423), .B(n2422), .Z(n2621) );
  XNOR U5976 ( .A(x[688]), .B(y[688]), .Z(n2427) );
  XNOR U5977 ( .A(x[686]), .B(y[686]), .Z(n2425) );
  XOR U5978 ( .A(x[1454]), .B(y[1454]), .Z(n2424) );
  XNOR U5979 ( .A(n2425), .B(n2424), .Z(n2426) );
  XOR U5980 ( .A(n2427), .B(n2426), .Z(n2618) );
  XNOR U5981 ( .A(x[589]), .B(y[589]), .Z(n923) );
  XOR U5982 ( .A(x[1597]), .B(y[1597]), .Z(n922) );
  XNOR U5983 ( .A(n923), .B(n922), .Z(n924) );
  XNOR U5984 ( .A(x[595]), .B(y[595]), .Z(n4655) );
  XOR U5985 ( .A(x[597]), .B(y[597]), .Z(n4654) );
  XNOR U5986 ( .A(n4655), .B(n4654), .Z(n925) );
  XOR U5987 ( .A(n924), .B(n925), .Z(n2619) );
  XNOR U5988 ( .A(n2618), .B(n2619), .Z(n2620) );
  XNOR U5989 ( .A(n2621), .B(n2620), .Z(n3685) );
  XOR U5990 ( .A(n3686), .B(n3685), .Z(n1323) );
  XNOR U5991 ( .A(n1322), .B(n1323), .Z(n1324) );
  XOR U5992 ( .A(n1325), .B(n1324), .Z(n1356) );
  XOR U5993 ( .A(n1357), .B(n1356), .Z(n1359) );
  XNOR U5994 ( .A(x[730]), .B(y[730]), .Z(n2305) );
  XNOR U5995 ( .A(x[726]), .B(y[726]), .Z(n2303) );
  XOR U5996 ( .A(x[1446]), .B(y[1446]), .Z(n2302) );
  XNOR U5997 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U5998 ( .A(n2305), .B(n2304), .Z(n936) );
  XNOR U5999 ( .A(x[736]), .B(y[736]), .Z(n2273) );
  XNOR U6000 ( .A(x[734]), .B(y[734]), .Z(n2271) );
  XOR U6001 ( .A(x[1114]), .B(y[1114]), .Z(n2270) );
  XNOR U6002 ( .A(n2271), .B(n2270), .Z(n2272) );
  XNOR U6003 ( .A(n2273), .B(n2272), .Z(n934) );
  XNOR U6004 ( .A(x[740]), .B(y[740]), .Z(n2269) );
  XNOR U6005 ( .A(x[738]), .B(y[738]), .Z(n2267) );
  XOR U6006 ( .A(x[1444]), .B(y[1444]), .Z(n2266) );
  XNOR U6007 ( .A(n2267), .B(n2266), .Z(n2268) );
  XNOR U6008 ( .A(n2269), .B(n2268), .Z(n935) );
  XNOR U6009 ( .A(n934), .B(n935), .Z(n937) );
  XNOR U6010 ( .A(n936), .B(n937), .Z(n3642) );
  XNOR U6011 ( .A(x[744]), .B(y[744]), .Z(n3786) );
  XNOR U6012 ( .A(x[742]), .B(y[742]), .Z(n3784) );
  XOR U6013 ( .A(x[1118]), .B(y[1118]), .Z(n3783) );
  XNOR U6014 ( .A(n3784), .B(n3783), .Z(n3785) );
  XOR U6015 ( .A(n3786), .B(n3785), .Z(n2615) );
  XNOR U6016 ( .A(x[752]), .B(y[752]), .Z(n3782) );
  XNOR U6017 ( .A(x[748]), .B(y[748]), .Z(n3780) );
  XOR U6018 ( .A(x[1442]), .B(y[1442]), .Z(n3779) );
  XNOR U6019 ( .A(n3780), .B(n3779), .Z(n3781) );
  XOR U6020 ( .A(n3782), .B(n3781), .Z(n2612) );
  XNOR U6021 ( .A(x[329]), .B(y[329]), .Z(n2791) );
  XNOR U6022 ( .A(x[331]), .B(y[331]), .Z(n2789) );
  XOR U6023 ( .A(x[332]), .B(y[332]), .Z(n2788) );
  XNOR U6024 ( .A(n2789), .B(n2788), .Z(n2790) );
  XNOR U6025 ( .A(n2791), .B(n2790), .Z(n2613) );
  XNOR U6026 ( .A(n2612), .B(n2613), .Z(n2614) );
  XOR U6027 ( .A(n2615), .B(n2614), .Z(n3641) );
  XOR U6028 ( .A(n3642), .B(n3641), .Z(n3644) );
  XNOR U6029 ( .A(x[756]), .B(y[756]), .Z(n3764) );
  XNOR U6030 ( .A(x[754]), .B(y[754]), .Z(n3762) );
  XOR U6031 ( .A(x[1122]), .B(y[1122]), .Z(n3761) );
  XNOR U6032 ( .A(n3762), .B(n3761), .Z(n3763) );
  XOR U6033 ( .A(n3764), .B(n3763), .Z(n2609) );
  XNOR U6034 ( .A(x[760]), .B(y[760]), .Z(n3760) );
  XNOR U6035 ( .A(x[758]), .B(y[758]), .Z(n3758) );
  XOR U6036 ( .A(x[1440]), .B(y[1440]), .Z(n3757) );
  XNOR U6037 ( .A(n3758), .B(n3757), .Z(n3759) );
  XOR U6038 ( .A(n3760), .B(n3759), .Z(n2606) );
  XNOR U6039 ( .A(x[309]), .B(y[309]), .Z(n2795) );
  XNOR U6040 ( .A(x[313]), .B(y[313]), .Z(n2793) );
  XOR U6041 ( .A(x[317]), .B(y[317]), .Z(n2792) );
  XNOR U6042 ( .A(n2793), .B(n2792), .Z(n2794) );
  XNOR U6043 ( .A(n2795), .B(n2794), .Z(n2607) );
  XNOR U6044 ( .A(n2606), .B(n2607), .Z(n2608) );
  XNOR U6045 ( .A(n2609), .B(n2608), .Z(n3643) );
  XNOR U6046 ( .A(n3644), .B(n3643), .Z(n1265) );
  XNOR U6047 ( .A(x[796]), .B(y[796]), .Z(n3213) );
  XNOR U6048 ( .A(x[794]), .B(y[794]), .Z(n3211) );
  XOR U6049 ( .A(x[1138]), .B(y[1138]), .Z(n3210) );
  XNOR U6050 ( .A(n3211), .B(n3210), .Z(n3212) );
  XOR U6051 ( .A(n3213), .B(n3212), .Z(n2061) );
  XNOR U6052 ( .A(x[802]), .B(y[802]), .Z(n2013) );
  XNOR U6053 ( .A(x[798]), .B(y[798]), .Z(n2011) );
  XOR U6054 ( .A(x[1432]), .B(y[1432]), .Z(n2010) );
  XNOR U6055 ( .A(n2011), .B(n2010), .Z(n2012) );
  XOR U6056 ( .A(n2013), .B(n2012), .Z(n2058) );
  XNOR U6057 ( .A(x[257]), .B(y[257]), .Z(n3021) );
  XNOR U6058 ( .A(x[259]), .B(y[259]), .Z(n3019) );
  XOR U6059 ( .A(x[263]), .B(y[263]), .Z(n3018) );
  XNOR U6060 ( .A(n3019), .B(n3018), .Z(n3020) );
  XNOR U6061 ( .A(n3021), .B(n3020), .Z(n2059) );
  XNOR U6062 ( .A(n2058), .B(n2059), .Z(n2060) );
  XNOR U6063 ( .A(n2061), .B(n2060), .Z(n2161) );
  XNOR U6064 ( .A(x[1330]), .B(y[1330]), .Z(n4691) );
  XNOR U6065 ( .A(x[1328]), .B(y[1328]), .Z(n4689) );
  XOR U6066 ( .A(x[1338]), .B(y[1338]), .Z(n4688) );
  XNOR U6067 ( .A(n4689), .B(n4688), .Z(n4690) );
  XOR U6068 ( .A(n4691), .B(n4690), .Z(n1837) );
  XNOR U6069 ( .A(x[1350]), .B(y[1350]), .Z(n4687) );
  XNOR U6070 ( .A(x[1344]), .B(y[1344]), .Z(n4685) );
  XOR U6071 ( .A(x[1348]), .B(y[1348]), .Z(n4684) );
  XNOR U6072 ( .A(n4685), .B(n4684), .Z(n4686) );
  XOR U6073 ( .A(n4687), .B(n4686), .Z(n1834) );
  XNOR U6074 ( .A(x[1352]), .B(y[1352]), .Z(n4683) );
  XNOR U6075 ( .A(x[1332]), .B(y[1332]), .Z(n4681) );
  XOR U6076 ( .A(x[1336]), .B(y[1336]), .Z(n4680) );
  XNOR U6077 ( .A(n4681), .B(n4680), .Z(n4682) );
  XNOR U6078 ( .A(n4683), .B(n4682), .Z(n1835) );
  XNOR U6079 ( .A(n1834), .B(n1835), .Z(n1836) );
  XOR U6080 ( .A(n1837), .B(n1836), .Z(n2160) );
  XOR U6081 ( .A(n2161), .B(n2160), .Z(n2163) );
  XNOR U6082 ( .A(x[808]), .B(y[808]), .Z(n885) );
  XNOR U6083 ( .A(x[806]), .B(y[806]), .Z(n883) );
  XOR U6084 ( .A(x[1142]), .B(y[1142]), .Z(n882) );
  XNOR U6085 ( .A(n883), .B(n882), .Z(n884) );
  XOR U6086 ( .A(n885), .B(n884), .Z(n1059) );
  XNOR U6087 ( .A(x[812]), .B(y[812]), .Z(n881) );
  XNOR U6088 ( .A(x[810]), .B(y[810]), .Z(n879) );
  XOR U6089 ( .A(x[1430]), .B(y[1430]), .Z(n878) );
  XNOR U6090 ( .A(n879), .B(n878), .Z(n880) );
  XOR U6091 ( .A(n881), .B(n880), .Z(n1056) );
  XNOR U6092 ( .A(x[241]), .B(y[241]), .Z(n3003) );
  XNOR U6093 ( .A(x[243]), .B(y[243]), .Z(n3001) );
  XNOR U6094 ( .A(x[428]), .B(y[428]), .Z(n3000) );
  XNOR U6095 ( .A(n3001), .B(n3000), .Z(n3002) );
  XOR U6096 ( .A(n3003), .B(n3002), .Z(n1057) );
  XNOR U6097 ( .A(n1056), .B(n1057), .Z(n1058) );
  XNOR U6098 ( .A(n1059), .B(n1058), .Z(n2162) );
  XNOR U6099 ( .A(n2163), .B(n2162), .Z(n1262) );
  XNOR U6100 ( .A(x[766]), .B(y[766]), .Z(n2029) );
  XNOR U6101 ( .A(x[762]), .B(y[762]), .Z(n2027) );
  XOR U6102 ( .A(x[1126]), .B(y[1126]), .Z(n2026) );
  XNOR U6103 ( .A(n2027), .B(n2026), .Z(n2028) );
  XOR U6104 ( .A(n2029), .B(n2028), .Z(n2633) );
  XNOR U6105 ( .A(x[776]), .B(y[776]), .Z(n2017) );
  XNOR U6106 ( .A(x[774]), .B(y[774]), .Z(n2015) );
  XOR U6107 ( .A(x[1130]), .B(y[1130]), .Z(n2014) );
  XNOR U6108 ( .A(n2015), .B(n2014), .Z(n2016) );
  XOR U6109 ( .A(n2017), .B(n2016), .Z(n2630) );
  XNOR U6110 ( .A(x[772]), .B(y[772]), .Z(n2025) );
  XNOR U6111 ( .A(x[770]), .B(y[770]), .Z(n2023) );
  XOR U6112 ( .A(x[1438]), .B(y[1438]), .Z(n2022) );
  XNOR U6113 ( .A(n2023), .B(n2022), .Z(n2024) );
  XNOR U6114 ( .A(n2025), .B(n2024), .Z(n2631) );
  XNOR U6115 ( .A(n2630), .B(n2631), .Z(n2632) );
  XNOR U6116 ( .A(n2633), .B(n2632), .Z(n2107) );
  XNOR U6117 ( .A(x[572]), .B(y[572]), .Z(n2173) );
  XNOR U6118 ( .A(x[570]), .B(y[570]), .Z(n2171) );
  XOR U6119 ( .A(x[854]), .B(y[854]), .Z(n2170) );
  XNOR U6120 ( .A(n2171), .B(n2170), .Z(n2172) );
  XOR U6121 ( .A(n2173), .B(n2172), .Z(n4707) );
  XNOR U6122 ( .A(x[576]), .B(y[576]), .Z(n4653) );
  XNOR U6123 ( .A(x[574]), .B(y[574]), .Z(n4651) );
  XOR U6124 ( .A(x[858]), .B(y[858]), .Z(n4650) );
  XNOR U6125 ( .A(n4651), .B(n4650), .Z(n4652) );
  XOR U6126 ( .A(n4653), .B(n4652), .Z(n4704) );
  XNOR U6127 ( .A(x[1340]), .B(y[1340]), .Z(n4659) );
  XNOR U6128 ( .A(x[1334]), .B(y[1334]), .Z(n4657) );
  XOR U6129 ( .A(x[1346]), .B(y[1346]), .Z(n4656) );
  XNOR U6130 ( .A(n4657), .B(n4656), .Z(n4658) );
  XNOR U6131 ( .A(n4659), .B(n4658), .Z(n4705) );
  XNOR U6132 ( .A(n4704), .B(n4705), .Z(n4706) );
  XOR U6133 ( .A(n4707), .B(n4706), .Z(n2106) );
  XOR U6134 ( .A(n2107), .B(n2106), .Z(n2109) );
  XNOR U6135 ( .A(x[780]), .B(y[780]), .Z(n2699) );
  XNOR U6136 ( .A(x[778]), .B(y[778]), .Z(n2697) );
  XOR U6137 ( .A(x[1436]), .B(y[1436]), .Z(n2696) );
  XNOR U6138 ( .A(n2697), .B(n2696), .Z(n2698) );
  XOR U6139 ( .A(n2699), .B(n2698), .Z(n2085) );
  XNOR U6140 ( .A(x[792]), .B(y[792]), .Z(n3125) );
  XNOR U6141 ( .A(x[790]), .B(y[790]), .Z(n3123) );
  XNOR U6142 ( .A(x[1434]), .B(y[1434]), .Z(n3122) );
  XNOR U6143 ( .A(n3123), .B(n3122), .Z(n3124) );
  XNOR U6144 ( .A(n3125), .B(n3124), .Z(n2082) );
  XNOR U6145 ( .A(x[788]), .B(y[788]), .Z(n2733) );
  XNOR U6146 ( .A(x[784]), .B(y[784]), .Z(n2731) );
  XOR U6147 ( .A(x[1134]), .B(y[1134]), .Z(n2730) );
  XNOR U6148 ( .A(n2731), .B(n2730), .Z(n2732) );
  XNOR U6149 ( .A(n2733), .B(n2732), .Z(n2083) );
  XNOR U6150 ( .A(n2082), .B(n2083), .Z(n2084) );
  XNOR U6151 ( .A(n2085), .B(n2084), .Z(n2108) );
  XOR U6152 ( .A(n2109), .B(n2108), .Z(n1263) );
  XNOR U6153 ( .A(n1262), .B(n1263), .Z(n1264) );
  XNOR U6154 ( .A(n1265), .B(n1264), .Z(n1358) );
  XOR U6155 ( .A(n1359), .B(n1358), .Z(n1173) );
  XNOR U6156 ( .A(n1172), .B(n1173), .Z(n1174) );
  XOR U6157 ( .A(n1175), .B(n1174), .Z(n804) );
  XOR U6158 ( .A(n805), .B(n804), .Z(o[0]) );
  NANDN U6159 ( .A(n803), .B(n802), .Z(n807) );
  OR U6160 ( .A(n805), .B(n804), .Z(n806) );
  NAND U6161 ( .A(n807), .B(n806), .Z(n6747) );
  NAND U6162 ( .A(n809), .B(n808), .Z(n813) );
  NANDN U6163 ( .A(n811), .B(n810), .Z(n812) );
  NAND U6164 ( .A(n813), .B(n812), .Z(n4966) );
  NANDN U6165 ( .A(n815), .B(n814), .Z(n819) );
  NAND U6166 ( .A(n817), .B(n816), .Z(n818) );
  NAND U6167 ( .A(n819), .B(n818), .Z(n6776) );
  NANDN U6168 ( .A(n821), .B(n820), .Z(n825) );
  NAND U6169 ( .A(n823), .B(n822), .Z(n824) );
  AND U6170 ( .A(n825), .B(n824), .Z(n6777) );
  XNOR U6171 ( .A(n6776), .B(n6777), .Z(n6778) );
  NANDN U6172 ( .A(n827), .B(n826), .Z(n831) );
  NAND U6173 ( .A(n829), .B(n828), .Z(n830) );
  NAND U6174 ( .A(n831), .B(n830), .Z(n6901) );
  OR U6175 ( .A(n837), .B(n836), .Z(n841) );
  NANDN U6176 ( .A(n839), .B(n838), .Z(n840) );
  NAND U6177 ( .A(n841), .B(n840), .Z(n5438) );
  OR U6178 ( .A(n843), .B(n842), .Z(n847) );
  NANDN U6179 ( .A(n845), .B(n844), .Z(n846) );
  NAND U6180 ( .A(n847), .B(n846), .Z(n5441) );
  XOR U6181 ( .A(n5440), .B(n5441), .Z(n6898) );
  XNOR U6182 ( .A(n6021), .B(n6022), .Z(n6899) );
  XNOR U6183 ( .A(n6898), .B(n6899), .Z(n6900) );
  XOR U6184 ( .A(n6901), .B(n6900), .Z(n7145) );
  XNOR U6185 ( .A(n5780), .B(n5779), .Z(n5781) );
  XOR U6186 ( .A(n5781), .B(n5782), .Z(n7121) );
  OR U6187 ( .A(n873), .B(n872), .Z(n877) );
  NANDN U6188 ( .A(n875), .B(n874), .Z(n876) );
  NAND U6189 ( .A(n877), .B(n876), .Z(n5493) );
  XOR U6190 ( .A(n5494), .B(n5495), .Z(n7118) );
  XNOR U6191 ( .A(n5979), .B(n5980), .Z(n7119) );
  XNOR U6192 ( .A(n7118), .B(n7119), .Z(n7120) );
  XNOR U6193 ( .A(n7121), .B(n7120), .Z(n7142) );
  XOR U6194 ( .A(n5608), .B(n5609), .Z(n7133) );
  XOR U6195 ( .A(n5991), .B(n5992), .Z(n7130) );
  XNOR U6196 ( .A(n5387), .B(n5386), .Z(n7131) );
  XNOR U6197 ( .A(n7130), .B(n7131), .Z(n7132) );
  XOR U6198 ( .A(n7133), .B(n7132), .Z(n7143) );
  XNOR U6199 ( .A(n7142), .B(n7143), .Z(n7144) );
  XNOR U6200 ( .A(n7145), .B(n7144), .Z(n5416) );
  OR U6201 ( .A(n935), .B(n934), .Z(n939) );
  OR U6202 ( .A(n937), .B(n936), .Z(n938) );
  NAND U6203 ( .A(n939), .B(n938), .Z(n5137) );
  NANDN U6204 ( .A(n941), .B(n940), .Z(n945) );
  OR U6205 ( .A(n943), .B(n942), .Z(n944) );
  NAND U6206 ( .A(n945), .B(n944), .Z(n5134) );
  XNOR U6207 ( .A(n5263), .B(n5262), .Z(n5264) );
  OR U6208 ( .A(n955), .B(n954), .Z(n959) );
  NANDN U6209 ( .A(n957), .B(n956), .Z(n958) );
  NAND U6210 ( .A(n959), .B(n958), .Z(n5265) );
  XOR U6211 ( .A(n5264), .B(n5265), .Z(n5998) );
  OR U6212 ( .A(n965), .B(n964), .Z(n969) );
  NANDN U6213 ( .A(n967), .B(n966), .Z(n968) );
  AND U6214 ( .A(n969), .B(n968), .Z(n5773) );
  XNOR U6215 ( .A(n5774), .B(n5773), .Z(n5775) );
  OR U6216 ( .A(n971), .B(n970), .Z(n975) );
  NANDN U6217 ( .A(n973), .B(n972), .Z(n974) );
  NAND U6218 ( .A(n975), .B(n974), .Z(n5776) );
  XOR U6219 ( .A(n5775), .B(n5776), .Z(n5995) );
  OR U6220 ( .A(n977), .B(n976), .Z(n981) );
  NAND U6221 ( .A(n979), .B(n978), .Z(n980) );
  NAND U6222 ( .A(n981), .B(n980), .Z(n5996) );
  XNOR U6223 ( .A(n5995), .B(n5996), .Z(n5997) );
  XOR U6224 ( .A(n5998), .B(n5997), .Z(n5135) );
  XNOR U6225 ( .A(n5134), .B(n5135), .Z(n5136) );
  XNOR U6226 ( .A(n5137), .B(n5136), .Z(n5414) );
  XOR U6227 ( .A(n5414), .B(n5415), .Z(n5417) );
  XNOR U6228 ( .A(n5416), .B(n5417), .Z(n6779) );
  XNOR U6229 ( .A(n6778), .B(n6779), .Z(n6790) );
  XNOR U6230 ( .A(n5577), .B(n5576), .Z(n5578) );
  XOR U6231 ( .A(n5578), .B(n5579), .Z(n7208) );
  XNOR U6232 ( .A(n5565), .B(n5564), .Z(n5566) );
  XNOR U6233 ( .A(n5566), .B(n5567), .Z(n7206) );
  OR U6234 ( .A(n1011), .B(n1010), .Z(n1015) );
  NAND U6235 ( .A(n1013), .B(n1012), .Z(n1014) );
  NAND U6236 ( .A(n1015), .B(n1014), .Z(n7207) );
  XOR U6237 ( .A(n7208), .B(n7209), .Z(n6931) );
  OR U6238 ( .A(n1021), .B(n1020), .Z(n1025) );
  NANDN U6239 ( .A(n1023), .B(n1022), .Z(n1024) );
  AND U6240 ( .A(n1025), .B(n1024), .Z(n5600) );
  XNOR U6241 ( .A(n5601), .B(n5600), .Z(n5602) );
  XOR U6242 ( .A(n5602), .B(n5603), .Z(n5217) );
  XNOR U6243 ( .A(n6698), .B(n6697), .Z(n6699) );
  OR U6244 ( .A(n1039), .B(n1038), .Z(n1043) );
  NANDN U6245 ( .A(n1041), .B(n1040), .Z(n1042) );
  NAND U6246 ( .A(n1043), .B(n1042), .Z(n6700) );
  XOR U6247 ( .A(n6699), .B(n6700), .Z(n5214) );
  NANDN U6248 ( .A(n1045), .B(n1044), .Z(n1049) );
  NAND U6249 ( .A(n1047), .B(n1046), .Z(n1048) );
  NAND U6250 ( .A(n1049), .B(n1048), .Z(n5215) );
  XNOR U6251 ( .A(n5214), .B(n5215), .Z(n5216) );
  XNOR U6252 ( .A(n5217), .B(n5216), .Z(n6928) );
  NANDN U6253 ( .A(n1051), .B(n1050), .Z(n1055) );
  NAND U6254 ( .A(n1053), .B(n1052), .Z(n1054) );
  NAND U6255 ( .A(n1055), .B(n1054), .Z(n6929) );
  XNOR U6256 ( .A(n6928), .B(n6929), .Z(n6930) );
  XOR U6257 ( .A(n6931), .B(n6930), .Z(n5131) );
  NANDN U6258 ( .A(n1057), .B(n1056), .Z(n1061) );
  NAND U6259 ( .A(n1059), .B(n1058), .Z(n1060) );
  NAND U6260 ( .A(n1061), .B(n1060), .Z(n6913) );
  NANDN U6261 ( .A(n1063), .B(n1062), .Z(n1067) );
  NAND U6262 ( .A(n1065), .B(n1064), .Z(n1066) );
  NAND U6263 ( .A(n1067), .B(n1066), .Z(n6911) );
  NANDN U6264 ( .A(n1069), .B(n1068), .Z(n1073) );
  NAND U6265 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U6266 ( .A(n1073), .B(n1072), .Z(n6910) );
  XNOR U6267 ( .A(n6911), .B(n6910), .Z(n6912) );
  XNOR U6268 ( .A(n6913), .B(n6912), .Z(n6940) );
  XNOR U6269 ( .A(n5257), .B(n5256), .Z(n5258) );
  XOR U6270 ( .A(n5258), .B(n5259), .Z(n6959) );
  OR U6271 ( .A(n1087), .B(n1086), .Z(n1091) );
  NANDN U6272 ( .A(n1089), .B(n1088), .Z(n1090) );
  NAND U6273 ( .A(n1091), .B(n1090), .Z(n5924) );
  OR U6274 ( .A(n1093), .B(n1092), .Z(n1097) );
  NANDN U6275 ( .A(n1095), .B(n1094), .Z(n1096) );
  NAND U6276 ( .A(n1097), .B(n1096), .Z(n5923) );
  OR U6277 ( .A(n1099), .B(n1098), .Z(n1103) );
  NANDN U6278 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U6279 ( .A(n1103), .B(n1102), .Z(n5926) );
  XOR U6280 ( .A(n5925), .B(n5926), .Z(n6956) );
  XNOR U6281 ( .A(n5614), .B(n5615), .Z(n6957) );
  XNOR U6282 ( .A(n6956), .B(n6957), .Z(n6958) );
  XOR U6283 ( .A(n6959), .B(n6958), .Z(n6941) );
  XOR U6284 ( .A(n6940), .B(n6941), .Z(n6942) );
  OR U6285 ( .A(n1117), .B(n1116), .Z(n1121) );
  NANDN U6286 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U6287 ( .A(n1121), .B(n1120), .Z(n6704) );
  OR U6288 ( .A(n1123), .B(n1122), .Z(n1127) );
  NANDN U6289 ( .A(n1125), .B(n1124), .Z(n1126) );
  NAND U6290 ( .A(n1127), .B(n1126), .Z(n6703) );
  OR U6291 ( .A(n1129), .B(n1128), .Z(n1133) );
  NANDN U6292 ( .A(n1131), .B(n1130), .Z(n1132) );
  NAND U6293 ( .A(n1133), .B(n1132), .Z(n6706) );
  XOR U6294 ( .A(n6705), .B(n6706), .Z(n6953) );
  XOR U6295 ( .A(n6027), .B(n6028), .Z(n6950) );
  OR U6296 ( .A(n1147), .B(n1146), .Z(n1151) );
  NANDN U6297 ( .A(n1149), .B(n1148), .Z(n1150) );
  NAND U6298 ( .A(n1151), .B(n1150), .Z(n5391) );
  OR U6299 ( .A(n1157), .B(n1156), .Z(n1161) );
  NANDN U6300 ( .A(n1159), .B(n1158), .Z(n1160) );
  NAND U6301 ( .A(n1161), .B(n1160), .Z(n5393) );
  XNOR U6302 ( .A(n5392), .B(n5393), .Z(n6951) );
  XNOR U6303 ( .A(n6950), .B(n6951), .Z(n6952) );
  XOR U6304 ( .A(n6953), .B(n6952), .Z(n6943) );
  XOR U6305 ( .A(n6942), .B(n6943), .Z(n5128) );
  NAND U6306 ( .A(n1163), .B(n1162), .Z(n1167) );
  NAND U6307 ( .A(n1165), .B(n1164), .Z(n1166) );
  AND U6308 ( .A(n1167), .B(n1166), .Z(n5129) );
  XOR U6309 ( .A(n5128), .B(n5129), .Z(n5130) );
  XNOR U6310 ( .A(n5131), .B(n5130), .Z(n6788) );
  XOR U6311 ( .A(n6788), .B(n6789), .Z(n6791) );
  XNOR U6312 ( .A(n6790), .B(n6791), .Z(n4964) );
  NANDN U6313 ( .A(n1173), .B(n1172), .Z(n1177) );
  NAND U6314 ( .A(n1175), .B(n1174), .Z(n1176) );
  NAND U6315 ( .A(n1177), .B(n1176), .Z(n4965) );
  XOR U6316 ( .A(n4964), .B(n4965), .Z(n4967) );
  XOR U6317 ( .A(n4966), .B(n4967), .Z(n6746) );
  XNOR U6318 ( .A(n6747), .B(n6746), .Z(n6749) );
  NANDN U6319 ( .A(n1179), .B(n1178), .Z(n1183) );
  NANDN U6320 ( .A(n1181), .B(n1180), .Z(n1182) );
  NAND U6321 ( .A(n1183), .B(n1182), .Z(n6830) );
  NANDN U6322 ( .A(n1185), .B(n1184), .Z(n1189) );
  NAND U6323 ( .A(n1187), .B(n1186), .Z(n1188) );
  NAND U6324 ( .A(n1189), .B(n1188), .Z(n6829) );
  NANDN U6325 ( .A(n1195), .B(n1194), .Z(n1199) );
  NAND U6326 ( .A(n1197), .B(n1196), .Z(n1198) );
  NAND U6327 ( .A(n1199), .B(n1198), .Z(n5471) );
  XNOR U6328 ( .A(n6079), .B(n6080), .Z(n5468) );
  NANDN U6329 ( .A(n1213), .B(n1212), .Z(n1217) );
  NAND U6330 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U6331 ( .A(n1217), .B(n1216), .Z(n5469) );
  XOR U6332 ( .A(n5471), .B(n5470), .Z(n5059) );
  XOR U6333 ( .A(n5058), .B(n5059), .Z(n5060) );
  OR U6334 ( .A(n1219), .B(n1218), .Z(n1223) );
  NANDN U6335 ( .A(n1221), .B(n1220), .Z(n1222) );
  NAND U6336 ( .A(n1223), .B(n1222), .Z(n6632) );
  OR U6337 ( .A(n1229), .B(n1228), .Z(n1233) );
  NANDN U6338 ( .A(n1231), .B(n1230), .Z(n1232) );
  NAND U6339 ( .A(n1233), .B(n1232), .Z(n6634) );
  XOR U6340 ( .A(n6633), .B(n6634), .Z(n5805) );
  OR U6341 ( .A(n1235), .B(n1234), .Z(n1239) );
  NANDN U6342 ( .A(n1237), .B(n1236), .Z(n1238) );
  NAND U6343 ( .A(n1239), .B(n1238), .Z(n6638) );
  OR U6344 ( .A(n1241), .B(n1240), .Z(n1245) );
  NANDN U6345 ( .A(n1243), .B(n1242), .Z(n1244) );
  NAND U6346 ( .A(n1245), .B(n1244), .Z(n6637) );
  OR U6347 ( .A(n1247), .B(n1246), .Z(n1251) );
  NANDN U6348 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U6349 ( .A(n1251), .B(n1250), .Z(n6640) );
  XNOR U6350 ( .A(n6639), .B(n6640), .Z(n5803) );
  OR U6351 ( .A(n1253), .B(n1252), .Z(n1257) );
  NAND U6352 ( .A(n1255), .B(n1254), .Z(n1256) );
  NAND U6353 ( .A(n1257), .B(n1256), .Z(n5804) );
  XOR U6354 ( .A(n5805), .B(n5806), .Z(n5061) );
  XNOR U6355 ( .A(n5060), .B(n5061), .Z(n6828) );
  XNOR U6356 ( .A(n6829), .B(n6828), .Z(n6831) );
  XNOR U6357 ( .A(n6830), .B(n6831), .Z(n5835) );
  NANDN U6358 ( .A(n1263), .B(n1262), .Z(n1267) );
  NAND U6359 ( .A(n1265), .B(n1264), .Z(n1266) );
  NAND U6360 ( .A(n1267), .B(n1266), .Z(n6823) );
  NANDN U6361 ( .A(n1269), .B(n1268), .Z(n1273) );
  OR U6362 ( .A(n1271), .B(n1270), .Z(n1272) );
  NAND U6363 ( .A(n1273), .B(n1272), .Z(n7108) );
  NANDN U6364 ( .A(n1275), .B(n1274), .Z(n1279) );
  NAND U6365 ( .A(n1277), .B(n1276), .Z(n1278) );
  NAND U6366 ( .A(n1279), .B(n1278), .Z(n6971) );
  OR U6367 ( .A(n1281), .B(n1280), .Z(n1285) );
  OR U6368 ( .A(n1283), .B(n1282), .Z(n1284) );
  NAND U6369 ( .A(n1285), .B(n1284), .Z(n6144) );
  OR U6370 ( .A(n1287), .B(n1286), .Z(n1291) );
  OR U6371 ( .A(n1289), .B(n1288), .Z(n1290) );
  AND U6372 ( .A(n1291), .B(n1290), .Z(n6143) );
  XNOR U6373 ( .A(n6144), .B(n6143), .Z(n6145) );
  OR U6374 ( .A(n1293), .B(n1292), .Z(n1297) );
  OR U6375 ( .A(n1295), .B(n1294), .Z(n1296) );
  NAND U6376 ( .A(n1297), .B(n1296), .Z(n6146) );
  XOR U6377 ( .A(n6145), .B(n6146), .Z(n6968) );
  NANDN U6378 ( .A(n1299), .B(n1298), .Z(n1303) );
  NAND U6379 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U6380 ( .A(n1303), .B(n1302), .Z(n6969) );
  XNOR U6381 ( .A(n6968), .B(n6969), .Z(n6970) );
  XOR U6382 ( .A(n6971), .B(n6970), .Z(n7109) );
  XOR U6383 ( .A(n7108), .B(n7109), .Z(n7110) );
  OR U6384 ( .A(n1305), .B(n1304), .Z(n1309) );
  NAND U6385 ( .A(n1307), .B(n1306), .Z(n1308) );
  NAND U6386 ( .A(n1309), .B(n1308), .Z(n5155) );
  OR U6387 ( .A(n1311), .B(n1310), .Z(n1315) );
  NANDN U6388 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U6389 ( .A(n1315), .B(n1314), .Z(n5153) );
  OR U6390 ( .A(n1317), .B(n1316), .Z(n1321) );
  NAND U6391 ( .A(n1319), .B(n1318), .Z(n1320) );
  AND U6392 ( .A(n1321), .B(n1320), .Z(n5152) );
  XNOR U6393 ( .A(n5153), .B(n5152), .Z(n5154) );
  XOR U6394 ( .A(n5155), .B(n5154), .Z(n7111) );
  XNOR U6395 ( .A(n7110), .B(n7111), .Z(n6822) );
  XNOR U6396 ( .A(n6823), .B(n6822), .Z(n6825) );
  XNOR U6397 ( .A(n6824), .B(n6825), .Z(n5833) );
  NANDN U6398 ( .A(n1323), .B(n1322), .Z(n1327) );
  NAND U6399 ( .A(n1325), .B(n1324), .Z(n1326) );
  NAND U6400 ( .A(n1327), .B(n1326), .Z(n6837) );
  NANDN U6401 ( .A(n1329), .B(n1328), .Z(n1333) );
  OR U6402 ( .A(n1331), .B(n1330), .Z(n1332) );
  NAND U6403 ( .A(n1333), .B(n1332), .Z(n7087) );
  OR U6404 ( .A(n1335), .B(n1334), .Z(n1339) );
  NAND U6405 ( .A(n1337), .B(n1336), .Z(n1338) );
  NAND U6406 ( .A(n1339), .B(n1338), .Z(n7084) );
  XNOR U6407 ( .A(n7084), .B(n7085), .Z(n7086) );
  XNOR U6408 ( .A(n7087), .B(n7086), .Z(n6834) );
  NAND U6409 ( .A(n1345), .B(n1344), .Z(n1349) );
  NAND U6410 ( .A(n1347), .B(n1346), .Z(n1348) );
  NAND U6411 ( .A(n1349), .B(n1348), .Z(n6835) );
  XNOR U6412 ( .A(n6834), .B(n6835), .Z(n6836) );
  XOR U6413 ( .A(n6837), .B(n6836), .Z(n5834) );
  XNOR U6414 ( .A(n5833), .B(n5834), .Z(n5836) );
  XNOR U6415 ( .A(n5835), .B(n5836), .Z(n7251) );
  NAND U6416 ( .A(n1351), .B(n1350), .Z(n1355) );
  NAND U6417 ( .A(n1353), .B(n1352), .Z(n1354) );
  NAND U6418 ( .A(n1355), .B(n1354), .Z(n7248) );
  NANDN U6419 ( .A(n1357), .B(n1356), .Z(n1361) );
  OR U6420 ( .A(n1359), .B(n1358), .Z(n1360) );
  NAND U6421 ( .A(n1361), .B(n1360), .Z(n7249) );
  XNOR U6422 ( .A(n7248), .B(n7249), .Z(n7250) );
  XOR U6423 ( .A(n7251), .B(n7250), .Z(n6795) );
  NANDN U6424 ( .A(n1363), .B(n1362), .Z(n1367) );
  OR U6425 ( .A(n1365), .B(n1364), .Z(n1366) );
  NAND U6426 ( .A(n1367), .B(n1366), .Z(n6843) );
  OR U6427 ( .A(n1369), .B(n1368), .Z(n1373) );
  NANDN U6428 ( .A(n1371), .B(n1370), .Z(n1372) );
  NAND U6429 ( .A(n1373), .B(n1372), .Z(n6840) );
  OR U6430 ( .A(n1375), .B(n1374), .Z(n1379) );
  NANDN U6431 ( .A(n1377), .B(n1376), .Z(n1378) );
  NAND U6432 ( .A(n1379), .B(n1378), .Z(n6541) );
  XOR U6433 ( .A(n6542), .B(n6543), .Z(n6362) );
  OR U6434 ( .A(n1389), .B(n1388), .Z(n1393) );
  NANDN U6435 ( .A(n1391), .B(n1390), .Z(n1392) );
  NAND U6436 ( .A(n1393), .B(n1392), .Z(n7237) );
  XNOR U6437 ( .A(n7237), .B(n7236), .Z(n7238) );
  XNOR U6438 ( .A(n7238), .B(n7239), .Z(n6359) );
  OR U6439 ( .A(n1403), .B(n1402), .Z(n1407) );
  NANDN U6440 ( .A(n1405), .B(n1404), .Z(n1406) );
  NAND U6441 ( .A(n1407), .B(n1406), .Z(n6360) );
  XOR U6442 ( .A(n6362), .B(n6361), .Z(n6841) );
  XNOR U6443 ( .A(n6840), .B(n6841), .Z(n6842) );
  XNOR U6444 ( .A(n6843), .B(n6842), .Z(n5109) );
  NANDN U6445 ( .A(n1409), .B(n1408), .Z(n1413) );
  OR U6446 ( .A(n1411), .B(n1410), .Z(n1412) );
  NAND U6447 ( .A(n1413), .B(n1412), .Z(n5143) );
  OR U6448 ( .A(n1423), .B(n1422), .Z(n1427) );
  NANDN U6449 ( .A(n1425), .B(n1424), .Z(n1426) );
  AND U6450 ( .A(n1427), .B(n1426), .Z(n5304) );
  XNOR U6451 ( .A(n5305), .B(n5304), .Z(n5306) );
  OR U6452 ( .A(n1429), .B(n1428), .Z(n1433) );
  NANDN U6453 ( .A(n1431), .B(n1430), .Z(n1432) );
  NAND U6454 ( .A(n1433), .B(n1432), .Z(n5307) );
  XOR U6455 ( .A(n5306), .B(n5307), .Z(n7191) );
  NANDN U6456 ( .A(n1435), .B(n1434), .Z(n1439) );
  NAND U6457 ( .A(n1437), .B(n1436), .Z(n1438) );
  NAND U6458 ( .A(n1439), .B(n1438), .Z(n7189) );
  NANDN U6459 ( .A(n1441), .B(n1440), .Z(n1445) );
  NAND U6460 ( .A(n1443), .B(n1442), .Z(n1444) );
  AND U6461 ( .A(n1445), .B(n1444), .Z(n7188) );
  XNOR U6462 ( .A(n7189), .B(n7188), .Z(n7190) );
  XOR U6463 ( .A(n7191), .B(n7190), .Z(n5141) );
  XNOR U6464 ( .A(n5140), .B(n5141), .Z(n5142) );
  XNOR U6465 ( .A(n5143), .B(n5142), .Z(n5107) );
  NANDN U6466 ( .A(n1447), .B(n1446), .Z(n1451) );
  OR U6467 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U6468 ( .A(n1451), .B(n1450), .Z(n6849) );
  OR U6469 ( .A(n1453), .B(n1452), .Z(n1457) );
  NANDN U6470 ( .A(n1455), .B(n1454), .Z(n1456) );
  NAND U6471 ( .A(n1457), .B(n1456), .Z(n6300) );
  OR U6472 ( .A(n1459), .B(n1458), .Z(n1463) );
  NANDN U6473 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U6474 ( .A(n1463), .B(n1462), .Z(n6299) );
  XNOR U6475 ( .A(n6300), .B(n6299), .Z(n6301) );
  OR U6476 ( .A(n1465), .B(n1464), .Z(n1469) );
  NANDN U6477 ( .A(n1467), .B(n1466), .Z(n1468) );
  NAND U6478 ( .A(n1469), .B(n1468), .Z(n6302) );
  XNOR U6479 ( .A(n6301), .B(n6302), .Z(n6922) );
  OR U6480 ( .A(n1471), .B(n1470), .Z(n1475) );
  NAND U6481 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U6482 ( .A(n1475), .B(n1474), .Z(n6923) );
  NANDN U6483 ( .A(n1477), .B(n1476), .Z(n1481) );
  NAND U6484 ( .A(n1479), .B(n1478), .Z(n1480) );
  AND U6485 ( .A(n1481), .B(n1480), .Z(n6925) );
  XNOR U6486 ( .A(n6924), .B(n6925), .Z(n6847) );
  OR U6487 ( .A(n1483), .B(n1482), .Z(n1487) );
  NANDN U6488 ( .A(n1485), .B(n1484), .Z(n1486) );
  AND U6489 ( .A(n1487), .B(n1486), .Z(n6846) );
  XNOR U6490 ( .A(n6847), .B(n6846), .Z(n6848) );
  XNOR U6491 ( .A(n6849), .B(n6848), .Z(n5106) );
  XOR U6492 ( .A(n5107), .B(n5106), .Z(n5108) );
  XOR U6493 ( .A(n5109), .B(n5108), .Z(n5183) );
  NANDN U6494 ( .A(n1489), .B(n1488), .Z(n1493) );
  NAND U6495 ( .A(n1491), .B(n1490), .Z(n1492) );
  NAND U6496 ( .A(n1493), .B(n1492), .Z(n7263) );
  OR U6497 ( .A(n1499), .B(n1498), .Z(n1503) );
  NANDN U6498 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U6499 ( .A(n1503), .B(n1502), .Z(n6209) );
  XNOR U6500 ( .A(n6210), .B(n6209), .Z(n6211) );
  XOR U6501 ( .A(n6211), .B(n6212), .Z(n5193) );
  NANDN U6502 ( .A(n1509), .B(n1508), .Z(n1513) );
  NAND U6503 ( .A(n1511), .B(n1510), .Z(n1512) );
  NAND U6504 ( .A(n1513), .B(n1512), .Z(n5191) );
  NANDN U6505 ( .A(n1515), .B(n1514), .Z(n1519) );
  NAND U6506 ( .A(n1517), .B(n1516), .Z(n1518) );
  AND U6507 ( .A(n1519), .B(n1518), .Z(n5190) );
  XNOR U6508 ( .A(n5191), .B(n5190), .Z(n5192) );
  XNOR U6509 ( .A(n5193), .B(n5192), .Z(n5826) );
  OR U6510 ( .A(n1525), .B(n1524), .Z(n1529) );
  NANDN U6511 ( .A(n1527), .B(n1526), .Z(n1528) );
  AND U6512 ( .A(n1529), .B(n1528), .Z(n6245) );
  XNOR U6513 ( .A(n6246), .B(n6245), .Z(n6247) );
  OR U6514 ( .A(n1531), .B(n1530), .Z(n1535) );
  NANDN U6515 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U6516 ( .A(n1535), .B(n1534), .Z(n6248) );
  XOR U6517 ( .A(n6247), .B(n6248), .Z(n5736) );
  OR U6518 ( .A(n1537), .B(n1536), .Z(n1541) );
  NAND U6519 ( .A(n1539), .B(n1538), .Z(n1540) );
  NAND U6520 ( .A(n1541), .B(n1540), .Z(n5737) );
  XNOR U6521 ( .A(n5736), .B(n5737), .Z(n5738) );
  NANDN U6522 ( .A(n1543), .B(n1542), .Z(n1547) );
  NAND U6523 ( .A(n1545), .B(n1544), .Z(n1546) );
  AND U6524 ( .A(n1547), .B(n1546), .Z(n5739) );
  XNOR U6525 ( .A(n5738), .B(n5739), .Z(n5823) );
  NANDN U6526 ( .A(n1549), .B(n1548), .Z(n1553) );
  NAND U6527 ( .A(n1551), .B(n1550), .Z(n1552) );
  NAND U6528 ( .A(n1553), .B(n1552), .Z(n5149) );
  OR U6529 ( .A(n1555), .B(n1554), .Z(n1559) );
  NAND U6530 ( .A(n1557), .B(n1556), .Z(n1558) );
  NAND U6531 ( .A(n1559), .B(n1558), .Z(n5147) );
  NANDN U6532 ( .A(n1561), .B(n1560), .Z(n1565) );
  NAND U6533 ( .A(n1563), .B(n1562), .Z(n1564) );
  AND U6534 ( .A(n1565), .B(n1564), .Z(n5146) );
  XNOR U6535 ( .A(n5147), .B(n5146), .Z(n5148) );
  XOR U6536 ( .A(n5149), .B(n5148), .Z(n5824) );
  XOR U6537 ( .A(n5823), .B(n5824), .Z(n5825) );
  XOR U6538 ( .A(n5826), .B(n5825), .Z(n7260) );
  XNOR U6539 ( .A(n5299), .B(n5298), .Z(n5300) );
  OR U6540 ( .A(n1575), .B(n1574), .Z(n1579) );
  NANDN U6541 ( .A(n1577), .B(n1576), .Z(n1578) );
  NAND U6542 ( .A(n1579), .B(n1578), .Z(n5301) );
  XOR U6543 ( .A(n5300), .B(n5301), .Z(n6221) );
  XNOR U6544 ( .A(n5335), .B(n5334), .Z(n5336) );
  XNOR U6545 ( .A(n5336), .B(n5337), .Z(n6222) );
  XNOR U6546 ( .A(n6221), .B(n6222), .Z(n6223) );
  NANDN U6547 ( .A(n1593), .B(n1592), .Z(n1597) );
  NAND U6548 ( .A(n1595), .B(n1594), .Z(n1596) );
  NAND U6549 ( .A(n1597), .B(n1596), .Z(n6224) );
  XOR U6550 ( .A(n6223), .B(n6224), .Z(n5501) );
  OR U6551 ( .A(n1599), .B(n1598), .Z(n1603) );
  NANDN U6552 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U6553 ( .A(n1603), .B(n1602), .Z(n6529) );
  OR U6554 ( .A(n1605), .B(n1604), .Z(n1609) );
  NANDN U6555 ( .A(n1607), .B(n1606), .Z(n1608) );
  AND U6556 ( .A(n1609), .B(n1608), .Z(n6528) );
  XNOR U6557 ( .A(n6529), .B(n6528), .Z(n6530) );
  XOR U6558 ( .A(n6530), .B(n6531), .Z(n5944) );
  OR U6559 ( .A(n1615), .B(n1614), .Z(n1619) );
  NANDN U6560 ( .A(n1617), .B(n1616), .Z(n1618) );
  NAND U6561 ( .A(n1619), .B(n1618), .Z(n6523) );
  XNOR U6562 ( .A(n6523), .B(n6522), .Z(n6524) );
  OR U6563 ( .A(n1625), .B(n1624), .Z(n1629) );
  NANDN U6564 ( .A(n1627), .B(n1626), .Z(n1628) );
  NAND U6565 ( .A(n1629), .B(n1628), .Z(n6525) );
  XOR U6566 ( .A(n6524), .B(n6525), .Z(n5941) );
  OR U6567 ( .A(n1631), .B(n1630), .Z(n1635) );
  NANDN U6568 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U6569 ( .A(n1635), .B(n1634), .Z(n7042) );
  XNOR U6570 ( .A(n7042), .B(n7041), .Z(n7043) );
  XNOR U6571 ( .A(n7043), .B(n7044), .Z(n5942) );
  XNOR U6572 ( .A(n5941), .B(n5942), .Z(n5943) );
  XNOR U6573 ( .A(n5944), .B(n5943), .Z(n5498) );
  NANDN U6574 ( .A(n1645), .B(n1644), .Z(n1649) );
  OR U6575 ( .A(n1647), .B(n1646), .Z(n1648) );
  AND U6576 ( .A(n1649), .B(n1648), .Z(n5499) );
  XNOR U6577 ( .A(n5498), .B(n5499), .Z(n5500) );
  XNOR U6578 ( .A(n5501), .B(n5500), .Z(n7261) );
  XNOR U6579 ( .A(n7260), .B(n7261), .Z(n7262) );
  XNOR U6580 ( .A(n7263), .B(n7262), .Z(n5180) );
  OR U6581 ( .A(n1651), .B(n1650), .Z(n1655) );
  NANDN U6582 ( .A(n1653), .B(n1652), .Z(n1654) );
  NAND U6583 ( .A(n1655), .B(n1654), .Z(n5239) );
  OR U6584 ( .A(n1657), .B(n1656), .Z(n1661) );
  NANDN U6585 ( .A(n1659), .B(n1658), .Z(n1660) );
  AND U6586 ( .A(n1661), .B(n1660), .Z(n5238) );
  XNOR U6587 ( .A(n5239), .B(n5238), .Z(n5240) );
  OR U6588 ( .A(n1663), .B(n1662), .Z(n1667) );
  NANDN U6589 ( .A(n1665), .B(n1664), .Z(n1666) );
  NAND U6590 ( .A(n1667), .B(n1666), .Z(n5241) );
  XOR U6591 ( .A(n5240), .B(n5241), .Z(n5402) );
  OR U6592 ( .A(n1669), .B(n1668), .Z(n1673) );
  NAND U6593 ( .A(n1671), .B(n1670), .Z(n1672) );
  NAND U6594 ( .A(n1673), .B(n1672), .Z(n5403) );
  XNOR U6595 ( .A(n5402), .B(n5403), .Z(n5404) );
  NANDN U6596 ( .A(n1675), .B(n1674), .Z(n1679) );
  NAND U6597 ( .A(n1677), .B(n1676), .Z(n1678) );
  AND U6598 ( .A(n1679), .B(n1678), .Z(n5405) );
  XNOR U6599 ( .A(n5404), .B(n5405), .Z(n5588) );
  NANDN U6600 ( .A(n1681), .B(n1680), .Z(n1685) );
  NAND U6601 ( .A(n1683), .B(n1682), .Z(n1684) );
  NAND U6602 ( .A(n1685), .B(n1684), .Z(n7221) );
  OR U6603 ( .A(n1691), .B(n1690), .Z(n1695) );
  NANDN U6604 ( .A(n1693), .B(n1692), .Z(n1694) );
  AND U6605 ( .A(n1695), .B(n1694), .Z(n5208) );
  XNOR U6606 ( .A(n5209), .B(n5208), .Z(n5210) );
  XOR U6607 ( .A(n5210), .B(n5211), .Z(n7218) );
  NANDN U6608 ( .A(n1701), .B(n1700), .Z(n1705) );
  NAND U6609 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U6610 ( .A(n1705), .B(n1704), .Z(n7219) );
  XNOR U6611 ( .A(n7218), .B(n7219), .Z(n7220) );
  XOR U6612 ( .A(n7221), .B(n7220), .Z(n5589) );
  XOR U6613 ( .A(n5588), .B(n5589), .Z(n5590) );
  OR U6614 ( .A(n1707), .B(n1706), .Z(n1711) );
  NANDN U6615 ( .A(n1709), .B(n1708), .Z(n1710) );
  NAND U6616 ( .A(n1711), .B(n1710), .Z(n6294) );
  XNOR U6617 ( .A(n6294), .B(n6293), .Z(n6295) );
  XOR U6618 ( .A(n6295), .B(n6296), .Z(n6278) );
  XOR U6619 ( .A(n5312), .B(n5313), .Z(n6275) );
  NANDN U6620 ( .A(n1733), .B(n1732), .Z(n1737) );
  NAND U6621 ( .A(n1735), .B(n1734), .Z(n1736) );
  NAND U6622 ( .A(n1737), .B(n1736), .Z(n6276) );
  XNOR U6623 ( .A(n6275), .B(n6276), .Z(n6277) );
  XNOR U6624 ( .A(n6278), .B(n6277), .Z(n5591) );
  XOR U6625 ( .A(n5590), .B(n5591), .Z(n6861) );
  OR U6626 ( .A(n1747), .B(n1746), .Z(n1751) );
  OR U6627 ( .A(n1749), .B(n1748), .Z(n1750) );
  NAND U6628 ( .A(n1751), .B(n1750), .Z(n5518) );
  OR U6629 ( .A(n1753), .B(n1752), .Z(n1757) );
  OR U6630 ( .A(n1755), .B(n1754), .Z(n1756) );
  AND U6631 ( .A(n1757), .B(n1756), .Z(n5519) );
  XNOR U6632 ( .A(n5518), .B(n5519), .Z(n5520) );
  XNOR U6633 ( .A(n5521), .B(n5520), .Z(n5618) );
  XNOR U6634 ( .A(n5619), .B(n5618), .Z(n5620) );
  NANDN U6635 ( .A(n1759), .B(n1758), .Z(n1763) );
  NAND U6636 ( .A(n1761), .B(n1760), .Z(n1762) );
  NAND U6637 ( .A(n1763), .B(n1762), .Z(n5621) );
  XOR U6638 ( .A(n5620), .B(n5621), .Z(n6046) );
  NANDN U6639 ( .A(n1765), .B(n1764), .Z(n1769) );
  NAND U6640 ( .A(n1767), .B(n1766), .Z(n1768) );
  NAND U6641 ( .A(n1769), .B(n1768), .Z(n5381) );
  XNOR U6642 ( .A(n5233), .B(n5232), .Z(n5234) );
  XNOR U6643 ( .A(n5234), .B(n5235), .Z(n5378) );
  OR U6644 ( .A(n1783), .B(n1782), .Z(n1787) );
  NANDN U6645 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U6646 ( .A(n1787), .B(n1786), .Z(n5379) );
  XOR U6647 ( .A(n5381), .B(n5380), .Z(n6043) );
  NANDN U6648 ( .A(n1789), .B(n1788), .Z(n1793) );
  NAND U6649 ( .A(n1791), .B(n1790), .Z(n1792) );
  NAND U6650 ( .A(n1793), .B(n1792), .Z(n6595) );
  NANDN U6651 ( .A(n1795), .B(n1794), .Z(n1799) );
  NAND U6652 ( .A(n1797), .B(n1796), .Z(n1798) );
  NAND U6653 ( .A(n1799), .B(n1798), .Z(n6594) );
  NANDN U6654 ( .A(n1801), .B(n1800), .Z(n1805) );
  NAND U6655 ( .A(n1803), .B(n1802), .Z(n1804) );
  NAND U6656 ( .A(n1805), .B(n1804), .Z(n6597) );
  XNOR U6657 ( .A(n6596), .B(n6597), .Z(n6044) );
  XNOR U6658 ( .A(n6043), .B(n6044), .Z(n6045) );
  XNOR U6659 ( .A(n6046), .B(n6045), .Z(n6859) );
  OR U6660 ( .A(n1807), .B(n1806), .Z(n1811) );
  OR U6661 ( .A(n1809), .B(n1808), .Z(n1810) );
  NAND U6662 ( .A(n1811), .B(n1810), .Z(n6192) );
  OR U6663 ( .A(n1813), .B(n1812), .Z(n1817) );
  OR U6664 ( .A(n1815), .B(n1814), .Z(n1816) );
  AND U6665 ( .A(n1817), .B(n1816), .Z(n6191) );
  XNOR U6666 ( .A(n6192), .B(n6191), .Z(n6193) );
  XOR U6667 ( .A(n6193), .B(n6194), .Z(n5229) );
  XNOR U6668 ( .A(n6160), .B(n6159), .Z(n6161) );
  XOR U6669 ( .A(n6161), .B(n6162), .Z(n5226) );
  NANDN U6670 ( .A(n1835), .B(n1834), .Z(n1839) );
  NAND U6671 ( .A(n1837), .B(n1836), .Z(n1838) );
  NAND U6672 ( .A(n1839), .B(n1838), .Z(n5227) );
  XNOR U6673 ( .A(n5226), .B(n5227), .Z(n5228) );
  XNOR U6674 ( .A(n5229), .B(n5228), .Z(n6230) );
  NANDN U6675 ( .A(n1841), .B(n1840), .Z(n1845) );
  NAND U6676 ( .A(n1843), .B(n1842), .Z(n1844) );
  NAND U6677 ( .A(n1845), .B(n1844), .Z(n5477) );
  XNOR U6678 ( .A(n6084), .B(n6083), .Z(n6085) );
  XOR U6679 ( .A(n6085), .B(n6086), .Z(n5474) );
  NANDN U6680 ( .A(n1859), .B(n1858), .Z(n1863) );
  NAND U6681 ( .A(n1861), .B(n1860), .Z(n1862) );
  NAND U6682 ( .A(n1863), .B(n1862), .Z(n5475) );
  XNOR U6683 ( .A(n5474), .B(n5475), .Z(n5476) );
  XOR U6684 ( .A(n5477), .B(n5476), .Z(n6227) );
  OR U6685 ( .A(n1865), .B(n1864), .Z(n1869) );
  NAND U6686 ( .A(n1867), .B(n1866), .Z(n1868) );
  NAND U6687 ( .A(n1869), .B(n1868), .Z(n6016) );
  XNOR U6688 ( .A(n5397), .B(n5396), .Z(n5398) );
  XOR U6689 ( .A(n5398), .B(n5399), .Z(n6013) );
  NANDN U6690 ( .A(n1883), .B(n1882), .Z(n1887) );
  NAND U6691 ( .A(n1885), .B(n1884), .Z(n1886) );
  NAND U6692 ( .A(n1887), .B(n1886), .Z(n6014) );
  XNOR U6693 ( .A(n6013), .B(n6014), .Z(n6015) );
  XNOR U6694 ( .A(n6016), .B(n6015), .Z(n6228) );
  XNOR U6695 ( .A(n6227), .B(n6228), .Z(n6229) );
  XOR U6696 ( .A(n6230), .B(n6229), .Z(n6858) );
  XNOR U6697 ( .A(n6859), .B(n6858), .Z(n6860) );
  XNOR U6698 ( .A(n6861), .B(n6860), .Z(n5181) );
  XNOR U6699 ( .A(n5180), .B(n5181), .Z(n5182) );
  XOR U6700 ( .A(n5183), .B(n5182), .Z(n6792) );
  NANDN U6701 ( .A(n1889), .B(n1888), .Z(n1893) );
  OR U6702 ( .A(n1891), .B(n1890), .Z(n1892) );
  NAND U6703 ( .A(n1893), .B(n1892), .Z(n7117) );
  XNOR U6704 ( .A(n5786), .B(n5785), .Z(n5787) );
  XOR U6705 ( .A(n5787), .B(n5788), .Z(n7161) );
  XNOR U6706 ( .A(n5269), .B(n5268), .Z(n5270) );
  XOR U6707 ( .A(n5270), .B(n5271), .Z(n7158) );
  NANDN U6708 ( .A(n1919), .B(n1918), .Z(n1923) );
  NAND U6709 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U6710 ( .A(n1923), .B(n1922), .Z(n7159) );
  XNOR U6711 ( .A(n7158), .B(n7159), .Z(n7160) );
  XNOR U6712 ( .A(n7161), .B(n7160), .Z(n7114) );
  NANDN U6713 ( .A(n1925), .B(n1924), .Z(n1929) );
  OR U6714 ( .A(n1927), .B(n1926), .Z(n1928) );
  AND U6715 ( .A(n1929), .B(n1928), .Z(n7115) );
  XNOR U6716 ( .A(n7114), .B(n7115), .Z(n7116) );
  XNOR U6717 ( .A(n7117), .B(n7116), .Z(n7170) );
  NANDN U6718 ( .A(n1931), .B(n1930), .Z(n1935) );
  NAND U6719 ( .A(n1933), .B(n1932), .Z(n1934) );
  NAND U6720 ( .A(n1935), .B(n1934), .Z(n6719) );
  OR U6721 ( .A(n1941), .B(n1940), .Z(n1945) );
  NANDN U6722 ( .A(n1943), .B(n1942), .Z(n1944) );
  NAND U6723 ( .A(n1945), .B(n1944), .Z(n5863) );
  OR U6724 ( .A(n1947), .B(n1946), .Z(n1951) );
  NANDN U6725 ( .A(n1949), .B(n1948), .Z(n1950) );
  NAND U6726 ( .A(n1951), .B(n1950), .Z(n5866) );
  XOR U6727 ( .A(n5865), .B(n5866), .Z(n6716) );
  NANDN U6728 ( .A(n1953), .B(n1952), .Z(n1957) );
  NAND U6729 ( .A(n1955), .B(n1954), .Z(n1956) );
  NAND U6730 ( .A(n1957), .B(n1956), .Z(n6717) );
  XNOR U6731 ( .A(n6716), .B(n6717), .Z(n6718) );
  XOR U6732 ( .A(n6719), .B(n6718), .Z(n5711) );
  OR U6733 ( .A(n1967), .B(n1966), .Z(n1971) );
  NANDN U6734 ( .A(n1969), .B(n1968), .Z(n1970) );
  NAND U6735 ( .A(n1971), .B(n1970), .Z(n7233) );
  XOR U6736 ( .A(n7232), .B(n7233), .Z(n6651) );
  OR U6737 ( .A(n1973), .B(n1972), .Z(n1977) );
  NANDN U6738 ( .A(n1975), .B(n1974), .Z(n1976) );
  NAND U6739 ( .A(n1977), .B(n1976), .Z(n6999) );
  XNOR U6740 ( .A(n6999), .B(n6998), .Z(n7000) );
  XNOR U6741 ( .A(n7000), .B(n7001), .Z(n6649) );
  NANDN U6742 ( .A(n1987), .B(n1986), .Z(n1991) );
  NAND U6743 ( .A(n1989), .B(n1988), .Z(n1990) );
  NAND U6744 ( .A(n1991), .B(n1990), .Z(n6650) );
  XOR U6745 ( .A(n6651), .B(n6652), .Z(n5708) );
  NANDN U6746 ( .A(n1993), .B(n1992), .Z(n1997) );
  NANDN U6747 ( .A(n1995), .B(n1994), .Z(n1996) );
  AND U6748 ( .A(n1997), .B(n1996), .Z(n5709) );
  XNOR U6749 ( .A(n5708), .B(n5709), .Z(n5710) );
  XOR U6750 ( .A(n5711), .B(n5710), .Z(n7171) );
  XOR U6751 ( .A(n7170), .B(n7171), .Z(n7172) );
  OR U6752 ( .A(n1999), .B(n1998), .Z(n2003) );
  NANDN U6753 ( .A(n2001), .B(n2000), .Z(n2002) );
  NAND U6754 ( .A(n2003), .B(n2002), .Z(n5699) );
  OR U6755 ( .A(n2005), .B(n2004), .Z(n2009) );
  NANDN U6756 ( .A(n2007), .B(n2006), .Z(n2008) );
  NAND U6757 ( .A(n2009), .B(n2008), .Z(n6336) );
  XOR U6758 ( .A(n6337), .B(n6338), .Z(n6500) );
  XNOR U6759 ( .A(n6378), .B(n6377), .Z(n6379) );
  XOR U6760 ( .A(n6379), .B(n6380), .Z(n6497) );
  OR U6761 ( .A(n2031), .B(n2030), .Z(n2035) );
  NANDN U6762 ( .A(n2033), .B(n2032), .Z(n2034) );
  NAND U6763 ( .A(n2035), .B(n2034), .Z(n6098) );
  OR U6764 ( .A(n2037), .B(n2036), .Z(n2041) );
  NANDN U6765 ( .A(n2039), .B(n2038), .Z(n2040) );
  NAND U6766 ( .A(n2041), .B(n2040), .Z(n6096) );
  XOR U6767 ( .A(n6096), .B(n6095), .Z(n6097) );
  XNOR U6768 ( .A(n6098), .B(n6097), .Z(n6498) );
  XNOR U6769 ( .A(n6497), .B(n6498), .Z(n6499) );
  XNOR U6770 ( .A(n6500), .B(n6499), .Z(n5697) );
  OR U6771 ( .A(n2047), .B(n2046), .Z(n2051) );
  NANDN U6772 ( .A(n2049), .B(n2048), .Z(n2050) );
  AND U6773 ( .A(n2051), .B(n2050), .Z(n5696) );
  XNOR U6774 ( .A(n5697), .B(n5696), .Z(n5698) );
  XOR U6775 ( .A(n5699), .B(n5698), .Z(n7173) );
  XNOR U6776 ( .A(n7172), .B(n7173), .Z(n6785) );
  OR U6777 ( .A(n2053), .B(n2052), .Z(n2057) );
  NAND U6778 ( .A(n2055), .B(n2054), .Z(n2056) );
  NAND U6779 ( .A(n2057), .B(n2056), .Z(n6917) );
  NANDN U6780 ( .A(n2059), .B(n2058), .Z(n2063) );
  NAND U6781 ( .A(n2061), .B(n2060), .Z(n2062) );
  AND U6782 ( .A(n2063), .B(n2062), .Z(n6916) );
  XNOR U6783 ( .A(n6917), .B(n6916), .Z(n6918) );
  OR U6784 ( .A(n2065), .B(n2064), .Z(n2069) );
  NANDN U6785 ( .A(n2067), .B(n2066), .Z(n2068) );
  NAND U6786 ( .A(n2069), .B(n2068), .Z(n6919) );
  XOR U6787 ( .A(n6918), .B(n6919), .Z(n7139) );
  OR U6788 ( .A(n2071), .B(n2070), .Z(n2075) );
  NAND U6789 ( .A(n2073), .B(n2072), .Z(n2074) );
  NAND U6790 ( .A(n2075), .B(n2074), .Z(n7185) );
  OR U6791 ( .A(n2077), .B(n2076), .Z(n2081) );
  NAND U6792 ( .A(n2079), .B(n2078), .Z(n2080) );
  NAND U6793 ( .A(n2081), .B(n2080), .Z(n7183) );
  NANDN U6794 ( .A(n2083), .B(n2082), .Z(n2087) );
  NAND U6795 ( .A(n2085), .B(n2084), .Z(n2086) );
  AND U6796 ( .A(n2087), .B(n2086), .Z(n7182) );
  XNOR U6797 ( .A(n7183), .B(n7182), .Z(n7184) );
  XOR U6798 ( .A(n7185), .B(n7184), .Z(n7136) );
  NANDN U6799 ( .A(n2089), .B(n2088), .Z(n2093) );
  NANDN U6800 ( .A(n2091), .B(n2090), .Z(n2092) );
  NAND U6801 ( .A(n2093), .B(n2092), .Z(n7177) );
  OR U6802 ( .A(n2095), .B(n2094), .Z(n2099) );
  NANDN U6803 ( .A(n2097), .B(n2096), .Z(n2098) );
  AND U6804 ( .A(n2099), .B(n2098), .Z(n7176) );
  XNOR U6805 ( .A(n7177), .B(n7176), .Z(n7178) );
  OR U6806 ( .A(n2101), .B(n2100), .Z(n2105) );
  NANDN U6807 ( .A(n2103), .B(n2102), .Z(n2104) );
  NAND U6808 ( .A(n2105), .B(n2104), .Z(n7179) );
  XNOR U6809 ( .A(n7178), .B(n7179), .Z(n7137) );
  XNOR U6810 ( .A(n7136), .B(n7137), .Z(n7138) );
  XNOR U6811 ( .A(n7139), .B(n7138), .Z(n6503) );
  NANDN U6812 ( .A(n2107), .B(n2106), .Z(n2111) );
  OR U6813 ( .A(n2109), .B(n2108), .Z(n2110) );
  NAND U6814 ( .A(n2111), .B(n2110), .Z(n5695) );
  OR U6815 ( .A(n2113), .B(n2112), .Z(n2117) );
  NANDN U6816 ( .A(n2115), .B(n2114), .Z(n2116) );
  NAND U6817 ( .A(n2117), .B(n2116), .Z(n6601) );
  OR U6818 ( .A(n2119), .B(n2118), .Z(n2123) );
  NANDN U6819 ( .A(n2121), .B(n2120), .Z(n2122) );
  NAND U6820 ( .A(n2123), .B(n2122), .Z(n6600) );
  OR U6821 ( .A(n2125), .B(n2124), .Z(n2129) );
  NANDN U6822 ( .A(n2127), .B(n2126), .Z(n2128) );
  NAND U6823 ( .A(n2129), .B(n2128), .Z(n6603) );
  XOR U6824 ( .A(n6602), .B(n6603), .Z(n5368) );
  OR U6825 ( .A(n2131), .B(n2130), .Z(n2135) );
  NANDN U6826 ( .A(n2133), .B(n2132), .Z(n2134) );
  NAND U6827 ( .A(n2135), .B(n2134), .Z(n5203) );
  OR U6828 ( .A(n2137), .B(n2136), .Z(n2141) );
  NANDN U6829 ( .A(n2139), .B(n2138), .Z(n2140) );
  AND U6830 ( .A(n2141), .B(n2140), .Z(n5202) );
  XNOR U6831 ( .A(n5203), .B(n5202), .Z(n5204) );
  OR U6832 ( .A(n2143), .B(n2142), .Z(n2147) );
  NANDN U6833 ( .A(n2145), .B(n2144), .Z(n2146) );
  NAND U6834 ( .A(n2147), .B(n2146), .Z(n5205) );
  XOR U6835 ( .A(n5204), .B(n5205), .Z(n5365) );
  OR U6836 ( .A(n2149), .B(n2148), .Z(n2153) );
  NANDN U6837 ( .A(n2151), .B(n2150), .Z(n2152) );
  NAND U6838 ( .A(n2153), .B(n2152), .Z(n5366) );
  XNOR U6839 ( .A(n5365), .B(n5366), .Z(n5367) );
  XNOR U6840 ( .A(n5368), .B(n5367), .Z(n5692) );
  NANDN U6841 ( .A(n2155), .B(n2154), .Z(n2159) );
  OR U6842 ( .A(n2157), .B(n2156), .Z(n2158) );
  AND U6843 ( .A(n2159), .B(n2158), .Z(n5693) );
  XNOR U6844 ( .A(n5692), .B(n5693), .Z(n5694) );
  XNOR U6845 ( .A(n5695), .B(n5694), .Z(n6504) );
  XOR U6846 ( .A(n6503), .B(n6504), .Z(n6505) );
  NANDN U6847 ( .A(n2161), .B(n2160), .Z(n2165) );
  OR U6848 ( .A(n2163), .B(n2162), .Z(n2164) );
  NAND U6849 ( .A(n2165), .B(n2164), .Z(n5659) );
  XNOR U6850 ( .A(n6056), .B(n6055), .Z(n6057) );
  XNOR U6851 ( .A(n6057), .B(n6058), .Z(n5374) );
  OR U6852 ( .A(n2179), .B(n2178), .Z(n2183) );
  NANDN U6853 ( .A(n2181), .B(n2180), .Z(n2182) );
  NAND U6854 ( .A(n2183), .B(n2182), .Z(n6987) );
  OR U6855 ( .A(n2185), .B(n2184), .Z(n2189) );
  NANDN U6856 ( .A(n2187), .B(n2186), .Z(n2188) );
  NAND U6857 ( .A(n2189), .B(n2188), .Z(n6986) );
  OR U6858 ( .A(n2191), .B(n2190), .Z(n2195) );
  NANDN U6859 ( .A(n2193), .B(n2192), .Z(n2194) );
  NAND U6860 ( .A(n2195), .B(n2194), .Z(n6989) );
  XOR U6861 ( .A(n6988), .B(n6989), .Z(n5371) );
  OR U6862 ( .A(n2197), .B(n2196), .Z(n2201) );
  NANDN U6863 ( .A(n2199), .B(n2198), .Z(n2200) );
  NAND U6864 ( .A(n2201), .B(n2200), .Z(n5372) );
  XNOR U6865 ( .A(n5371), .B(n5372), .Z(n5373) );
  XNOR U6866 ( .A(n5374), .B(n5373), .Z(n5657) );
  NANDN U6867 ( .A(n2203), .B(n2202), .Z(n2207) );
  OR U6868 ( .A(n2205), .B(n2204), .Z(n2206) );
  AND U6869 ( .A(n2207), .B(n2206), .Z(n5656) );
  XOR U6870 ( .A(n5657), .B(n5656), .Z(n5658) );
  XOR U6871 ( .A(n5659), .B(n5658), .Z(n6506) );
  XOR U6872 ( .A(n6505), .B(n6506), .Z(n6782) );
  NANDN U6873 ( .A(n2209), .B(n2208), .Z(n2213) );
  OR U6874 ( .A(n2211), .B(n2210), .Z(n2212) );
  NAND U6875 ( .A(n2213), .B(n2212), .Z(n4979) );
  NANDN U6876 ( .A(n2215), .B(n2214), .Z(n2219) );
  NAND U6877 ( .A(n2217), .B(n2216), .Z(n2218) );
  NAND U6878 ( .A(n2219), .B(n2218), .Z(n7167) );
  NANDN U6879 ( .A(n2221), .B(n2220), .Z(n2225) );
  NAND U6880 ( .A(n2223), .B(n2222), .Z(n2224) );
  NAND U6881 ( .A(n2225), .B(n2224), .Z(n7165) );
  NANDN U6882 ( .A(n2227), .B(n2226), .Z(n2231) );
  NAND U6883 ( .A(n2229), .B(n2228), .Z(n2230) );
  AND U6884 ( .A(n2231), .B(n2230), .Z(n7164) );
  XNOR U6885 ( .A(n7165), .B(n7164), .Z(n7166) );
  XNOR U6886 ( .A(n7167), .B(n7166), .Z(n4976) );
  XNOR U6887 ( .A(n6090), .B(n6089), .Z(n6091) );
  XOR U6888 ( .A(n6091), .B(n6092), .Z(n6513) );
  XNOR U6889 ( .A(n6060), .B(n6059), .Z(n6061) );
  XNOR U6890 ( .A(n6062), .B(n6061), .Z(n6510) );
  XOR U6891 ( .A(n6510), .B(n6511), .Z(n6512) );
  XOR U6892 ( .A(n6513), .B(n6512), .Z(n4977) );
  XOR U6893 ( .A(n4976), .B(n4977), .Z(n4978) );
  XOR U6894 ( .A(n4979), .B(n4978), .Z(n6740) );
  OR U6895 ( .A(n2261), .B(n2260), .Z(n2265) );
  NANDN U6896 ( .A(n2263), .B(n2262), .Z(n2264) );
  NAND U6897 ( .A(n2265), .B(n2264), .Z(n6326) );
  XNOR U6898 ( .A(n6390), .B(n6389), .Z(n6391) );
  XOR U6899 ( .A(n6391), .B(n6392), .Z(n6323) );
  OR U6900 ( .A(n2279), .B(n2278), .Z(n2283) );
  NAND U6901 ( .A(n2281), .B(n2280), .Z(n2282) );
  NAND U6902 ( .A(n2283), .B(n2282), .Z(n6324) );
  XNOR U6903 ( .A(n6323), .B(n6324), .Z(n6325) );
  XNOR U6904 ( .A(n6326), .B(n6325), .Z(n5652) );
  XNOR U6905 ( .A(n7005), .B(n7004), .Z(n7006) );
  OR U6906 ( .A(n2293), .B(n2292), .Z(n2297) );
  NANDN U6907 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U6908 ( .A(n2297), .B(n2296), .Z(n7007) );
  XOR U6909 ( .A(n7006), .B(n7007), .Z(n5854) );
  XNOR U6910 ( .A(n6420), .B(n6419), .Z(n6421) );
  XOR U6911 ( .A(n6421), .B(n6422), .Z(n5851) );
  OR U6912 ( .A(n2311), .B(n2310), .Z(n2315) );
  NAND U6913 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U6914 ( .A(n2315), .B(n2314), .Z(n5852) );
  XNOR U6915 ( .A(n5851), .B(n5852), .Z(n5853) );
  XOR U6916 ( .A(n5854), .B(n5853), .Z(n5653) );
  XOR U6917 ( .A(n5652), .B(n5653), .Z(n5654) );
  OR U6918 ( .A(n2317), .B(n2316), .Z(n2321) );
  NANDN U6919 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U6920 ( .A(n2321), .B(n2320), .Z(n7011) );
  XNOR U6921 ( .A(n7011), .B(n7010), .Z(n7012) );
  XOR U6922 ( .A(n7012), .B(n7013), .Z(n5875) );
  OR U6923 ( .A(n2331), .B(n2330), .Z(n2335) );
  NANDN U6924 ( .A(n2333), .B(n2332), .Z(n2334) );
  NAND U6925 ( .A(n2335), .B(n2334), .Z(n6434) );
  XNOR U6926 ( .A(n6431), .B(n6432), .Z(n6433) );
  XNOR U6927 ( .A(n6434), .B(n6433), .Z(n5876) );
  XNOR U6928 ( .A(n5875), .B(n5876), .Z(n5877) );
  XNOR U6929 ( .A(n6467), .B(n6468), .Z(n6469) );
  XOR U6930 ( .A(n6470), .B(n6469), .Z(n5878) );
  XOR U6931 ( .A(n5877), .B(n5878), .Z(n5655) );
  XOR U6932 ( .A(n5654), .B(n5655), .Z(n6741) );
  XNOR U6933 ( .A(n6740), .B(n6741), .Z(n6742) );
  OR U6934 ( .A(n2361), .B(n2360), .Z(n2365) );
  NANDN U6935 ( .A(n2363), .B(n2362), .Z(n2364) );
  AND U6936 ( .A(n2365), .B(n2364), .Z(n6661) );
  XNOR U6937 ( .A(n6662), .B(n6661), .Z(n6663) );
  OR U6938 ( .A(n2367), .B(n2366), .Z(n2371) );
  NANDN U6939 ( .A(n2369), .B(n2368), .Z(n2370) );
  NAND U6940 ( .A(n2371), .B(n2370), .Z(n6664) );
  XOR U6941 ( .A(n6663), .B(n6664), .Z(n6350) );
  OR U6942 ( .A(n2373), .B(n2372), .Z(n2377) );
  NANDN U6943 ( .A(n2375), .B(n2374), .Z(n2376) );
  NAND U6944 ( .A(n2377), .B(n2376), .Z(n6565) );
  OR U6945 ( .A(n2379), .B(n2378), .Z(n2383) );
  NANDN U6946 ( .A(n2381), .B(n2380), .Z(n2382) );
  AND U6947 ( .A(n2383), .B(n2382), .Z(n6564) );
  XNOR U6948 ( .A(n6565), .B(n6564), .Z(n6566) );
  XOR U6949 ( .A(n6566), .B(n6567), .Z(n6347) );
  OR U6950 ( .A(n2389), .B(n2388), .Z(n2393) );
  NANDN U6951 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U6952 ( .A(n2393), .B(n2392), .Z(n6132) );
  XNOR U6953 ( .A(n6132), .B(n6131), .Z(n6133) );
  XNOR U6954 ( .A(n6133), .B(n6134), .Z(n6348) );
  XNOR U6955 ( .A(n6347), .B(n6348), .Z(n6349) );
  XNOR U6956 ( .A(n6350), .B(n6349), .Z(n5665) );
  OR U6957 ( .A(n2407), .B(n2406), .Z(n2411) );
  OR U6958 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U6959 ( .A(n2411), .B(n2410), .Z(n5511) );
  XNOR U6960 ( .A(n5511), .B(n5510), .Z(n5512) );
  XNOR U6961 ( .A(n5513), .B(n5512), .Z(n5881) );
  XNOR U6962 ( .A(n6643), .B(n6644), .Z(n6645) );
  XNOR U6963 ( .A(n6646), .B(n6645), .Z(n5882) );
  XOR U6964 ( .A(n5881), .B(n5882), .Z(n5883) );
  OR U6965 ( .A(n2429), .B(n2428), .Z(n2433) );
  NANDN U6966 ( .A(n2431), .B(n2430), .Z(n2432) );
  NAND U6967 ( .A(n2433), .B(n2432), .Z(n6482) );
  XNOR U6968 ( .A(n6479), .B(n6480), .Z(n6481) );
  XNOR U6969 ( .A(n6482), .B(n6481), .Z(n5884) );
  XOR U6970 ( .A(n5883), .B(n5884), .Z(n5662) );
  OR U6971 ( .A(n2443), .B(n2442), .Z(n2447) );
  NANDN U6972 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U6973 ( .A(n2447), .B(n2446), .Z(n6102) );
  OR U6974 ( .A(n2449), .B(n2448), .Z(n2453) );
  NANDN U6975 ( .A(n2451), .B(n2450), .Z(n2452) );
  AND U6976 ( .A(n2453), .B(n2452), .Z(n6101) );
  XNOR U6977 ( .A(n6102), .B(n6101), .Z(n6103) );
  OR U6978 ( .A(n2455), .B(n2454), .Z(n2459) );
  NANDN U6979 ( .A(n2457), .B(n2456), .Z(n2458) );
  NAND U6980 ( .A(n2459), .B(n2458), .Z(n6104) );
  XOR U6981 ( .A(n6103), .B(n6104), .Z(n5905) );
  OR U6982 ( .A(n2461), .B(n2460), .Z(n2465) );
  NANDN U6983 ( .A(n2463), .B(n2462), .Z(n2464) );
  NAND U6984 ( .A(n2465), .B(n2464), .Z(n6688) );
  XNOR U6985 ( .A(n6685), .B(n6686), .Z(n6687) );
  XNOR U6986 ( .A(n6688), .B(n6687), .Z(n5906) );
  XNOR U6987 ( .A(n5905), .B(n5906), .Z(n5907) );
  XNOR U6988 ( .A(n6722), .B(n6723), .Z(n6724) );
  XNOR U6989 ( .A(n6725), .B(n6724), .Z(n5908) );
  XNOR U6990 ( .A(n5907), .B(n5908), .Z(n5663) );
  XNOR U6991 ( .A(n5662), .B(n5663), .Z(n5664) );
  XOR U6992 ( .A(n5665), .B(n5664), .Z(n6743) );
  XOR U6993 ( .A(n6742), .B(n6743), .Z(n6783) );
  XOR U6994 ( .A(n6782), .B(n6783), .Z(n6784) );
  XOR U6995 ( .A(n6785), .B(n6784), .Z(n6793) );
  XNOR U6996 ( .A(n6792), .B(n6793), .Z(n6794) );
  XOR U6997 ( .A(n6795), .B(n6794), .Z(n6889) );
  OR U6998 ( .A(n2491), .B(n2490), .Z(n2495) );
  NANDN U6999 ( .A(n2493), .B(n2492), .Z(n2494) );
  AND U7000 ( .A(n2495), .B(n2494), .Z(n5540) );
  XNOR U7001 ( .A(n5541), .B(n5540), .Z(n5542) );
  XOR U7002 ( .A(n5542), .B(n5543), .Z(n6197) );
  NANDN U7003 ( .A(n2501), .B(n2500), .Z(n2505) );
  NAND U7004 ( .A(n2503), .B(n2502), .Z(n2504) );
  NAND U7005 ( .A(n2505), .B(n2504), .Z(n6198) );
  XNOR U7006 ( .A(n6197), .B(n6198), .Z(n6199) );
  NANDN U7007 ( .A(n2507), .B(n2506), .Z(n2511) );
  NAND U7008 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U7009 ( .A(n2511), .B(n2510), .Z(n6200) );
  XNOR U7010 ( .A(n6199), .B(n6200), .Z(n7147) );
  OR U7011 ( .A(n2513), .B(n2512), .Z(n2517) );
  NANDN U7012 ( .A(n2515), .B(n2514), .Z(n2516) );
  NAND U7013 ( .A(n2517), .B(n2516), .Z(n5481) );
  OR U7014 ( .A(n2519), .B(n2518), .Z(n2523) );
  NANDN U7015 ( .A(n2521), .B(n2520), .Z(n2522) );
  AND U7016 ( .A(n2523), .B(n2522), .Z(n5480) );
  XNOR U7017 ( .A(n5481), .B(n5480), .Z(n5482) );
  OR U7018 ( .A(n2525), .B(n2524), .Z(n2529) );
  NANDN U7019 ( .A(n2527), .B(n2526), .Z(n2528) );
  NAND U7020 ( .A(n2529), .B(n2528), .Z(n5483) );
  XNOR U7021 ( .A(n5482), .B(n5483), .Z(n5594) );
  NANDN U7022 ( .A(n2531), .B(n2530), .Z(n2535) );
  NANDN U7023 ( .A(n2533), .B(n2532), .Z(n2534) );
  AND U7024 ( .A(n2535), .B(n2534), .Z(n5595) );
  OR U7025 ( .A(n2541), .B(n2540), .Z(n2545) );
  OR U7026 ( .A(n2543), .B(n2542), .Z(n2544) );
  AND U7027 ( .A(n2545), .B(n2544), .Z(n5816) );
  XNOR U7028 ( .A(n5815), .B(n5816), .Z(n5817) );
  OR U7029 ( .A(n2547), .B(n2546), .Z(n2551) );
  NANDN U7030 ( .A(n2549), .B(n2548), .Z(n2550) );
  AND U7031 ( .A(n2551), .B(n2550), .Z(n5818) );
  XNOR U7032 ( .A(n5817), .B(n5818), .Z(n5596) );
  XOR U7033 ( .A(n7147), .B(n7146), .Z(n7149) );
  OR U7034 ( .A(n2553), .B(n2552), .Z(n2557) );
  NANDN U7035 ( .A(n2555), .B(n2554), .Z(n2556) );
  NAND U7036 ( .A(n2557), .B(n2556), .Z(n6032) );
  OR U7037 ( .A(n2559), .B(n2558), .Z(n2563) );
  NANDN U7038 ( .A(n2561), .B(n2560), .Z(n2562) );
  AND U7039 ( .A(n2563), .B(n2562), .Z(n6031) );
  XNOR U7040 ( .A(n6032), .B(n6031), .Z(n6033) );
  OR U7041 ( .A(n2565), .B(n2564), .Z(n2569) );
  NANDN U7042 ( .A(n2567), .B(n2566), .Z(n2568) );
  NAND U7043 ( .A(n2569), .B(n2568), .Z(n6034) );
  XOR U7044 ( .A(n6033), .B(n6034), .Z(n6621) );
  OR U7045 ( .A(n2571), .B(n2570), .Z(n2575) );
  NANDN U7046 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U7047 ( .A(n2575), .B(n2574), .Z(n5984) );
  OR U7048 ( .A(n2577), .B(n2576), .Z(n2581) );
  NANDN U7049 ( .A(n2579), .B(n2578), .Z(n2580) );
  AND U7050 ( .A(n2581), .B(n2580), .Z(n5983) );
  XNOR U7051 ( .A(n5984), .B(n5983), .Z(n5985) );
  OR U7052 ( .A(n2583), .B(n2582), .Z(n2587) );
  NANDN U7053 ( .A(n2585), .B(n2584), .Z(n2586) );
  NAND U7054 ( .A(n2587), .B(n2586), .Z(n5986) );
  XNOR U7055 ( .A(n5985), .B(n5986), .Z(n6618) );
  OR U7056 ( .A(n2589), .B(n2588), .Z(n2593) );
  NANDN U7057 ( .A(n2591), .B(n2590), .Z(n2592) );
  NAND U7058 ( .A(n2593), .B(n2592), .Z(n6619) );
  XNOR U7059 ( .A(n6621), .B(n6620), .Z(n7148) );
  XNOR U7060 ( .A(n7149), .B(n7148), .Z(n5179) );
  NANDN U7061 ( .A(n2595), .B(n2594), .Z(n2599) );
  NAND U7062 ( .A(n2597), .B(n2596), .Z(n2598) );
  NAND U7063 ( .A(n2599), .B(n2598), .Z(n5177) );
  NANDN U7064 ( .A(n2601), .B(n2600), .Z(n2605) );
  NAND U7065 ( .A(n2603), .B(n2602), .Z(n2604) );
  NAND U7066 ( .A(n2605), .B(n2604), .Z(n7215) );
  NANDN U7067 ( .A(n2607), .B(n2606), .Z(n2611) );
  NAND U7068 ( .A(n2609), .B(n2608), .Z(n2610) );
  NAND U7069 ( .A(n2611), .B(n2610), .Z(n7213) );
  NANDN U7070 ( .A(n2613), .B(n2612), .Z(n2617) );
  NAND U7071 ( .A(n2615), .B(n2614), .Z(n2616) );
  AND U7072 ( .A(n2617), .B(n2616), .Z(n7212) );
  XNOR U7073 ( .A(n7213), .B(n7212), .Z(n7214) );
  XOR U7074 ( .A(n7215), .B(n7214), .Z(n6947) );
  NANDN U7075 ( .A(n2619), .B(n2618), .Z(n2623) );
  NAND U7076 ( .A(n2621), .B(n2620), .Z(n2622) );
  NAND U7077 ( .A(n2623), .B(n2622), .Z(n7203) );
  NANDN U7078 ( .A(n2625), .B(n2624), .Z(n2629) );
  NAND U7079 ( .A(n2627), .B(n2626), .Z(n2628) );
  NAND U7080 ( .A(n2629), .B(n2628), .Z(n7201) );
  NANDN U7081 ( .A(n2631), .B(n2630), .Z(n2635) );
  NAND U7082 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U7083 ( .A(n2635), .B(n2634), .Z(n7200) );
  XNOR U7084 ( .A(n7201), .B(n7200), .Z(n7202) );
  XOR U7085 ( .A(n7203), .B(n7202), .Z(n6944) );
  NANDN U7086 ( .A(n2637), .B(n2636), .Z(n2641) );
  NAND U7087 ( .A(n2639), .B(n2638), .Z(n2640) );
  NAND U7088 ( .A(n2641), .B(n2640), .Z(n7195) );
  NANDN U7089 ( .A(n2643), .B(n2642), .Z(n2647) );
  NAND U7090 ( .A(n2645), .B(n2644), .Z(n2646) );
  AND U7091 ( .A(n2647), .B(n2646), .Z(n7194) );
  XNOR U7092 ( .A(n7195), .B(n7194), .Z(n7196) );
  NANDN U7093 ( .A(n2649), .B(n2648), .Z(n2653) );
  NAND U7094 ( .A(n2651), .B(n2650), .Z(n2652) );
  NAND U7095 ( .A(n2653), .B(n2652), .Z(n7197) );
  XNOR U7096 ( .A(n7196), .B(n7197), .Z(n6945) );
  XNOR U7097 ( .A(n6944), .B(n6945), .Z(n6946) );
  XOR U7098 ( .A(n6947), .B(n6946), .Z(n5176) );
  XNOR U7099 ( .A(n5177), .B(n5176), .Z(n5178) );
  XNOR U7100 ( .A(n5179), .B(n5178), .Z(n5100) );
  NANDN U7101 ( .A(n2655), .B(n2654), .Z(n2659) );
  OR U7102 ( .A(n2657), .B(n2656), .Z(n2658) );
  AND U7103 ( .A(n2659), .B(n2658), .Z(n5101) );
  XOR U7104 ( .A(n5100), .B(n5101), .Z(n5103) );
  NANDN U7105 ( .A(n2661), .B(n2660), .Z(n2665) );
  NAND U7106 ( .A(n2663), .B(n2662), .Z(n2664) );
  NAND U7107 ( .A(n2665), .B(n2664), .Z(n5465) );
  NANDN U7108 ( .A(n2667), .B(n2666), .Z(n2671) );
  NAND U7109 ( .A(n2669), .B(n2668), .Z(n2670) );
  NAND U7110 ( .A(n2671), .B(n2670), .Z(n5462) );
  NANDN U7111 ( .A(n2673), .B(n2672), .Z(n2677) );
  OR U7112 ( .A(n2675), .B(n2674), .Z(n2676) );
  NAND U7113 ( .A(n2677), .B(n2676), .Z(n5848) );
  OR U7114 ( .A(n2679), .B(n2678), .Z(n2683) );
  NANDN U7115 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U7116 ( .A(n2683), .B(n2682), .Z(n5583) );
  OR U7117 ( .A(n2685), .B(n2684), .Z(n2689) );
  NANDN U7118 ( .A(n2687), .B(n2686), .Z(n2688) );
  AND U7119 ( .A(n2689), .B(n2688), .Z(n5582) );
  XNOR U7120 ( .A(n5583), .B(n5582), .Z(n5584) );
  OR U7121 ( .A(n2691), .B(n2690), .Z(n2695) );
  NANDN U7122 ( .A(n2693), .B(n2692), .Z(n2694) );
  NAND U7123 ( .A(n2695), .B(n2694), .Z(n5585) );
  XOR U7124 ( .A(n5584), .B(n5585), .Z(n5007) );
  XNOR U7125 ( .A(n5159), .B(n5158), .Z(n5160) );
  XOR U7126 ( .A(n5160), .B(n5161), .Z(n5004) );
  NANDN U7127 ( .A(n2709), .B(n2708), .Z(n2713) );
  NAND U7128 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U7129 ( .A(n2713), .B(n2712), .Z(n5005) );
  XNOR U7130 ( .A(n5004), .B(n5005), .Z(n5006) );
  XNOR U7131 ( .A(n5007), .B(n5006), .Z(n5845) );
  OR U7132 ( .A(n2719), .B(n2718), .Z(n2723) );
  NANDN U7133 ( .A(n2721), .B(n2720), .Z(n2722) );
  AND U7134 ( .A(n2723), .B(n2722), .Z(n5552) );
  XNOR U7135 ( .A(n5553), .B(n5552), .Z(n5554) );
  OR U7136 ( .A(n2725), .B(n2724), .Z(n2729) );
  NANDN U7137 ( .A(n2727), .B(n2726), .Z(n2728) );
  NAND U7138 ( .A(n2729), .B(n2728), .Z(n5555) );
  XOR U7139 ( .A(n5554), .B(n5555), .Z(n6907) );
  XNOR U7140 ( .A(n5165), .B(n5164), .Z(n5166) );
  XOR U7141 ( .A(n5166), .B(n5167), .Z(n6904) );
  OR U7142 ( .A(n2747), .B(n2746), .Z(n2751) );
  NANDN U7143 ( .A(n2749), .B(n2748), .Z(n2750) );
  AND U7144 ( .A(n2751), .B(n2750), .Z(n5558) );
  XNOR U7145 ( .A(n5559), .B(n5558), .Z(n5560) );
  OR U7146 ( .A(n2753), .B(n2752), .Z(n2757) );
  NANDN U7147 ( .A(n2755), .B(n2754), .Z(n2756) );
  NAND U7148 ( .A(n2757), .B(n2756), .Z(n5561) );
  XNOR U7149 ( .A(n5560), .B(n5561), .Z(n6905) );
  XNOR U7150 ( .A(n6904), .B(n6905), .Z(n6906) );
  XOR U7151 ( .A(n6907), .B(n6906), .Z(n5846) );
  XNOR U7152 ( .A(n5845), .B(n5846), .Z(n5847) );
  XOR U7153 ( .A(n5848), .B(n5847), .Z(n5463) );
  XNOR U7154 ( .A(n5462), .B(n5463), .Z(n5464) );
  XNOR U7155 ( .A(n5465), .B(n5464), .Z(n5102) );
  XNOR U7156 ( .A(n5103), .B(n5102), .Z(n4973) );
  NANDN U7157 ( .A(n2759), .B(n2758), .Z(n2763) );
  NAND U7158 ( .A(n2761), .B(n2760), .Z(n2762) );
  NAND U7159 ( .A(n2763), .B(n2762), .Z(n5085) );
  XOR U7160 ( .A(n7067), .B(n7068), .Z(n5082) );
  NANDN U7161 ( .A(n2777), .B(n2776), .Z(n2781) );
  NAND U7162 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U7163 ( .A(n2781), .B(n2780), .Z(n5083) );
  XNOR U7164 ( .A(n5082), .B(n5083), .Z(n5084) );
  XOR U7165 ( .A(n5085), .B(n5084), .Z(n5651) );
  OR U7166 ( .A(n2783), .B(n2782), .Z(n2787) );
  NANDN U7167 ( .A(n2785), .B(n2784), .Z(n2786) );
  NAND U7168 ( .A(n2787), .B(n2786), .Z(n6981) );
  XOR U7169 ( .A(n6982), .B(n6983), .Z(n5073) );
  NANDN U7170 ( .A(n2797), .B(n2796), .Z(n2801) );
  NAND U7171 ( .A(n2799), .B(n2798), .Z(n2800) );
  NAND U7172 ( .A(n2801), .B(n2800), .Z(n5071) );
  NANDN U7173 ( .A(n2803), .B(n2802), .Z(n2807) );
  NAND U7174 ( .A(n2805), .B(n2804), .Z(n2806) );
  AND U7175 ( .A(n2807), .B(n2806), .Z(n5070) );
  XNOR U7176 ( .A(n5071), .B(n5070), .Z(n5072) );
  XNOR U7177 ( .A(n5073), .B(n5072), .Z(n5648) );
  OR U7178 ( .A(n2809), .B(n2808), .Z(n2813) );
  NANDN U7179 ( .A(n2811), .B(n2810), .Z(n2812) );
  NAND U7180 ( .A(n2813), .B(n2812), .Z(n7048) );
  OR U7181 ( .A(n2815), .B(n2814), .Z(n2819) );
  NANDN U7182 ( .A(n2817), .B(n2816), .Z(n2818) );
  AND U7183 ( .A(n2819), .B(n2818), .Z(n7047) );
  XNOR U7184 ( .A(n7048), .B(n7047), .Z(n7049) );
  OR U7185 ( .A(n2821), .B(n2820), .Z(n2825) );
  NANDN U7186 ( .A(n2823), .B(n2822), .Z(n2824) );
  NAND U7187 ( .A(n2825), .B(n2824), .Z(n7050) );
  XOR U7188 ( .A(n7049), .B(n7050), .Z(n7290) );
  NANDN U7189 ( .A(n2827), .B(n2826), .Z(n2831) );
  NANDN U7190 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U7191 ( .A(n2831), .B(n2830), .Z(n7291) );
  XNOR U7192 ( .A(n7290), .B(n7291), .Z(n7292) );
  OR U7193 ( .A(n2833), .B(n2832), .Z(n2837) );
  NAND U7194 ( .A(n2835), .B(n2834), .Z(n2836) );
  NAND U7195 ( .A(n2837), .B(n2836), .Z(n7293) );
  XNOR U7196 ( .A(n7292), .B(n7293), .Z(n5649) );
  XNOR U7197 ( .A(n5648), .B(n5649), .Z(n5650) );
  XNOR U7198 ( .A(n5651), .B(n5650), .Z(n6137) );
  NANDN U7199 ( .A(n2839), .B(n2838), .Z(n2843) );
  OR U7200 ( .A(n2841), .B(n2840), .Z(n2842) );
  NAND U7201 ( .A(n2843), .B(n2842), .Z(n6855) );
  NANDN U7202 ( .A(n2845), .B(n2844), .Z(n2849) );
  NAND U7203 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U7204 ( .A(n2849), .B(n2848), .Z(n5049) );
  XOR U7205 ( .A(n7061), .B(n7062), .Z(n5046) );
  NANDN U7206 ( .A(n2863), .B(n2862), .Z(n2867) );
  NAND U7207 ( .A(n2865), .B(n2864), .Z(n2866) );
  NAND U7208 ( .A(n2867), .B(n2866), .Z(n5047) );
  XNOR U7209 ( .A(n5046), .B(n5047), .Z(n5048) );
  XOR U7210 ( .A(n5049), .B(n5048), .Z(n6852) );
  OR U7211 ( .A(n2869), .B(n2868), .Z(n2873) );
  NANDN U7212 ( .A(n2871), .B(n2870), .Z(n2872) );
  AND U7213 ( .A(n2873), .B(n2872), .Z(n6853) );
  XNOR U7214 ( .A(n6852), .B(n6853), .Z(n6854) );
  XOR U7215 ( .A(n6855), .B(n6854), .Z(n6138) );
  XOR U7216 ( .A(n6137), .B(n6138), .Z(n6140) );
  XOR U7217 ( .A(n6657), .B(n6658), .Z(n5067) );
  XOR U7218 ( .A(n6572), .B(n6573), .Z(n5064) );
  NANDN U7219 ( .A(n2899), .B(n2898), .Z(n2903) );
  NAND U7220 ( .A(n2901), .B(n2900), .Z(n2902) );
  NAND U7221 ( .A(n2903), .B(n2902), .Z(n5065) );
  XNOR U7222 ( .A(n5064), .B(n5065), .Z(n5066) );
  XNOR U7223 ( .A(n5067), .B(n5066), .Z(n5637) );
  XNOR U7224 ( .A(n6577), .B(n6576), .Z(n6578) );
  OR U7225 ( .A(n2913), .B(n2912), .Z(n2917) );
  NANDN U7226 ( .A(n2915), .B(n2914), .Z(n2916) );
  NAND U7227 ( .A(n2917), .B(n2916), .Z(n6579) );
  XOR U7228 ( .A(n6578), .B(n6579), .Z(n7269) );
  OR U7229 ( .A(n2919), .B(n2918), .Z(n2923) );
  NANDN U7230 ( .A(n2921), .B(n2920), .Z(n2922) );
  NAND U7231 ( .A(n2923), .B(n2922), .Z(n6559) );
  OR U7232 ( .A(n2925), .B(n2924), .Z(n2929) );
  NANDN U7233 ( .A(n2927), .B(n2926), .Z(n2928) );
  AND U7234 ( .A(n2929), .B(n2928), .Z(n6558) );
  XNOR U7235 ( .A(n6559), .B(n6558), .Z(n6560) );
  OR U7236 ( .A(n2931), .B(n2930), .Z(n2935) );
  NANDN U7237 ( .A(n2933), .B(n2932), .Z(n2934) );
  NAND U7238 ( .A(n2935), .B(n2934), .Z(n6561) );
  XOR U7239 ( .A(n6560), .B(n6561), .Z(n7266) );
  OR U7240 ( .A(n2937), .B(n2936), .Z(n2941) );
  NANDN U7241 ( .A(n2939), .B(n2938), .Z(n2940) );
  NAND U7242 ( .A(n2941), .B(n2940), .Z(n7267) );
  XNOR U7243 ( .A(n7266), .B(n7267), .Z(n7268) );
  XOR U7244 ( .A(n7269), .B(n7268), .Z(n5636) );
  XNOR U7245 ( .A(n5637), .B(n5636), .Z(n5638) );
  XOR U7246 ( .A(n6669), .B(n6670), .Z(n5079) );
  OR U7247 ( .A(n2955), .B(n2954), .Z(n2959) );
  NANDN U7248 ( .A(n2957), .B(n2956), .Z(n2958) );
  NAND U7249 ( .A(n2959), .B(n2958), .Z(n6674) );
  OR U7250 ( .A(n2965), .B(n2964), .Z(n2969) );
  NANDN U7251 ( .A(n2967), .B(n2966), .Z(n2968) );
  NAND U7252 ( .A(n2969), .B(n2968), .Z(n6676) );
  XOR U7253 ( .A(n6675), .B(n6676), .Z(n5076) );
  NANDN U7254 ( .A(n2971), .B(n2970), .Z(n2975) );
  NAND U7255 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U7256 ( .A(n2975), .B(n2974), .Z(n5077) );
  XNOR U7257 ( .A(n5076), .B(n5077), .Z(n5078) );
  XOR U7258 ( .A(n5079), .B(n5078), .Z(n5639) );
  XOR U7259 ( .A(n5638), .B(n5639), .Z(n6139) );
  XOR U7260 ( .A(n6140), .B(n6139), .Z(n7257) );
  NANDN U7261 ( .A(n2977), .B(n2976), .Z(n2981) );
  NAND U7262 ( .A(n2979), .B(n2978), .Z(n2980) );
  NAND U7263 ( .A(n2981), .B(n2980), .Z(n7099) );
  OR U7264 ( .A(n2983), .B(n2982), .Z(n2987) );
  NANDN U7265 ( .A(n2985), .B(n2984), .Z(n2986) );
  NAND U7266 ( .A(n2987), .B(n2986), .Z(n5287) );
  OR U7267 ( .A(n2989), .B(n2988), .Z(n2993) );
  NANDN U7268 ( .A(n2991), .B(n2990), .Z(n2992) );
  AND U7269 ( .A(n2993), .B(n2992), .Z(n5286) );
  XNOR U7270 ( .A(n5287), .B(n5286), .Z(n5288) );
  OR U7271 ( .A(n2995), .B(n2994), .Z(n2999) );
  NANDN U7272 ( .A(n2997), .B(n2996), .Z(n2998) );
  NAND U7273 ( .A(n2999), .B(n2998), .Z(n5289) );
  XOR U7274 ( .A(n5288), .B(n5289), .Z(n7097) );
  OR U7275 ( .A(n3001), .B(n3000), .Z(n3005) );
  OR U7276 ( .A(n3003), .B(n3002), .Z(n3004) );
  AND U7277 ( .A(n3005), .B(n3004), .Z(n5822) );
  OR U7278 ( .A(n3007), .B(n3006), .Z(n3011) );
  OR U7279 ( .A(n3009), .B(n3008), .Z(n3010) );
  NAND U7280 ( .A(n3011), .B(n3010), .Z(n5819) );
  OR U7281 ( .A(n3013), .B(n3012), .Z(n3017) );
  OR U7282 ( .A(n3015), .B(n3014), .Z(n3016) );
  AND U7283 ( .A(n3017), .B(n3016), .Z(n5820) );
  XNOR U7284 ( .A(n5819), .B(n5820), .Z(n5821) );
  XNOR U7285 ( .A(n5822), .B(n5821), .Z(n7096) );
  XNOR U7286 ( .A(n7097), .B(n7096), .Z(n7098) );
  XNOR U7287 ( .A(n7099), .B(n7098), .Z(n5914) );
  XNOR U7288 ( .A(n5451), .B(n5450), .Z(n5452) );
  XOR U7289 ( .A(n5452), .B(n5453), .Z(n7090) );
  NANDN U7290 ( .A(n3031), .B(n3030), .Z(n3035) );
  NAND U7291 ( .A(n3033), .B(n3032), .Z(n3034) );
  NAND U7292 ( .A(n3035), .B(n3034), .Z(n7091) );
  XNOR U7293 ( .A(n7090), .B(n7091), .Z(n7092) );
  OR U7294 ( .A(n3037), .B(n3036), .Z(n3041) );
  NANDN U7295 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U7296 ( .A(n3041), .B(n3040), .Z(n5549) );
  OR U7297 ( .A(n3043), .B(n3042), .Z(n3047) );
  NANDN U7298 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U7299 ( .A(n3047), .B(n3046), .Z(n5546) );
  OR U7300 ( .A(n3049), .B(n3048), .Z(n3053) );
  NANDN U7301 ( .A(n3051), .B(n3050), .Z(n3052) );
  AND U7302 ( .A(n3053), .B(n3052), .Z(n5547) );
  XNOR U7303 ( .A(n5546), .B(n5547), .Z(n5548) );
  XNOR U7304 ( .A(n5549), .B(n5548), .Z(n7093) );
  XOR U7305 ( .A(n7092), .B(n7093), .Z(n5911) );
  OR U7306 ( .A(n3055), .B(n3054), .Z(n3059) );
  NANDN U7307 ( .A(n3057), .B(n3056), .Z(n3058) );
  NAND U7308 ( .A(n3059), .B(n3058), .Z(n6692) );
  OR U7309 ( .A(n3061), .B(n3060), .Z(n3065) );
  NANDN U7310 ( .A(n3063), .B(n3062), .Z(n3064) );
  AND U7311 ( .A(n3065), .B(n3064), .Z(n6691) );
  XNOR U7312 ( .A(n6692), .B(n6691), .Z(n6693) );
  OR U7313 ( .A(n3067), .B(n3066), .Z(n3071) );
  NANDN U7314 ( .A(n3069), .B(n3068), .Z(n3070) );
  NAND U7315 ( .A(n3071), .B(n3070), .Z(n6694) );
  XOR U7316 ( .A(n6693), .B(n6694), .Z(n5001) );
  OR U7317 ( .A(n3077), .B(n3076), .Z(n3081) );
  NANDN U7318 ( .A(n3079), .B(n3078), .Z(n3080) );
  AND U7319 ( .A(n3081), .B(n3080), .Z(n5514) );
  XNOR U7320 ( .A(n5515), .B(n5514), .Z(n5516) );
  OR U7321 ( .A(n3083), .B(n3082), .Z(n3087) );
  NANDN U7322 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U7323 ( .A(n3087), .B(n3086), .Z(n5517) );
  XNOR U7324 ( .A(n5516), .B(n5517), .Z(n4999) );
  OR U7325 ( .A(n3089), .B(n3088), .Z(n3093) );
  NANDN U7326 ( .A(n3091), .B(n3090), .Z(n3092) );
  NAND U7327 ( .A(n3093), .B(n3092), .Z(n5571) );
  OR U7328 ( .A(n3095), .B(n3094), .Z(n3099) );
  NANDN U7329 ( .A(n3097), .B(n3096), .Z(n3098) );
  AND U7330 ( .A(n3099), .B(n3098), .Z(n5570) );
  XNOR U7331 ( .A(n5571), .B(n5570), .Z(n5572) );
  OR U7332 ( .A(n3101), .B(n3100), .Z(n3105) );
  NANDN U7333 ( .A(n3103), .B(n3102), .Z(n3104) );
  NAND U7334 ( .A(n3105), .B(n3104), .Z(n5573) );
  XNOR U7335 ( .A(n5572), .B(n5573), .Z(n4998) );
  XOR U7336 ( .A(n4999), .B(n4998), .Z(n5000) );
  XOR U7337 ( .A(n5001), .B(n5000), .Z(n5912) );
  XNOR U7338 ( .A(n5911), .B(n5912), .Z(n5913) );
  XNOR U7339 ( .A(n5914), .B(n5913), .Z(n5831) );
  OR U7340 ( .A(n3111), .B(n3110), .Z(n3115) );
  NANDN U7341 ( .A(n3113), .B(n3112), .Z(n3114) );
  NAND U7342 ( .A(n3115), .B(n3114), .Z(n5292) );
  OR U7343 ( .A(n3117), .B(n3116), .Z(n3121) );
  NANDN U7344 ( .A(n3119), .B(n3118), .Z(n3120) );
  NAND U7345 ( .A(n3121), .B(n3120), .Z(n5295) );
  XOR U7346 ( .A(n5294), .B(n5295), .Z(n5031) );
  OR U7347 ( .A(n3123), .B(n3122), .Z(n3127) );
  OR U7348 ( .A(n3125), .B(n3124), .Z(n3126) );
  NAND U7349 ( .A(n3127), .B(n3126), .Z(n5810) );
  OR U7350 ( .A(n3129), .B(n3128), .Z(n3133) );
  OR U7351 ( .A(n3131), .B(n3130), .Z(n3132) );
  NAND U7352 ( .A(n3133), .B(n3132), .Z(n5809) );
  OR U7353 ( .A(n3135), .B(n3134), .Z(n3139) );
  OR U7354 ( .A(n3137), .B(n3136), .Z(n3138) );
  NAND U7355 ( .A(n3139), .B(n3138), .Z(n5812) );
  XOR U7356 ( .A(n5811), .B(n5812), .Z(n5028) );
  XNOR U7357 ( .A(n5330), .B(n5331), .Z(n5029) );
  XNOR U7358 ( .A(n5028), .B(n5029), .Z(n5030) );
  XNOR U7359 ( .A(n5031), .B(n5030), .Z(n5423) );
  OR U7360 ( .A(n3153), .B(n3152), .Z(n3157) );
  NANDN U7361 ( .A(n3155), .B(n3154), .Z(n3156) );
  NAND U7362 ( .A(n3157), .B(n3156), .Z(n5535) );
  OR U7363 ( .A(n3159), .B(n3158), .Z(n3163) );
  NANDN U7364 ( .A(n3161), .B(n3160), .Z(n3162) );
  NAND U7365 ( .A(n3163), .B(n3162), .Z(n5534) );
  OR U7366 ( .A(n3165), .B(n3164), .Z(n3169) );
  NANDN U7367 ( .A(n3167), .B(n3166), .Z(n3168) );
  NAND U7368 ( .A(n3169), .B(n3168), .Z(n5537) );
  XOR U7369 ( .A(n5536), .B(n5537), .Z(n4992) );
  NANDN U7370 ( .A(n3171), .B(n3170), .Z(n3175) );
  NAND U7371 ( .A(n3173), .B(n3172), .Z(n3174) );
  NAND U7372 ( .A(n3175), .B(n3174), .Z(n4993) );
  XNOR U7373 ( .A(n4992), .B(n4993), .Z(n4994) );
  OR U7374 ( .A(n3177), .B(n3176), .Z(n3181) );
  NANDN U7375 ( .A(n3179), .B(n3178), .Z(n3180) );
  NAND U7376 ( .A(n3181), .B(n3180), .Z(n6218) );
  OR U7377 ( .A(n3183), .B(n3182), .Z(n3187) );
  NANDN U7378 ( .A(n3185), .B(n3184), .Z(n3186) );
  AND U7379 ( .A(n3187), .B(n3186), .Z(n6215) );
  OR U7380 ( .A(n3189), .B(n3188), .Z(n3193) );
  NANDN U7381 ( .A(n3191), .B(n3190), .Z(n3192) );
  AND U7382 ( .A(n3193), .B(n3192), .Z(n6216) );
  XNOR U7383 ( .A(n6218), .B(n6217), .Z(n4995) );
  XOR U7384 ( .A(n4994), .B(n4995), .Z(n5420) );
  OR U7385 ( .A(n3199), .B(n3198), .Z(n3203) );
  NANDN U7386 ( .A(n3201), .B(n3200), .Z(n3202) );
  NAND U7387 ( .A(n3203), .B(n3202), .Z(n6203) );
  OR U7388 ( .A(n3205), .B(n3204), .Z(n3209) );
  NANDN U7389 ( .A(n3207), .B(n3206), .Z(n3208) );
  NAND U7390 ( .A(n3209), .B(n3208), .Z(n6206) );
  XOR U7391 ( .A(n6205), .B(n6206), .Z(n4983) );
  OR U7392 ( .A(n3219), .B(n3218), .Z(n3223) );
  NANDN U7393 ( .A(n3221), .B(n3220), .Z(n3222) );
  NAND U7394 ( .A(n3223), .B(n3222), .Z(n5489) );
  XOR U7395 ( .A(n5488), .B(n5489), .Z(n4980) );
  OR U7396 ( .A(n3225), .B(n3224), .Z(n3229) );
  NANDN U7397 ( .A(n3227), .B(n3226), .Z(n3228) );
  NAND U7398 ( .A(n3229), .B(n3228), .Z(n5323) );
  OR U7399 ( .A(n3231), .B(n3230), .Z(n3235) );
  NANDN U7400 ( .A(n3233), .B(n3232), .Z(n3234) );
  NAND U7401 ( .A(n3235), .B(n3234), .Z(n5322) );
  OR U7402 ( .A(n3237), .B(n3236), .Z(n3241) );
  NANDN U7403 ( .A(n3239), .B(n3238), .Z(n3240) );
  NAND U7404 ( .A(n3241), .B(n3240), .Z(n5325) );
  XNOR U7405 ( .A(n5324), .B(n5325), .Z(n4981) );
  XNOR U7406 ( .A(n4980), .B(n4981), .Z(n4982) );
  XOR U7407 ( .A(n4983), .B(n4982), .Z(n5421) );
  XNOR U7408 ( .A(n5420), .B(n5421), .Z(n5422) );
  XNOR U7409 ( .A(n5423), .B(n5422), .Z(n5829) );
  NANDN U7410 ( .A(n3243), .B(n3242), .Z(n3247) );
  NAND U7411 ( .A(n3245), .B(n3244), .Z(n3246) );
  NAND U7412 ( .A(n3247), .B(n3246), .Z(n5037) );
  XOR U7413 ( .A(n5756), .B(n5757), .Z(n5034) );
  NANDN U7414 ( .A(n3261), .B(n3260), .Z(n3265) );
  NAND U7415 ( .A(n3263), .B(n3262), .Z(n3264) );
  NAND U7416 ( .A(n3265), .B(n3264), .Z(n5035) );
  XNOR U7417 ( .A(n5034), .B(n5035), .Z(n5036) );
  XOR U7418 ( .A(n5037), .B(n5036), .Z(n5733) );
  NANDN U7419 ( .A(n3267), .B(n3266), .Z(n3271) );
  NAND U7420 ( .A(n3269), .B(n3268), .Z(n3270) );
  NAND U7421 ( .A(n3271), .B(n3270), .Z(n5055) );
  IV U7422 ( .A(n3276), .Z(n3277) );
  OR U7423 ( .A(n3278), .B(n3277), .Z(n3282) );
  NANDN U7424 ( .A(n3280), .B(n3279), .Z(n3281) );
  NAND U7425 ( .A(n3282), .B(n3281), .Z(n5742) );
  XOR U7426 ( .A(n5744), .B(n5745), .Z(n5052) );
  NANDN U7427 ( .A(n3288), .B(n3287), .Z(n3292) );
  NAND U7428 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U7429 ( .A(n3292), .B(n3291), .Z(n5053) );
  XNOR U7430 ( .A(n5052), .B(n5053), .Z(n5054) );
  XOR U7431 ( .A(n5055), .B(n5054), .Z(n5730) );
  OR U7432 ( .A(n3298), .B(n3297), .Z(n3302) );
  NANDN U7433 ( .A(n3300), .B(n3299), .Z(n3301) );
  NAND U7434 ( .A(n3302), .B(n3301), .Z(n5196) );
  OR U7435 ( .A(n3304), .B(n3303), .Z(n3308) );
  NANDN U7436 ( .A(n3306), .B(n3305), .Z(n3307) );
  NAND U7437 ( .A(n3308), .B(n3307), .Z(n5199) );
  XOR U7438 ( .A(n5198), .B(n5199), .Z(n5025) );
  XOR U7439 ( .A(n6241), .B(n6242), .Z(n5022) );
  OR U7440 ( .A(n3322), .B(n3321), .Z(n3326) );
  NAND U7441 ( .A(n3324), .B(n3323), .Z(n3325) );
  NAND U7442 ( .A(n3326), .B(n3325), .Z(n5023) );
  XNOR U7443 ( .A(n5022), .B(n5023), .Z(n5024) );
  XOR U7444 ( .A(n5025), .B(n5024), .Z(n5731) );
  XNOR U7445 ( .A(n5730), .B(n5731), .Z(n5732) );
  XOR U7446 ( .A(n5733), .B(n5732), .Z(n5830) );
  XNOR U7447 ( .A(n5829), .B(n5830), .Z(n5832) );
  XNOR U7448 ( .A(n5831), .B(n5832), .Z(n7254) );
  NAND U7449 ( .A(n3328), .B(n3327), .Z(n3332) );
  NANDN U7450 ( .A(n3330), .B(n3329), .Z(n3331) );
  NAND U7451 ( .A(n3332), .B(n3331), .Z(n5411) );
  OR U7452 ( .A(n3342), .B(n3341), .Z(n3346) );
  NANDN U7453 ( .A(n3344), .B(n3343), .Z(n3345) );
  NAND U7454 ( .A(n3346), .B(n3345), .Z(n5349) );
  XOR U7455 ( .A(n5348), .B(n5349), .Z(n4986) );
  NANDN U7456 ( .A(n3348), .B(n3347), .Z(n3352) );
  NAND U7457 ( .A(n3350), .B(n3349), .Z(n3351) );
  NAND U7458 ( .A(n3352), .B(n3351), .Z(n4987) );
  XNOR U7459 ( .A(n4986), .B(n4987), .Z(n4988) );
  NANDN U7460 ( .A(n3354), .B(n3353), .Z(n3358) );
  NAND U7461 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U7462 ( .A(n3358), .B(n3357), .Z(n4989) );
  XNOR U7463 ( .A(n4988), .B(n4989), .Z(n5408) );
  NANDN U7464 ( .A(n3360), .B(n3359), .Z(n3364) );
  NAND U7465 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U7466 ( .A(n3364), .B(n3363), .Z(n5043) );
  OR U7467 ( .A(n3366), .B(n3365), .Z(n3370) );
  NANDN U7468 ( .A(n3368), .B(n3367), .Z(n3369) );
  NAND U7469 ( .A(n3370), .B(n3369), .Z(n5930) );
  XOR U7470 ( .A(n5931), .B(n5932), .Z(n5040) );
  NANDN U7471 ( .A(n3380), .B(n3379), .Z(n3384) );
  NAND U7472 ( .A(n3382), .B(n3381), .Z(n3383) );
  NAND U7473 ( .A(n3384), .B(n3383), .Z(n5041) );
  XNOR U7474 ( .A(n5040), .B(n5041), .Z(n5042) );
  XOR U7475 ( .A(n5043), .B(n5042), .Z(n5409) );
  XOR U7476 ( .A(n5408), .B(n5409), .Z(n5410) );
  XOR U7477 ( .A(n5411), .B(n5410), .Z(n5531) );
  OR U7478 ( .A(n3390), .B(n3389), .Z(n3394) );
  NANDN U7479 ( .A(n3392), .B(n3391), .Z(n3393) );
  NAND U7480 ( .A(n3394), .B(n3393), .Z(n5352) );
  OR U7481 ( .A(n3396), .B(n3395), .Z(n3400) );
  NANDN U7482 ( .A(n3398), .B(n3397), .Z(n3399) );
  NAND U7483 ( .A(n3400), .B(n3399), .Z(n5355) );
  XOR U7484 ( .A(n5354), .B(n5355), .Z(n5094) );
  NANDN U7485 ( .A(n3402), .B(n3401), .Z(n3406) );
  NAND U7486 ( .A(n3404), .B(n3403), .Z(n3405) );
  NAND U7487 ( .A(n3406), .B(n3405), .Z(n5095) );
  XNOR U7488 ( .A(n5094), .B(n5095), .Z(n5096) );
  NANDN U7489 ( .A(n3408), .B(n3407), .Z(n3412) );
  NAND U7490 ( .A(n3410), .B(n3409), .Z(n3411) );
  AND U7491 ( .A(n3412), .B(n3411), .Z(n5097) );
  XNOR U7492 ( .A(n5096), .B(n5097), .Z(n5220) );
  OR U7493 ( .A(n3414), .B(n3413), .Z(n3418) );
  NANDN U7494 ( .A(n3416), .B(n3415), .Z(n3417) );
  NAND U7495 ( .A(n3418), .B(n3417), .Z(n7299) );
  OR U7496 ( .A(n3420), .B(n3419), .Z(n3424) );
  NANDN U7497 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U7498 ( .A(n3424), .B(n3423), .Z(n5960) );
  XNOR U7499 ( .A(n5960), .B(n5959), .Z(n5961) );
  OR U7500 ( .A(n3430), .B(n3429), .Z(n3434) );
  NANDN U7501 ( .A(n3432), .B(n3431), .Z(n3433) );
  NAND U7502 ( .A(n3434), .B(n3433), .Z(n5962) );
  XNOR U7503 ( .A(n5961), .B(n5962), .Z(n7296) );
  OR U7504 ( .A(n3436), .B(n3435), .Z(n3440) );
  NAND U7505 ( .A(n3438), .B(n3437), .Z(n3439) );
  NAND U7506 ( .A(n3440), .B(n3439), .Z(n7297) );
  XOR U7507 ( .A(n7299), .B(n7298), .Z(n5221) );
  XOR U7508 ( .A(n5220), .B(n5221), .Z(n5222) );
  NANDN U7509 ( .A(n3442), .B(n3441), .Z(n3446) );
  NAND U7510 ( .A(n3444), .B(n3443), .Z(n3445) );
  NAND U7511 ( .A(n3446), .B(n3445), .Z(n7281) );
  OR U7512 ( .A(n3448), .B(n3447), .Z(n3452) );
  NANDN U7513 ( .A(n3450), .B(n3449), .Z(n3451) );
  NAND U7514 ( .A(n3452), .B(n3451), .Z(n5954) );
  OR U7515 ( .A(n3454), .B(n3453), .Z(n3458) );
  NANDN U7516 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U7517 ( .A(n3458), .B(n3457), .Z(n5953) );
  XOR U7518 ( .A(n5955), .B(n5956), .Z(n7278) );
  NANDN U7519 ( .A(n3464), .B(n3463), .Z(n3468) );
  NAND U7520 ( .A(n3466), .B(n3465), .Z(n3467) );
  NAND U7521 ( .A(n3468), .B(n3467), .Z(n7279) );
  XNOR U7522 ( .A(n7278), .B(n7279), .Z(n7280) );
  XOR U7523 ( .A(n7281), .B(n7280), .Z(n5223) );
  XOR U7524 ( .A(n5222), .B(n5223), .Z(n5528) );
  OR U7525 ( .A(n3470), .B(n3469), .Z(n3474) );
  NANDN U7526 ( .A(n3472), .B(n3471), .Z(n3473) );
  NAND U7527 ( .A(n3474), .B(n3473), .Z(n6535) );
  OR U7528 ( .A(n3476), .B(n3475), .Z(n3480) );
  NANDN U7529 ( .A(n3478), .B(n3477), .Z(n3479) );
  AND U7530 ( .A(n3480), .B(n3479), .Z(n6534) );
  XNOR U7531 ( .A(n6535), .B(n6534), .Z(n6536) );
  OR U7532 ( .A(n3482), .B(n3481), .Z(n3486) );
  NANDN U7533 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U7534 ( .A(n3486), .B(n3485), .Z(n6537) );
  XOR U7535 ( .A(n6536), .B(n6537), .Z(n7302) );
  OR U7536 ( .A(n3488), .B(n3487), .Z(n3492) );
  NANDN U7537 ( .A(n3490), .B(n3489), .Z(n3491) );
  NAND U7538 ( .A(n3492), .B(n3491), .Z(n6607) );
  OR U7539 ( .A(n3494), .B(n3493), .Z(n3498) );
  NANDN U7540 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U7541 ( .A(n3498), .B(n3497), .Z(n6606) );
  XNOR U7542 ( .A(n6607), .B(n6606), .Z(n6608) );
  OR U7543 ( .A(n3500), .B(n3499), .Z(n3504) );
  NANDN U7544 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U7545 ( .A(n3504), .B(n3503), .Z(n6609) );
  XNOR U7546 ( .A(n6608), .B(n6609), .Z(n7303) );
  XNOR U7547 ( .A(n7302), .B(n7303), .Z(n7304) );
  OR U7548 ( .A(n3506), .B(n3505), .Z(n3510) );
  NAND U7549 ( .A(n3508), .B(n3507), .Z(n3509) );
  NAND U7550 ( .A(n3510), .B(n3509), .Z(n7305) );
  XOR U7551 ( .A(n7304), .B(n7305), .Z(n5343) );
  OR U7552 ( .A(n3516), .B(n3515), .Z(n3520) );
  NANDN U7553 ( .A(n3518), .B(n3517), .Z(n3519) );
  NAND U7554 ( .A(n3520), .B(n3519), .Z(n6125) );
  XOR U7555 ( .A(n6127), .B(n6128), .Z(n7287) );
  OR U7556 ( .A(n3530), .B(n3529), .Z(n3534) );
  NANDN U7557 ( .A(n3532), .B(n3531), .Z(n3533) );
  NAND U7558 ( .A(n3534), .B(n3533), .Z(n5857) );
  OR U7559 ( .A(n3536), .B(n3535), .Z(n3540) );
  NANDN U7560 ( .A(n3538), .B(n3537), .Z(n3539) );
  NAND U7561 ( .A(n3540), .B(n3539), .Z(n5860) );
  XOR U7562 ( .A(n5859), .B(n5860), .Z(n7284) );
  NANDN U7563 ( .A(n3542), .B(n3541), .Z(n3546) );
  NAND U7564 ( .A(n3544), .B(n3543), .Z(n3545) );
  NAND U7565 ( .A(n3546), .B(n3545), .Z(n7285) );
  XNOR U7566 ( .A(n7284), .B(n7285), .Z(n7286) );
  XNOR U7567 ( .A(n7287), .B(n7286), .Z(n5340) );
  OR U7568 ( .A(n3552), .B(n3551), .Z(n3556) );
  NANDN U7569 ( .A(n3554), .B(n3553), .Z(n3555) );
  NAND U7570 ( .A(n3556), .B(n3555), .Z(n5887) );
  OR U7571 ( .A(n3558), .B(n3557), .Z(n3562) );
  NANDN U7572 ( .A(n3560), .B(n3559), .Z(n3561) );
  NAND U7573 ( .A(n3562), .B(n3561), .Z(n5890) );
  XOR U7574 ( .A(n5889), .B(n5890), .Z(n7275) );
  OR U7575 ( .A(n3564), .B(n3563), .Z(n3568) );
  NANDN U7576 ( .A(n3566), .B(n3565), .Z(n3567) );
  NAND U7577 ( .A(n3568), .B(n3567), .Z(n5900) );
  OR U7578 ( .A(n3570), .B(n3569), .Z(n3574) );
  NANDN U7579 ( .A(n3572), .B(n3571), .Z(n3573) );
  NAND U7580 ( .A(n3574), .B(n3573), .Z(n5899) );
  OR U7581 ( .A(n3576), .B(n3575), .Z(n3580) );
  NANDN U7582 ( .A(n3578), .B(n3577), .Z(n3579) );
  NAND U7583 ( .A(n3580), .B(n3579), .Z(n5902) );
  XOR U7584 ( .A(n5901), .B(n5902), .Z(n7272) );
  NANDN U7585 ( .A(n3582), .B(n3581), .Z(n3586) );
  NAND U7586 ( .A(n3584), .B(n3583), .Z(n3585) );
  NAND U7587 ( .A(n3586), .B(n3585), .Z(n7273) );
  XNOR U7588 ( .A(n7272), .B(n7273), .Z(n7274) );
  XOR U7589 ( .A(n7275), .B(n7274), .Z(n5341) );
  XNOR U7590 ( .A(n5340), .B(n5341), .Z(n5342) );
  XNOR U7591 ( .A(n5343), .B(n5342), .Z(n5529) );
  XNOR U7592 ( .A(n5528), .B(n5529), .Z(n5530) );
  XNOR U7593 ( .A(n5531), .B(n5530), .Z(n7255) );
  XNOR U7594 ( .A(n7254), .B(n7255), .Z(n7256) );
  XNOR U7595 ( .A(n7257), .B(n7256), .Z(n4971) );
  NANDN U7596 ( .A(n3588), .B(n3587), .Z(n3592) );
  NAND U7597 ( .A(n3590), .B(n3589), .Z(n3591) );
  NAND U7598 ( .A(n3592), .B(n3591), .Z(n6319) );
  NANDN U7599 ( .A(n3594), .B(n3593), .Z(n3598) );
  OR U7600 ( .A(n3596), .B(n3595), .Z(n3597) );
  NAND U7601 ( .A(n3598), .B(n3597), .Z(n5689) );
  OR U7602 ( .A(n3604), .B(n3603), .Z(n3608) );
  NANDN U7603 ( .A(n3606), .B(n3605), .Z(n3607) );
  NAND U7604 ( .A(n3608), .B(n3607), .Z(n6589) );
  OR U7605 ( .A(n3610), .B(n3609), .Z(n3614) );
  NANDN U7606 ( .A(n3612), .B(n3611), .Z(n3613) );
  AND U7607 ( .A(n3614), .B(n3613), .Z(n6588) );
  XNOR U7608 ( .A(n6589), .B(n6588), .Z(n6590) );
  OR U7609 ( .A(n3616), .B(n3615), .Z(n3620) );
  NANDN U7610 ( .A(n3618), .B(n3617), .Z(n3619) );
  NAND U7611 ( .A(n3620), .B(n3619), .Z(n6591) );
  XOR U7612 ( .A(n6590), .B(n6591), .Z(n5950) );
  OR U7613 ( .A(n3626), .B(n3625), .Z(n3630) );
  NANDN U7614 ( .A(n3628), .B(n3627), .Z(n3629) );
  AND U7615 ( .A(n3630), .B(n3629), .Z(n7016) );
  XNOR U7616 ( .A(n7017), .B(n7016), .Z(n7018) );
  XOR U7617 ( .A(n7018), .B(n7019), .Z(n5947) );
  NANDN U7618 ( .A(n3636), .B(n3635), .Z(n3640) );
  NAND U7619 ( .A(n3638), .B(n3637), .Z(n3639) );
  NAND U7620 ( .A(n3640), .B(n3639), .Z(n5948) );
  XNOR U7621 ( .A(n5947), .B(n5948), .Z(n5949) );
  XOR U7622 ( .A(n5950), .B(n5949), .Z(n5687) );
  XNOR U7623 ( .A(n5686), .B(n5687), .Z(n5688) );
  XNOR U7624 ( .A(n5689), .B(n5688), .Z(n5839) );
  NANDN U7625 ( .A(n3642), .B(n3641), .Z(n3646) );
  OR U7626 ( .A(n3644), .B(n3643), .Z(n3645) );
  NAND U7627 ( .A(n3646), .B(n3645), .Z(n5677) );
  OR U7628 ( .A(n3648), .B(n3647), .Z(n3652) );
  NANDN U7629 ( .A(n3650), .B(n3649), .Z(n3651) );
  NAND U7630 ( .A(n3652), .B(n3651), .Z(n6553) );
  XNOR U7631 ( .A(n6553), .B(n6552), .Z(n6554) );
  XOR U7632 ( .A(n6554), .B(n6555), .Z(n5974) );
  OR U7633 ( .A(n3666), .B(n3665), .Z(n3670) );
  NANDN U7634 ( .A(n3668), .B(n3667), .Z(n3669) );
  AND U7635 ( .A(n3670), .B(n3669), .Z(n7022) );
  XNOR U7636 ( .A(n7023), .B(n7022), .Z(n7024) );
  OR U7637 ( .A(n3672), .B(n3671), .Z(n3676) );
  NANDN U7638 ( .A(n3674), .B(n3673), .Z(n3675) );
  NAND U7639 ( .A(n3676), .B(n3675), .Z(n7025) );
  XOR U7640 ( .A(n7024), .B(n7025), .Z(n5971) );
  OR U7641 ( .A(n3678), .B(n3677), .Z(n3682) );
  NANDN U7642 ( .A(n3680), .B(n3679), .Z(n3681) );
  NAND U7643 ( .A(n3682), .B(n3681), .Z(n5972) );
  XNOR U7644 ( .A(n5971), .B(n5972), .Z(n5973) );
  XNOR U7645 ( .A(n5974), .B(n5973), .Z(n5674) );
  NANDN U7646 ( .A(n3684), .B(n3683), .Z(n3688) );
  OR U7647 ( .A(n3686), .B(n3685), .Z(n3687) );
  AND U7648 ( .A(n3688), .B(n3687), .Z(n5675) );
  XNOR U7649 ( .A(n5674), .B(n5675), .Z(n5676) );
  XOR U7650 ( .A(n5677), .B(n5676), .Z(n5840) );
  XOR U7651 ( .A(n5839), .B(n5840), .Z(n5842) );
  XNOR U7652 ( .A(n6583), .B(n6582), .Z(n6584) );
  OR U7653 ( .A(n3698), .B(n3697), .Z(n3702) );
  NANDN U7654 ( .A(n3700), .B(n3699), .Z(n3701) );
  NAND U7655 ( .A(n3702), .B(n3701), .Z(n6585) );
  XOR U7656 ( .A(n6584), .B(n6585), .Z(n6452) );
  OR U7657 ( .A(n3704), .B(n3703), .Z(n3708) );
  NANDN U7658 ( .A(n3706), .B(n3705), .Z(n3707) );
  NAND U7659 ( .A(n3708), .B(n3707), .Z(n6108) );
  OR U7660 ( .A(n3710), .B(n3709), .Z(n3714) );
  NANDN U7661 ( .A(n3712), .B(n3711), .Z(n3713) );
  AND U7662 ( .A(n3714), .B(n3713), .Z(n6107) );
  XNOR U7663 ( .A(n6108), .B(n6107), .Z(n6109) );
  XOR U7664 ( .A(n6109), .B(n6110), .Z(n6449) );
  NANDN U7665 ( .A(n3720), .B(n3719), .Z(n3724) );
  NANDN U7666 ( .A(n3722), .B(n3721), .Z(n3723) );
  AND U7667 ( .A(n3724), .B(n3723), .Z(n6450) );
  XNOR U7668 ( .A(n6449), .B(n6450), .Z(n6451) );
  XNOR U7669 ( .A(n6452), .B(n6451), .Z(n5682) );
  OR U7670 ( .A(n3726), .B(n3725), .Z(n3730) );
  NANDN U7671 ( .A(n3728), .B(n3727), .Z(n3729) );
  NAND U7672 ( .A(n3730), .B(n3729), .Z(n6330) );
  OR U7673 ( .A(n3736), .B(n3735), .Z(n3740) );
  NANDN U7674 ( .A(n3738), .B(n3737), .Z(n3739) );
  NAND U7675 ( .A(n3740), .B(n3739), .Z(n6332) );
  XOR U7676 ( .A(n6331), .B(n6332), .Z(n6473) );
  NANDN U7677 ( .A(n3742), .B(n3741), .Z(n3746) );
  NAND U7678 ( .A(n3744), .B(n3743), .Z(n3745) );
  NAND U7679 ( .A(n3746), .B(n3745), .Z(n6474) );
  XNOR U7680 ( .A(n6473), .B(n6474), .Z(n6475) );
  NANDN U7681 ( .A(n3748), .B(n3747), .Z(n3752) );
  NAND U7682 ( .A(n3750), .B(n3749), .Z(n3751) );
  AND U7683 ( .A(n3752), .B(n3751), .Z(n6476) );
  XNOR U7684 ( .A(n6475), .B(n6476), .Z(n5681) );
  XNOR U7685 ( .A(n6396), .B(n6395), .Z(n6397) );
  XOR U7686 ( .A(n6397), .B(n6398), .Z(n6446) );
  OR U7687 ( .A(n3766), .B(n3765), .Z(n3770) );
  NANDN U7688 ( .A(n3768), .B(n3767), .Z(n3769) );
  NAND U7689 ( .A(n3770), .B(n3769), .Z(n6547) );
  XOR U7690 ( .A(n6548), .B(n6549), .Z(n6443) );
  XNOR U7691 ( .A(n6366), .B(n6365), .Z(n6367) );
  XNOR U7692 ( .A(n6367), .B(n6368), .Z(n6444) );
  XNOR U7693 ( .A(n6443), .B(n6444), .Z(n6445) );
  XOR U7694 ( .A(n6446), .B(n6445), .Z(n5680) );
  XOR U7695 ( .A(n5681), .B(n5680), .Z(n5683) );
  XOR U7696 ( .A(n5682), .B(n5683), .Z(n5841) );
  XOR U7697 ( .A(n5842), .B(n5841), .Z(n6318) );
  OR U7698 ( .A(n3792), .B(n3791), .Z(n3796) );
  NANDN U7699 ( .A(n3794), .B(n3793), .Z(n3795) );
  NAND U7700 ( .A(n3796), .B(n3795), .Z(n6807) );
  OR U7701 ( .A(n3798), .B(n3797), .Z(n3802) );
  NANDN U7702 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U7703 ( .A(n3802), .B(n3801), .Z(n6804) );
  NANDN U7704 ( .A(n3804), .B(n3803), .Z(n3808) );
  NAND U7705 ( .A(n3806), .B(n3805), .Z(n3807) );
  NAND U7706 ( .A(n3808), .B(n3807), .Z(n7127) );
  OR U7707 ( .A(n3814), .B(n3813), .Z(n3818) );
  NANDN U7708 ( .A(n3816), .B(n3815), .Z(n3817) );
  NAND U7709 ( .A(n3818), .B(n3817), .Z(n6974) );
  OR U7710 ( .A(n3820), .B(n3819), .Z(n3824) );
  NANDN U7711 ( .A(n3822), .B(n3821), .Z(n3823) );
  NAND U7712 ( .A(n3824), .B(n3823), .Z(n6977) );
  XNOR U7713 ( .A(n6976), .B(n6977), .Z(n7124) );
  NANDN U7714 ( .A(n3826), .B(n3825), .Z(n3830) );
  NAND U7715 ( .A(n3828), .B(n3827), .Z(n3829) );
  NAND U7716 ( .A(n3830), .B(n3829), .Z(n7125) );
  XOR U7717 ( .A(n7127), .B(n7126), .Z(n6805) );
  XOR U7718 ( .A(n6804), .B(n6805), .Z(n6806) );
  XOR U7719 ( .A(n6807), .B(n6806), .Z(n6311) );
  IV U7720 ( .A(n3835), .Z(n3836) );
  OR U7721 ( .A(n3837), .B(n3836), .Z(n3841) );
  NANDN U7722 ( .A(n3839), .B(n3838), .Z(n3840) );
  NAND U7723 ( .A(n3841), .B(n3840), .Z(n6113) );
  XNOR U7724 ( .A(n6115), .B(n6116), .Z(n6710) );
  NANDN U7725 ( .A(n3847), .B(n3846), .Z(n3851) );
  NAND U7726 ( .A(n3849), .B(n3848), .Z(n3850) );
  NAND U7727 ( .A(n3851), .B(n3850), .Z(n6711) );
  NANDN U7728 ( .A(n3853), .B(n3852), .Z(n3857) );
  NAND U7729 ( .A(n3855), .B(n3854), .Z(n3856) );
  NAND U7730 ( .A(n3857), .B(n3856), .Z(n6713) );
  XOR U7731 ( .A(n6712), .B(n6713), .Z(n6767) );
  NANDN U7732 ( .A(n3859), .B(n3858), .Z(n3863) );
  NAND U7733 ( .A(n3861), .B(n3860), .Z(n3862) );
  NAND U7734 ( .A(n3863), .B(n3862), .Z(n6965) );
  XNOR U7735 ( .A(n6614), .B(n6615), .Z(n6962) );
  NANDN U7736 ( .A(n3877), .B(n3876), .Z(n3881) );
  NAND U7737 ( .A(n3879), .B(n3878), .Z(n3880) );
  NAND U7738 ( .A(n3881), .B(n3880), .Z(n6963) );
  XOR U7739 ( .A(n6965), .B(n6964), .Z(n6764) );
  XOR U7740 ( .A(n7030), .B(n7031), .Z(n6895) );
  NANDN U7741 ( .A(n3895), .B(n3894), .Z(n3899) );
  NAND U7742 ( .A(n3897), .B(n3896), .Z(n3898) );
  NAND U7743 ( .A(n3899), .B(n3898), .Z(n6893) );
  NANDN U7744 ( .A(n3901), .B(n3900), .Z(n3905) );
  NAND U7745 ( .A(n3903), .B(n3902), .Z(n3904) );
  NAND U7746 ( .A(n3905), .B(n3904), .Z(n6892) );
  XOR U7747 ( .A(n6895), .B(n6894), .Z(n6765) );
  XNOR U7748 ( .A(n6764), .B(n6765), .Z(n6766) );
  XNOR U7749 ( .A(n6767), .B(n6766), .Z(n6312) );
  XNOR U7750 ( .A(n6311), .B(n6312), .Z(n6313) );
  XNOR U7751 ( .A(n6120), .B(n6119), .Z(n6121) );
  XOR U7752 ( .A(n6121), .B(n6122), .Z(n5010) );
  OR U7753 ( .A(n3923), .B(n3922), .Z(n3927) );
  NANDN U7754 ( .A(n3925), .B(n3924), .Z(n3926) );
  NAND U7755 ( .A(n3927), .B(n3926), .Z(n5011) );
  XNOR U7756 ( .A(n5010), .B(n5011), .Z(n5012) );
  XOR U7757 ( .A(n5013), .B(n5012), .Z(n6883) );
  NANDN U7758 ( .A(n3929), .B(n3928), .Z(n3933) );
  NAND U7759 ( .A(n3931), .B(n3930), .Z(n3932) );
  NAND U7760 ( .A(n3933), .B(n3932), .Z(n7105) );
  XNOR U7761 ( .A(n7054), .B(n7053), .Z(n7055) );
  OR U7762 ( .A(n3943), .B(n3942), .Z(n3947) );
  NANDN U7763 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U7764 ( .A(n3947), .B(n3946), .Z(n7056) );
  XNOR U7765 ( .A(n7055), .B(n7056), .Z(n7102) );
  NANDN U7766 ( .A(n3949), .B(n3948), .Z(n3953) );
  NAND U7767 ( .A(n3951), .B(n3950), .Z(n3952) );
  NAND U7768 ( .A(n3953), .B(n3952), .Z(n7103) );
  XOR U7769 ( .A(n7105), .B(n7104), .Z(n6880) );
  NANDN U7770 ( .A(n3955), .B(n3954), .Z(n3959) );
  NAND U7771 ( .A(n3957), .B(n3956), .Z(n3958) );
  NAND U7772 ( .A(n3959), .B(n3958), .Z(n5091) );
  OR U7773 ( .A(n3961), .B(n3960), .Z(n3965) );
  NANDN U7774 ( .A(n3963), .B(n3962), .Z(n3964) );
  NAND U7775 ( .A(n3965), .B(n3964), .Z(n7072) );
  OR U7776 ( .A(n3967), .B(n3966), .Z(n3971) );
  NANDN U7777 ( .A(n3969), .B(n3968), .Z(n3970) );
  NAND U7778 ( .A(n3971), .B(n3970), .Z(n7071) );
  OR U7779 ( .A(n3973), .B(n3972), .Z(n3977) );
  NANDN U7780 ( .A(n3975), .B(n3974), .Z(n3976) );
  NAND U7781 ( .A(n3977), .B(n3976), .Z(n7074) );
  XOR U7782 ( .A(n7073), .B(n7074), .Z(n5088) );
  NANDN U7783 ( .A(n3979), .B(n3978), .Z(n3983) );
  NAND U7784 ( .A(n3981), .B(n3980), .Z(n3982) );
  NAND U7785 ( .A(n3983), .B(n3982), .Z(n5089) );
  XNOR U7786 ( .A(n5088), .B(n5089), .Z(n5090) );
  XNOR U7787 ( .A(n5091), .B(n5090), .Z(n6881) );
  XNOR U7788 ( .A(n6880), .B(n6881), .Z(n6882) );
  XOR U7789 ( .A(n6883), .B(n6882), .Z(n6314) );
  XOR U7790 ( .A(n6313), .B(n6314), .Z(n6317) );
  XNOR U7791 ( .A(n6318), .B(n6317), .Z(n6320) );
  XNOR U7792 ( .A(n6319), .B(n6320), .Z(n4970) );
  XNOR U7793 ( .A(n4971), .B(n4970), .Z(n4972) );
  XNOR U7794 ( .A(n4973), .B(n4972), .Z(n6887) );
  OR U7795 ( .A(n3985), .B(n3984), .Z(n3989) );
  NANDN U7796 ( .A(n3987), .B(n3986), .Z(n3988) );
  NAND U7797 ( .A(n3989), .B(n3988), .Z(n6870) );
  OR U7798 ( .A(n3991), .B(n3990), .Z(n3995) );
  NANDN U7799 ( .A(n3993), .B(n3992), .Z(n3994) );
  NAND U7800 ( .A(n3995), .B(n3994), .Z(n6869) );
  OR U7801 ( .A(n3997), .B(n3996), .Z(n4001) );
  NANDN U7802 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U7803 ( .A(n4001), .B(n4000), .Z(n7225) );
  XOR U7804 ( .A(n7226), .B(n7227), .Z(n6410) );
  OR U7805 ( .A(n4011), .B(n4010), .Z(n4015) );
  NANDN U7806 ( .A(n4013), .B(n4012), .Z(n4014) );
  NAND U7807 ( .A(n4015), .B(n4014), .Z(n6050) );
  XOR U7808 ( .A(n6050), .B(n6049), .Z(n6051) );
  XNOR U7809 ( .A(n6051), .B(n6052), .Z(n6407) );
  OR U7810 ( .A(n4025), .B(n4024), .Z(n4029) );
  NANDN U7811 ( .A(n4027), .B(n4026), .Z(n4028) );
  NAND U7812 ( .A(n4029), .B(n4028), .Z(n6408) );
  XOR U7813 ( .A(n6407), .B(n6408), .Z(n6409) );
  XOR U7814 ( .A(n6410), .B(n6409), .Z(n6868) );
  XOR U7815 ( .A(n6869), .B(n6868), .Z(n6871) );
  XNOR U7816 ( .A(n6870), .B(n6871), .Z(n5110) );
  OR U7817 ( .A(n4031), .B(n4030), .Z(n4035) );
  NANDN U7818 ( .A(n4033), .B(n4032), .Z(n4034) );
  NAND U7819 ( .A(n4035), .B(n4034), .Z(n6877) );
  OR U7820 ( .A(n4037), .B(n4036), .Z(n4041) );
  NAND U7821 ( .A(n4039), .B(n4038), .Z(n4040) );
  NAND U7822 ( .A(n4041), .B(n4040), .Z(n6354) );
  OR U7823 ( .A(n4043), .B(n4042), .Z(n4047) );
  NANDN U7824 ( .A(n4045), .B(n4044), .Z(n4046) );
  NAND U7825 ( .A(n4047), .B(n4046), .Z(n6353) );
  NANDN U7826 ( .A(n4049), .B(n4048), .Z(n4053) );
  NAND U7827 ( .A(n4051), .B(n4050), .Z(n4052) );
  AND U7828 ( .A(n4053), .B(n4052), .Z(n6356) );
  XNOR U7829 ( .A(n6355), .B(n6356), .Z(n6875) );
  OR U7830 ( .A(n4055), .B(n4054), .Z(n4059) );
  NANDN U7831 ( .A(n4057), .B(n4056), .Z(n4058) );
  AND U7832 ( .A(n4059), .B(n4058), .Z(n6874) );
  XNOR U7833 ( .A(n6875), .B(n6874), .Z(n6876) );
  XNOR U7834 ( .A(n6877), .B(n6876), .Z(n5111) );
  XNOR U7835 ( .A(n5110), .B(n5111), .Z(n5112) );
  OR U7836 ( .A(n4061), .B(n4060), .Z(n4065) );
  NANDN U7837 ( .A(n4063), .B(n4062), .Z(n4064) );
  NAND U7838 ( .A(n4065), .B(n4064), .Z(n6813) );
  NANDN U7839 ( .A(n4067), .B(n4066), .Z(n4071) );
  NAND U7840 ( .A(n4069), .B(n4068), .Z(n4070) );
  NAND U7841 ( .A(n4071), .B(n4070), .Z(n6386) );
  NANDN U7842 ( .A(n4073), .B(n4072), .Z(n4077) );
  NANDN U7843 ( .A(n4075), .B(n4074), .Z(n4076) );
  AND U7844 ( .A(n4077), .B(n4076), .Z(n6383) );
  NANDN U7845 ( .A(n4079), .B(n4078), .Z(n4083) );
  NAND U7846 ( .A(n4081), .B(n4080), .Z(n4082) );
  NAND U7847 ( .A(n4083), .B(n4082), .Z(n6384) );
  XOR U7848 ( .A(n6386), .B(n6385), .Z(n6810) );
  OR U7849 ( .A(n4085), .B(n4084), .Z(n4089) );
  NANDN U7850 ( .A(n4087), .B(n4086), .Z(n4088) );
  AND U7851 ( .A(n4089), .B(n4088), .Z(n6811) );
  XNOR U7852 ( .A(n6810), .B(n6811), .Z(n6812) );
  XNOR U7853 ( .A(n6813), .B(n6812), .Z(n5113) );
  XOR U7854 ( .A(n5112), .B(n5113), .Z(n5187) );
  NANDN U7855 ( .A(n4095), .B(n4094), .Z(n4099) );
  OR U7856 ( .A(n4097), .B(n4096), .Z(n4098) );
  NAND U7857 ( .A(n4099), .B(n4098), .Z(n5705) );
  OR U7858 ( .A(n4101), .B(n4100), .Z(n4105) );
  NANDN U7859 ( .A(n4103), .B(n4102), .Z(n4104) );
  NAND U7860 ( .A(n4105), .B(n4104), .Z(n5702) );
  OR U7861 ( .A(n4111), .B(n4110), .Z(n4115) );
  NANDN U7862 ( .A(n4113), .B(n4112), .Z(n4114) );
  AND U7863 ( .A(n4115), .B(n4114), .Z(n5316) );
  XNOR U7864 ( .A(n5317), .B(n5316), .Z(n5318) );
  OR U7865 ( .A(n4117), .B(n4116), .Z(n4121) );
  NANDN U7866 ( .A(n4119), .B(n4118), .Z(n4120) );
  NAND U7867 ( .A(n4121), .B(n4120), .Z(n5319) );
  XOR U7868 ( .A(n5318), .B(n5319), .Z(n5919) );
  XNOR U7869 ( .A(n6288), .B(n6287), .Z(n6289) );
  OR U7870 ( .A(n4131), .B(n4130), .Z(n4135) );
  NANDN U7871 ( .A(n4133), .B(n4132), .Z(n4134) );
  NAND U7872 ( .A(n4135), .B(n4134), .Z(n6290) );
  XNOR U7873 ( .A(n6289), .B(n6290), .Z(n5917) );
  OR U7874 ( .A(n4137), .B(n4136), .Z(n4141) );
  NAND U7875 ( .A(n4139), .B(n4138), .Z(n4140) );
  NAND U7876 ( .A(n4141), .B(n4140), .Z(n5918) );
  XOR U7877 ( .A(n5919), .B(n5920), .Z(n5703) );
  XOR U7878 ( .A(n5702), .B(n5703), .Z(n5704) );
  XOR U7879 ( .A(n5705), .B(n5704), .Z(n6934) );
  NANDN U7880 ( .A(n4147), .B(n4146), .Z(n4151) );
  OR U7881 ( .A(n4149), .B(n4148), .Z(n4150) );
  NAND U7882 ( .A(n4151), .B(n4150), .Z(n5668) );
  OR U7883 ( .A(n4153), .B(n4152), .Z(n4157) );
  NANDN U7884 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U7885 ( .A(n4157), .B(n4156), .Z(n6414) );
  OR U7886 ( .A(n4159), .B(n4158), .Z(n4163) );
  NANDN U7887 ( .A(n4161), .B(n4160), .Z(n4162) );
  AND U7888 ( .A(n4163), .B(n4162), .Z(n6413) );
  XNOR U7889 ( .A(n6414), .B(n6413), .Z(n6415) );
  OR U7890 ( .A(n4165), .B(n4164), .Z(n4169) );
  NAND U7891 ( .A(n4167), .B(n4166), .Z(n4168) );
  NAND U7892 ( .A(n4169), .B(n4168), .Z(n6416) );
  XNOR U7893 ( .A(n6415), .B(n6416), .Z(n5669) );
  XNOR U7894 ( .A(n5668), .B(n5669), .Z(n5670) );
  XNOR U7895 ( .A(n5671), .B(n5670), .Z(n6935) );
  XNOR U7896 ( .A(n6934), .B(n6935), .Z(n6936) );
  XOR U7897 ( .A(n6937), .B(n6936), .Z(n5184) );
  OR U7898 ( .A(n4171), .B(n4170), .Z(n4175) );
  NANDN U7899 ( .A(n4173), .B(n4172), .Z(n4174) );
  NAND U7900 ( .A(n4175), .B(n4174), .Z(n6755) );
  OR U7901 ( .A(n4177), .B(n4176), .Z(n4181) );
  NAND U7902 ( .A(n4179), .B(n4178), .Z(n4180) );
  NAND U7903 ( .A(n4181), .B(n4180), .Z(n6752) );
  NANDN U7904 ( .A(n4183), .B(n4182), .Z(n4187) );
  NAND U7905 ( .A(n4185), .B(n4184), .Z(n4186) );
  NAND U7906 ( .A(n4187), .B(n4186), .Z(n6438) );
  NANDN U7907 ( .A(n4189), .B(n4188), .Z(n4193) );
  NAND U7908 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND U7909 ( .A(n4193), .B(n4192), .Z(n6437) );
  NANDN U7910 ( .A(n4195), .B(n4194), .Z(n4199) );
  NAND U7911 ( .A(n4197), .B(n4196), .Z(n4198) );
  NAND U7912 ( .A(n4199), .B(n4198), .Z(n6440) );
  XNOR U7913 ( .A(n6439), .B(n6440), .Z(n6753) );
  XNOR U7914 ( .A(n6752), .B(n6753), .Z(n6754) );
  XNOR U7915 ( .A(n6755), .B(n6754), .Z(n5118) );
  OR U7916 ( .A(n4201), .B(n4200), .Z(n4205) );
  NANDN U7917 ( .A(n4203), .B(n4202), .Z(n4204) );
  NAND U7918 ( .A(n4205), .B(n4204), .Z(n6761) );
  OR U7919 ( .A(n4207), .B(n4206), .Z(n4211) );
  NANDN U7920 ( .A(n4209), .B(n4208), .Z(n4210) );
  NAND U7921 ( .A(n4211), .B(n4210), .Z(n6758) );
  XOR U7922 ( .A(n6186), .B(n6185), .Z(n6187) );
  XNOR U7923 ( .A(n6187), .B(n6188), .Z(n6628) );
  XOR U7924 ( .A(n6064), .B(n6063), .Z(n6065) );
  XNOR U7925 ( .A(n6065), .B(n6066), .Z(n6625) );
  NANDN U7926 ( .A(n4237), .B(n4236), .Z(n4241) );
  NAND U7927 ( .A(n4239), .B(n4238), .Z(n4240) );
  NAND U7928 ( .A(n4241), .B(n4240), .Z(n6626) );
  XOR U7929 ( .A(n6625), .B(n6626), .Z(n6627) );
  XNOR U7930 ( .A(n6628), .B(n6627), .Z(n6759) );
  XNOR U7931 ( .A(n6758), .B(n6759), .Z(n6760) );
  XNOR U7932 ( .A(n6761), .B(n6760), .Z(n5117) );
  OR U7933 ( .A(n4243), .B(n4242), .Z(n4247) );
  NANDN U7934 ( .A(n4245), .B(n4244), .Z(n4246) );
  NAND U7935 ( .A(n4247), .B(n4246), .Z(n6819) );
  NANDN U7936 ( .A(n4249), .B(n4248), .Z(n4253) );
  NAND U7937 ( .A(n4251), .B(n4250), .Z(n4252) );
  NAND U7938 ( .A(n4253), .B(n4252), .Z(n7155) );
  NANDN U7939 ( .A(n4255), .B(n4254), .Z(n4259) );
  NAND U7940 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U7941 ( .A(n4259), .B(n4258), .Z(n7153) );
  XOR U7942 ( .A(n7155), .B(n7154), .Z(n6816) );
  OR U7943 ( .A(n4265), .B(n4264), .Z(n4269) );
  NANDN U7944 ( .A(n4267), .B(n4266), .Z(n4268) );
  AND U7945 ( .A(n4269), .B(n4268), .Z(n6817) );
  XNOR U7946 ( .A(n6816), .B(n6817), .Z(n6818) );
  XOR U7947 ( .A(n6819), .B(n6818), .Z(n5116) );
  XOR U7948 ( .A(n5117), .B(n5116), .Z(n5119) );
  XOR U7949 ( .A(n5118), .B(n5119), .Z(n5185) );
  XNOR U7950 ( .A(n5184), .B(n5185), .Z(n5186) );
  XNOR U7951 ( .A(n5187), .B(n5186), .Z(n7245) );
  OR U7952 ( .A(n4271), .B(n4270), .Z(n4275) );
  NAND U7953 ( .A(n4273), .B(n4272), .Z(n4274) );
  NAND U7954 ( .A(n4275), .B(n4274), .Z(n6865) );
  XOR U7955 ( .A(n6493), .B(n6494), .Z(n5799) );
  XNOR U7956 ( .A(n6487), .B(n6488), .Z(n5797) );
  NANDN U7957 ( .A(n4301), .B(n4300), .Z(n4305) );
  NAND U7958 ( .A(n4303), .B(n4302), .Z(n4304) );
  NAND U7959 ( .A(n4305), .B(n4304), .Z(n5798) );
  XOR U7960 ( .A(n5799), .B(n5800), .Z(n5019) );
  OR U7961 ( .A(n4307), .B(n4306), .Z(n4311) );
  NANDN U7962 ( .A(n4309), .B(n4308), .Z(n4310) );
  NAND U7963 ( .A(n4311), .B(n4310), .Z(n5016) );
  XNOR U7964 ( .A(n5016), .B(n5017), .Z(n5018) );
  XOR U7965 ( .A(n5019), .B(n5018), .Z(n6862) );
  NANDN U7966 ( .A(n4317), .B(n4316), .Z(n4321) );
  NAND U7967 ( .A(n4319), .B(n4318), .Z(n4320) );
  AND U7968 ( .A(n4321), .B(n4320), .Z(n6863) );
  XNOR U7969 ( .A(n6862), .B(n6863), .Z(n6864) );
  XNOR U7970 ( .A(n6865), .B(n6864), .Z(n5720) );
  NANDN U7971 ( .A(n4323), .B(n4322), .Z(n4327) );
  NAND U7972 ( .A(n4325), .B(n4324), .Z(n4326) );
  NAND U7973 ( .A(n4327), .B(n4326), .Z(n5721) );
  XNOR U7974 ( .A(n5720), .B(n5721), .Z(n5722) );
  XNOR U7975 ( .A(n6462), .B(n6461), .Z(n6463) );
  XOR U7976 ( .A(n6463), .B(n6464), .Z(n5280) );
  NANDN U7977 ( .A(n4341), .B(n4340), .Z(n4345) );
  NAND U7978 ( .A(n4343), .B(n4342), .Z(n4344) );
  NAND U7979 ( .A(n4345), .B(n4344), .Z(n5281) );
  XNOR U7980 ( .A(n5280), .B(n5281), .Z(n5282) );
  XNOR U7981 ( .A(n6425), .B(n6426), .Z(n6427) );
  XNOR U7982 ( .A(n6428), .B(n6427), .Z(n5283) );
  XOR U7983 ( .A(n5282), .B(n5283), .Z(n5647) );
  OR U7984 ( .A(n4359), .B(n4358), .Z(n4363) );
  NANDN U7985 ( .A(n4361), .B(n4360), .Z(n4362) );
  NAND U7986 ( .A(n4363), .B(n4362), .Z(n6402) );
  OR U7987 ( .A(n4365), .B(n4364), .Z(n4369) );
  NANDN U7988 ( .A(n4367), .B(n4366), .Z(n4368) );
  NAND U7989 ( .A(n4369), .B(n4368), .Z(n6401) );
  OR U7990 ( .A(n4371), .B(n4370), .Z(n4375) );
  NANDN U7991 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U7992 ( .A(n4375), .B(n4374), .Z(n6404) );
  XOR U7993 ( .A(n6403), .B(n6404), .Z(n5277) );
  OR U7994 ( .A(n4377), .B(n4376), .Z(n4381) );
  NANDN U7995 ( .A(n4379), .B(n4378), .Z(n4380) );
  NAND U7996 ( .A(n4381), .B(n4380), .Z(n6372) );
  OR U7997 ( .A(n4383), .B(n4382), .Z(n4387) );
  NANDN U7998 ( .A(n4385), .B(n4384), .Z(n4386) );
  NAND U7999 ( .A(n4387), .B(n4386), .Z(n6371) );
  OR U8000 ( .A(n4389), .B(n4388), .Z(n4393) );
  NANDN U8001 ( .A(n4391), .B(n4390), .Z(n4392) );
  NAND U8002 ( .A(n4393), .B(n4392), .Z(n6374) );
  XOR U8003 ( .A(n6373), .B(n6374), .Z(n5274) );
  OR U8004 ( .A(n4395), .B(n4394), .Z(n4399) );
  NAND U8005 ( .A(n4397), .B(n4396), .Z(n4398) );
  NAND U8006 ( .A(n4399), .B(n4398), .Z(n5275) );
  XNOR U8007 ( .A(n5274), .B(n5275), .Z(n5276) );
  XNOR U8008 ( .A(n5277), .B(n5276), .Z(n5644) );
  NANDN U8009 ( .A(n4401), .B(n4400), .Z(n4405) );
  OR U8010 ( .A(n4403), .B(n4402), .Z(n4404) );
  AND U8011 ( .A(n4405), .B(n4404), .Z(n5645) );
  XNOR U8012 ( .A(n5644), .B(n5645), .Z(n5646) );
  XNOR U8013 ( .A(n5647), .B(n5646), .Z(n7311) );
  OR U8014 ( .A(n4407), .B(n4406), .Z(n4411) );
  NANDN U8015 ( .A(n4409), .B(n4408), .Z(n4410) );
  NAND U8016 ( .A(n4411), .B(n4410), .Z(n6456) );
  OR U8017 ( .A(n4413), .B(n4412), .Z(n4417) );
  NANDN U8018 ( .A(n4415), .B(n4414), .Z(n4416) );
  AND U8019 ( .A(n4417), .B(n4416), .Z(n6455) );
  XNOR U8020 ( .A(n6456), .B(n6455), .Z(n6457) );
  XOR U8021 ( .A(n6457), .B(n6458), .Z(n6995) );
  OR U8022 ( .A(n4423), .B(n4422), .Z(n4427) );
  NAND U8023 ( .A(n4425), .B(n4424), .Z(n4426) );
  NAND U8024 ( .A(n4427), .B(n4426), .Z(n6993) );
  OR U8025 ( .A(n4429), .B(n4428), .Z(n4433) );
  NAND U8026 ( .A(n4431), .B(n4430), .Z(n4432) );
  AND U8027 ( .A(n4433), .B(n4432), .Z(n6992) );
  XNOR U8028 ( .A(n6993), .B(n6992), .Z(n6994) );
  XNOR U8029 ( .A(n6995), .B(n6994), .Z(n5627) );
  XNOR U8030 ( .A(n5870), .B(n5869), .Z(n5871) );
  XOR U8031 ( .A(n5871), .B(n5872), .Z(n5794) );
  OR U8032 ( .A(n4447), .B(n4446), .Z(n4451) );
  NAND U8033 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U8034 ( .A(n4451), .B(n4450), .Z(n5792) );
  OR U8035 ( .A(n4453), .B(n4452), .Z(n4457) );
  NAND U8036 ( .A(n4455), .B(n4454), .Z(n4456) );
  AND U8037 ( .A(n4457), .B(n4456), .Z(n5791) );
  XNOR U8038 ( .A(n5792), .B(n5791), .Z(n5793) );
  XNOR U8039 ( .A(n5794), .B(n5793), .Z(n5624) );
  NANDN U8040 ( .A(n4459), .B(n4458), .Z(n4463) );
  OR U8041 ( .A(n4461), .B(n4460), .Z(n4462) );
  AND U8042 ( .A(n4463), .B(n4462), .Z(n5625) );
  XNOR U8043 ( .A(n5624), .B(n5625), .Z(n5626) );
  XOR U8044 ( .A(n5627), .B(n5626), .Z(n7308) );
  OR U8045 ( .A(n4465), .B(n4464), .Z(n4469) );
  OR U8046 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U8047 ( .A(n4469), .B(n4468), .Z(n7309) );
  XOR U8048 ( .A(n7308), .B(n7309), .Z(n7310) );
  XOR U8049 ( .A(n7311), .B(n7310), .Z(n5723) );
  XOR U8050 ( .A(n5722), .B(n5723), .Z(n7242) );
  NANDN U8051 ( .A(n4471), .B(n4470), .Z(n4475) );
  NAND U8052 ( .A(n4473), .B(n4472), .Z(n4474) );
  NAND U8053 ( .A(n4475), .B(n4474), .Z(n5717) );
  NAND U8054 ( .A(n4477), .B(n4476), .Z(n4481) );
  NAND U8055 ( .A(n4479), .B(n4478), .Z(n4480) );
  NAND U8056 ( .A(n4481), .B(n4480), .Z(n5715) );
  OR U8057 ( .A(n4483), .B(n4482), .Z(n4487) );
  NAND U8058 ( .A(n4485), .B(n4484), .Z(n4486) );
  NAND U8059 ( .A(n4487), .B(n4486), .Z(n5770) );
  OR U8060 ( .A(n4489), .B(n4488), .Z(n4493) );
  NANDN U8061 ( .A(n4491), .B(n4490), .Z(n4492) );
  NAND U8062 ( .A(n4493), .B(n4492), .Z(n6342) );
  OR U8063 ( .A(n4495), .B(n4494), .Z(n4499) );
  NANDN U8064 ( .A(n4497), .B(n4496), .Z(n4498) );
  AND U8065 ( .A(n4499), .B(n4498), .Z(n6341) );
  XNOR U8066 ( .A(n6342), .B(n6341), .Z(n6343) );
  OR U8067 ( .A(n4501), .B(n4500), .Z(n4505) );
  NANDN U8068 ( .A(n4503), .B(n4502), .Z(n4504) );
  NAND U8069 ( .A(n4505), .B(n4504), .Z(n6344) );
  XOR U8070 ( .A(n6343), .B(n6344), .Z(n5767) );
  OR U8071 ( .A(n4507), .B(n4506), .Z(n4511) );
  NAND U8072 ( .A(n4509), .B(n4508), .Z(n4510) );
  NAND U8073 ( .A(n4511), .B(n4510), .Z(n5768) );
  XNOR U8074 ( .A(n5767), .B(n5768), .Z(n5769) );
  XNOR U8075 ( .A(n5770), .B(n5769), .Z(n5640) );
  OR U8076 ( .A(n4513), .B(n4512), .Z(n4517) );
  NANDN U8077 ( .A(n4515), .B(n4514), .Z(n4516) );
  NAND U8078 ( .A(n4517), .B(n4516), .Z(n5435) );
  OR U8079 ( .A(n4519), .B(n4518), .Z(n4523) );
  NANDN U8080 ( .A(n4521), .B(n4520), .Z(n4522) );
  NAND U8081 ( .A(n4523), .B(n4522), .Z(n5433) );
  NANDN U8082 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U8083 ( .A(n4527), .B(n4526), .Z(n4528) );
  AND U8084 ( .A(n4529), .B(n4528), .Z(n5432) );
  XNOR U8085 ( .A(n5433), .B(n5432), .Z(n5434) );
  XOR U8086 ( .A(n5435), .B(n5434), .Z(n5641) );
  XNOR U8087 ( .A(n5640), .B(n5641), .Z(n5642) );
  OR U8088 ( .A(n4531), .B(n4530), .Z(n4535) );
  NANDN U8089 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U8090 ( .A(n4535), .B(n4534), .Z(n6680) );
  OR U8091 ( .A(n4537), .B(n4536), .Z(n4541) );
  NANDN U8092 ( .A(n4539), .B(n4538), .Z(n4540) );
  NAND U8093 ( .A(n4541), .B(n4540), .Z(n6679) );
  OR U8094 ( .A(n4543), .B(n4542), .Z(n4547) );
  NANDN U8095 ( .A(n4545), .B(n4544), .Z(n4546) );
  NAND U8096 ( .A(n4547), .B(n4546), .Z(n6682) );
  XOR U8097 ( .A(n6681), .B(n6682), .Z(n5764) );
  OR U8098 ( .A(n4549), .B(n4548), .Z(n4553) );
  NANDN U8099 ( .A(n4551), .B(n4550), .Z(n4552) );
  NAND U8100 ( .A(n4553), .B(n4552), .Z(n6264) );
  XNOR U8101 ( .A(n6264), .B(n6263), .Z(n6265) );
  XOR U8102 ( .A(n6265), .B(n6266), .Z(n5761) );
  OR U8103 ( .A(n4563), .B(n4562), .Z(n4567) );
  NANDN U8104 ( .A(n4565), .B(n4564), .Z(n4566) );
  NAND U8105 ( .A(n4567), .B(n4566), .Z(n6735) );
  OR U8106 ( .A(n4569), .B(n4568), .Z(n4573) );
  NANDN U8107 ( .A(n4571), .B(n4570), .Z(n4572) );
  AND U8108 ( .A(n4573), .B(n4572), .Z(n6734) );
  XNOR U8109 ( .A(n6735), .B(n6734), .Z(n6736) );
  OR U8110 ( .A(n4575), .B(n4574), .Z(n4579) );
  NANDN U8111 ( .A(n4577), .B(n4576), .Z(n4578) );
  NAND U8112 ( .A(n4579), .B(n4578), .Z(n6737) );
  XNOR U8113 ( .A(n6736), .B(n6737), .Z(n5762) );
  XNOR U8114 ( .A(n5761), .B(n5762), .Z(n5763) );
  XOR U8115 ( .A(n5764), .B(n5763), .Z(n5643) );
  XOR U8116 ( .A(n5642), .B(n5643), .Z(n5714) );
  XNOR U8117 ( .A(n5715), .B(n5714), .Z(n5716) );
  XNOR U8118 ( .A(n5717), .B(n5716), .Z(n5125) );
  NANDN U8119 ( .A(n4585), .B(n4584), .Z(n4589) );
  NAND U8120 ( .A(n4587), .B(n4586), .Z(n4588) );
  NAND U8121 ( .A(n4589), .B(n4588), .Z(n6004) );
  OR U8122 ( .A(n4591), .B(n4590), .Z(n4595) );
  NANDN U8123 ( .A(n4593), .B(n4592), .Z(n4594) );
  NAND U8124 ( .A(n4595), .B(n4594), .Z(n5749) );
  OR U8125 ( .A(n4597), .B(n4596), .Z(n4601) );
  NANDN U8126 ( .A(n4599), .B(n4598), .Z(n4600) );
  NAND U8127 ( .A(n4601), .B(n4600), .Z(n5748) );
  OR U8128 ( .A(n4603), .B(n4602), .Z(n4607) );
  NANDN U8129 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U8130 ( .A(n4607), .B(n4606), .Z(n5751) );
  XOR U8131 ( .A(n5750), .B(n5751), .Z(n6001) );
  NANDN U8132 ( .A(n4609), .B(n4608), .Z(n4613) );
  NAND U8133 ( .A(n4611), .B(n4610), .Z(n4612) );
  NAND U8134 ( .A(n4613), .B(n4612), .Z(n6002) );
  XNOR U8135 ( .A(n6001), .B(n6002), .Z(n6003) );
  XOR U8136 ( .A(n6004), .B(n6003), .Z(n6306) );
  XOR U8137 ( .A(n6305), .B(n6306), .Z(n6307) );
  NANDN U8138 ( .A(n4615), .B(n4614), .Z(n4619) );
  NAND U8139 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U8140 ( .A(n4619), .B(n4618), .Z(n5525) );
  XNOR U8141 ( .A(n6729), .B(n6728), .Z(n6730) );
  XOR U8142 ( .A(n6730), .B(n6731), .Z(n5522) );
  OR U8143 ( .A(n4641), .B(n4640), .Z(n4645) );
  OR U8144 ( .A(n4643), .B(n4642), .Z(n4644) );
  AND U8145 ( .A(n4645), .B(n4644), .Z(n6073) );
  XNOR U8146 ( .A(n6074), .B(n6073), .Z(n6075) );
  XNOR U8147 ( .A(n6076), .B(n6075), .Z(n5523) );
  XNOR U8148 ( .A(n5522), .B(n5523), .Z(n5524) );
  XOR U8149 ( .A(n5525), .B(n5524), .Z(n6308) );
  XOR U8150 ( .A(n6307), .B(n6308), .Z(n6801) );
  XNOR U8151 ( .A(n6165), .B(n6166), .Z(n6167) );
  XNOR U8152 ( .A(n6178), .B(n6177), .Z(n6168) );
  XOR U8153 ( .A(n6167), .B(n6168), .Z(n6173) );
  XNOR U8154 ( .A(n6171), .B(n6172), .Z(n6174) );
  XOR U8155 ( .A(n6173), .B(n6174), .Z(n5253) );
  XNOR U8156 ( .A(n6180), .B(n6179), .Z(n6181) );
  XNOR U8157 ( .A(n6181), .B(n6182), .Z(n5251) );
  XNOR U8158 ( .A(n6150), .B(n6149), .Z(n6151) );
  XOR U8159 ( .A(n6151), .B(n6152), .Z(n5250) );
  XNOR U8160 ( .A(n5251), .B(n5250), .Z(n5252) );
  XOR U8161 ( .A(n5253), .B(n5252), .Z(n6040) );
  NANDN U8162 ( .A(n4693), .B(n4692), .Z(n4697) );
  NAND U8163 ( .A(n4695), .B(n4694), .Z(n4696) );
  NAND U8164 ( .A(n4697), .B(n4696), .Z(n7081) );
  NANDN U8165 ( .A(n4699), .B(n4698), .Z(n4703) );
  NAND U8166 ( .A(n4701), .B(n4700), .Z(n4702) );
  NAND U8167 ( .A(n4703), .B(n4702), .Z(n7078) );
  NANDN U8168 ( .A(n4705), .B(n4704), .Z(n4709) );
  NAND U8169 ( .A(n4707), .B(n4706), .Z(n4708) );
  AND U8170 ( .A(n4709), .B(n4708), .Z(n7079) );
  XNOR U8171 ( .A(n7078), .B(n7079), .Z(n7080) );
  XNOR U8172 ( .A(n7081), .B(n7080), .Z(n6037) );
  XOR U8173 ( .A(n5446), .B(n5447), .Z(n7038) );
  OR U8174 ( .A(n4723), .B(n4722), .Z(n4727) );
  NANDN U8175 ( .A(n4725), .B(n4724), .Z(n4726) );
  NAND U8176 ( .A(n4727), .B(n4726), .Z(n5171) );
  OR U8177 ( .A(n4729), .B(n4728), .Z(n4733) );
  NANDN U8178 ( .A(n4731), .B(n4730), .Z(n4732) );
  NAND U8179 ( .A(n4733), .B(n4732), .Z(n5170) );
  XOR U8180 ( .A(n5172), .B(n5173), .Z(n7035) );
  NANDN U8181 ( .A(n4739), .B(n4738), .Z(n4743) );
  NAND U8182 ( .A(n4741), .B(n4740), .Z(n4742) );
  NAND U8183 ( .A(n4743), .B(n4742), .Z(n7036) );
  XNOR U8184 ( .A(n7035), .B(n7036), .Z(n7037) );
  XNOR U8185 ( .A(n7038), .B(n7037), .Z(n6038) );
  XNOR U8186 ( .A(n6037), .B(n6038), .Z(n6039) );
  XOR U8187 ( .A(n6040), .B(n6039), .Z(n6798) );
  OR U8188 ( .A(n4745), .B(n4744), .Z(n4749) );
  NAND U8189 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U8190 ( .A(n4749), .B(n4748), .Z(n5429) );
  OR U8191 ( .A(n4751), .B(n4750), .Z(n4755) );
  NANDN U8192 ( .A(n4753), .B(n4752), .Z(n4754) );
  NAND U8193 ( .A(n4755), .B(n4754), .Z(n6258) );
  OR U8194 ( .A(n4757), .B(n4756), .Z(n4761) );
  NANDN U8195 ( .A(n4759), .B(n4758), .Z(n4760) );
  AND U8196 ( .A(n4761), .B(n4760), .Z(n6257) );
  XNOR U8197 ( .A(n6258), .B(n6257), .Z(n6259) );
  OR U8198 ( .A(n4763), .B(n4762), .Z(n4767) );
  NANDN U8199 ( .A(n4765), .B(n4764), .Z(n4766) );
  NAND U8200 ( .A(n4767), .B(n4766), .Z(n6260) );
  XOR U8201 ( .A(n6259), .B(n6260), .Z(n5426) );
  NANDN U8202 ( .A(n4769), .B(n4768), .Z(n4773) );
  NAND U8203 ( .A(n4771), .B(n4770), .Z(n4772) );
  NAND U8204 ( .A(n4773), .B(n4772), .Z(n5427) );
  XNOR U8205 ( .A(n5426), .B(n5427), .Z(n5428) );
  XOR U8206 ( .A(n5429), .B(n5428), .Z(n5459) );
  NANDN U8207 ( .A(n4775), .B(n4774), .Z(n4779) );
  NAND U8208 ( .A(n4777), .B(n4776), .Z(n4778) );
  NAND U8209 ( .A(n4779), .B(n4778), .Z(n6236) );
  XNOR U8210 ( .A(n6270), .B(n6269), .Z(n6271) );
  XOR U8211 ( .A(n6271), .B(n6272), .Z(n6233) );
  NANDN U8212 ( .A(n4793), .B(n4792), .Z(n4797) );
  NAND U8213 ( .A(n4795), .B(n4794), .Z(n4796) );
  NAND U8214 ( .A(n4797), .B(n4796), .Z(n6234) );
  XNOR U8215 ( .A(n6233), .B(n6234), .Z(n6235) );
  XOR U8216 ( .A(n6236), .B(n6235), .Z(n5456) );
  OR U8217 ( .A(n4799), .B(n4798), .Z(n4803) );
  NANDN U8218 ( .A(n4801), .B(n4800), .Z(n4802) );
  NAND U8219 ( .A(n4803), .B(n4802), .Z(n5894) );
  OR U8220 ( .A(n4809), .B(n4808), .Z(n4813) );
  NANDN U8221 ( .A(n4811), .B(n4810), .Z(n4812) );
  NAND U8222 ( .A(n4813), .B(n4812), .Z(n5896) );
  XOR U8223 ( .A(n5895), .B(n5896), .Z(n5507) );
  OR U8224 ( .A(n4819), .B(n4818), .Z(n4823) );
  NANDN U8225 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U8226 ( .A(n4823), .B(n4822), .Z(n5935) );
  XOR U8227 ( .A(n5937), .B(n5938), .Z(n5504) );
  NANDN U8228 ( .A(n4829), .B(n4828), .Z(n4833) );
  NAND U8229 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U8230 ( .A(n4833), .B(n4832), .Z(n5505) );
  XNOR U8231 ( .A(n5504), .B(n5505), .Z(n5506) );
  XOR U8232 ( .A(n5507), .B(n5506), .Z(n5457) );
  XNOR U8233 ( .A(n5456), .B(n5457), .Z(n5458) );
  XNOR U8234 ( .A(n5459), .B(n5458), .Z(n6799) );
  XOR U8235 ( .A(n6798), .B(n6799), .Z(n6800) );
  XNOR U8236 ( .A(n6801), .B(n6800), .Z(n5123) );
  NANDN U8237 ( .A(n4835), .B(n4834), .Z(n4839) );
  NAND U8238 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U8239 ( .A(n4839), .B(n4838), .Z(n6771) );
  OR U8240 ( .A(n4841), .B(n4840), .Z(n4845) );
  OR U8241 ( .A(n4843), .B(n4842), .Z(n4844) );
  NAND U8242 ( .A(n4845), .B(n4844), .Z(n6070) );
  XNOR U8243 ( .A(n6070), .B(n6069), .Z(n6071) );
  OR U8244 ( .A(n4851), .B(n4850), .Z(n4855) );
  OR U8245 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U8246 ( .A(n4855), .B(n4854), .Z(n6072) );
  XNOR U8247 ( .A(n6071), .B(n6072), .Z(n6519) );
  OR U8248 ( .A(n4857), .B(n4856), .Z(n4861) );
  OR U8249 ( .A(n4859), .B(n4858), .Z(n4860) );
  NAND U8250 ( .A(n4861), .B(n4860), .Z(n6156) );
  XNOR U8251 ( .A(n6156), .B(n6155), .Z(n6157) );
  XNOR U8252 ( .A(n6157), .B(n6158), .Z(n6516) );
  NANDN U8253 ( .A(n4871), .B(n4870), .Z(n4875) );
  NAND U8254 ( .A(n4873), .B(n4872), .Z(n4874) );
  NAND U8255 ( .A(n4875), .B(n4874), .Z(n6517) );
  XOR U8256 ( .A(n6516), .B(n6517), .Z(n6518) );
  XNOR U8257 ( .A(n6519), .B(n6518), .Z(n5726) );
  OR U8258 ( .A(n4881), .B(n4880), .Z(n4885) );
  NANDN U8259 ( .A(n4883), .B(n4882), .Z(n4884) );
  AND U8260 ( .A(n4885), .B(n4884), .Z(n5965) );
  XNOR U8261 ( .A(n5966), .B(n5965), .Z(n5967) );
  OR U8262 ( .A(n4887), .B(n4886), .Z(n4891) );
  NANDN U8263 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U8264 ( .A(n4891), .B(n4890), .Z(n5968) );
  XOR U8265 ( .A(n5967), .B(n5968), .Z(n6010) );
  OR U8266 ( .A(n4897), .B(n4896), .Z(n4901) );
  NANDN U8267 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U8268 ( .A(n4901), .B(n4900), .Z(n5358) );
  OR U8269 ( .A(n4903), .B(n4902), .Z(n4907) );
  NANDN U8270 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U8271 ( .A(n4907), .B(n4906), .Z(n5361) );
  XOR U8272 ( .A(n5360), .B(n5361), .Z(n6007) );
  OR U8273 ( .A(n4909), .B(n4908), .Z(n4913) );
  NANDN U8274 ( .A(n4911), .B(n4910), .Z(n4912) );
  NAND U8275 ( .A(n4913), .B(n4912), .Z(n6008) );
  XNOR U8276 ( .A(n6007), .B(n6008), .Z(n6009) );
  XOR U8277 ( .A(n6010), .B(n6009), .Z(n5727) );
  XOR U8278 ( .A(n5726), .B(n5727), .Z(n5728) );
  OR U8279 ( .A(n4919), .B(n4918), .Z(n4923) );
  NANDN U8280 ( .A(n4921), .B(n4920), .Z(n4922) );
  NAND U8281 ( .A(n4923), .B(n4922), .Z(n6251) );
  XOR U8282 ( .A(n6253), .B(n6254), .Z(n6284) );
  XNOR U8283 ( .A(n5245), .B(n5244), .Z(n5246) );
  XOR U8284 ( .A(n5246), .B(n5247), .Z(n6281) );
  NANDN U8285 ( .A(n4941), .B(n4940), .Z(n4945) );
  NAND U8286 ( .A(n4943), .B(n4942), .Z(n4944) );
  NAND U8287 ( .A(n4945), .B(n4944), .Z(n6282) );
  XNOR U8288 ( .A(n6281), .B(n6282), .Z(n6283) );
  XOR U8289 ( .A(n6284), .B(n6283), .Z(n5729) );
  XOR U8290 ( .A(n5728), .B(n5729), .Z(n6770) );
  XNOR U8291 ( .A(n6771), .B(n6770), .Z(n6772) );
  NANDN U8292 ( .A(n4947), .B(n4946), .Z(n4951) );
  OR U8293 ( .A(n4949), .B(n4948), .Z(n4950) );
  NAND U8294 ( .A(n4951), .B(n4950), .Z(n5633) );
  NANDN U8295 ( .A(n4953), .B(n4952), .Z(n4957) );
  OR U8296 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U8297 ( .A(n4957), .B(n4956), .Z(n5631) );
  NANDN U8298 ( .A(n4959), .B(n4958), .Z(n4963) );
  OR U8299 ( .A(n4961), .B(n4960), .Z(n4962) );
  AND U8300 ( .A(n4963), .B(n4962), .Z(n5630) );
  XNOR U8301 ( .A(n5631), .B(n5630), .Z(n5632) );
  XOR U8302 ( .A(n5633), .B(n5632), .Z(n6773) );
  XOR U8303 ( .A(n6772), .B(n6773), .Z(n5122) );
  XOR U8304 ( .A(n5123), .B(n5122), .Z(n5124) );
  XOR U8305 ( .A(n5125), .B(n5124), .Z(n7243) );
  XNOR U8306 ( .A(n7242), .B(n7243), .Z(n7244) );
  XNOR U8307 ( .A(n7245), .B(n7244), .Z(n6886) );
  XNOR U8308 ( .A(n6887), .B(n6886), .Z(n6888) );
  XOR U8309 ( .A(n6889), .B(n6888), .Z(n6748) );
  XOR U8310 ( .A(n6749), .B(n6748), .Z(o[1]) );
  NANDN U8311 ( .A(n4965), .B(n4964), .Z(n4969) );
  OR U8312 ( .A(n4967), .B(n4966), .Z(n4968) );
  NAND U8313 ( .A(n4969), .B(n4968), .Z(n8297) );
  NANDN U8314 ( .A(n4971), .B(n4970), .Z(n4975) );
  NAND U8315 ( .A(n4973), .B(n4972), .Z(n4974) );
  NAND U8316 ( .A(n4975), .B(n4974), .Z(n8294) );
  NANDN U8317 ( .A(n4981), .B(n4980), .Z(n4985) );
  NAND U8318 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U8319 ( .A(n4985), .B(n4984), .Z(n8135) );
  NANDN U8320 ( .A(n4987), .B(n4986), .Z(n4991) );
  NAND U8321 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U8322 ( .A(n4991), .B(n4990), .Z(n8133) );
  NANDN U8323 ( .A(n4993), .B(n4992), .Z(n4997) );
  NANDN U8324 ( .A(n4995), .B(n4994), .Z(n4996) );
  AND U8325 ( .A(n4997), .B(n4996), .Z(n8132) );
  XNOR U8326 ( .A(n8133), .B(n8132), .Z(n8134) );
  XOR U8327 ( .A(n8135), .B(n8134), .Z(n8012) );
  OR U8328 ( .A(n4999), .B(n4998), .Z(n5003) );
  NAND U8329 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U8330 ( .A(n5003), .B(n5002), .Z(n7743) );
  NANDN U8331 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U8332 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U8333 ( .A(n5009), .B(n5008), .Z(n7740) );
  NANDN U8334 ( .A(n5011), .B(n5010), .Z(n5015) );
  NANDN U8335 ( .A(n5013), .B(n5012), .Z(n5014) );
  AND U8336 ( .A(n5015), .B(n5014), .Z(n7741) );
  XNOR U8337 ( .A(n7740), .B(n7741), .Z(n7742) );
  XNOR U8338 ( .A(n7743), .B(n7742), .Z(n8013) );
  XNOR U8339 ( .A(n8012), .B(n8013), .Z(n8014) );
  XNOR U8340 ( .A(n8015), .B(n8014), .Z(n7901) );
  NANDN U8341 ( .A(n5017), .B(n5016), .Z(n5021) );
  NAND U8342 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U8343 ( .A(n5021), .B(n5020), .Z(n8427) );
  NANDN U8344 ( .A(n5023), .B(n5022), .Z(n5027) );
  NAND U8345 ( .A(n5025), .B(n5024), .Z(n5026) );
  NAND U8346 ( .A(n5027), .B(n5026), .Z(n7827) );
  NANDN U8347 ( .A(n5029), .B(n5028), .Z(n5033) );
  NAND U8348 ( .A(n5031), .B(n5030), .Z(n5032) );
  NAND U8349 ( .A(n5033), .B(n5032), .Z(n7825) );
  NANDN U8350 ( .A(n5035), .B(n5034), .Z(n5039) );
  NANDN U8351 ( .A(n5037), .B(n5036), .Z(n5038) );
  NAND U8352 ( .A(n5039), .B(n5038), .Z(n7824) );
  XNOR U8353 ( .A(n7827), .B(n7826), .Z(n8426) );
  XNOR U8354 ( .A(n8427), .B(n8426), .Z(n8428) );
  NANDN U8355 ( .A(n5041), .B(n5040), .Z(n5045) );
  NANDN U8356 ( .A(n5043), .B(n5042), .Z(n5044) );
  NAND U8357 ( .A(n5045), .B(n5044), .Z(n7833) );
  NANDN U8358 ( .A(n5047), .B(n5046), .Z(n5051) );
  NANDN U8359 ( .A(n5049), .B(n5048), .Z(n5050) );
  NAND U8360 ( .A(n5051), .B(n5050), .Z(n7831) );
  NANDN U8361 ( .A(n5053), .B(n5052), .Z(n5057) );
  NANDN U8362 ( .A(n5055), .B(n5054), .Z(n5056) );
  NAND U8363 ( .A(n5057), .B(n5056), .Z(n7830) );
  XOR U8364 ( .A(n7833), .B(n7832), .Z(n8429) );
  XNOR U8365 ( .A(n8428), .B(n8429), .Z(n7898) );
  OR U8366 ( .A(n5059), .B(n5058), .Z(n5063) );
  NANDN U8367 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U8368 ( .A(n5063), .B(n5062), .Z(n8355) );
  NANDN U8369 ( .A(n5065), .B(n5064), .Z(n5069) );
  NAND U8370 ( .A(n5067), .B(n5066), .Z(n5068) );
  NAND U8371 ( .A(n5069), .B(n5068), .Z(n8087) );
  NANDN U8372 ( .A(n5071), .B(n5070), .Z(n5075) );
  NAND U8373 ( .A(n5073), .B(n5072), .Z(n5074) );
  NAND U8374 ( .A(n5075), .B(n5074), .Z(n8085) );
  NANDN U8375 ( .A(n5077), .B(n5076), .Z(n5081) );
  NAND U8376 ( .A(n5079), .B(n5078), .Z(n5080) );
  NAND U8377 ( .A(n5081), .B(n5080), .Z(n8084) );
  XOR U8378 ( .A(n8087), .B(n8086), .Z(n8352) );
  NANDN U8379 ( .A(n5083), .B(n5082), .Z(n5087) );
  NANDN U8380 ( .A(n5085), .B(n5084), .Z(n5086) );
  NAND U8381 ( .A(n5087), .B(n5086), .Z(n8205) );
  NANDN U8382 ( .A(n5089), .B(n5088), .Z(n5093) );
  NANDN U8383 ( .A(n5091), .B(n5090), .Z(n5092) );
  AND U8384 ( .A(n5093), .B(n5092), .Z(n8202) );
  NANDN U8385 ( .A(n5095), .B(n5094), .Z(n5099) );
  NAND U8386 ( .A(n5097), .B(n5096), .Z(n5098) );
  AND U8387 ( .A(n5099), .B(n5098), .Z(n8203) );
  XNOR U8388 ( .A(n8205), .B(n8204), .Z(n8353) );
  XNOR U8389 ( .A(n8352), .B(n8353), .Z(n8354) );
  XNOR U8390 ( .A(n8355), .B(n8354), .Z(n7899) );
  XNOR U8391 ( .A(n7898), .B(n7899), .Z(n7900) );
  XOR U8392 ( .A(n7901), .B(n7900), .Z(n8441) );
  NANDN U8393 ( .A(n5101), .B(n5100), .Z(n5105) );
  OR U8394 ( .A(n5103), .B(n5102), .Z(n5104) );
  NAND U8395 ( .A(n5105), .B(n5104), .Z(n8438) );
  NANDN U8396 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U8397 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U8398 ( .A(n5115), .B(n5114), .Z(n7806) );
  NANDN U8399 ( .A(n5117), .B(n5116), .Z(n5121) );
  OR U8400 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U8401 ( .A(n5121), .B(n5120), .Z(n7807) );
  XNOR U8402 ( .A(n7806), .B(n7807), .Z(n7808) );
  XOR U8403 ( .A(n7809), .B(n7808), .Z(n8439) );
  XOR U8404 ( .A(n8438), .B(n8439), .Z(n8440) );
  XNOR U8405 ( .A(n8441), .B(n8440), .Z(n8295) );
  XNOR U8406 ( .A(n8294), .B(n8295), .Z(n8296) );
  XOR U8407 ( .A(n8297), .B(n8296), .Z(n7699) );
  NAND U8408 ( .A(n5123), .B(n5122), .Z(n5127) );
  NANDN U8409 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U8410 ( .A(n5127), .B(n5126), .Z(n7693) );
  NAND U8411 ( .A(n5129), .B(n5128), .Z(n5133) );
  NANDN U8412 ( .A(n5131), .B(n5130), .Z(n5132) );
  NAND U8413 ( .A(n5133), .B(n5132), .Z(n7503) );
  NANDN U8414 ( .A(n5135), .B(n5134), .Z(n5139) );
  NAND U8415 ( .A(n5137), .B(n5136), .Z(n5138) );
  NAND U8416 ( .A(n5139), .B(n5138), .Z(n7632) );
  NANDN U8417 ( .A(n5141), .B(n5140), .Z(n5145) );
  NAND U8418 ( .A(n5143), .B(n5142), .Z(n5144) );
  NAND U8419 ( .A(n5145), .B(n5144), .Z(n7631) );
  NANDN U8420 ( .A(n5147), .B(n5146), .Z(n5151) );
  NANDN U8421 ( .A(n5149), .B(n5148), .Z(n5150) );
  NAND U8422 ( .A(n5151), .B(n5150), .Z(n7839) );
  NANDN U8423 ( .A(n5153), .B(n5152), .Z(n5157) );
  NANDN U8424 ( .A(n5155), .B(n5154), .Z(n5156) );
  NAND U8425 ( .A(n5157), .B(n5156), .Z(n7836) );
  NANDN U8426 ( .A(n5159), .B(n5158), .Z(n5163) );
  NANDN U8427 ( .A(n5161), .B(n5160), .Z(n5162) );
  NAND U8428 ( .A(n5163), .B(n5162), .Z(n8393) );
  NANDN U8429 ( .A(n5165), .B(n5164), .Z(n5169) );
  NANDN U8430 ( .A(n5167), .B(n5166), .Z(n5168) );
  NAND U8431 ( .A(n5169), .B(n5168), .Z(n8390) );
  OR U8432 ( .A(n5171), .B(n5170), .Z(n5175) );
  NANDN U8433 ( .A(n5173), .B(n5172), .Z(n5174) );
  AND U8434 ( .A(n5175), .B(n5174), .Z(n8391) );
  XNOR U8435 ( .A(n8390), .B(n8391), .Z(n8392) );
  XOR U8436 ( .A(n8393), .B(n8392), .Z(n7837) );
  XNOR U8437 ( .A(n7836), .B(n7837), .Z(n7838) );
  XOR U8438 ( .A(n7839), .B(n7838), .Z(n7630) );
  XOR U8439 ( .A(n7631), .B(n7630), .Z(n7633) );
  XOR U8440 ( .A(n7632), .B(n7633), .Z(n7502) );
  XNOR U8441 ( .A(n7503), .B(n7502), .Z(n7505) );
  XNOR U8442 ( .A(n7505), .B(n7504), .Z(n7692) );
  XNOR U8443 ( .A(n7693), .B(n7692), .Z(n7695) );
  XOR U8444 ( .A(n7695), .B(n7694), .Z(n7593) );
  NANDN U8445 ( .A(n5185), .B(n5184), .Z(n5189) );
  NAND U8446 ( .A(n5187), .B(n5186), .Z(n5188) );
  NAND U8447 ( .A(n5189), .B(n5188), .Z(n7637) );
  NANDN U8448 ( .A(n5191), .B(n5190), .Z(n5195) );
  NAND U8449 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U8450 ( .A(n5195), .B(n5194), .Z(n8227) );
  OR U8451 ( .A(n5197), .B(n5196), .Z(n5201) );
  NANDN U8452 ( .A(n5199), .B(n5198), .Z(n5200) );
  NAND U8453 ( .A(n5201), .B(n5200), .Z(n8265) );
  NANDN U8454 ( .A(n5203), .B(n5202), .Z(n5207) );
  NANDN U8455 ( .A(n5205), .B(n5204), .Z(n5206) );
  NAND U8456 ( .A(n5207), .B(n5206), .Z(n8262) );
  NANDN U8457 ( .A(n5209), .B(n5208), .Z(n5213) );
  NANDN U8458 ( .A(n5211), .B(n5210), .Z(n5212) );
  AND U8459 ( .A(n5213), .B(n5212), .Z(n8263) );
  XNOR U8460 ( .A(n8262), .B(n8263), .Z(n8264) );
  XOR U8461 ( .A(n8265), .B(n8264), .Z(n8226) );
  XOR U8462 ( .A(n8227), .B(n8226), .Z(n8229) );
  NANDN U8463 ( .A(n5215), .B(n5214), .Z(n5219) );
  NAND U8464 ( .A(n5217), .B(n5216), .Z(n5218) );
  NAND U8465 ( .A(n5219), .B(n5218), .Z(n8228) );
  XNOR U8466 ( .A(n8229), .B(n8228), .Z(n7655) );
  OR U8467 ( .A(n5221), .B(n5220), .Z(n5225) );
  NANDN U8468 ( .A(n5223), .B(n5222), .Z(n5224) );
  NAND U8469 ( .A(n5225), .B(n5224), .Z(n7652) );
  NANDN U8470 ( .A(n5227), .B(n5226), .Z(n5231) );
  NAND U8471 ( .A(n5229), .B(n5228), .Z(n5230) );
  NAND U8472 ( .A(n5231), .B(n5230), .Z(n8281) );
  NANDN U8473 ( .A(n5233), .B(n5232), .Z(n5237) );
  NANDN U8474 ( .A(n5235), .B(n5234), .Z(n5236) );
  NAND U8475 ( .A(n5237), .B(n5236), .Z(n8153) );
  NANDN U8476 ( .A(n5239), .B(n5238), .Z(n5243) );
  NANDN U8477 ( .A(n5241), .B(n5240), .Z(n5242) );
  NAND U8478 ( .A(n5243), .B(n5242), .Z(n8150) );
  NANDN U8479 ( .A(n5245), .B(n5244), .Z(n5249) );
  NANDN U8480 ( .A(n5247), .B(n5246), .Z(n5248) );
  AND U8481 ( .A(n5249), .B(n5248), .Z(n8151) );
  XNOR U8482 ( .A(n8150), .B(n8151), .Z(n8152) );
  XNOR U8483 ( .A(n8153), .B(n8152), .Z(n8278) );
  NANDN U8484 ( .A(n5251), .B(n5250), .Z(n5255) );
  NANDN U8485 ( .A(n5253), .B(n5252), .Z(n5254) );
  NAND U8486 ( .A(n5255), .B(n5254), .Z(n8279) );
  XNOR U8487 ( .A(n8278), .B(n8279), .Z(n8280) );
  XNOR U8488 ( .A(n8281), .B(n8280), .Z(n7653) );
  XNOR U8489 ( .A(n7652), .B(n7653), .Z(n7654) );
  XNOR U8490 ( .A(n7655), .B(n7654), .Z(n7414) );
  NANDN U8491 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U8492 ( .A(n5259), .B(n5258), .Z(n5260) );
  NAND U8493 ( .A(n5261), .B(n5260), .Z(n8387) );
  NANDN U8494 ( .A(n5263), .B(n5262), .Z(n5267) );
  NANDN U8495 ( .A(n5265), .B(n5264), .Z(n5266) );
  NAND U8496 ( .A(n5267), .B(n5266), .Z(n8384) );
  NANDN U8497 ( .A(n5269), .B(n5268), .Z(n5273) );
  NANDN U8498 ( .A(n5271), .B(n5270), .Z(n5272) );
  AND U8499 ( .A(n5273), .B(n5272), .Z(n8385) );
  XNOR U8500 ( .A(n8384), .B(n8385), .Z(n8386) );
  XNOR U8501 ( .A(n8387), .B(n8386), .Z(n8329) );
  NANDN U8502 ( .A(n5275), .B(n5274), .Z(n5279) );
  NAND U8503 ( .A(n5277), .B(n5276), .Z(n5278) );
  AND U8504 ( .A(n5279), .B(n5278), .Z(n8328) );
  XNOR U8505 ( .A(n8329), .B(n8328), .Z(n8330) );
  NANDN U8506 ( .A(n5281), .B(n5280), .Z(n5285) );
  NANDN U8507 ( .A(n5283), .B(n5282), .Z(n5284) );
  NAND U8508 ( .A(n5285), .B(n5284), .Z(n8331) );
  XOR U8509 ( .A(n8330), .B(n8331), .Z(n7667) );
  NANDN U8510 ( .A(n5287), .B(n5286), .Z(n5291) );
  NANDN U8511 ( .A(n5289), .B(n5288), .Z(n5290) );
  NAND U8512 ( .A(n5291), .B(n5290), .Z(n7444) );
  OR U8513 ( .A(n5293), .B(n5292), .Z(n5297) );
  NANDN U8514 ( .A(n5295), .B(n5294), .Z(n5296) );
  AND U8515 ( .A(n5297), .B(n5296), .Z(n7442) );
  NANDN U8516 ( .A(n5299), .B(n5298), .Z(n5303) );
  NANDN U8517 ( .A(n5301), .B(n5300), .Z(n5302) );
  AND U8518 ( .A(n5303), .B(n5302), .Z(n7443) );
  XOR U8519 ( .A(n7444), .B(n7445), .Z(n8271) );
  NANDN U8520 ( .A(n5305), .B(n5304), .Z(n5309) );
  NANDN U8521 ( .A(n5307), .B(n5306), .Z(n5308) );
  NAND U8522 ( .A(n5309), .B(n5308), .Z(n7383) );
  OR U8523 ( .A(n5311), .B(n5310), .Z(n5315) );
  NANDN U8524 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U8525 ( .A(n5315), .B(n5314), .Z(n7380) );
  NANDN U8526 ( .A(n5317), .B(n5316), .Z(n5321) );
  NANDN U8527 ( .A(n5319), .B(n5318), .Z(n5320) );
  AND U8528 ( .A(n5321), .B(n5320), .Z(n7381) );
  XNOR U8529 ( .A(n7380), .B(n7381), .Z(n7382) );
  XNOR U8530 ( .A(n7383), .B(n7382), .Z(n8268) );
  OR U8531 ( .A(n5323), .B(n5322), .Z(n5327) );
  NANDN U8532 ( .A(n5325), .B(n5324), .Z(n5326) );
  NAND U8533 ( .A(n5327), .B(n5326), .Z(n7529) );
  OR U8534 ( .A(n5329), .B(n5328), .Z(n5333) );
  NANDN U8535 ( .A(n5331), .B(n5330), .Z(n5332) );
  AND U8536 ( .A(n5333), .B(n5332), .Z(n7526) );
  NANDN U8537 ( .A(n5335), .B(n5334), .Z(n5339) );
  NANDN U8538 ( .A(n5337), .B(n5336), .Z(n5338) );
  AND U8539 ( .A(n5339), .B(n5338), .Z(n7527) );
  XOR U8540 ( .A(n7529), .B(n7528), .Z(n8269) );
  XNOR U8541 ( .A(n8268), .B(n8269), .Z(n8270) );
  XOR U8542 ( .A(n8271), .B(n8270), .Z(n7664) );
  NANDN U8543 ( .A(n5341), .B(n5340), .Z(n5345) );
  NAND U8544 ( .A(n5343), .B(n5342), .Z(n5344) );
  AND U8545 ( .A(n5345), .B(n5344), .Z(n7665) );
  XOR U8546 ( .A(n7664), .B(n7665), .Z(n7666) );
  XOR U8547 ( .A(n7667), .B(n7666), .Z(n7415) );
  XNOR U8548 ( .A(n7414), .B(n7415), .Z(n7416) );
  OR U8549 ( .A(n5347), .B(n5346), .Z(n5351) );
  NANDN U8550 ( .A(n5349), .B(n5348), .Z(n5350) );
  NAND U8551 ( .A(n5351), .B(n5350), .Z(n7553) );
  IV U8552 ( .A(n7553), .Z(n7555) );
  OR U8553 ( .A(n5353), .B(n5352), .Z(n5357) );
  NANDN U8554 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U8555 ( .A(n5357), .B(n5356), .Z(n7557) );
  OR U8556 ( .A(n5359), .B(n5358), .Z(n5363) );
  NANDN U8557 ( .A(n5361), .B(n5360), .Z(n5362) );
  AND U8558 ( .A(n5363), .B(n5362), .Z(n7554) );
  XOR U8559 ( .A(n7557), .B(n7554), .Z(n5364) );
  XNOR U8560 ( .A(n7555), .B(n5364), .Z(n7923) );
  NANDN U8561 ( .A(n5366), .B(n5365), .Z(n5370) );
  NAND U8562 ( .A(n5368), .B(n5367), .Z(n5369) );
  AND U8563 ( .A(n5370), .B(n5369), .Z(n7922) );
  NANDN U8564 ( .A(n5372), .B(n5371), .Z(n5376) );
  NANDN U8565 ( .A(n5374), .B(n5373), .Z(n5375) );
  NAND U8566 ( .A(n5376), .B(n5375), .Z(n7924) );
  XOR U8567 ( .A(n7922), .B(n7924), .Z(n5377) );
  XOR U8568 ( .A(n7923), .B(n5377), .Z(n7660) );
  OR U8569 ( .A(n5379), .B(n5378), .Z(n5383) );
  NANDN U8570 ( .A(n5381), .B(n5380), .Z(n5382) );
  NAND U8571 ( .A(n5383), .B(n5382), .Z(n8056) );
  OR U8572 ( .A(n5385), .B(n5384), .Z(n5389) );
  NAND U8573 ( .A(n5387), .B(n5386), .Z(n5388) );
  NAND U8574 ( .A(n5389), .B(n5388), .Z(n7797) );
  OR U8575 ( .A(n5391), .B(n5390), .Z(n5395) );
  NANDN U8576 ( .A(n5393), .B(n5392), .Z(n5394) );
  NAND U8577 ( .A(n5395), .B(n5394), .Z(n7794) );
  NANDN U8578 ( .A(n5397), .B(n5396), .Z(n5401) );
  NANDN U8579 ( .A(n5399), .B(n5398), .Z(n5400) );
  AND U8580 ( .A(n5401), .B(n5400), .Z(n7795) );
  XNOR U8581 ( .A(n7794), .B(n7795), .Z(n7796) );
  XNOR U8582 ( .A(n7797), .B(n7796), .Z(n8054) );
  NANDN U8583 ( .A(n5403), .B(n5402), .Z(n5407) );
  NAND U8584 ( .A(n5405), .B(n5404), .Z(n5406) );
  AND U8585 ( .A(n5407), .B(n5406), .Z(n8055) );
  XOR U8586 ( .A(n8056), .B(n8057), .Z(n7658) );
  OR U8587 ( .A(n5409), .B(n5408), .Z(n5413) );
  NANDN U8588 ( .A(n5411), .B(n5410), .Z(n5412) );
  NAND U8589 ( .A(n5413), .B(n5412), .Z(n7659) );
  XOR U8590 ( .A(n7658), .B(n7659), .Z(n7661) );
  XNOR U8591 ( .A(n7660), .B(n7661), .Z(n7417) );
  XOR U8592 ( .A(n7416), .B(n7417), .Z(n7636) );
  XNOR U8593 ( .A(n7637), .B(n7636), .Z(n7638) );
  NANDN U8594 ( .A(n5415), .B(n5414), .Z(n5419) );
  NANDN U8595 ( .A(n5417), .B(n5416), .Z(n5418) );
  NAND U8596 ( .A(n5419), .B(n5418), .Z(n7584) );
  NANDN U8597 ( .A(n5421), .B(n5420), .Z(n5425) );
  NAND U8598 ( .A(n5423), .B(n5422), .Z(n5424) );
  NAND U8599 ( .A(n5425), .B(n5424), .Z(n7679) );
  NANDN U8600 ( .A(n5427), .B(n5426), .Z(n5431) );
  NANDN U8601 ( .A(n5429), .B(n5428), .Z(n5430) );
  NAND U8602 ( .A(n5431), .B(n5430), .Z(n7953) );
  NANDN U8603 ( .A(n5433), .B(n5432), .Z(n5437) );
  NANDN U8604 ( .A(n5435), .B(n5434), .Z(n5436) );
  NAND U8605 ( .A(n5437), .B(n5436), .Z(n7950) );
  OR U8606 ( .A(n5439), .B(n5438), .Z(n5443) );
  NANDN U8607 ( .A(n5441), .B(n5440), .Z(n5442) );
  NAND U8608 ( .A(n5443), .B(n5442), .Z(n7791) );
  OR U8609 ( .A(n5445), .B(n5444), .Z(n5449) );
  NANDN U8610 ( .A(n5447), .B(n5446), .Z(n5448) );
  NAND U8611 ( .A(n5449), .B(n5448), .Z(n7788) );
  NANDN U8612 ( .A(n5451), .B(n5450), .Z(n5455) );
  NANDN U8613 ( .A(n5453), .B(n5452), .Z(n5454) );
  AND U8614 ( .A(n5455), .B(n5454), .Z(n7789) );
  XNOR U8615 ( .A(n7788), .B(n7789), .Z(n7790) );
  XOR U8616 ( .A(n7791), .B(n7790), .Z(n7951) );
  XNOR U8617 ( .A(n7950), .B(n7951), .Z(n7952) );
  XNOR U8618 ( .A(n7953), .B(n7952), .Z(n7676) );
  NANDN U8619 ( .A(n5457), .B(n5456), .Z(n5461) );
  NAND U8620 ( .A(n5459), .B(n5458), .Z(n5460) );
  AND U8621 ( .A(n5461), .B(n5460), .Z(n7677) );
  XNOR U8622 ( .A(n7676), .B(n7677), .Z(n7678) );
  XNOR U8623 ( .A(n7679), .B(n7678), .Z(n7585) );
  XOR U8624 ( .A(n7584), .B(n7585), .Z(n7586) );
  NANDN U8625 ( .A(n5463), .B(n5462), .Z(n5467) );
  NAND U8626 ( .A(n5465), .B(n5464), .Z(n5466) );
  AND U8627 ( .A(n5467), .B(n5466), .Z(n7587) );
  XOR U8628 ( .A(n7586), .B(n7587), .Z(n7639) );
  XOR U8629 ( .A(n7638), .B(n7639), .Z(n7590) );
  OR U8630 ( .A(n5469), .B(n5468), .Z(n5473) );
  NANDN U8631 ( .A(n5471), .B(n5470), .Z(n5472) );
  NAND U8632 ( .A(n5473), .B(n5472), .Z(n7475) );
  NANDN U8633 ( .A(n5475), .B(n5474), .Z(n5479) );
  NANDN U8634 ( .A(n5477), .B(n5476), .Z(n5478) );
  NAND U8635 ( .A(n5479), .B(n5478), .Z(n7472) );
  NANDN U8636 ( .A(n5481), .B(n5480), .Z(n5485) );
  NANDN U8637 ( .A(n5483), .B(n5482), .Z(n5484) );
  NAND U8638 ( .A(n5485), .B(n5484), .Z(n7785) );
  OR U8639 ( .A(n5487), .B(n5486), .Z(n5491) );
  NANDN U8640 ( .A(n5489), .B(n5488), .Z(n5490) );
  NAND U8641 ( .A(n5491), .B(n5490), .Z(n7782) );
  OR U8642 ( .A(n5493), .B(n5492), .Z(n5497) );
  NANDN U8643 ( .A(n5495), .B(n5494), .Z(n5496) );
  AND U8644 ( .A(n5497), .B(n5496), .Z(n7783) );
  XNOR U8645 ( .A(n7782), .B(n7783), .Z(n7784) );
  XOR U8646 ( .A(n7785), .B(n7784), .Z(n7473) );
  XNOR U8647 ( .A(n7472), .B(n7473), .Z(n7474) );
  XNOR U8648 ( .A(n7475), .B(n7474), .Z(n8184) );
  NANDN U8649 ( .A(n5499), .B(n5498), .Z(n5503) );
  NAND U8650 ( .A(n5501), .B(n5500), .Z(n5502) );
  AND U8651 ( .A(n5503), .B(n5502), .Z(n8185) );
  XOR U8652 ( .A(n8184), .B(n8185), .Z(n8187) );
  NANDN U8653 ( .A(n5505), .B(n5504), .Z(n5509) );
  NAND U8654 ( .A(n5507), .B(n5506), .Z(n5508) );
  NAND U8655 ( .A(n5509), .B(n5508), .Z(n7746) );
  XNOR U8656 ( .A(n8408), .B(n8409), .Z(n8411) );
  XNOR U8657 ( .A(n8410), .B(n8411), .Z(n7747) );
  XOR U8658 ( .A(n7746), .B(n7747), .Z(n7748) );
  NANDN U8659 ( .A(n5523), .B(n5522), .Z(n5527) );
  NANDN U8660 ( .A(n5525), .B(n5524), .Z(n5526) );
  AND U8661 ( .A(n5527), .B(n5526), .Z(n7749) );
  XNOR U8662 ( .A(n7748), .B(n7749), .Z(n8186) );
  XNOR U8663 ( .A(n8187), .B(n8186), .Z(n7983) );
  NANDN U8664 ( .A(n5529), .B(n5528), .Z(n5533) );
  NAND U8665 ( .A(n5531), .B(n5530), .Z(n5532) );
  NAND U8666 ( .A(n5533), .B(n5532), .Z(n7981) );
  OR U8667 ( .A(n5535), .B(n5534), .Z(n5539) );
  NANDN U8668 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U8669 ( .A(n5539), .B(n5538), .Z(n7484) );
  NANDN U8670 ( .A(n5541), .B(n5540), .Z(n5545) );
  NANDN U8671 ( .A(n5543), .B(n5542), .Z(n5544) );
  AND U8672 ( .A(n5545), .B(n5544), .Z(n7485) );
  NANDN U8673 ( .A(n5547), .B(n5546), .Z(n5551) );
  NAND U8674 ( .A(n5549), .B(n5548), .Z(n5550) );
  AND U8675 ( .A(n5551), .B(n5550), .Z(n7487) );
  XNOR U8676 ( .A(n7486), .B(n7487), .Z(n8245) );
  NANDN U8677 ( .A(n5553), .B(n5552), .Z(n5557) );
  NANDN U8678 ( .A(n5555), .B(n5554), .Z(n5556) );
  NAND U8679 ( .A(n5557), .B(n5556), .Z(n8337) );
  NANDN U8680 ( .A(n5559), .B(n5558), .Z(n5563) );
  NANDN U8681 ( .A(n5561), .B(n5560), .Z(n5562) );
  NAND U8682 ( .A(n5563), .B(n5562), .Z(n8334) );
  NANDN U8683 ( .A(n5565), .B(n5564), .Z(n5569) );
  NANDN U8684 ( .A(n5567), .B(n5566), .Z(n5568) );
  AND U8685 ( .A(n5569), .B(n5568), .Z(n8335) );
  XNOR U8686 ( .A(n8334), .B(n8335), .Z(n8336) );
  XOR U8687 ( .A(n8337), .B(n8336), .Z(n8244) );
  XOR U8688 ( .A(n8245), .B(n8244), .Z(n8247) );
  NANDN U8689 ( .A(n5571), .B(n5570), .Z(n5575) );
  NANDN U8690 ( .A(n5573), .B(n5572), .Z(n5574) );
  NAND U8691 ( .A(n5575), .B(n5574), .Z(n7731) );
  NANDN U8692 ( .A(n5577), .B(n5576), .Z(n5581) );
  NANDN U8693 ( .A(n5579), .B(n5578), .Z(n5580) );
  NAND U8694 ( .A(n5581), .B(n5580), .Z(n7728) );
  NANDN U8695 ( .A(n5583), .B(n5582), .Z(n5587) );
  NANDN U8696 ( .A(n5585), .B(n5584), .Z(n5586) );
  AND U8697 ( .A(n5587), .B(n5586), .Z(n7729) );
  XNOR U8698 ( .A(n7728), .B(n7729), .Z(n7730) );
  XNOR U8699 ( .A(n7731), .B(n7730), .Z(n8246) );
  XNOR U8700 ( .A(n8247), .B(n8246), .Z(n8211) );
  OR U8701 ( .A(n5589), .B(n5588), .Z(n5593) );
  NANDN U8702 ( .A(n5591), .B(n5590), .Z(n5592) );
  NAND U8703 ( .A(n5593), .B(n5592), .Z(n8208) );
  OR U8704 ( .A(n5595), .B(n5594), .Z(n5599) );
  NANDN U8705 ( .A(n5597), .B(n5596), .Z(n5598) );
  NAND U8706 ( .A(n5599), .B(n5598), .Z(n7463) );
  NANDN U8707 ( .A(n5601), .B(n5600), .Z(n5605) );
  NANDN U8708 ( .A(n5603), .B(n5602), .Z(n5604) );
  NAND U8709 ( .A(n5605), .B(n5604), .Z(n7713) );
  OR U8710 ( .A(n5607), .B(n5606), .Z(n5611) );
  NANDN U8711 ( .A(n5609), .B(n5608), .Z(n5610) );
  NAND U8712 ( .A(n5611), .B(n5610), .Z(n7710) );
  OR U8713 ( .A(n5613), .B(n5612), .Z(n5617) );
  NANDN U8714 ( .A(n5615), .B(n5614), .Z(n5616) );
  AND U8715 ( .A(n5617), .B(n5616), .Z(n7711) );
  XNOR U8716 ( .A(n7710), .B(n7711), .Z(n7712) );
  XNOR U8717 ( .A(n7713), .B(n7712), .Z(n7460) );
  NANDN U8718 ( .A(n5619), .B(n5618), .Z(n5623) );
  NANDN U8719 ( .A(n5621), .B(n5620), .Z(n5622) );
  AND U8720 ( .A(n5623), .B(n5622), .Z(n7461) );
  XNOR U8721 ( .A(n7460), .B(n7461), .Z(n7462) );
  XNOR U8722 ( .A(n7463), .B(n7462), .Z(n8209) );
  XNOR U8723 ( .A(n8208), .B(n8209), .Z(n8210) );
  XOR U8724 ( .A(n8211), .B(n8210), .Z(n7980) );
  XNOR U8725 ( .A(n7981), .B(n7980), .Z(n7982) );
  XNOR U8726 ( .A(n7983), .B(n7982), .Z(n8434) );
  NANDN U8727 ( .A(n5625), .B(n5624), .Z(n5629) );
  NAND U8728 ( .A(n5627), .B(n5626), .Z(n5628) );
  NAND U8729 ( .A(n5629), .B(n5628), .Z(n7673) );
  NANDN U8730 ( .A(n5631), .B(n5630), .Z(n5635) );
  NANDN U8731 ( .A(n5633), .B(n5632), .Z(n5634) );
  NAND U8732 ( .A(n5635), .B(n5634), .Z(n7670) );
  XNOR U8733 ( .A(n7670), .B(n7671), .Z(n7672) );
  XOR U8734 ( .A(n7673), .B(n7672), .Z(n7334) );
  XNOR U8735 ( .A(n7619), .B(n7618), .Z(n7620) );
  XNOR U8736 ( .A(n7621), .B(n7620), .Z(n7333) );
  OR U8737 ( .A(n5657), .B(n5656), .Z(n5661) );
  NAND U8738 ( .A(n5659), .B(n5658), .Z(n5660) );
  NAND U8739 ( .A(n5661), .B(n5660), .Z(n7467) );
  XNOR U8740 ( .A(n7466), .B(n7467), .Z(n7468) );
  NANDN U8741 ( .A(n5663), .B(n5662), .Z(n5667) );
  NAND U8742 ( .A(n5665), .B(n5664), .Z(n5666) );
  AND U8743 ( .A(n5667), .B(n5666), .Z(n7469) );
  XOR U8744 ( .A(n7468), .B(n7469), .Z(n7332) );
  XOR U8745 ( .A(n7333), .B(n7332), .Z(n7335) );
  XNOR U8746 ( .A(n7334), .B(n7335), .Z(n8433) );
  NANDN U8747 ( .A(n5669), .B(n5668), .Z(n5673) );
  NAND U8748 ( .A(n5671), .B(n5670), .Z(n5672) );
  NAND U8749 ( .A(n5673), .B(n5672), .Z(n7541) );
  NANDN U8750 ( .A(n5675), .B(n5674), .Z(n5679) );
  NAND U8751 ( .A(n5677), .B(n5676), .Z(n5678) );
  NAND U8752 ( .A(n5679), .B(n5678), .Z(n7538) );
  NANDN U8753 ( .A(n5681), .B(n5680), .Z(n5685) );
  OR U8754 ( .A(n5683), .B(n5682), .Z(n5684) );
  NAND U8755 ( .A(n5685), .B(n5684), .Z(n7539) );
  XNOR U8756 ( .A(n7538), .B(n7539), .Z(n7540) );
  XNOR U8757 ( .A(n7541), .B(n7540), .Z(n7991) );
  NANDN U8758 ( .A(n5687), .B(n5686), .Z(n5691) );
  NAND U8759 ( .A(n5689), .B(n5688), .Z(n5690) );
  NAND U8760 ( .A(n5691), .B(n5690), .Z(n7989) );
  XNOR U8761 ( .A(n7989), .B(n7988), .Z(n7990) );
  XOR U8762 ( .A(n7991), .B(n7990), .Z(n7879) );
  NANDN U8763 ( .A(n5697), .B(n5696), .Z(n5701) );
  NANDN U8764 ( .A(n5699), .B(n5698), .Z(n5700) );
  NAND U8765 ( .A(n5701), .B(n5700), .Z(n7341) );
  OR U8766 ( .A(n5703), .B(n5702), .Z(n5707) );
  NANDN U8767 ( .A(n5705), .B(n5704), .Z(n5706) );
  NAND U8768 ( .A(n5707), .B(n5706), .Z(n7338) );
  NANDN U8769 ( .A(n5709), .B(n5708), .Z(n5713) );
  NAND U8770 ( .A(n5711), .B(n5710), .Z(n5712) );
  NAND U8771 ( .A(n5713), .B(n5712), .Z(n7339) );
  XNOR U8772 ( .A(n7338), .B(n7339), .Z(n7340) );
  XNOR U8773 ( .A(n7341), .B(n7340), .Z(n7876) );
  NANDN U8774 ( .A(n5715), .B(n5714), .Z(n5719) );
  NAND U8775 ( .A(n5717), .B(n5716), .Z(n5718) );
  NAND U8776 ( .A(n5719), .B(n5718), .Z(n7877) );
  XNOR U8777 ( .A(n7876), .B(n7877), .Z(n7878) );
  XNOR U8778 ( .A(n7879), .B(n7878), .Z(n8432) );
  XNOR U8779 ( .A(n8433), .B(n8432), .Z(n8435) );
  XOR U8780 ( .A(n8434), .B(n8435), .Z(n7591) );
  XNOR U8781 ( .A(n7590), .B(n7591), .Z(n7592) );
  XNOR U8782 ( .A(n7593), .B(n7592), .Z(n7698) );
  XNOR U8783 ( .A(n7699), .B(n7698), .Z(n7701) );
  NANDN U8784 ( .A(n5721), .B(n5720), .Z(n5725) );
  NAND U8785 ( .A(n5723), .B(n5722), .Z(n5724) );
  NAND U8786 ( .A(n5725), .B(n5724), .Z(n8452) );
  NANDN U8787 ( .A(n5731), .B(n5730), .Z(n5735) );
  NAND U8788 ( .A(n5733), .B(n5732), .Z(n5734) );
  NAND U8789 ( .A(n5735), .B(n5734), .Z(n7647) );
  XNOR U8790 ( .A(n7646), .B(n7647), .Z(n7648) );
  NANDN U8791 ( .A(n5737), .B(n5736), .Z(n5741) );
  NAND U8792 ( .A(n5739), .B(n5738), .Z(n5740) );
  NAND U8793 ( .A(n5741), .B(n5740), .Z(n8165) );
  OR U8794 ( .A(n5743), .B(n5742), .Z(n5747) );
  NANDN U8795 ( .A(n5745), .B(n5744), .Z(n5746) );
  NAND U8796 ( .A(n5747), .B(n5746), .Z(n7552) );
  OR U8797 ( .A(n5749), .B(n5748), .Z(n5753) );
  NANDN U8798 ( .A(n5751), .B(n5750), .Z(n5752) );
  AND U8799 ( .A(n5753), .B(n5752), .Z(n7551) );
  OR U8800 ( .A(n5755), .B(n5754), .Z(n5759) );
  NANDN U8801 ( .A(n5757), .B(n5756), .Z(n5758) );
  AND U8802 ( .A(n5759), .B(n5758), .Z(n7550) );
  XNOR U8803 ( .A(n7551), .B(n7550), .Z(n5760) );
  XNOR U8804 ( .A(n7552), .B(n5760), .Z(n8163) );
  NANDN U8805 ( .A(n5762), .B(n5761), .Z(n5766) );
  NAND U8806 ( .A(n5764), .B(n5763), .Z(n5765) );
  AND U8807 ( .A(n5766), .B(n5765), .Z(n8162) );
  XNOR U8808 ( .A(n8165), .B(n8164), .Z(n7649) );
  XOR U8809 ( .A(n7648), .B(n7649), .Z(n7845) );
  NANDN U8810 ( .A(n5768), .B(n5767), .Z(n5772) );
  NANDN U8811 ( .A(n5770), .B(n5769), .Z(n5771) );
  NAND U8812 ( .A(n5772), .B(n5771), .Z(n7563) );
  NANDN U8813 ( .A(n5774), .B(n5773), .Z(n5778) );
  NANDN U8814 ( .A(n5776), .B(n5775), .Z(n5777) );
  NAND U8815 ( .A(n5778), .B(n5777), .Z(n8399) );
  NANDN U8816 ( .A(n5780), .B(n5779), .Z(n5784) );
  NANDN U8817 ( .A(n5782), .B(n5781), .Z(n5783) );
  NAND U8818 ( .A(n5784), .B(n5783), .Z(n8396) );
  NANDN U8819 ( .A(n5786), .B(n5785), .Z(n5790) );
  NANDN U8820 ( .A(n5788), .B(n5787), .Z(n5789) );
  AND U8821 ( .A(n5790), .B(n5789), .Z(n8397) );
  XNOR U8822 ( .A(n8396), .B(n8397), .Z(n8398) );
  XNOR U8823 ( .A(n8399), .B(n8398), .Z(n7560) );
  NANDN U8824 ( .A(n5792), .B(n5791), .Z(n5796) );
  NAND U8825 ( .A(n5794), .B(n5793), .Z(n5795) );
  AND U8826 ( .A(n5796), .B(n5795), .Z(n7561) );
  XNOR U8827 ( .A(n7560), .B(n7561), .Z(n7562) );
  XNOR U8828 ( .A(n7563), .B(n7562), .Z(n7627) );
  OR U8829 ( .A(n5798), .B(n5797), .Z(n5802) );
  NANDN U8830 ( .A(n5800), .B(n5799), .Z(n5801) );
  NAND U8831 ( .A(n5802), .B(n5801), .Z(n8191) );
  OR U8832 ( .A(n5804), .B(n5803), .Z(n5808) );
  NANDN U8833 ( .A(n5806), .B(n5805), .Z(n5807) );
  AND U8834 ( .A(n5808), .B(n5807), .Z(n8190) );
  XNOR U8835 ( .A(n8191), .B(n8190), .Z(n8192) );
  OR U8836 ( .A(n5810), .B(n5809), .Z(n5814) );
  NANDN U8837 ( .A(n5812), .B(n5811), .Z(n5813) );
  NAND U8838 ( .A(n5814), .B(n5813), .Z(n8402) );
  XNOR U8839 ( .A(n8402), .B(n8403), .Z(n8404) );
  XNOR U8840 ( .A(n8404), .B(n8405), .Z(n8193) );
  XOR U8841 ( .A(n8192), .B(n8193), .Z(n7624) );
  OR U8842 ( .A(n5824), .B(n5823), .Z(n5828) );
  NANDN U8843 ( .A(n5826), .B(n5825), .Z(n5827) );
  AND U8844 ( .A(n5828), .B(n5827), .Z(n7625) );
  XNOR U8845 ( .A(n7624), .B(n7625), .Z(n7626) );
  XOR U8846 ( .A(n7627), .B(n7626), .Z(n7842) );
  XNOR U8847 ( .A(n7842), .B(n7843), .Z(n7844) );
  XNOR U8848 ( .A(n7845), .B(n7844), .Z(n8451) );
  OR U8849 ( .A(n5834), .B(n5833), .Z(n5838) );
  OR U8850 ( .A(n5836), .B(n5835), .Z(n5837) );
  AND U8851 ( .A(n5838), .B(n5837), .Z(n8450) );
  XOR U8852 ( .A(n8451), .B(n8450), .Z(n8453) );
  XNOR U8853 ( .A(n8452), .B(n8453), .Z(n8290) );
  NANDN U8854 ( .A(n5840), .B(n5839), .Z(n5844) );
  NANDN U8855 ( .A(n5842), .B(n5841), .Z(n5843) );
  NAND U8856 ( .A(n5844), .B(n5843), .Z(n8215) );
  NANDN U8857 ( .A(n5846), .B(n5845), .Z(n5850) );
  NAND U8858 ( .A(n5848), .B(n5847), .Z(n5849) );
  NAND U8859 ( .A(n5850), .B(n5849), .Z(n8069) );
  NANDN U8860 ( .A(n5852), .B(n5851), .Z(n5856) );
  NAND U8861 ( .A(n5854), .B(n5853), .Z(n5855) );
  NAND U8862 ( .A(n5856), .B(n5855), .Z(n7857) );
  OR U8863 ( .A(n5858), .B(n5857), .Z(n5862) );
  NANDN U8864 ( .A(n5860), .B(n5859), .Z(n5861) );
  NAND U8865 ( .A(n5862), .B(n5861), .Z(n7725) );
  OR U8866 ( .A(n5864), .B(n5863), .Z(n5868) );
  NANDN U8867 ( .A(n5866), .B(n5865), .Z(n5867) );
  NAND U8868 ( .A(n5868), .B(n5867), .Z(n7722) );
  NANDN U8869 ( .A(n5870), .B(n5869), .Z(n5874) );
  NANDN U8870 ( .A(n5872), .B(n5871), .Z(n5873) );
  AND U8871 ( .A(n5874), .B(n5873), .Z(n7723) );
  XNOR U8872 ( .A(n7722), .B(n7723), .Z(n7724) );
  XNOR U8873 ( .A(n7725), .B(n7724), .Z(n7854) );
  NANDN U8874 ( .A(n5876), .B(n5875), .Z(n5880) );
  NAND U8875 ( .A(n5878), .B(n5877), .Z(n5879) );
  AND U8876 ( .A(n5880), .B(n5879), .Z(n7855) );
  XNOR U8877 ( .A(n7854), .B(n7855), .Z(n7856) );
  XNOR U8878 ( .A(n7857), .B(n7856), .Z(n8066) );
  OR U8879 ( .A(n5882), .B(n5881), .Z(n5886) );
  NANDN U8880 ( .A(n5884), .B(n5883), .Z(n5885) );
  NAND U8881 ( .A(n5886), .B(n5885), .Z(n7869) );
  OR U8882 ( .A(n5888), .B(n5887), .Z(n5892) );
  NANDN U8883 ( .A(n5890), .B(n5889), .Z(n5891) );
  NAND U8884 ( .A(n5892), .B(n5891), .Z(n7767) );
  OR U8885 ( .A(n5894), .B(n5893), .Z(n5898) );
  NANDN U8886 ( .A(n5896), .B(n5895), .Z(n5897) );
  NAND U8887 ( .A(n5898), .B(n5897), .Z(n7764) );
  OR U8888 ( .A(n5900), .B(n5899), .Z(n5904) );
  NANDN U8889 ( .A(n5902), .B(n5901), .Z(n5903) );
  AND U8890 ( .A(n5904), .B(n5903), .Z(n7765) );
  XNOR U8891 ( .A(n7764), .B(n7765), .Z(n7766) );
  XNOR U8892 ( .A(n7767), .B(n7766), .Z(n7866) );
  NANDN U8893 ( .A(n5906), .B(n5905), .Z(n5910) );
  NANDN U8894 ( .A(n5908), .B(n5907), .Z(n5909) );
  AND U8895 ( .A(n5910), .B(n5909), .Z(n7867) );
  XNOR U8896 ( .A(n7866), .B(n7867), .Z(n7868) );
  XNOR U8897 ( .A(n7869), .B(n7868), .Z(n8067) );
  XOR U8898 ( .A(n8066), .B(n8067), .Z(n8068) );
  XNOR U8899 ( .A(n8069), .B(n8068), .Z(n8214) );
  XNOR U8900 ( .A(n8215), .B(n8214), .Z(n8216) );
  NANDN U8901 ( .A(n5912), .B(n5911), .Z(n5916) );
  NAND U8902 ( .A(n5914), .B(n5913), .Z(n5915) );
  NAND U8903 ( .A(n5916), .B(n5915), .Z(n8181) );
  OR U8904 ( .A(n5918), .B(n5917), .Z(n5922) );
  NANDN U8905 ( .A(n5920), .B(n5919), .Z(n5921) );
  NAND U8906 ( .A(n5922), .B(n5921), .Z(n8043) );
  OR U8907 ( .A(n5924), .B(n5923), .Z(n5928) );
  NANDN U8908 ( .A(n5926), .B(n5925), .Z(n5927) );
  NAND U8909 ( .A(n5928), .B(n5927), .Z(n7755) );
  OR U8910 ( .A(n5930), .B(n5929), .Z(n5934) );
  NANDN U8911 ( .A(n5932), .B(n5931), .Z(n5933) );
  NAND U8912 ( .A(n5934), .B(n5933), .Z(n7752) );
  OR U8913 ( .A(n5936), .B(n5935), .Z(n5940) );
  NANDN U8914 ( .A(n5938), .B(n5937), .Z(n5939) );
  AND U8915 ( .A(n5940), .B(n5939), .Z(n7753) );
  XNOR U8916 ( .A(n7752), .B(n7753), .Z(n7754) );
  XOR U8917 ( .A(n7755), .B(n7754), .Z(n8042) );
  XOR U8918 ( .A(n8043), .B(n8042), .Z(n8045) );
  NANDN U8919 ( .A(n5942), .B(n5941), .Z(n5946) );
  NAND U8920 ( .A(n5944), .B(n5943), .Z(n5945) );
  NAND U8921 ( .A(n5946), .B(n5945), .Z(n8044) );
  XNOR U8922 ( .A(n8045), .B(n8044), .Z(n8178) );
  NANDN U8923 ( .A(n5948), .B(n5947), .Z(n5952) );
  NAND U8924 ( .A(n5950), .B(n5949), .Z(n5951) );
  NAND U8925 ( .A(n5952), .B(n5951), .Z(n8039) );
  OR U8926 ( .A(n5954), .B(n5953), .Z(n5958) );
  NANDN U8927 ( .A(n5956), .B(n5955), .Z(n5957) );
  NAND U8928 ( .A(n5958), .B(n5957), .Z(n7719) );
  NANDN U8929 ( .A(n5960), .B(n5959), .Z(n5964) );
  NANDN U8930 ( .A(n5962), .B(n5961), .Z(n5963) );
  NAND U8931 ( .A(n5964), .B(n5963), .Z(n7716) );
  NANDN U8932 ( .A(n5966), .B(n5965), .Z(n5970) );
  NANDN U8933 ( .A(n5968), .B(n5967), .Z(n5969) );
  AND U8934 ( .A(n5970), .B(n5969), .Z(n7717) );
  XNOR U8935 ( .A(n7716), .B(n7717), .Z(n7718) );
  XNOR U8936 ( .A(n7719), .B(n7718), .Z(n8036) );
  NANDN U8937 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U8938 ( .A(n5974), .B(n5973), .Z(n5975) );
  AND U8939 ( .A(n5976), .B(n5975), .Z(n8037) );
  XNOR U8940 ( .A(n8036), .B(n8037), .Z(n8038) );
  XNOR U8941 ( .A(n8039), .B(n8038), .Z(n8179) );
  XNOR U8942 ( .A(n8178), .B(n8179), .Z(n8180) );
  XOR U8943 ( .A(n8181), .B(n8180), .Z(n8217) );
  XNOR U8944 ( .A(n8216), .B(n8217), .Z(n7689) );
  OR U8945 ( .A(n5978), .B(n5977), .Z(n5982) );
  NANDN U8946 ( .A(n5980), .B(n5979), .Z(n5981) );
  NAND U8947 ( .A(n5982), .B(n5981), .Z(n7707) );
  NANDN U8948 ( .A(n5984), .B(n5983), .Z(n5988) );
  NANDN U8949 ( .A(n5986), .B(n5985), .Z(n5987) );
  NAND U8950 ( .A(n5988), .B(n5987), .Z(n7704) );
  OR U8951 ( .A(n5990), .B(n5989), .Z(n5994) );
  NANDN U8952 ( .A(n5992), .B(n5991), .Z(n5993) );
  AND U8953 ( .A(n5994), .B(n5993), .Z(n7705) );
  XNOR U8954 ( .A(n7704), .B(n7705), .Z(n7706) );
  XNOR U8955 ( .A(n7707), .B(n7706), .Z(n7515) );
  NANDN U8956 ( .A(n5996), .B(n5995), .Z(n6000) );
  NAND U8957 ( .A(n5998), .B(n5997), .Z(n5999) );
  NAND U8958 ( .A(n6000), .B(n5999), .Z(n7514) );
  NANDN U8959 ( .A(n6002), .B(n6001), .Z(n6006) );
  NANDN U8960 ( .A(n6004), .B(n6003), .Z(n6005) );
  AND U8961 ( .A(n6006), .B(n6005), .Z(n7517) );
  XNOR U8962 ( .A(n7516), .B(n7517), .Z(n7814) );
  NANDN U8963 ( .A(n6008), .B(n6007), .Z(n6012) );
  NAND U8964 ( .A(n6010), .B(n6009), .Z(n6011) );
  NAND U8965 ( .A(n6012), .B(n6011), .Z(n7510) );
  NANDN U8966 ( .A(n6014), .B(n6013), .Z(n6018) );
  NANDN U8967 ( .A(n6016), .B(n6015), .Z(n6017) );
  AND U8968 ( .A(n6018), .B(n6017), .Z(n7508) );
  OR U8969 ( .A(n6020), .B(n6019), .Z(n6024) );
  NANDN U8970 ( .A(n6022), .B(n6021), .Z(n6023) );
  NAND U8971 ( .A(n6024), .B(n6023), .Z(n7547) );
  OR U8972 ( .A(n6026), .B(n6025), .Z(n6030) );
  NANDN U8973 ( .A(n6028), .B(n6027), .Z(n6029) );
  AND U8974 ( .A(n6030), .B(n6029), .Z(n7544) );
  NANDN U8975 ( .A(n6032), .B(n6031), .Z(n6036) );
  NANDN U8976 ( .A(n6034), .B(n6033), .Z(n6035) );
  AND U8977 ( .A(n6036), .B(n6035), .Z(n7545) );
  XOR U8978 ( .A(n7547), .B(n7546), .Z(n7509) );
  XOR U8979 ( .A(n7510), .B(n7511), .Z(n7812) );
  NANDN U8980 ( .A(n6038), .B(n6037), .Z(n6042) );
  NAND U8981 ( .A(n6040), .B(n6039), .Z(n6041) );
  NAND U8982 ( .A(n6042), .B(n6041), .Z(n7813) );
  XOR U8983 ( .A(n7812), .B(n7813), .Z(n7815) );
  XNOR U8984 ( .A(n7814), .B(n7815), .Z(n7421) );
  NANDN U8985 ( .A(n6044), .B(n6043), .Z(n6048) );
  NAND U8986 ( .A(n6046), .B(n6045), .Z(n6047) );
  NAND U8987 ( .A(n6048), .B(n6047), .Z(n7819) );
  OR U8988 ( .A(n6050), .B(n6049), .Z(n6054) );
  NANDN U8989 ( .A(n6052), .B(n6051), .Z(n6053) );
  NAND U8990 ( .A(n6054), .B(n6053), .Z(n8123) );
  XNOR U8991 ( .A(n8120), .B(n8121), .Z(n8122) );
  XNOR U8992 ( .A(n8123), .B(n8122), .Z(n7387) );
  OR U8993 ( .A(n6064), .B(n6063), .Z(n6068) );
  NANDN U8994 ( .A(n6066), .B(n6065), .Z(n6067) );
  NAND U8995 ( .A(n6068), .B(n6067), .Z(n8129) );
  XNOR U8996 ( .A(n8126), .B(n8127), .Z(n8128) );
  XOR U8997 ( .A(n8129), .B(n8128), .Z(n7386) );
  XNOR U8998 ( .A(n7387), .B(n7386), .Z(n7388) );
  OR U8999 ( .A(n6078), .B(n6077), .Z(n6082) );
  NANDN U9000 ( .A(n6080), .B(n6079), .Z(n6081) );
  NAND U9001 ( .A(n6082), .B(n6081), .Z(n7359) );
  NANDN U9002 ( .A(n6084), .B(n6083), .Z(n6088) );
  NANDN U9003 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U9004 ( .A(n6088), .B(n6087), .Z(n7356) );
  NANDN U9005 ( .A(n6090), .B(n6089), .Z(n6094) );
  NANDN U9006 ( .A(n6092), .B(n6091), .Z(n6093) );
  AND U9007 ( .A(n6094), .B(n6093), .Z(n7357) );
  XNOR U9008 ( .A(n7356), .B(n7357), .Z(n7358) );
  XOR U9009 ( .A(n7359), .B(n7358), .Z(n7389) );
  XOR U9010 ( .A(n7388), .B(n7389), .Z(n7818) );
  XNOR U9011 ( .A(n7819), .B(n7818), .Z(n7821) );
  OR U9012 ( .A(n6096), .B(n6095), .Z(n6100) );
  NANDN U9013 ( .A(n6098), .B(n6097), .Z(n6099) );
  NAND U9014 ( .A(n6100), .B(n6099), .Z(n7800) );
  NANDN U9015 ( .A(n6102), .B(n6101), .Z(n6106) );
  NANDN U9016 ( .A(n6104), .B(n6103), .Z(n6105) );
  NAND U9017 ( .A(n6106), .B(n6105), .Z(n7575) );
  NANDN U9018 ( .A(n6108), .B(n6107), .Z(n6112) );
  NANDN U9019 ( .A(n6110), .B(n6109), .Z(n6111) );
  AND U9020 ( .A(n6112), .B(n6111), .Z(n7572) );
  OR U9021 ( .A(n6114), .B(n6113), .Z(n6118) );
  NANDN U9022 ( .A(n6116), .B(n6115), .Z(n6117) );
  AND U9023 ( .A(n6118), .B(n6117), .Z(n7573) );
  XNOR U9024 ( .A(n7575), .B(n7574), .Z(n7801) );
  XNOR U9025 ( .A(n7800), .B(n7801), .Z(n7802) );
  NANDN U9026 ( .A(n6120), .B(n6119), .Z(n6124) );
  NANDN U9027 ( .A(n6122), .B(n6121), .Z(n6123) );
  NAND U9028 ( .A(n6124), .B(n6123), .Z(n7522) );
  OR U9029 ( .A(n6126), .B(n6125), .Z(n6130) );
  NANDN U9030 ( .A(n6128), .B(n6127), .Z(n6129) );
  AND U9031 ( .A(n6130), .B(n6129), .Z(n7520) );
  NANDN U9032 ( .A(n6132), .B(n6131), .Z(n6136) );
  NANDN U9033 ( .A(n6134), .B(n6133), .Z(n6135) );
  AND U9034 ( .A(n6136), .B(n6135), .Z(n7521) );
  XOR U9035 ( .A(n7522), .B(n7523), .Z(n7803) );
  XNOR U9036 ( .A(n7802), .B(n7803), .Z(n7820) );
  XOR U9037 ( .A(n7821), .B(n7820), .Z(n7418) );
  NANDN U9038 ( .A(n6138), .B(n6137), .Z(n6142) );
  NANDN U9039 ( .A(n6140), .B(n6139), .Z(n6141) );
  AND U9040 ( .A(n6142), .B(n6141), .Z(n7419) );
  XNOR U9041 ( .A(n7418), .B(n7419), .Z(n7420) );
  XNOR U9042 ( .A(n7421), .B(n7420), .Z(n7687) );
  NANDN U9043 ( .A(n6144), .B(n6143), .Z(n6148) );
  NANDN U9044 ( .A(n6146), .B(n6145), .Z(n6147) );
  NAND U9045 ( .A(n6148), .B(n6147), .Z(n7399) );
  NANDN U9046 ( .A(n6150), .B(n6149), .Z(n6154) );
  NAND U9047 ( .A(n6152), .B(n6151), .Z(n6153) );
  AND U9048 ( .A(n6154), .B(n6153), .Z(n7396) );
  XNOR U9049 ( .A(n7399), .B(n7398), .Z(n7779) );
  NANDN U9050 ( .A(n6160), .B(n6159), .Z(n6164) );
  NANDN U9051 ( .A(n6162), .B(n6161), .Z(n6163) );
  NAND U9052 ( .A(n6164), .B(n6163), .Z(n8372) );
  NANDN U9053 ( .A(n6166), .B(n6165), .Z(n6170) );
  NAND U9054 ( .A(n6168), .B(n6167), .Z(n6169) );
  NAND U9055 ( .A(n6170), .B(n6169), .Z(n8373) );
  XNOR U9056 ( .A(n8372), .B(n8373), .Z(n8374) );
  NANDN U9057 ( .A(n6172), .B(n6171), .Z(n6176) );
  NAND U9058 ( .A(n6174), .B(n6173), .Z(n6175) );
  AND U9059 ( .A(n6176), .B(n6175), .Z(n8375) );
  XNOR U9060 ( .A(n8374), .B(n8375), .Z(n7776) );
  NANDN U9061 ( .A(n6178), .B(n6177), .Z(n8365) );
  NANDN U9062 ( .A(n6180), .B(n6179), .Z(n6184) );
  NAND U9063 ( .A(n6182), .B(n6181), .Z(n6183) );
  NAND U9064 ( .A(n6184), .B(n6183), .Z(n8364) );
  XNOR U9065 ( .A(n8365), .B(n8364), .Z(n7404) );
  OR U9066 ( .A(n6186), .B(n6185), .Z(n6190) );
  NANDN U9067 ( .A(n6188), .B(n6187), .Z(n6189) );
  AND U9068 ( .A(n6190), .B(n6189), .Z(n7402) );
  NANDN U9069 ( .A(n6192), .B(n6191), .Z(n6196) );
  NANDN U9070 ( .A(n6194), .B(n6193), .Z(n6195) );
  AND U9071 ( .A(n6196), .B(n6195), .Z(n7403) );
  XOR U9072 ( .A(n7404), .B(n7405), .Z(n7777) );
  XOR U9073 ( .A(n7776), .B(n7777), .Z(n7778) );
  XOR U9074 ( .A(n7779), .B(n7778), .Z(n7935) );
  NANDN U9075 ( .A(n6198), .B(n6197), .Z(n6202) );
  NAND U9076 ( .A(n6200), .B(n6199), .Z(n6201) );
  NAND U9077 ( .A(n6202), .B(n6201), .Z(n8241) );
  OR U9078 ( .A(n6204), .B(n6203), .Z(n6208) );
  NANDN U9079 ( .A(n6206), .B(n6205), .Z(n6207) );
  NAND U9080 ( .A(n6208), .B(n6207), .Z(n8256) );
  NANDN U9081 ( .A(n6210), .B(n6209), .Z(n6214) );
  NANDN U9082 ( .A(n6212), .B(n6211), .Z(n6213) );
  AND U9083 ( .A(n6214), .B(n6213), .Z(n8257) );
  XNOR U9084 ( .A(n8256), .B(n8257), .Z(n8258) );
  OR U9085 ( .A(n6216), .B(n6215), .Z(n6220) );
  NAND U9086 ( .A(n6218), .B(n6217), .Z(n6219) );
  NAND U9087 ( .A(n6220), .B(n6219), .Z(n8259) );
  XOR U9088 ( .A(n8258), .B(n8259), .Z(n8238) );
  NANDN U9089 ( .A(n6222), .B(n6221), .Z(n6226) );
  NANDN U9090 ( .A(n6224), .B(n6223), .Z(n6225) );
  AND U9091 ( .A(n6226), .B(n6225), .Z(n8239) );
  XNOR U9092 ( .A(n8238), .B(n8239), .Z(n8240) );
  XNOR U9093 ( .A(n8241), .B(n8240), .Z(n7933) );
  NANDN U9094 ( .A(n6228), .B(n6227), .Z(n6232) );
  NAND U9095 ( .A(n6230), .B(n6229), .Z(n6231) );
  AND U9096 ( .A(n6232), .B(n6231), .Z(n7932) );
  XNOR U9097 ( .A(n7933), .B(n7932), .Z(n7934) );
  XNOR U9098 ( .A(n7935), .B(n7934), .Z(n8223) );
  NANDN U9099 ( .A(n6234), .B(n6233), .Z(n6238) );
  NANDN U9100 ( .A(n6236), .B(n6235), .Z(n6237) );
  NAND U9101 ( .A(n6238), .B(n6237), .Z(n8275) );
  OR U9102 ( .A(n6240), .B(n6239), .Z(n6244) );
  NANDN U9103 ( .A(n6242), .B(n6241), .Z(n6243) );
  NAND U9104 ( .A(n6244), .B(n6243), .Z(n7377) );
  NANDN U9105 ( .A(n6246), .B(n6245), .Z(n6250) );
  NANDN U9106 ( .A(n6248), .B(n6247), .Z(n6249) );
  NAND U9107 ( .A(n6250), .B(n6249), .Z(n7374) );
  OR U9108 ( .A(n6252), .B(n6251), .Z(n6256) );
  NANDN U9109 ( .A(n6254), .B(n6253), .Z(n6255) );
  AND U9110 ( .A(n6256), .B(n6255), .Z(n7375) );
  XNOR U9111 ( .A(n7374), .B(n7375), .Z(n7376) );
  XNOR U9112 ( .A(n7377), .B(n7376), .Z(n8272) );
  NANDN U9113 ( .A(n6258), .B(n6257), .Z(n6262) );
  NANDN U9114 ( .A(n6260), .B(n6259), .Z(n6261) );
  NAND U9115 ( .A(n6262), .B(n6261), .Z(n7347) );
  NANDN U9116 ( .A(n6264), .B(n6263), .Z(n6268) );
  NANDN U9117 ( .A(n6266), .B(n6265), .Z(n6267) );
  NAND U9118 ( .A(n6268), .B(n6267), .Z(n7344) );
  NANDN U9119 ( .A(n6270), .B(n6269), .Z(n6274) );
  NANDN U9120 ( .A(n6272), .B(n6271), .Z(n6273) );
  AND U9121 ( .A(n6274), .B(n6273), .Z(n7345) );
  XNOR U9122 ( .A(n7344), .B(n7345), .Z(n7346) );
  XOR U9123 ( .A(n7347), .B(n7346), .Z(n8273) );
  XNOR U9124 ( .A(n8272), .B(n8273), .Z(n8274) );
  XNOR U9125 ( .A(n8275), .B(n8274), .Z(n8075) );
  NANDN U9126 ( .A(n6276), .B(n6275), .Z(n6280) );
  NAND U9127 ( .A(n6278), .B(n6277), .Z(n6279) );
  NAND U9128 ( .A(n6280), .B(n6279), .Z(n7365) );
  NANDN U9129 ( .A(n6282), .B(n6281), .Z(n6286) );
  NAND U9130 ( .A(n6284), .B(n6283), .Z(n6285) );
  NAND U9131 ( .A(n6286), .B(n6285), .Z(n7362) );
  NANDN U9132 ( .A(n6288), .B(n6287), .Z(n6292) );
  NANDN U9133 ( .A(n6290), .B(n6289), .Z(n6291) );
  NAND U9134 ( .A(n6292), .B(n6291), .Z(n7568) );
  NANDN U9135 ( .A(n6294), .B(n6293), .Z(n6298) );
  NANDN U9136 ( .A(n6296), .B(n6295), .Z(n6297) );
  AND U9137 ( .A(n6298), .B(n6297), .Z(n7566) );
  NANDN U9138 ( .A(n6300), .B(n6299), .Z(n6304) );
  NANDN U9139 ( .A(n6302), .B(n6301), .Z(n6303) );
  AND U9140 ( .A(n6304), .B(n6303), .Z(n7567) );
  XOR U9141 ( .A(n7568), .B(n7569), .Z(n7363) );
  XOR U9142 ( .A(n7362), .B(n7363), .Z(n7364) );
  XOR U9143 ( .A(n7365), .B(n7364), .Z(n8072) );
  OR U9144 ( .A(n6306), .B(n6305), .Z(n6310) );
  NANDN U9145 ( .A(n6308), .B(n6307), .Z(n6309) );
  AND U9146 ( .A(n6310), .B(n6309), .Z(n8073) );
  XNOR U9147 ( .A(n8072), .B(n8073), .Z(n8074) );
  XOR U9148 ( .A(n8075), .B(n8074), .Z(n8220) );
  NANDN U9149 ( .A(n6312), .B(n6311), .Z(n6316) );
  NAND U9150 ( .A(n6314), .B(n6313), .Z(n6315) );
  AND U9151 ( .A(n6316), .B(n6315), .Z(n8221) );
  XNOR U9152 ( .A(n8220), .B(n8221), .Z(n8222) );
  XOR U9153 ( .A(n8223), .B(n8222), .Z(n7686) );
  XOR U9154 ( .A(n7687), .B(n7686), .Z(n7688) );
  XNOR U9155 ( .A(n7689), .B(n7688), .Z(n8291) );
  XNOR U9156 ( .A(n8290), .B(n8291), .Z(n8292) );
  NAND U9157 ( .A(n6318), .B(n6317), .Z(n6322) );
  NANDN U9158 ( .A(n6320), .B(n6319), .Z(n6321) );
  NAND U9159 ( .A(n6322), .B(n6321), .Z(n7680) );
  NANDN U9160 ( .A(n6324), .B(n6323), .Z(n6328) );
  NANDN U9161 ( .A(n6326), .B(n6325), .Z(n6327) );
  NAND U9162 ( .A(n6328), .B(n6327), .Z(n8009) );
  OR U9163 ( .A(n6330), .B(n6329), .Z(n6334) );
  NANDN U9164 ( .A(n6332), .B(n6331), .Z(n6333) );
  NAND U9165 ( .A(n6334), .B(n6333), .Z(n7737) );
  OR U9166 ( .A(n6336), .B(n6335), .Z(n6340) );
  NANDN U9167 ( .A(n6338), .B(n6337), .Z(n6339) );
  NAND U9168 ( .A(n6340), .B(n6339), .Z(n7734) );
  NANDN U9169 ( .A(n6342), .B(n6341), .Z(n6346) );
  NANDN U9170 ( .A(n6344), .B(n6343), .Z(n6345) );
  AND U9171 ( .A(n6346), .B(n6345), .Z(n7735) );
  XNOR U9172 ( .A(n7734), .B(n7735), .Z(n7736) );
  XNOR U9173 ( .A(n7737), .B(n7736), .Z(n8006) );
  NANDN U9174 ( .A(n6348), .B(n6347), .Z(n6352) );
  NAND U9175 ( .A(n6350), .B(n6349), .Z(n6351) );
  AND U9176 ( .A(n6352), .B(n6351), .Z(n8007) );
  XNOR U9177 ( .A(n8006), .B(n8007), .Z(n8008) );
  XNOR U9178 ( .A(n8009), .B(n8008), .Z(n7941) );
  OR U9179 ( .A(n6354), .B(n6353), .Z(n6358) );
  NAND U9180 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U9181 ( .A(n6358), .B(n6357), .Z(n7996) );
  OR U9182 ( .A(n6360), .B(n6359), .Z(n6364) );
  NAND U9183 ( .A(n6362), .B(n6361), .Z(n6363) );
  NAND U9184 ( .A(n6364), .B(n6363), .Z(n7995) );
  NANDN U9185 ( .A(n6366), .B(n6365), .Z(n6370) );
  NANDN U9186 ( .A(n6368), .B(n6367), .Z(n6369) );
  NAND U9187 ( .A(n6370), .B(n6369), .Z(n8349) );
  OR U9188 ( .A(n6372), .B(n6371), .Z(n6376) );
  NANDN U9189 ( .A(n6374), .B(n6373), .Z(n6375) );
  NAND U9190 ( .A(n6376), .B(n6375), .Z(n8346) );
  NANDN U9191 ( .A(n6378), .B(n6377), .Z(n6382) );
  NANDN U9192 ( .A(n6380), .B(n6379), .Z(n6381) );
  AND U9193 ( .A(n6382), .B(n6381), .Z(n8347) );
  XNOR U9194 ( .A(n8346), .B(n8347), .Z(n8348) );
  XOR U9195 ( .A(n8349), .B(n8348), .Z(n7994) );
  XOR U9196 ( .A(n7995), .B(n7994), .Z(n7997) );
  XNOR U9197 ( .A(n7996), .B(n7997), .Z(n7938) );
  OR U9198 ( .A(n6384), .B(n6383), .Z(n6388) );
  NANDN U9199 ( .A(n6386), .B(n6385), .Z(n6387) );
  NAND U9200 ( .A(n6388), .B(n6387), .Z(n8111) );
  NANDN U9201 ( .A(n6390), .B(n6389), .Z(n6394) );
  NANDN U9202 ( .A(n6392), .B(n6391), .Z(n6393) );
  NAND U9203 ( .A(n6394), .B(n6393), .Z(n8343) );
  NANDN U9204 ( .A(n6396), .B(n6395), .Z(n6400) );
  NANDN U9205 ( .A(n6398), .B(n6397), .Z(n6399) );
  NAND U9206 ( .A(n6400), .B(n6399), .Z(n8340) );
  OR U9207 ( .A(n6402), .B(n6401), .Z(n6406) );
  NANDN U9208 ( .A(n6404), .B(n6403), .Z(n6405) );
  AND U9209 ( .A(n6406), .B(n6405), .Z(n8341) );
  XNOR U9210 ( .A(n8340), .B(n8341), .Z(n8342) );
  XNOR U9211 ( .A(n8343), .B(n8342), .Z(n8108) );
  OR U9212 ( .A(n6408), .B(n6407), .Z(n6412) );
  NAND U9213 ( .A(n6410), .B(n6409), .Z(n6411) );
  AND U9214 ( .A(n6412), .B(n6411), .Z(n8109) );
  XNOR U9215 ( .A(n8108), .B(n8109), .Z(n8110) );
  XNOR U9216 ( .A(n8111), .B(n8110), .Z(n7939) );
  XNOR U9217 ( .A(n7938), .B(n7939), .Z(n7940) );
  XOR U9218 ( .A(n7941), .B(n7940), .Z(n7912) );
  NANDN U9219 ( .A(n6414), .B(n6413), .Z(n6418) );
  NANDN U9220 ( .A(n6416), .B(n6415), .Z(n6417) );
  NAND U9221 ( .A(n6418), .B(n6417), .Z(n8002) );
  NANDN U9222 ( .A(n6420), .B(n6419), .Z(n6424) );
  NANDN U9223 ( .A(n6422), .B(n6421), .Z(n6423) );
  NAND U9224 ( .A(n6424), .B(n6423), .Z(n8366) );
  NANDN U9225 ( .A(n6426), .B(n6425), .Z(n6430) );
  NAND U9226 ( .A(n6428), .B(n6427), .Z(n6429) );
  NAND U9227 ( .A(n6430), .B(n6429), .Z(n8367) );
  XNOR U9228 ( .A(n8366), .B(n8367), .Z(n8368) );
  NANDN U9229 ( .A(n6432), .B(n6431), .Z(n6436) );
  NAND U9230 ( .A(n6434), .B(n6433), .Z(n6435) );
  NAND U9231 ( .A(n6436), .B(n6435), .Z(n8369) );
  XNOR U9232 ( .A(n8368), .B(n8369), .Z(n8000) );
  OR U9233 ( .A(n6438), .B(n6437), .Z(n6442) );
  NANDN U9234 ( .A(n6440), .B(n6439), .Z(n6441) );
  AND U9235 ( .A(n6442), .B(n6441), .Z(n8001) );
  XOR U9236 ( .A(n8002), .B(n8003), .Z(n7603) );
  NANDN U9237 ( .A(n6444), .B(n6443), .Z(n6448) );
  NAND U9238 ( .A(n6446), .B(n6445), .Z(n6447) );
  NAND U9239 ( .A(n6448), .B(n6447), .Z(n8033) );
  NANDN U9240 ( .A(n6450), .B(n6449), .Z(n6454) );
  NAND U9241 ( .A(n6452), .B(n6451), .Z(n6453) );
  NAND U9242 ( .A(n6454), .B(n6453), .Z(n8031) );
  NANDN U9243 ( .A(n6456), .B(n6455), .Z(n6460) );
  NANDN U9244 ( .A(n6458), .B(n6457), .Z(n6459) );
  NAND U9245 ( .A(n6460), .B(n6459), .Z(n8358) );
  NANDN U9246 ( .A(n6462), .B(n6461), .Z(n6466) );
  NANDN U9247 ( .A(n6464), .B(n6463), .Z(n6465) );
  AND U9248 ( .A(n6466), .B(n6465), .Z(n8359) );
  XNOR U9249 ( .A(n8358), .B(n8359), .Z(n8360) );
  NANDN U9250 ( .A(n6468), .B(n6467), .Z(n6472) );
  NAND U9251 ( .A(n6470), .B(n6469), .Z(n6471) );
  AND U9252 ( .A(n6472), .B(n6471), .Z(n8361) );
  XOR U9253 ( .A(n8360), .B(n8361), .Z(n8030) );
  XNOR U9254 ( .A(n8031), .B(n8030), .Z(n8032) );
  XNOR U9255 ( .A(n8033), .B(n8032), .Z(n7602) );
  XOR U9256 ( .A(n7603), .B(n7602), .Z(n7604) );
  NANDN U9257 ( .A(n6474), .B(n6473), .Z(n6478) );
  NAND U9258 ( .A(n6476), .B(n6475), .Z(n6477) );
  NAND U9259 ( .A(n6478), .B(n6477), .Z(n8105) );
  NANDN U9260 ( .A(n6480), .B(n6479), .Z(n6484) );
  NAND U9261 ( .A(n6482), .B(n6481), .Z(n6483) );
  AND U9262 ( .A(n6484), .B(n6483), .Z(n7393) );
  OR U9263 ( .A(n6486), .B(n6485), .Z(n6490) );
  NANDN U9264 ( .A(n6488), .B(n6487), .Z(n6489) );
  NAND U9265 ( .A(n6490), .B(n6489), .Z(n7391) );
  OR U9266 ( .A(n6492), .B(n6491), .Z(n6496) );
  NANDN U9267 ( .A(n6494), .B(n6493), .Z(n6495) );
  NAND U9268 ( .A(n6496), .B(n6495), .Z(n7390) );
  XOR U9269 ( .A(n7391), .B(n7390), .Z(n7392) );
  XNOR U9270 ( .A(n7393), .B(n7392), .Z(n8103) );
  NANDN U9271 ( .A(n6498), .B(n6497), .Z(n6502) );
  NAND U9272 ( .A(n6500), .B(n6499), .Z(n6501) );
  NAND U9273 ( .A(n6502), .B(n6501), .Z(n8102) );
  XOR U9274 ( .A(n8103), .B(n8102), .Z(n8104) );
  XOR U9275 ( .A(n8105), .B(n8104), .Z(n7605) );
  XOR U9276 ( .A(n7604), .B(n7605), .Z(n7910) );
  OR U9277 ( .A(n6504), .B(n6503), .Z(n6508) );
  NAND U9278 ( .A(n6506), .B(n6505), .Z(n6507) );
  AND U9279 ( .A(n6508), .B(n6507), .Z(n7911) );
  XOR U9280 ( .A(n7910), .B(n7911), .Z(n6509) );
  XNOR U9281 ( .A(n7912), .B(n6509), .Z(n7681) );
  XNOR U9282 ( .A(n7680), .B(n7681), .Z(n7682) );
  OR U9283 ( .A(n6511), .B(n6510), .Z(n6515) );
  NAND U9284 ( .A(n6513), .B(n6512), .Z(n6514) );
  NAND U9285 ( .A(n6515), .B(n6514), .Z(n7918) );
  OR U9286 ( .A(n6517), .B(n6516), .Z(n6521) );
  NANDN U9287 ( .A(n6519), .B(n6518), .Z(n6520) );
  NAND U9288 ( .A(n6521), .B(n6520), .Z(n7917) );
  NANDN U9289 ( .A(n6523), .B(n6522), .Z(n6527) );
  NANDN U9290 ( .A(n6525), .B(n6524), .Z(n6526) );
  NAND U9291 ( .A(n6527), .B(n6526), .Z(n8147) );
  NANDN U9292 ( .A(n6529), .B(n6528), .Z(n6533) );
  NANDN U9293 ( .A(n6531), .B(n6530), .Z(n6532) );
  NAND U9294 ( .A(n6533), .B(n6532), .Z(n8144) );
  NANDN U9295 ( .A(n6535), .B(n6534), .Z(n6539) );
  NANDN U9296 ( .A(n6537), .B(n6536), .Z(n6538) );
  AND U9297 ( .A(n6539), .B(n6538), .Z(n8145) );
  XNOR U9298 ( .A(n8144), .B(n8145), .Z(n8146) );
  XOR U9299 ( .A(n8147), .B(n8146), .Z(n7916) );
  XOR U9300 ( .A(n7917), .B(n7916), .Z(n7919) );
  XOR U9301 ( .A(n7918), .B(n7919), .Z(n7915) );
  OR U9302 ( .A(n6541), .B(n6540), .Z(n6545) );
  NANDN U9303 ( .A(n6543), .B(n6542), .Z(n6544) );
  NAND U9304 ( .A(n6545), .B(n6544), .Z(n7581) );
  OR U9305 ( .A(n6547), .B(n6546), .Z(n6551) );
  NANDN U9306 ( .A(n6549), .B(n6548), .Z(n6550) );
  NAND U9307 ( .A(n6551), .B(n6550), .Z(n7578) );
  NANDN U9308 ( .A(n6553), .B(n6552), .Z(n6557) );
  NANDN U9309 ( .A(n6555), .B(n6554), .Z(n6556) );
  AND U9310 ( .A(n6557), .B(n6556), .Z(n7579) );
  XNOR U9311 ( .A(n7578), .B(n7579), .Z(n7580) );
  XNOR U9312 ( .A(n7581), .B(n7580), .Z(n8158) );
  NANDN U9313 ( .A(n6559), .B(n6558), .Z(n6563) );
  NANDN U9314 ( .A(n6561), .B(n6560), .Z(n6562) );
  NAND U9315 ( .A(n6563), .B(n6562), .Z(n7433) );
  NANDN U9316 ( .A(n6565), .B(n6564), .Z(n6569) );
  NANDN U9317 ( .A(n6567), .B(n6566), .Z(n6568) );
  NAND U9318 ( .A(n6569), .B(n6568), .Z(n7430) );
  OR U9319 ( .A(n6571), .B(n6570), .Z(n6575) );
  NANDN U9320 ( .A(n6573), .B(n6572), .Z(n6574) );
  AND U9321 ( .A(n6575), .B(n6574), .Z(n7431) );
  XNOR U9322 ( .A(n7430), .B(n7431), .Z(n7432) );
  XNOR U9323 ( .A(n7433), .B(n7432), .Z(n8157) );
  NANDN U9324 ( .A(n6577), .B(n6576), .Z(n6581) );
  NANDN U9325 ( .A(n6579), .B(n6578), .Z(n6580) );
  NAND U9326 ( .A(n6581), .B(n6580), .Z(n7371) );
  NANDN U9327 ( .A(n6583), .B(n6582), .Z(n6587) );
  NANDN U9328 ( .A(n6585), .B(n6584), .Z(n6586) );
  NAND U9329 ( .A(n6587), .B(n6586), .Z(n7368) );
  NANDN U9330 ( .A(n6589), .B(n6588), .Z(n6593) );
  NANDN U9331 ( .A(n6591), .B(n6590), .Z(n6592) );
  AND U9332 ( .A(n6593), .B(n6592), .Z(n7369) );
  XNOR U9333 ( .A(n7368), .B(n7369), .Z(n7370) );
  XOR U9334 ( .A(n7371), .B(n7370), .Z(n8156) );
  XOR U9335 ( .A(n8157), .B(n8156), .Z(n8159) );
  XNOR U9336 ( .A(n8158), .B(n8159), .Z(n7913) );
  OR U9337 ( .A(n6595), .B(n6594), .Z(n6599) );
  NANDN U9338 ( .A(n6597), .B(n6596), .Z(n6598) );
  NAND U9339 ( .A(n6599), .B(n6598), .Z(n8171) );
  OR U9340 ( .A(n6601), .B(n6600), .Z(n6605) );
  NANDN U9341 ( .A(n6603), .B(n6602), .Z(n6604) );
  NAND U9342 ( .A(n6605), .B(n6604), .Z(n7439) );
  NANDN U9343 ( .A(n6607), .B(n6606), .Z(n6611) );
  NANDN U9344 ( .A(n6609), .B(n6608), .Z(n6610) );
  NAND U9345 ( .A(n6611), .B(n6610), .Z(n7436) );
  OR U9346 ( .A(n6613), .B(n6612), .Z(n6617) );
  NANDN U9347 ( .A(n6615), .B(n6614), .Z(n6616) );
  AND U9348 ( .A(n6617), .B(n6616), .Z(n7437) );
  XNOR U9349 ( .A(n7436), .B(n7437), .Z(n7438) );
  XNOR U9350 ( .A(n7439), .B(n7438), .Z(n8169) );
  OR U9351 ( .A(n6619), .B(n6618), .Z(n6623) );
  NAND U9352 ( .A(n6621), .B(n6620), .Z(n6622) );
  AND U9353 ( .A(n6623), .B(n6622), .Z(n8168) );
  XNOR U9354 ( .A(n8169), .B(n8168), .Z(n8170) );
  XNOR U9355 ( .A(n8171), .B(n8170), .Z(n7914) );
  XOR U9356 ( .A(n7913), .B(n7914), .Z(n6624) );
  XNOR U9357 ( .A(n7915), .B(n6624), .Z(n7887) );
  OR U9358 ( .A(n6626), .B(n6625), .Z(n6630) );
  NANDN U9359 ( .A(n6628), .B(n6627), .Z(n6629) );
  NAND U9360 ( .A(n6630), .B(n6629), .Z(n7863) );
  OR U9361 ( .A(n6632), .B(n6631), .Z(n6636) );
  NANDN U9362 ( .A(n6634), .B(n6633), .Z(n6635) );
  NAND U9363 ( .A(n6636), .B(n6635), .Z(n7499) );
  OR U9364 ( .A(n6638), .B(n6637), .Z(n6642) );
  NANDN U9365 ( .A(n6640), .B(n6639), .Z(n6641) );
  NAND U9366 ( .A(n6642), .B(n6641), .Z(n7496) );
  NANDN U9367 ( .A(n6644), .B(n6643), .Z(n6648) );
  NAND U9368 ( .A(n6646), .B(n6645), .Z(n6647) );
  NAND U9369 ( .A(n6648), .B(n6647), .Z(n7497) );
  XNOR U9370 ( .A(n7496), .B(n7497), .Z(n7498) );
  XNOR U9371 ( .A(n7499), .B(n7498), .Z(n7861) );
  OR U9372 ( .A(n6650), .B(n6649), .Z(n6654) );
  NANDN U9373 ( .A(n6652), .B(n6651), .Z(n6653) );
  AND U9374 ( .A(n6654), .B(n6653), .Z(n7860) );
  XNOR U9375 ( .A(n7861), .B(n7860), .Z(n7862) );
  XOR U9376 ( .A(n7863), .B(n7862), .Z(n7931) );
  OR U9377 ( .A(n6656), .B(n6655), .Z(n6660) );
  NANDN U9378 ( .A(n6658), .B(n6657), .Z(n6659) );
  NAND U9379 ( .A(n6660), .B(n6659), .Z(n7353) );
  NANDN U9380 ( .A(n6662), .B(n6661), .Z(n6666) );
  NANDN U9381 ( .A(n6664), .B(n6663), .Z(n6665) );
  NAND U9382 ( .A(n6666), .B(n6665), .Z(n7350) );
  OR U9383 ( .A(n6668), .B(n6667), .Z(n6672) );
  NANDN U9384 ( .A(n6670), .B(n6669), .Z(n6671) );
  AND U9385 ( .A(n6672), .B(n6671), .Z(n7351) );
  XNOR U9386 ( .A(n7350), .B(n7351), .Z(n7352) );
  XOR U9387 ( .A(n7353), .B(n7352), .Z(n7927) );
  OR U9388 ( .A(n6674), .B(n6673), .Z(n6678) );
  NANDN U9389 ( .A(n6676), .B(n6675), .Z(n6677) );
  NAND U9390 ( .A(n6678), .B(n6677), .Z(n7490) );
  OR U9391 ( .A(n6680), .B(n6679), .Z(n6684) );
  NANDN U9392 ( .A(n6682), .B(n6681), .Z(n6683) );
  AND U9393 ( .A(n6684), .B(n6683), .Z(n7491) );
  XNOR U9394 ( .A(n7490), .B(n7491), .Z(n7492) );
  NANDN U9395 ( .A(n6686), .B(n6685), .Z(n6690) );
  NAND U9396 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U9397 ( .A(n6690), .B(n6689), .Z(n7493) );
  XNOR U9398 ( .A(n7492), .B(n7493), .Z(n7925) );
  NANDN U9399 ( .A(n6692), .B(n6691), .Z(n6696) );
  NANDN U9400 ( .A(n6694), .B(n6693), .Z(n6695) );
  NAND U9401 ( .A(n6696), .B(n6695), .Z(n7761) );
  NANDN U9402 ( .A(n6698), .B(n6697), .Z(n6702) );
  NANDN U9403 ( .A(n6700), .B(n6699), .Z(n6701) );
  NAND U9404 ( .A(n6702), .B(n6701), .Z(n7758) );
  OR U9405 ( .A(n6704), .B(n6703), .Z(n6708) );
  NANDN U9406 ( .A(n6706), .B(n6705), .Z(n6707) );
  AND U9407 ( .A(n6708), .B(n6707), .Z(n7759) );
  XNOR U9408 ( .A(n7758), .B(n7759), .Z(n7760) );
  XNOR U9409 ( .A(n7761), .B(n7760), .Z(n7926) );
  XOR U9410 ( .A(n7925), .B(n7926), .Z(n6709) );
  XOR U9411 ( .A(n7927), .B(n6709), .Z(n7928) );
  OR U9412 ( .A(n6711), .B(n6710), .Z(n6715) );
  NANDN U9413 ( .A(n6713), .B(n6712), .Z(n6714) );
  NAND U9414 ( .A(n6715), .B(n6714), .Z(n8099) );
  NANDN U9415 ( .A(n6717), .B(n6716), .Z(n6721) );
  NANDN U9416 ( .A(n6719), .B(n6718), .Z(n6720) );
  NAND U9417 ( .A(n6721), .B(n6720), .Z(n8096) );
  NANDN U9418 ( .A(n6723), .B(n6722), .Z(n6727) );
  NAND U9419 ( .A(n6725), .B(n6724), .Z(n6726) );
  NAND U9420 ( .A(n6727), .B(n6726), .Z(n8117) );
  NANDN U9421 ( .A(n6729), .B(n6728), .Z(n6733) );
  NANDN U9422 ( .A(n6731), .B(n6730), .Z(n6732) );
  AND U9423 ( .A(n6733), .B(n6732), .Z(n8114) );
  NANDN U9424 ( .A(n6735), .B(n6734), .Z(n6739) );
  NANDN U9425 ( .A(n6737), .B(n6736), .Z(n6738) );
  AND U9426 ( .A(n6739), .B(n6738), .Z(n8115) );
  XOR U9427 ( .A(n8114), .B(n8115), .Z(n8116) );
  XNOR U9428 ( .A(n8117), .B(n8116), .Z(n8097) );
  XNOR U9429 ( .A(n8096), .B(n8097), .Z(n8098) );
  XNOR U9430 ( .A(n8099), .B(n8098), .Z(n7929) );
  XNOR U9431 ( .A(n7928), .B(n7929), .Z(n7930) );
  XNOR U9432 ( .A(n7931), .B(n7930), .Z(n7884) );
  NANDN U9433 ( .A(n6741), .B(n6740), .Z(n6745) );
  NAND U9434 ( .A(n6743), .B(n6742), .Z(n6744) );
  AND U9435 ( .A(n6745), .B(n6744), .Z(n7885) );
  XNOR U9436 ( .A(n7884), .B(n7885), .Z(n7886) );
  XNOR U9437 ( .A(n7887), .B(n7886), .Z(n7683) );
  XNOR U9438 ( .A(n7682), .B(n7683), .Z(n8293) );
  XOR U9439 ( .A(n8292), .B(n8293), .Z(n7700) );
  XNOR U9440 ( .A(n7701), .B(n7700), .Z(n7315) );
  NAND U9441 ( .A(n6747), .B(n6746), .Z(n6751) );
  OR U9442 ( .A(n6749), .B(n6748), .Z(n6750) );
  AND U9443 ( .A(n6751), .B(n6750), .Z(n7314) );
  XOR U9444 ( .A(n7315), .B(n7314), .Z(n7316) );
  NANDN U9445 ( .A(n6753), .B(n6752), .Z(n6757) );
  NAND U9446 ( .A(n6755), .B(n6754), .Z(n6756) );
  NAND U9447 ( .A(n6757), .B(n6756), .Z(n8423) );
  NANDN U9448 ( .A(n6759), .B(n6758), .Z(n6763) );
  NAND U9449 ( .A(n6761), .B(n6760), .Z(n6762) );
  NAND U9450 ( .A(n6763), .B(n6762), .Z(n8421) );
  NANDN U9451 ( .A(n6765), .B(n6764), .Z(n6769) );
  NAND U9452 ( .A(n6767), .B(n6766), .Z(n6768) );
  AND U9453 ( .A(n6769), .B(n6768), .Z(n8420) );
  XNOR U9454 ( .A(n8421), .B(n8420), .Z(n8422) );
  XOR U9455 ( .A(n8423), .B(n8422), .Z(n7640) );
  NAND U9456 ( .A(n6771), .B(n6770), .Z(n6775) );
  OR U9457 ( .A(n6773), .B(n6772), .Z(n6774) );
  NAND U9458 ( .A(n6775), .B(n6774), .Z(n7641) );
  XNOR U9459 ( .A(n7640), .B(n7641), .Z(n7642) );
  NANDN U9460 ( .A(n6777), .B(n6776), .Z(n6781) );
  NAND U9461 ( .A(n6779), .B(n6778), .Z(n6780) );
  NAND U9462 ( .A(n6781), .B(n6780), .Z(n7643) );
  XOR U9463 ( .A(n7642), .B(n7643), .Z(n8309) );
  NAND U9464 ( .A(n6783), .B(n6782), .Z(n6787) );
  NAND U9465 ( .A(n6785), .B(n6784), .Z(n6786) );
  NAND U9466 ( .A(n6787), .B(n6786), .Z(n8307) );
  XNOR U9467 ( .A(n8307), .B(n8306), .Z(n8308) );
  XNOR U9468 ( .A(n8309), .B(n8308), .Z(n7329) );
  NANDN U9469 ( .A(n6793), .B(n6792), .Z(n6797) );
  NAND U9470 ( .A(n6795), .B(n6794), .Z(n6796) );
  NAND U9471 ( .A(n6797), .B(n6796), .Z(n7327) );
  OR U9472 ( .A(n6799), .B(n6798), .Z(n6803) );
  NAND U9473 ( .A(n6801), .B(n6800), .Z(n6802) );
  NAND U9474 ( .A(n6803), .B(n6802), .Z(n7599) );
  OR U9475 ( .A(n6805), .B(n6804), .Z(n6809) );
  NANDN U9476 ( .A(n6807), .B(n6806), .Z(n6808) );
  NAND U9477 ( .A(n6809), .B(n6808), .Z(n8414) );
  NANDN U9478 ( .A(n6811), .B(n6810), .Z(n6815) );
  NAND U9479 ( .A(n6813), .B(n6812), .Z(n6814) );
  NAND U9480 ( .A(n6815), .B(n6814), .Z(n8415) );
  XNOR U9481 ( .A(n8414), .B(n8415), .Z(n8416) );
  NANDN U9482 ( .A(n6817), .B(n6816), .Z(n6821) );
  NAND U9483 ( .A(n6819), .B(n6818), .Z(n6820) );
  NAND U9484 ( .A(n6821), .B(n6820), .Z(n8417) );
  XOR U9485 ( .A(n8416), .B(n8417), .Z(n7596) );
  NAND U9486 ( .A(n6823), .B(n6822), .Z(n6827) );
  NANDN U9487 ( .A(n6825), .B(n6824), .Z(n6826) );
  NAND U9488 ( .A(n6827), .B(n6826), .Z(n7597) );
  XNOR U9489 ( .A(n7596), .B(n7597), .Z(n7598) );
  XNOR U9490 ( .A(n7599), .B(n7598), .Z(n8446) );
  NAND U9491 ( .A(n6829), .B(n6828), .Z(n6833) );
  NANDN U9492 ( .A(n6831), .B(n6830), .Z(n6832) );
  NAND U9493 ( .A(n6833), .B(n6832), .Z(n8321) );
  NANDN U9494 ( .A(n6835), .B(n6834), .Z(n6839) );
  NAND U9495 ( .A(n6837), .B(n6836), .Z(n6838) );
  NAND U9496 ( .A(n6839), .B(n6838), .Z(n8319) );
  NANDN U9497 ( .A(n6841), .B(n6840), .Z(n6845) );
  NAND U9498 ( .A(n6843), .B(n6842), .Z(n6844) );
  NAND U9499 ( .A(n6845), .B(n6844), .Z(n7609) );
  NANDN U9500 ( .A(n6847), .B(n6846), .Z(n6851) );
  NANDN U9501 ( .A(n6849), .B(n6848), .Z(n6850) );
  NAND U9502 ( .A(n6851), .B(n6850), .Z(n7606) );
  NANDN U9503 ( .A(n6853), .B(n6852), .Z(n6857) );
  NAND U9504 ( .A(n6855), .B(n6854), .Z(n6856) );
  NAND U9505 ( .A(n6857), .B(n6856), .Z(n7607) );
  XNOR U9506 ( .A(n7606), .B(n7607), .Z(n7608) );
  XNOR U9507 ( .A(n7609), .B(n7608), .Z(n8318) );
  XOR U9508 ( .A(n8319), .B(n8318), .Z(n8320) );
  XNOR U9509 ( .A(n8321), .B(n8320), .Z(n8444) );
  NAND U9510 ( .A(n6863), .B(n6862), .Z(n6867) );
  OR U9511 ( .A(n6865), .B(n6864), .Z(n6866) );
  NAND U9512 ( .A(n6867), .B(n6866), .Z(n7424) );
  NANDN U9513 ( .A(n6869), .B(n6868), .Z(n6873) );
  OR U9514 ( .A(n6871), .B(n6870), .Z(n6872) );
  NAND U9515 ( .A(n6873), .B(n6872), .Z(n7615) );
  NANDN U9516 ( .A(n6875), .B(n6874), .Z(n6879) );
  NANDN U9517 ( .A(n6877), .B(n6876), .Z(n6878) );
  NAND U9518 ( .A(n6879), .B(n6878), .Z(n7612) );
  NANDN U9519 ( .A(n6881), .B(n6880), .Z(n6885) );
  NAND U9520 ( .A(n6883), .B(n6882), .Z(n6884) );
  NAND U9521 ( .A(n6885), .B(n6884), .Z(n7613) );
  XNOR U9522 ( .A(n7612), .B(n7613), .Z(n7614) );
  XOR U9523 ( .A(n7615), .B(n7614), .Z(n7425) );
  XNOR U9524 ( .A(n7424), .B(n7425), .Z(n7426) );
  XNOR U9525 ( .A(n7427), .B(n7426), .Z(n8445) );
  XOR U9526 ( .A(n8444), .B(n8445), .Z(n8447) );
  XOR U9527 ( .A(n8446), .B(n8447), .Z(n7326) );
  XNOR U9528 ( .A(n7327), .B(n7326), .Z(n7328) );
  XNOR U9529 ( .A(n7329), .B(n7328), .Z(n8303) );
  OR U9530 ( .A(n6887), .B(n6886), .Z(n6891) );
  OR U9531 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U9532 ( .A(n6891), .B(n6890), .Z(n8300) );
  OR U9533 ( .A(n6893), .B(n6892), .Z(n6897) );
  NAND U9534 ( .A(n6895), .B(n6894), .Z(n6896) );
  NAND U9535 ( .A(n6897), .B(n6896), .Z(n7773) );
  NANDN U9536 ( .A(n6899), .B(n6898), .Z(n6903) );
  NANDN U9537 ( .A(n6901), .B(n6900), .Z(n6902) );
  NAND U9538 ( .A(n6903), .B(n6902), .Z(n7770) );
  NANDN U9539 ( .A(n6905), .B(n6904), .Z(n6909) );
  NAND U9540 ( .A(n6907), .B(n6906), .Z(n6908) );
  AND U9541 ( .A(n6909), .B(n6908), .Z(n7771) );
  XNOR U9542 ( .A(n7770), .B(n7771), .Z(n7772) );
  XNOR U9543 ( .A(n7773), .B(n7772), .Z(n7873) );
  NANDN U9544 ( .A(n6911), .B(n6910), .Z(n6915) );
  NANDN U9545 ( .A(n6913), .B(n6912), .Z(n6914) );
  NAND U9546 ( .A(n6915), .B(n6914), .Z(n7947) );
  NANDN U9547 ( .A(n6917), .B(n6916), .Z(n6921) );
  NANDN U9548 ( .A(n6919), .B(n6918), .Z(n6920) );
  AND U9549 ( .A(n6921), .B(n6920), .Z(n7944) );
  OR U9550 ( .A(n6923), .B(n6922), .Z(n6927) );
  NAND U9551 ( .A(n6925), .B(n6924), .Z(n6926) );
  AND U9552 ( .A(n6927), .B(n6926), .Z(n7945) );
  XNOR U9553 ( .A(n7947), .B(n7946), .Z(n7871) );
  NANDN U9554 ( .A(n6929), .B(n6928), .Z(n6933) );
  NAND U9555 ( .A(n6931), .B(n6930), .Z(n6932) );
  AND U9556 ( .A(n6933), .B(n6932), .Z(n7870) );
  XNOR U9557 ( .A(n7871), .B(n7870), .Z(n7872) );
  XOR U9558 ( .A(n7873), .B(n7872), .Z(n7883) );
  NANDN U9559 ( .A(n6935), .B(n6934), .Z(n6939) );
  NANDN U9560 ( .A(n6937), .B(n6936), .Z(n6938) );
  AND U9561 ( .A(n6939), .B(n6938), .Z(n7880) );
  NANDN U9562 ( .A(n6945), .B(n6944), .Z(n6949) );
  NAND U9563 ( .A(n6947), .B(n6946), .Z(n6948) );
  NAND U9564 ( .A(n6949), .B(n6948), .Z(n7969) );
  NANDN U9565 ( .A(n6951), .B(n6950), .Z(n6955) );
  NAND U9566 ( .A(n6953), .B(n6952), .Z(n6954) );
  NAND U9567 ( .A(n6955), .B(n6954), .Z(n8093) );
  NANDN U9568 ( .A(n6957), .B(n6956), .Z(n6961) );
  NAND U9569 ( .A(n6959), .B(n6958), .Z(n6960) );
  NAND U9570 ( .A(n6961), .B(n6960), .Z(n8090) );
  OR U9571 ( .A(n6963), .B(n6962), .Z(n6967) );
  NANDN U9572 ( .A(n6965), .B(n6964), .Z(n6966) );
  AND U9573 ( .A(n6967), .B(n6966), .Z(n8091) );
  XNOR U9574 ( .A(n8090), .B(n8091), .Z(n8092) );
  XOR U9575 ( .A(n8093), .B(n8092), .Z(n7968) );
  XNOR U9576 ( .A(n7969), .B(n7968), .Z(n7970) );
  XOR U9577 ( .A(n7971), .B(n7970), .Z(n7881) );
  XOR U9578 ( .A(n7880), .B(n7881), .Z(n7882) );
  XOR U9579 ( .A(n7883), .B(n7882), .Z(n7985) );
  NANDN U9580 ( .A(n6969), .B(n6968), .Z(n6973) );
  NANDN U9581 ( .A(n6971), .B(n6970), .Z(n6972) );
  AND U9582 ( .A(n6973), .B(n6972), .Z(n8050) );
  OR U9583 ( .A(n6975), .B(n6974), .Z(n6979) );
  NANDN U9584 ( .A(n6977), .B(n6976), .Z(n6978) );
  NAND U9585 ( .A(n6979), .B(n6978), .Z(n7535) );
  OR U9586 ( .A(n6981), .B(n6980), .Z(n6985) );
  NANDN U9587 ( .A(n6983), .B(n6982), .Z(n6984) );
  NAND U9588 ( .A(n6985), .B(n6984), .Z(n7532) );
  OR U9589 ( .A(n6987), .B(n6986), .Z(n6991) );
  NANDN U9590 ( .A(n6989), .B(n6988), .Z(n6990) );
  AND U9591 ( .A(n6991), .B(n6990), .Z(n7533) );
  XNOR U9592 ( .A(n7532), .B(n7533), .Z(n7534) );
  XNOR U9593 ( .A(n7535), .B(n7534), .Z(n8048) );
  NANDN U9594 ( .A(n6993), .B(n6992), .Z(n6997) );
  NAND U9595 ( .A(n6995), .B(n6994), .Z(n6996) );
  AND U9596 ( .A(n6997), .B(n6996), .Z(n8049) );
  XOR U9597 ( .A(n8048), .B(n8049), .Z(n8051) );
  NANDN U9598 ( .A(n6999), .B(n6998), .Z(n7003) );
  NANDN U9599 ( .A(n7001), .B(n7000), .Z(n7002) );
  NAND U9600 ( .A(n7003), .B(n7002), .Z(n8140) );
  NANDN U9601 ( .A(n7005), .B(n7004), .Z(n7009) );
  NANDN U9602 ( .A(n7007), .B(n7006), .Z(n7008) );
  AND U9603 ( .A(n7009), .B(n7008), .Z(n8138) );
  NANDN U9604 ( .A(n7011), .B(n7010), .Z(n7015) );
  NANDN U9605 ( .A(n7013), .B(n7012), .Z(n7014) );
  AND U9606 ( .A(n7015), .B(n7014), .Z(n8139) );
  XOR U9607 ( .A(n8140), .B(n8141), .Z(n8381) );
  NANDN U9608 ( .A(n7017), .B(n7016), .Z(n7021) );
  NANDN U9609 ( .A(n7019), .B(n7018), .Z(n7020) );
  NAND U9610 ( .A(n7021), .B(n7020), .Z(n7456) );
  NANDN U9611 ( .A(n7023), .B(n7022), .Z(n7027) );
  NANDN U9612 ( .A(n7025), .B(n7024), .Z(n7026) );
  NAND U9613 ( .A(n7027), .B(n7026), .Z(n7454) );
  OR U9614 ( .A(n7029), .B(n7028), .Z(n7033) );
  NANDN U9615 ( .A(n7031), .B(n7030), .Z(n7032) );
  NAND U9616 ( .A(n7033), .B(n7032), .Z(n7455) );
  XNOR U9617 ( .A(n7454), .B(n7455), .Z(n7034) );
  XOR U9618 ( .A(n7456), .B(n7034), .Z(n8378) );
  NANDN U9619 ( .A(n7036), .B(n7035), .Z(n7040) );
  NAND U9620 ( .A(n7038), .B(n7037), .Z(n7039) );
  NAND U9621 ( .A(n7040), .B(n7039), .Z(n8379) );
  XOR U9622 ( .A(n8378), .B(n8379), .Z(n8380) );
  XOR U9623 ( .A(n8381), .B(n8380), .Z(n8019) );
  NANDN U9624 ( .A(n7042), .B(n7041), .Z(n7046) );
  NANDN U9625 ( .A(n7044), .B(n7043), .Z(n7045) );
  NAND U9626 ( .A(n7046), .B(n7045), .Z(n7450) );
  NANDN U9627 ( .A(n7048), .B(n7047), .Z(n7052) );
  NANDN U9628 ( .A(n7050), .B(n7049), .Z(n7051) );
  AND U9629 ( .A(n7052), .B(n7051), .Z(n7448) );
  NANDN U9630 ( .A(n7054), .B(n7053), .Z(n7058) );
  NANDN U9631 ( .A(n7056), .B(n7055), .Z(n7057) );
  AND U9632 ( .A(n7058), .B(n7057), .Z(n7449) );
  XOR U9633 ( .A(n7450), .B(n7451), .Z(n7411) );
  OR U9634 ( .A(n7060), .B(n7059), .Z(n7064) );
  NANDN U9635 ( .A(n7062), .B(n7061), .Z(n7063) );
  NAND U9636 ( .A(n7064), .B(n7063), .Z(n7459) );
  OR U9637 ( .A(n7066), .B(n7065), .Z(n7070) );
  NANDN U9638 ( .A(n7068), .B(n7067), .Z(n7069) );
  NAND U9639 ( .A(n7070), .B(n7069), .Z(n7457) );
  OR U9640 ( .A(n7072), .B(n7071), .Z(n7076) );
  NANDN U9641 ( .A(n7074), .B(n7073), .Z(n7075) );
  NAND U9642 ( .A(n7076), .B(n7075), .Z(n7458) );
  XNOR U9643 ( .A(n7457), .B(n7458), .Z(n7077) );
  XOR U9644 ( .A(n7459), .B(n7077), .Z(n7408) );
  NANDN U9645 ( .A(n7079), .B(n7078), .Z(n7083) );
  NAND U9646 ( .A(n7081), .B(n7080), .Z(n7082) );
  AND U9647 ( .A(n7083), .B(n7082), .Z(n7409) );
  XOR U9648 ( .A(n7408), .B(n7409), .Z(n7410) );
  XOR U9649 ( .A(n7411), .B(n7410), .Z(n8018) );
  XOR U9650 ( .A(n8019), .B(n8018), .Z(n8020) );
  XOR U9651 ( .A(n8021), .B(n8020), .Z(n7897) );
  NANDN U9652 ( .A(n7085), .B(n7084), .Z(n7089) );
  NAND U9653 ( .A(n7087), .B(n7086), .Z(n7088) );
  NAND U9654 ( .A(n7089), .B(n7088), .Z(n8177) );
  NANDN U9655 ( .A(n7091), .B(n7090), .Z(n7095) );
  NANDN U9656 ( .A(n7093), .B(n7092), .Z(n7094) );
  NAND U9657 ( .A(n7095), .B(n7094), .Z(n7481) );
  NAND U9658 ( .A(n7097), .B(n7096), .Z(n7101) );
  OR U9659 ( .A(n7099), .B(n7098), .Z(n7100) );
  NAND U9660 ( .A(n7101), .B(n7100), .Z(n7478) );
  OR U9661 ( .A(n7103), .B(n7102), .Z(n7107) );
  NANDN U9662 ( .A(n7105), .B(n7104), .Z(n7106) );
  AND U9663 ( .A(n7107), .B(n7106), .Z(n7479) );
  XNOR U9664 ( .A(n7478), .B(n7479), .Z(n7480) );
  XNOR U9665 ( .A(n7481), .B(n7480), .Z(n8174) );
  OR U9666 ( .A(n7109), .B(n7108), .Z(n7113) );
  NANDN U9667 ( .A(n7111), .B(n7110), .Z(n7112) );
  NAND U9668 ( .A(n7113), .B(n7112), .Z(n8175) );
  XNOR U9669 ( .A(n8174), .B(n8175), .Z(n8176) );
  XNOR U9670 ( .A(n8177), .B(n8176), .Z(n7895) );
  NANDN U9671 ( .A(n7119), .B(n7118), .Z(n7123) );
  NAND U9672 ( .A(n7121), .B(n7120), .Z(n7122) );
  NAND U9673 ( .A(n7123), .B(n7122), .Z(n8325) );
  OR U9674 ( .A(n7125), .B(n7124), .Z(n7129) );
  NANDN U9675 ( .A(n7127), .B(n7126), .Z(n7128) );
  NAND U9676 ( .A(n7129), .B(n7128), .Z(n8322) );
  NANDN U9677 ( .A(n7131), .B(n7130), .Z(n7135) );
  NAND U9678 ( .A(n7133), .B(n7132), .Z(n7134) );
  AND U9679 ( .A(n7135), .B(n7134), .Z(n8323) );
  XNOR U9680 ( .A(n8322), .B(n8323), .Z(n8324) );
  XNOR U9681 ( .A(n8325), .B(n8324), .Z(n7963) );
  NANDN U9682 ( .A(n7137), .B(n7136), .Z(n7141) );
  NAND U9683 ( .A(n7139), .B(n7138), .Z(n7140) );
  AND U9684 ( .A(n7141), .B(n7140), .Z(n7962) );
  XNOR U9685 ( .A(n7963), .B(n7962), .Z(n7964) );
  XNOR U9686 ( .A(n7965), .B(n7964), .Z(n7894) );
  XOR U9687 ( .A(n7895), .B(n7894), .Z(n7896) );
  XNOR U9688 ( .A(n7897), .B(n7896), .Z(n7984) );
  XNOR U9689 ( .A(n7985), .B(n7984), .Z(n7986) );
  NANDN U9690 ( .A(n7147), .B(n7146), .Z(n7151) );
  OR U9691 ( .A(n7149), .B(n7148), .Z(n7150) );
  NAND U9692 ( .A(n7151), .B(n7150), .Z(n7848) );
  OR U9693 ( .A(n7153), .B(n7152), .Z(n7157) );
  NANDN U9694 ( .A(n7155), .B(n7154), .Z(n7156) );
  NAND U9695 ( .A(n7157), .B(n7156), .Z(n7959) );
  NANDN U9696 ( .A(n7159), .B(n7158), .Z(n7163) );
  NAND U9697 ( .A(n7161), .B(n7160), .Z(n7162) );
  AND U9698 ( .A(n7163), .B(n7162), .Z(n7956) );
  NANDN U9699 ( .A(n7165), .B(n7164), .Z(n7169) );
  NANDN U9700 ( .A(n7167), .B(n7166), .Z(n7168) );
  AND U9701 ( .A(n7169), .B(n7168), .Z(n7957) );
  XNOR U9702 ( .A(n7959), .B(n7958), .Z(n7849) );
  XNOR U9703 ( .A(n7848), .B(n7849), .Z(n7850) );
  XOR U9704 ( .A(n7851), .B(n7850), .Z(n7891) );
  NANDN U9705 ( .A(n7171), .B(n7170), .Z(n7175) );
  OR U9706 ( .A(n7173), .B(n7172), .Z(n7174) );
  AND U9707 ( .A(n7175), .B(n7174), .Z(n7889) );
  NANDN U9708 ( .A(n7177), .B(n7176), .Z(n7181) );
  NANDN U9709 ( .A(n7179), .B(n7178), .Z(n7180) );
  NAND U9710 ( .A(n7181), .B(n7180), .Z(n8235) );
  NANDN U9711 ( .A(n7183), .B(n7182), .Z(n7187) );
  NANDN U9712 ( .A(n7185), .B(n7184), .Z(n7186) );
  NAND U9713 ( .A(n7187), .B(n7186), .Z(n8232) );
  NANDN U9714 ( .A(n7189), .B(n7188), .Z(n7193) );
  NAND U9715 ( .A(n7191), .B(n7190), .Z(n7192) );
  AND U9716 ( .A(n7193), .B(n7192), .Z(n8233) );
  XNOR U9717 ( .A(n8232), .B(n8233), .Z(n8234) );
  XNOR U9718 ( .A(n8235), .B(n8234), .Z(n8024) );
  NANDN U9719 ( .A(n7195), .B(n7194), .Z(n7199) );
  NANDN U9720 ( .A(n7197), .B(n7196), .Z(n7198) );
  NAND U9721 ( .A(n7199), .B(n7198), .Z(n8062) );
  NANDN U9722 ( .A(n7201), .B(n7200), .Z(n7205) );
  NANDN U9723 ( .A(n7203), .B(n7202), .Z(n7204) );
  AND U9724 ( .A(n7205), .B(n7204), .Z(n8060) );
  OR U9725 ( .A(n7207), .B(n7206), .Z(n7211) );
  NANDN U9726 ( .A(n7209), .B(n7208), .Z(n7210) );
  AND U9727 ( .A(n7211), .B(n7210), .Z(n8061) );
  XOR U9728 ( .A(n8062), .B(n8063), .Z(n8025) );
  XOR U9729 ( .A(n8024), .B(n8025), .Z(n8026) );
  NANDN U9730 ( .A(n7213), .B(n7212), .Z(n7217) );
  NANDN U9731 ( .A(n7215), .B(n7214), .Z(n7216) );
  NAND U9732 ( .A(n7217), .B(n7216), .Z(n8287) );
  NANDN U9733 ( .A(n7219), .B(n7218), .Z(n7223) );
  NANDN U9734 ( .A(n7221), .B(n7220), .Z(n7222) );
  NAND U9735 ( .A(n7223), .B(n7222), .Z(n8284) );
  OR U9736 ( .A(n7225), .B(n7224), .Z(n7229) );
  NANDN U9737 ( .A(n7227), .B(n7226), .Z(n7228) );
  NAND U9738 ( .A(n7229), .B(n7228), .Z(n8253) );
  OR U9739 ( .A(n7231), .B(n7230), .Z(n7235) );
  NANDN U9740 ( .A(n7233), .B(n7232), .Z(n7234) );
  NAND U9741 ( .A(n7235), .B(n7234), .Z(n8250) );
  NANDN U9742 ( .A(n7237), .B(n7236), .Z(n7241) );
  NANDN U9743 ( .A(n7239), .B(n7238), .Z(n7240) );
  AND U9744 ( .A(n7241), .B(n7240), .Z(n8251) );
  XNOR U9745 ( .A(n8250), .B(n8251), .Z(n8252) );
  XOR U9746 ( .A(n8253), .B(n8252), .Z(n8285) );
  XNOR U9747 ( .A(n8284), .B(n8285), .Z(n8286) );
  XOR U9748 ( .A(n8287), .B(n8286), .Z(n8027) );
  XOR U9749 ( .A(n8026), .B(n8027), .Z(n7888) );
  XNOR U9750 ( .A(n7889), .B(n7888), .Z(n7890) );
  XOR U9751 ( .A(n7891), .B(n7890), .Z(n7987) );
  XOR U9752 ( .A(n7986), .B(n7987), .Z(n7323) );
  NANDN U9753 ( .A(n7243), .B(n7242), .Z(n7247) );
  NANDN U9754 ( .A(n7245), .B(n7244), .Z(n7246) );
  NAND U9755 ( .A(n7247), .B(n7246), .Z(n7321) );
  NANDN U9756 ( .A(n7249), .B(n7248), .Z(n7253) );
  NANDN U9757 ( .A(n7251), .B(n7250), .Z(n7252) );
  NAND U9758 ( .A(n7253), .B(n7252), .Z(n8315) );
  NANDN U9759 ( .A(n7255), .B(n7254), .Z(n7259) );
  NAND U9760 ( .A(n7257), .B(n7256), .Z(n7258) );
  NAND U9761 ( .A(n7259), .B(n7258), .Z(n8312) );
  NANDN U9762 ( .A(n7261), .B(n7260), .Z(n7265) );
  NANDN U9763 ( .A(n7263), .B(n7262), .Z(n7264) );
  NAND U9764 ( .A(n7265), .B(n7264), .Z(n7907) );
  NANDN U9765 ( .A(n7267), .B(n7266), .Z(n7271) );
  NAND U9766 ( .A(n7269), .B(n7268), .Z(n7270) );
  NAND U9767 ( .A(n7271), .B(n7270), .Z(n7977) );
  NANDN U9768 ( .A(n7273), .B(n7272), .Z(n7277) );
  NAND U9769 ( .A(n7275), .B(n7274), .Z(n7276) );
  NAND U9770 ( .A(n7277), .B(n7276), .Z(n8079) );
  NANDN U9771 ( .A(n7279), .B(n7278), .Z(n7283) );
  NANDN U9772 ( .A(n7281), .B(n7280), .Z(n7282) );
  AND U9773 ( .A(n7283), .B(n7282), .Z(n8078) );
  XNOR U9774 ( .A(n8079), .B(n8078), .Z(n8080) );
  NANDN U9775 ( .A(n7285), .B(n7284), .Z(n7289) );
  NAND U9776 ( .A(n7287), .B(n7286), .Z(n7288) );
  NAND U9777 ( .A(n7289), .B(n7288), .Z(n8081) );
  XOR U9778 ( .A(n8080), .B(n8081), .Z(n7974) );
  NANDN U9779 ( .A(n7291), .B(n7290), .Z(n7295) );
  NANDN U9780 ( .A(n7293), .B(n7292), .Z(n7294) );
  NAND U9781 ( .A(n7295), .B(n7294), .Z(n8199) );
  OR U9782 ( .A(n7297), .B(n7296), .Z(n7301) );
  NANDN U9783 ( .A(n7299), .B(n7298), .Z(n7300) );
  NAND U9784 ( .A(n7301), .B(n7300), .Z(n8196) );
  NANDN U9785 ( .A(n7303), .B(n7302), .Z(n7307) );
  NANDN U9786 ( .A(n7305), .B(n7304), .Z(n7306) );
  AND U9787 ( .A(n7307), .B(n7306), .Z(n8197) );
  XNOR U9788 ( .A(n8196), .B(n8197), .Z(n8198) );
  XNOR U9789 ( .A(n8199), .B(n8198), .Z(n7975) );
  XNOR U9790 ( .A(n7974), .B(n7975), .Z(n7976) );
  XNOR U9791 ( .A(n7977), .B(n7976), .Z(n7904) );
  OR U9792 ( .A(n7309), .B(n7308), .Z(n7313) );
  NAND U9793 ( .A(n7311), .B(n7310), .Z(n7312) );
  NAND U9794 ( .A(n7313), .B(n7312), .Z(n7905) );
  XNOR U9795 ( .A(n7904), .B(n7905), .Z(n7906) );
  XNOR U9796 ( .A(n7907), .B(n7906), .Z(n8313) );
  XNOR U9797 ( .A(n8312), .B(n8313), .Z(n8314) );
  XOR U9798 ( .A(n8315), .B(n8314), .Z(n7320) );
  XNOR U9799 ( .A(n7321), .B(n7320), .Z(n7322) );
  XNOR U9800 ( .A(n7323), .B(n7322), .Z(n8301) );
  XOR U9801 ( .A(n8300), .B(n8301), .Z(n8302) );
  XNOR U9802 ( .A(n8303), .B(n8302), .Z(n7317) );
  XNOR U9803 ( .A(n7316), .B(n7317), .Z(o[2]) );
  OR U9804 ( .A(n7315), .B(n7314), .Z(n7319) );
  NANDN U9805 ( .A(n7317), .B(n7316), .Z(n7318) );
  NAND U9806 ( .A(n7319), .B(n7318), .Z(n8456) );
  NANDN U9807 ( .A(n7321), .B(n7320), .Z(n7325) );
  NAND U9808 ( .A(n7323), .B(n7322), .Z(n7324) );
  NAND U9809 ( .A(n7325), .B(n7324), .Z(n8882) );
  NANDN U9810 ( .A(n7327), .B(n7326), .Z(n7331) );
  NAND U9811 ( .A(n7329), .B(n7328), .Z(n7330) );
  AND U9812 ( .A(n7331), .B(n7330), .Z(n8883) );
  XNOR U9813 ( .A(n8882), .B(n8883), .Z(n8884) );
  NANDN U9814 ( .A(n7333), .B(n7332), .Z(n7337) );
  OR U9815 ( .A(n7335), .B(n7334), .Z(n7336) );
  NAND U9816 ( .A(n7337), .B(n7336), .Z(n8708) );
  NANDN U9817 ( .A(n7339), .B(n7338), .Z(n7343) );
  NAND U9818 ( .A(n7341), .B(n7340), .Z(n7342) );
  NAND U9819 ( .A(n7343), .B(n7342), .Z(n8542) );
  NANDN U9820 ( .A(n7345), .B(n7344), .Z(n7349) );
  NAND U9821 ( .A(n7347), .B(n7346), .Z(n7348) );
  NAND U9822 ( .A(n7349), .B(n7348), .Z(n8831) );
  NANDN U9823 ( .A(n7351), .B(n7350), .Z(n7355) );
  NAND U9824 ( .A(n7353), .B(n7352), .Z(n7354) );
  NAND U9825 ( .A(n7355), .B(n7354), .Z(n8829) );
  NANDN U9826 ( .A(n7357), .B(n7356), .Z(n7361) );
  NAND U9827 ( .A(n7359), .B(n7358), .Z(n7360) );
  NAND U9828 ( .A(n7361), .B(n7360), .Z(n8828) );
  XOR U9829 ( .A(n8831), .B(n8830), .Z(n8512) );
  OR U9830 ( .A(n7363), .B(n7362), .Z(n7367) );
  NANDN U9831 ( .A(n7365), .B(n7364), .Z(n7366) );
  AND U9832 ( .A(n7367), .B(n7366), .Z(n8510) );
  NANDN U9833 ( .A(n7369), .B(n7368), .Z(n7373) );
  NAND U9834 ( .A(n7371), .B(n7370), .Z(n7372) );
  NAND U9835 ( .A(n7373), .B(n7372), .Z(n8921) );
  NANDN U9836 ( .A(n7375), .B(n7374), .Z(n7379) );
  NAND U9837 ( .A(n7377), .B(n7376), .Z(n7378) );
  AND U9838 ( .A(n7379), .B(n7378), .Z(n8918) );
  NANDN U9839 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U9840 ( .A(n7383), .B(n7382), .Z(n7384) );
  AND U9841 ( .A(n7385), .B(n7384), .Z(n8919) );
  XNOR U9842 ( .A(n8921), .B(n8920), .Z(n8511) );
  XOR U9843 ( .A(n8512), .B(n8513), .Z(n8543) );
  XOR U9844 ( .A(n8542), .B(n8543), .Z(n8544) );
  OR U9845 ( .A(n7391), .B(n7390), .Z(n7395) );
  NANDN U9846 ( .A(n7393), .B(n7392), .Z(n7394) );
  NAND U9847 ( .A(n7395), .B(n7394), .Z(n8848) );
  OR U9848 ( .A(n7397), .B(n7396), .Z(n7401) );
  NAND U9849 ( .A(n7399), .B(n7398), .Z(n7400) );
  NAND U9850 ( .A(n7401), .B(n7400), .Z(n8847) );
  OR U9851 ( .A(n7403), .B(n7402), .Z(n7407) );
  NANDN U9852 ( .A(n7405), .B(n7404), .Z(n7406) );
  NAND U9853 ( .A(n7407), .B(n7406), .Z(n8846) );
  XOR U9854 ( .A(n8848), .B(n8849), .Z(n8480) );
  NAND U9855 ( .A(n7409), .B(n7408), .Z(n7413) );
  NAND U9856 ( .A(n7411), .B(n7410), .Z(n7412) );
  NAND U9857 ( .A(n7413), .B(n7412), .Z(n8481) );
  XOR U9858 ( .A(n8480), .B(n8481), .Z(n8483) );
  XOR U9859 ( .A(n8482), .B(n8483), .Z(n8545) );
  XNOR U9860 ( .A(n8544), .B(n8545), .Z(n8709) );
  XNOR U9861 ( .A(n8708), .B(n8709), .Z(n8710) );
  XOR U9862 ( .A(n8710), .B(n8711), .Z(n9028) );
  NANDN U9863 ( .A(n7419), .B(n7418), .Z(n7423) );
  NAND U9864 ( .A(n7421), .B(n7420), .Z(n7422) );
  NAND U9865 ( .A(n7423), .B(n7422), .Z(n8861) );
  NANDN U9866 ( .A(n7425), .B(n7424), .Z(n7429) );
  NAND U9867 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U9868 ( .A(n7429), .B(n7428), .Z(n8858) );
  NANDN U9869 ( .A(n7431), .B(n7430), .Z(n7435) );
  NAND U9870 ( .A(n7433), .B(n7432), .Z(n7434) );
  NAND U9871 ( .A(n7435), .B(n7434), .Z(n8606) );
  NANDN U9872 ( .A(n7437), .B(n7436), .Z(n7441) );
  NAND U9873 ( .A(n7439), .B(n7438), .Z(n7440) );
  NAND U9874 ( .A(n7441), .B(n7440), .Z(n8604) );
  OR U9875 ( .A(n7443), .B(n7442), .Z(n7447) );
  NANDN U9876 ( .A(n7445), .B(n7444), .Z(n7446) );
  AND U9877 ( .A(n7447), .B(n7446), .Z(n8603) );
  XNOR U9878 ( .A(n8604), .B(n8603), .Z(n8605) );
  XOR U9879 ( .A(n8606), .B(n8605), .Z(n8939) );
  OR U9880 ( .A(n7449), .B(n7448), .Z(n7453) );
  NANDN U9881 ( .A(n7451), .B(n7450), .Z(n7452) );
  NAND U9882 ( .A(n7453), .B(n7452), .Z(n8612) );
  XOR U9883 ( .A(n8610), .B(n8609), .Z(n8611) );
  XOR U9884 ( .A(n8612), .B(n8611), .Z(n8936) );
  NANDN U9885 ( .A(n7461), .B(n7460), .Z(n7465) );
  NAND U9886 ( .A(n7463), .B(n7462), .Z(n7464) );
  NAND U9887 ( .A(n7465), .B(n7464), .Z(n8937) );
  XNOR U9888 ( .A(n8936), .B(n8937), .Z(n8938) );
  XNOR U9889 ( .A(n8939), .B(n8938), .Z(n8704) );
  NANDN U9890 ( .A(n7467), .B(n7466), .Z(n7471) );
  NAND U9891 ( .A(n7469), .B(n7468), .Z(n7470) );
  NAND U9892 ( .A(n7471), .B(n7470), .Z(n8703) );
  NANDN U9893 ( .A(n7473), .B(n7472), .Z(n7477) );
  NAND U9894 ( .A(n7475), .B(n7474), .Z(n7476) );
  NAND U9895 ( .A(n7477), .B(n7476), .Z(n8560) );
  NANDN U9896 ( .A(n7479), .B(n7478), .Z(n7483) );
  NAND U9897 ( .A(n7481), .B(n7480), .Z(n7482) );
  AND U9898 ( .A(n7483), .B(n7482), .Z(n8561) );
  XNOR U9899 ( .A(n8560), .B(n8561), .Z(n8562) );
  OR U9900 ( .A(n7485), .B(n7484), .Z(n7489) );
  NAND U9901 ( .A(n7487), .B(n7486), .Z(n7488) );
  NAND U9902 ( .A(n7489), .B(n7488), .Z(n8489) );
  NANDN U9903 ( .A(n7491), .B(n7490), .Z(n7495) );
  NANDN U9904 ( .A(n7493), .B(n7492), .Z(n7494) );
  NAND U9905 ( .A(n7495), .B(n7494), .Z(n8487) );
  NANDN U9906 ( .A(n7497), .B(n7496), .Z(n7501) );
  NAND U9907 ( .A(n7499), .B(n7498), .Z(n7500) );
  AND U9908 ( .A(n7501), .B(n7500), .Z(n8486) );
  XNOR U9909 ( .A(n8487), .B(n8486), .Z(n8488) );
  XOR U9910 ( .A(n8489), .B(n8488), .Z(n8563) );
  XNOR U9911 ( .A(n8562), .B(n8563), .Z(n8702) );
  XNOR U9912 ( .A(n8703), .B(n8702), .Z(n8705) );
  XOR U9913 ( .A(n8704), .B(n8705), .Z(n8859) );
  XOR U9914 ( .A(n8858), .B(n8859), .Z(n8860) );
  XNOR U9915 ( .A(n8861), .B(n8860), .Z(n9026) );
  NAND U9916 ( .A(n7503), .B(n7502), .Z(n7507) );
  NANDN U9917 ( .A(n7505), .B(n7504), .Z(n7506) );
  NAND U9918 ( .A(n7507), .B(n7506), .Z(n8761) );
  OR U9919 ( .A(n7509), .B(n7508), .Z(n7513) );
  NANDN U9920 ( .A(n7511), .B(n7510), .Z(n7512) );
  NAND U9921 ( .A(n7513), .B(n7512), .Z(n8900) );
  OR U9922 ( .A(n7515), .B(n7514), .Z(n7519) );
  NAND U9923 ( .A(n7517), .B(n7516), .Z(n7518) );
  NAND U9924 ( .A(n7519), .B(n7518), .Z(n8901) );
  XNOR U9925 ( .A(n8900), .B(n8901), .Z(n8902) );
  OR U9926 ( .A(n7521), .B(n7520), .Z(n7525) );
  NANDN U9927 ( .A(n7523), .B(n7522), .Z(n7524) );
  NAND U9928 ( .A(n7525), .B(n7524), .Z(n8495) );
  OR U9929 ( .A(n7527), .B(n7526), .Z(n7531) );
  NAND U9930 ( .A(n7529), .B(n7528), .Z(n7530) );
  NAND U9931 ( .A(n7531), .B(n7530), .Z(n8493) );
  NANDN U9932 ( .A(n7533), .B(n7532), .Z(n7537) );
  NAND U9933 ( .A(n7535), .B(n7534), .Z(n7536) );
  AND U9934 ( .A(n7537), .B(n7536), .Z(n8492) );
  XNOR U9935 ( .A(n8493), .B(n8492), .Z(n8494) );
  XOR U9936 ( .A(n8495), .B(n8494), .Z(n8903) );
  XOR U9937 ( .A(n8902), .B(n8903), .Z(n8696) );
  NANDN U9938 ( .A(n7539), .B(n7538), .Z(n7543) );
  NAND U9939 ( .A(n7541), .B(n7540), .Z(n7542) );
  AND U9940 ( .A(n7543), .B(n7542), .Z(n8697) );
  XNOR U9941 ( .A(n8696), .B(n8697), .Z(n8698) );
  OR U9942 ( .A(n7545), .B(n7544), .Z(n7549) );
  NAND U9943 ( .A(n7547), .B(n7546), .Z(n7548) );
  NAND U9944 ( .A(n7549), .B(n7548), .Z(n8618) );
  NANDN U9945 ( .A(n7553), .B(n7554), .Z(n7559) );
  NOR U9946 ( .A(n7555), .B(n7554), .Z(n7556) );
  OR U9947 ( .A(n7557), .B(n7556), .Z(n7558) );
  NAND U9948 ( .A(n7559), .B(n7558), .Z(n8616) );
  XOR U9949 ( .A(n8615), .B(n8616), .Z(n8617) );
  XOR U9950 ( .A(n8618), .B(n8617), .Z(n8924) );
  NANDN U9951 ( .A(n7561), .B(n7560), .Z(n7565) );
  NAND U9952 ( .A(n7563), .B(n7562), .Z(n7564) );
  NAND U9953 ( .A(n7565), .B(n7564), .Z(n8925) );
  XNOR U9954 ( .A(n8924), .B(n8925), .Z(n8926) );
  OR U9955 ( .A(n7567), .B(n7566), .Z(n7571) );
  NANDN U9956 ( .A(n7569), .B(n7568), .Z(n7570) );
  NAND U9957 ( .A(n7571), .B(n7570), .Z(n8909) );
  OR U9958 ( .A(n7573), .B(n7572), .Z(n7577) );
  NAND U9959 ( .A(n7575), .B(n7574), .Z(n7576) );
  NAND U9960 ( .A(n7577), .B(n7576), .Z(n8906) );
  NANDN U9961 ( .A(n7579), .B(n7578), .Z(n7583) );
  NAND U9962 ( .A(n7581), .B(n7580), .Z(n7582) );
  AND U9963 ( .A(n7583), .B(n7582), .Z(n8907) );
  XNOR U9964 ( .A(n8906), .B(n8907), .Z(n8908) );
  XOR U9965 ( .A(n8909), .B(n8908), .Z(n8927) );
  XOR U9966 ( .A(n8926), .B(n8927), .Z(n8699) );
  XNOR U9967 ( .A(n8698), .B(n8699), .Z(n8758) );
  OR U9968 ( .A(n7585), .B(n7584), .Z(n7589) );
  NAND U9969 ( .A(n7587), .B(n7586), .Z(n7588) );
  NAND U9970 ( .A(n7589), .B(n7588), .Z(n8759) );
  XNOR U9971 ( .A(n8758), .B(n8759), .Z(n8760) );
  XOR U9972 ( .A(n8761), .B(n8760), .Z(n9027) );
  XOR U9973 ( .A(n9026), .B(n9027), .Z(n9029) );
  XNOR U9974 ( .A(n9028), .B(n9029), .Z(n8885) );
  XNOR U9975 ( .A(n8884), .B(n8885), .Z(n8871) );
  NANDN U9976 ( .A(n7591), .B(n7590), .Z(n7595) );
  NAND U9977 ( .A(n7593), .B(n7592), .Z(n7594) );
  NAND U9978 ( .A(n7595), .B(n7594), .Z(n8889) );
  NANDN U9979 ( .A(n7597), .B(n7596), .Z(n7601) );
  NAND U9980 ( .A(n7599), .B(n7598), .Z(n7600) );
  NAND U9981 ( .A(n7601), .B(n7600), .Z(n8770) );
  NANDN U9982 ( .A(n7607), .B(n7606), .Z(n7611) );
  NANDN U9983 ( .A(n7609), .B(n7608), .Z(n7610) );
  NAND U9984 ( .A(n7611), .B(n7610), .Z(n8672) );
  NANDN U9985 ( .A(n7613), .B(n7612), .Z(n7617) );
  NAND U9986 ( .A(n7615), .B(n7614), .Z(n7616) );
  AND U9987 ( .A(n7617), .B(n7616), .Z(n8671) );
  XNOR U9988 ( .A(n8672), .B(n8671), .Z(n8673) );
  XNOR U9989 ( .A(n8674), .B(n8673), .Z(n8768) );
  NANDN U9990 ( .A(n7619), .B(n7618), .Z(n7623) );
  NAND U9991 ( .A(n7621), .B(n7620), .Z(n7622) );
  NAND U9992 ( .A(n7623), .B(n7622), .Z(n8743) );
  NANDN U9993 ( .A(n7625), .B(n7624), .Z(n7629) );
  NANDN U9994 ( .A(n7627), .B(n7626), .Z(n7628) );
  NAND U9995 ( .A(n7629), .B(n7628), .Z(n8741) );
  NANDN U9996 ( .A(n7631), .B(n7630), .Z(n7635) );
  OR U9997 ( .A(n7633), .B(n7632), .Z(n7634) );
  AND U9998 ( .A(n7635), .B(n7634), .Z(n8740) );
  XNOR U9999 ( .A(n8741), .B(n8740), .Z(n8742) );
  XNOR U10000 ( .A(n8743), .B(n8742), .Z(n8769) );
  XOR U10001 ( .A(n8768), .B(n8769), .Z(n8771) );
  XNOR U10002 ( .A(n8770), .B(n8771), .Z(n8780) );
  XNOR U10003 ( .A(n8780), .B(n8781), .Z(n8782) );
  NANDN U10004 ( .A(n7641), .B(n7640), .Z(n7645) );
  NANDN U10005 ( .A(n7643), .B(n7642), .Z(n7644) );
  NAND U10006 ( .A(n7645), .B(n7644), .Z(n8680) );
  NANDN U10007 ( .A(n7647), .B(n7646), .Z(n7651) );
  NANDN U10008 ( .A(n7649), .B(n7648), .Z(n7650) );
  NAND U10009 ( .A(n7651), .B(n7650), .Z(n8662) );
  NANDN U10010 ( .A(n7653), .B(n7652), .Z(n7657) );
  NAND U10011 ( .A(n7655), .B(n7654), .Z(n7656) );
  NAND U10012 ( .A(n7657), .B(n7656), .Z(n8659) );
  NANDN U10013 ( .A(n7659), .B(n7658), .Z(n7663) );
  NANDN U10014 ( .A(n7661), .B(n7660), .Z(n7662) );
  NAND U10015 ( .A(n7663), .B(n7662), .Z(n8660) );
  XNOR U10016 ( .A(n8659), .B(n8660), .Z(n8661) );
  XNOR U10017 ( .A(n8662), .B(n8661), .Z(n8677) );
  NAND U10018 ( .A(n7665), .B(n7664), .Z(n7669) );
  NAND U10019 ( .A(n7667), .B(n7666), .Z(n7668) );
  NAND U10020 ( .A(n7669), .B(n7668), .Z(n8752) );
  NANDN U10021 ( .A(n7671), .B(n7670), .Z(n7675) );
  NANDN U10022 ( .A(n7673), .B(n7672), .Z(n7674) );
  AND U10023 ( .A(n7675), .B(n7674), .Z(n8753) );
  XNOR U10024 ( .A(n8752), .B(n8753), .Z(n8754) );
  XNOR U10025 ( .A(n8754), .B(n8755), .Z(n8678) );
  XNOR U10026 ( .A(n8677), .B(n8678), .Z(n8679) );
  XNOR U10027 ( .A(n8680), .B(n8679), .Z(n8783) );
  XNOR U10028 ( .A(n8782), .B(n8783), .Z(n8888) );
  XOR U10029 ( .A(n8889), .B(n8888), .Z(n8890) );
  NANDN U10030 ( .A(n7681), .B(n7680), .Z(n7685) );
  NANDN U10031 ( .A(n7683), .B(n7682), .Z(n7684) );
  NAND U10032 ( .A(n7685), .B(n7684), .Z(n8727) );
  NAND U10033 ( .A(n7687), .B(n7686), .Z(n7691) );
  NAND U10034 ( .A(n7689), .B(n7688), .Z(n7690) );
  NAND U10035 ( .A(n7691), .B(n7690), .Z(n8724) );
  NAND U10036 ( .A(n7693), .B(n7692), .Z(n7697) );
  NANDN U10037 ( .A(n7695), .B(n7694), .Z(n7696) );
  NAND U10038 ( .A(n7697), .B(n7696), .Z(n8725) );
  XNOR U10039 ( .A(n8724), .B(n8725), .Z(n8726) );
  XNOR U10040 ( .A(n8727), .B(n8726), .Z(n8891) );
  XOR U10041 ( .A(n8890), .B(n8891), .Z(n8870) );
  XOR U10042 ( .A(n8871), .B(n8870), .Z(n8872) );
  OR U10043 ( .A(n7699), .B(n7698), .Z(n7703) );
  NANDN U10044 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U10045 ( .A(n7703), .B(n7702), .Z(n8873) );
  XNOR U10046 ( .A(n8872), .B(n8873), .Z(n8457) );
  XNOR U10047 ( .A(n8456), .B(n8457), .Z(n8458) );
  NANDN U10048 ( .A(n7705), .B(n7704), .Z(n7709) );
  NAND U10049 ( .A(n7707), .B(n7706), .Z(n7708) );
  NAND U10050 ( .A(n7709), .B(n7708), .Z(n8622) );
  NANDN U10051 ( .A(n7711), .B(n7710), .Z(n7715) );
  NAND U10052 ( .A(n7713), .B(n7712), .Z(n7714) );
  NAND U10053 ( .A(n7715), .B(n7714), .Z(n8621) );
  NANDN U10054 ( .A(n7717), .B(n7716), .Z(n7721) );
  NAND U10055 ( .A(n7719), .B(n7718), .Z(n7720) );
  NAND U10056 ( .A(n7721), .B(n7720), .Z(n8624) );
  XOR U10057 ( .A(n8623), .B(n8624), .Z(n9000) );
  NANDN U10058 ( .A(n7723), .B(n7722), .Z(n7727) );
  NAND U10059 ( .A(n7725), .B(n7724), .Z(n7726) );
  NAND U10060 ( .A(n7727), .B(n7726), .Z(n8975) );
  NANDN U10061 ( .A(n7729), .B(n7728), .Z(n7733) );
  NAND U10062 ( .A(n7731), .B(n7730), .Z(n7732) );
  NAND U10063 ( .A(n7733), .B(n7732), .Z(n8973) );
  NANDN U10064 ( .A(n7735), .B(n7734), .Z(n7739) );
  NAND U10065 ( .A(n7737), .B(n7736), .Z(n7738) );
  NAND U10066 ( .A(n7739), .B(n7738), .Z(n8972) );
  XNOR U10067 ( .A(n8975), .B(n8974), .Z(n8998) );
  NANDN U10068 ( .A(n7741), .B(n7740), .Z(n7745) );
  NAND U10069 ( .A(n7743), .B(n7742), .Z(n7744) );
  NAND U10070 ( .A(n7745), .B(n7744), .Z(n8999) );
  XOR U10071 ( .A(n9000), .B(n9001), .Z(n8541) );
  OR U10072 ( .A(n7747), .B(n7746), .Z(n7751) );
  NAND U10073 ( .A(n7749), .B(n7748), .Z(n7750) );
  NAND U10074 ( .A(n7751), .B(n7750), .Z(n8574) );
  NANDN U10075 ( .A(n7753), .B(n7752), .Z(n7757) );
  NAND U10076 ( .A(n7755), .B(n7754), .Z(n7756) );
  NAND U10077 ( .A(n7757), .B(n7756), .Z(n8825) );
  NANDN U10078 ( .A(n7759), .B(n7758), .Z(n7763) );
  NAND U10079 ( .A(n7761), .B(n7760), .Z(n7762) );
  NAND U10080 ( .A(n7763), .B(n7762), .Z(n8823) );
  NANDN U10081 ( .A(n7765), .B(n7764), .Z(n7769) );
  NAND U10082 ( .A(n7767), .B(n7766), .Z(n7768) );
  NAND U10083 ( .A(n7769), .B(n7768), .Z(n8822) );
  XNOR U10084 ( .A(n8825), .B(n8824), .Z(n8572) );
  NANDN U10085 ( .A(n7771), .B(n7770), .Z(n7775) );
  NAND U10086 ( .A(n7773), .B(n7772), .Z(n7774) );
  NAND U10087 ( .A(n7775), .B(n7774), .Z(n8573) );
  XOR U10088 ( .A(n8574), .B(n8575), .Z(n8539) );
  OR U10089 ( .A(n7777), .B(n7776), .Z(n7781) );
  NANDN U10090 ( .A(n7779), .B(n7778), .Z(n7780) );
  NAND U10091 ( .A(n7781), .B(n7780), .Z(n8477) );
  NANDN U10092 ( .A(n7783), .B(n7782), .Z(n7787) );
  NAND U10093 ( .A(n7785), .B(n7784), .Z(n7786) );
  NAND U10094 ( .A(n7787), .B(n7786), .Z(n8914) );
  NANDN U10095 ( .A(n7789), .B(n7788), .Z(n7793) );
  NAND U10096 ( .A(n7791), .B(n7790), .Z(n7792) );
  AND U10097 ( .A(n7793), .B(n7792), .Z(n8912) );
  NANDN U10098 ( .A(n7795), .B(n7794), .Z(n7799) );
  NANDN U10099 ( .A(n7797), .B(n7796), .Z(n7798) );
  AND U10100 ( .A(n7799), .B(n7798), .Z(n8913) );
  XOR U10101 ( .A(n8914), .B(n8915), .Z(n8474) );
  NANDN U10102 ( .A(n7801), .B(n7800), .Z(n7805) );
  NANDN U10103 ( .A(n7803), .B(n7802), .Z(n7804) );
  NAND U10104 ( .A(n7805), .B(n7804), .Z(n8475) );
  XNOR U10105 ( .A(n8474), .B(n8475), .Z(n8476) );
  XNOR U10106 ( .A(n8477), .B(n8476), .Z(n8538) );
  XOR U10107 ( .A(n8539), .B(n8538), .Z(n8540) );
  XOR U10108 ( .A(n8541), .B(n8540), .Z(n8763) );
  NANDN U10109 ( .A(n7807), .B(n7806), .Z(n7811) );
  NANDN U10110 ( .A(n7809), .B(n7808), .Z(n7810) );
  AND U10111 ( .A(n7811), .B(n7810), .Z(n8762) );
  XOR U10112 ( .A(n8763), .B(n8762), .Z(n8764) );
  NANDN U10113 ( .A(n7813), .B(n7812), .Z(n7817) );
  OR U10114 ( .A(n7815), .B(n7814), .Z(n7816) );
  NAND U10115 ( .A(n7817), .B(n7816), .Z(n8668) );
  NAND U10116 ( .A(n7819), .B(n7818), .Z(n7823) );
  NANDN U10117 ( .A(n7821), .B(n7820), .Z(n7822) );
  NAND U10118 ( .A(n7823), .B(n7822), .Z(n8665) );
  OR U10119 ( .A(n7825), .B(n7824), .Z(n7829) );
  NANDN U10120 ( .A(n7827), .B(n7826), .Z(n7828) );
  NAND U10121 ( .A(n7829), .B(n7828), .Z(n8593) );
  OR U10122 ( .A(n7831), .B(n7830), .Z(n7835) );
  NANDN U10123 ( .A(n7833), .B(n7832), .Z(n7834) );
  AND U10124 ( .A(n7835), .B(n7834), .Z(n8590) );
  NANDN U10125 ( .A(n7837), .B(n7836), .Z(n7841) );
  NAND U10126 ( .A(n7839), .B(n7838), .Z(n7840) );
  NAND U10127 ( .A(n7841), .B(n7840), .Z(n8591) );
  XNOR U10128 ( .A(n8593), .B(n8592), .Z(n8666) );
  XNOR U10129 ( .A(n8665), .B(n8666), .Z(n8667) );
  XOR U10130 ( .A(n8668), .B(n8667), .Z(n8765) );
  XOR U10131 ( .A(n8764), .B(n8765), .Z(n8866) );
  NANDN U10132 ( .A(n7843), .B(n7842), .Z(n7847) );
  NAND U10133 ( .A(n7845), .B(n7844), .Z(n7846) );
  NAND U10134 ( .A(n7847), .B(n7846), .Z(n8640) );
  NANDN U10135 ( .A(n7849), .B(n7848), .Z(n7853) );
  NANDN U10136 ( .A(n7851), .B(n7850), .Z(n7852) );
  NAND U10137 ( .A(n7853), .B(n7852), .Z(n8992) );
  NANDN U10138 ( .A(n7855), .B(n7854), .Z(n7859) );
  NAND U10139 ( .A(n7857), .B(n7856), .Z(n7858) );
  NAND U10140 ( .A(n7859), .B(n7858), .Z(n8951) );
  NANDN U10141 ( .A(n7861), .B(n7860), .Z(n7865) );
  NANDN U10142 ( .A(n7863), .B(n7862), .Z(n7864) );
  AND U10143 ( .A(n7865), .B(n7864), .Z(n8948) );
  XOR U10144 ( .A(n8951), .B(n8950), .Z(n8993) );
  XOR U10145 ( .A(n8992), .B(n8993), .Z(n8994) );
  NANDN U10146 ( .A(n7871), .B(n7870), .Z(n7875) );
  NANDN U10147 ( .A(n7873), .B(n7872), .Z(n7874) );
  NAND U10148 ( .A(n7875), .B(n7874), .Z(n8995) );
  XOR U10149 ( .A(n8994), .B(n8995), .Z(n8637) );
  XNOR U10150 ( .A(n8637), .B(n8638), .Z(n8639) );
  XOR U10151 ( .A(n8640), .B(n8639), .Z(n8864) );
  NANDN U10152 ( .A(n7889), .B(n7888), .Z(n7893) );
  NANDN U10153 ( .A(n7891), .B(n7890), .Z(n7892) );
  NAND U10154 ( .A(n7893), .B(n7892), .Z(n8529) );
  XNOR U10155 ( .A(n8528), .B(n8529), .Z(n8530) );
  XNOR U10156 ( .A(n8531), .B(n8530), .Z(n8865) );
  XNOR U10157 ( .A(n8864), .B(n8865), .Z(n8867) );
  XOR U10158 ( .A(n8866), .B(n8867), .Z(n8464) );
  NANDN U10159 ( .A(n7899), .B(n7898), .Z(n7903) );
  NANDN U10160 ( .A(n7901), .B(n7900), .Z(n7902) );
  NAND U10161 ( .A(n7903), .B(n7902), .Z(n8737) );
  NANDN U10162 ( .A(n7905), .B(n7904), .Z(n7909) );
  NAND U10163 ( .A(n7907), .B(n7906), .Z(n7908) );
  NAND U10164 ( .A(n7909), .B(n7908), .Z(n8557) );
  NANDN U10165 ( .A(n7917), .B(n7916), .Z(n7921) );
  OR U10166 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U10167 ( .A(n7921), .B(n7920), .Z(n8969) );
  XOR U10168 ( .A(n8966), .B(n8967), .Z(n8968) );
  XOR U10169 ( .A(n8969), .B(n8968), .Z(n8930) );
  XOR U10170 ( .A(n8931), .B(n8930), .Z(n8933) );
  XOR U10171 ( .A(n8933), .B(n8932), .Z(n8555) );
  XNOR U10172 ( .A(n8554), .B(n8555), .Z(n8556) );
  XNOR U10173 ( .A(n8557), .B(n8556), .Z(n8736) );
  XOR U10174 ( .A(n8737), .B(n8736), .Z(n8738) );
  XNOR U10175 ( .A(n8739), .B(n8738), .Z(n8717) );
  NANDN U10176 ( .A(n7933), .B(n7932), .Z(n7937) );
  NAND U10177 ( .A(n7935), .B(n7934), .Z(n7936) );
  NAND U10178 ( .A(n7937), .B(n7936), .Z(n8793) );
  NANDN U10179 ( .A(n7939), .B(n7938), .Z(n7943) );
  NANDN U10180 ( .A(n7941), .B(n7940), .Z(n7942) );
  AND U10181 ( .A(n7943), .B(n7942), .Z(n8792) );
  XNOR U10182 ( .A(n8793), .B(n8792), .Z(n8794) );
  OR U10183 ( .A(n7945), .B(n7944), .Z(n7949) );
  NAND U10184 ( .A(n7947), .B(n7946), .Z(n7948) );
  NAND U10185 ( .A(n7949), .B(n7948), .Z(n8801) );
  NANDN U10186 ( .A(n7951), .B(n7950), .Z(n7955) );
  NAND U10187 ( .A(n7953), .B(n7952), .Z(n7954) );
  NAND U10188 ( .A(n7955), .B(n7954), .Z(n8799) );
  OR U10189 ( .A(n7957), .B(n7956), .Z(n7961) );
  NAND U10190 ( .A(n7959), .B(n7958), .Z(n7960) );
  AND U10191 ( .A(n7961), .B(n7960), .Z(n8798) );
  XNOR U10192 ( .A(n8799), .B(n8798), .Z(n8800) );
  XOR U10193 ( .A(n8801), .B(n8800), .Z(n8795) );
  XOR U10194 ( .A(n8794), .B(n8795), .Z(n8551) );
  NANDN U10195 ( .A(n7963), .B(n7962), .Z(n7967) );
  NANDN U10196 ( .A(n7965), .B(n7964), .Z(n7966) );
  NAND U10197 ( .A(n7967), .B(n7966), .Z(n8507) );
  NANDN U10198 ( .A(n7969), .B(n7968), .Z(n7973) );
  NAND U10199 ( .A(n7971), .B(n7970), .Z(n7972) );
  NAND U10200 ( .A(n7973), .B(n7972), .Z(n8505) );
  NANDN U10201 ( .A(n7975), .B(n7974), .Z(n7979) );
  NAND U10202 ( .A(n7977), .B(n7976), .Z(n7978) );
  AND U10203 ( .A(n7979), .B(n7978), .Z(n8504) );
  XNOR U10204 ( .A(n8505), .B(n8504), .Z(n8506) );
  XOR U10205 ( .A(n8507), .B(n8506), .Z(n8548) );
  XNOR U10206 ( .A(n8548), .B(n8549), .Z(n8550) );
  XNOR U10207 ( .A(n8551), .B(n8550), .Z(n8714) );
  XNOR U10208 ( .A(n8714), .B(n8715), .Z(n8716) );
  XOR U10209 ( .A(n8717), .B(n8716), .Z(n8462) );
  NANDN U10210 ( .A(n7989), .B(n7988), .Z(n7993) );
  NAND U10211 ( .A(n7991), .B(n7990), .Z(n7992) );
  NAND U10212 ( .A(n7993), .B(n7992), .Z(n8636) );
  NANDN U10213 ( .A(n7995), .B(n7994), .Z(n7999) );
  OR U10214 ( .A(n7997), .B(n7996), .Z(n7998) );
  NAND U10215 ( .A(n7999), .B(n7998), .Z(n8813) );
  OR U10216 ( .A(n8001), .B(n8000), .Z(n8005) );
  NANDN U10217 ( .A(n8003), .B(n8002), .Z(n8004) );
  NAND U10218 ( .A(n8005), .B(n8004), .Z(n8811) );
  NANDN U10219 ( .A(n8007), .B(n8006), .Z(n8011) );
  NAND U10220 ( .A(n8009), .B(n8008), .Z(n8010) );
  AND U10221 ( .A(n8011), .B(n8010), .Z(n8810) );
  XNOR U10222 ( .A(n8811), .B(n8810), .Z(n8812) );
  XNOR U10223 ( .A(n8813), .B(n8812), .Z(n8633) );
  NANDN U10224 ( .A(n8013), .B(n8012), .Z(n8017) );
  NAND U10225 ( .A(n8015), .B(n8014), .Z(n8016) );
  AND U10226 ( .A(n8017), .B(n8016), .Z(n8634) );
  XNOR U10227 ( .A(n8633), .B(n8634), .Z(n8635) );
  XNOR U10228 ( .A(n8636), .B(n8635), .Z(n8789) );
  OR U10229 ( .A(n8019), .B(n8018), .Z(n8023) );
  NAND U10230 ( .A(n8021), .B(n8020), .Z(n8022) );
  NAND U10231 ( .A(n8023), .B(n8022), .Z(n8957) );
  OR U10232 ( .A(n8025), .B(n8024), .Z(n8029) );
  NAND U10233 ( .A(n8027), .B(n8026), .Z(n8028) );
  NAND U10234 ( .A(n8029), .B(n8028), .Z(n8955) );
  NANDN U10235 ( .A(n8031), .B(n8030), .Z(n8035) );
  NANDN U10236 ( .A(n8033), .B(n8032), .Z(n8034) );
  NAND U10237 ( .A(n8035), .B(n8034), .Z(n8855) );
  NANDN U10238 ( .A(n8037), .B(n8036), .Z(n8041) );
  NAND U10239 ( .A(n8039), .B(n8038), .Z(n8040) );
  AND U10240 ( .A(n8041), .B(n8040), .Z(n8852) );
  NANDN U10241 ( .A(n8043), .B(n8042), .Z(n8047) );
  OR U10242 ( .A(n8045), .B(n8044), .Z(n8046) );
  NAND U10243 ( .A(n8047), .B(n8046), .Z(n8853) );
  XNOR U10244 ( .A(n8855), .B(n8854), .Z(n8954) );
  XNOR U10245 ( .A(n8955), .B(n8954), .Z(n8956) );
  XNOR U10246 ( .A(n8957), .B(n8956), .Z(n8787) );
  NANDN U10247 ( .A(n8049), .B(n8048), .Z(n8053) );
  OR U10248 ( .A(n8051), .B(n8050), .Z(n8052) );
  NAND U10249 ( .A(n8053), .B(n8052), .Z(n8525) );
  OR U10250 ( .A(n8055), .B(n8054), .Z(n8059) );
  NANDN U10251 ( .A(n8057), .B(n8056), .Z(n8058) );
  NAND U10252 ( .A(n8059), .B(n8058), .Z(n8523) );
  OR U10253 ( .A(n8061), .B(n8060), .Z(n8065) );
  NANDN U10254 ( .A(n8063), .B(n8062), .Z(n8064) );
  NAND U10255 ( .A(n8065), .B(n8064), .Z(n8522) );
  XNOR U10256 ( .A(n8525), .B(n8524), .Z(n9024) );
  OR U10257 ( .A(n8067), .B(n8066), .Z(n8071) );
  NANDN U10258 ( .A(n8069), .B(n8068), .Z(n8070) );
  NAND U10259 ( .A(n8071), .B(n8070), .Z(n9023) );
  NANDN U10260 ( .A(n8073), .B(n8072), .Z(n8077) );
  NANDN U10261 ( .A(n8075), .B(n8074), .Z(n8076) );
  AND U10262 ( .A(n8077), .B(n8076), .Z(n9022) );
  XNOR U10263 ( .A(n9023), .B(n9022), .Z(n9025) );
  XOR U10264 ( .A(n9024), .B(n9025), .Z(n8786) );
  XOR U10265 ( .A(n8787), .B(n8786), .Z(n8788) );
  XOR U10266 ( .A(n8789), .B(n8788), .Z(n8894) );
  NANDN U10267 ( .A(n8079), .B(n8078), .Z(n8083) );
  NANDN U10268 ( .A(n8081), .B(n8080), .Z(n8082) );
  NAND U10269 ( .A(n8083), .B(n8082), .Z(n8569) );
  OR U10270 ( .A(n8085), .B(n8084), .Z(n8089) );
  NANDN U10271 ( .A(n8087), .B(n8086), .Z(n8088) );
  AND U10272 ( .A(n8089), .B(n8088), .Z(n8566) );
  NANDN U10273 ( .A(n8091), .B(n8090), .Z(n8095) );
  NAND U10274 ( .A(n8093), .B(n8092), .Z(n8094) );
  NAND U10275 ( .A(n8095), .B(n8094), .Z(n8567) );
  XNOR U10276 ( .A(n8569), .B(n8568), .Z(n8690) );
  NANDN U10277 ( .A(n8097), .B(n8096), .Z(n8101) );
  NAND U10278 ( .A(n8099), .B(n8098), .Z(n8100) );
  NAND U10279 ( .A(n8101), .B(n8100), .Z(n8807) );
  OR U10280 ( .A(n8103), .B(n8102), .Z(n8107) );
  NANDN U10281 ( .A(n8105), .B(n8104), .Z(n8106) );
  AND U10282 ( .A(n8107), .B(n8106), .Z(n8804) );
  NANDN U10283 ( .A(n8109), .B(n8108), .Z(n8113) );
  NAND U10284 ( .A(n8111), .B(n8110), .Z(n8112) );
  NAND U10285 ( .A(n8113), .B(n8112), .Z(n8805) );
  XOR U10286 ( .A(n8807), .B(n8806), .Z(n8691) );
  XOR U10287 ( .A(n8690), .B(n8691), .Z(n8692) );
  OR U10288 ( .A(n8115), .B(n8114), .Z(n8119) );
  NANDN U10289 ( .A(n8117), .B(n8116), .Z(n8118) );
  NAND U10290 ( .A(n8119), .B(n8118), .Z(n8843) );
  NANDN U10291 ( .A(n8121), .B(n8120), .Z(n8125) );
  NAND U10292 ( .A(n8123), .B(n8122), .Z(n8124) );
  NAND U10293 ( .A(n8125), .B(n8124), .Z(n8841) );
  NANDN U10294 ( .A(n8127), .B(n8126), .Z(n8131) );
  NAND U10295 ( .A(n8129), .B(n8128), .Z(n8130) );
  NAND U10296 ( .A(n8131), .B(n8130), .Z(n8840) );
  XOR U10297 ( .A(n8843), .B(n8842), .Z(n8581) );
  NANDN U10298 ( .A(n8133), .B(n8132), .Z(n8137) );
  NANDN U10299 ( .A(n8135), .B(n8134), .Z(n8136) );
  AND U10300 ( .A(n8137), .B(n8136), .Z(n8578) );
  OR U10301 ( .A(n8139), .B(n8138), .Z(n8143) );
  NANDN U10302 ( .A(n8141), .B(n8140), .Z(n8142) );
  NAND U10303 ( .A(n8143), .B(n8142), .Z(n8817) );
  NANDN U10304 ( .A(n8145), .B(n8144), .Z(n8149) );
  NAND U10305 ( .A(n8147), .B(n8146), .Z(n8148) );
  NAND U10306 ( .A(n8149), .B(n8148), .Z(n8816) );
  NANDN U10307 ( .A(n8151), .B(n8150), .Z(n8155) );
  NAND U10308 ( .A(n8153), .B(n8152), .Z(n8154) );
  NAND U10309 ( .A(n8155), .B(n8154), .Z(n8819) );
  XNOR U10310 ( .A(n8818), .B(n8819), .Z(n8579) );
  XNOR U10311 ( .A(n8581), .B(n8580), .Z(n8693) );
  XOR U10312 ( .A(n8692), .B(n8693), .Z(n8777) );
  NANDN U10313 ( .A(n8157), .B(n8156), .Z(n8161) );
  OR U10314 ( .A(n8159), .B(n8158), .Z(n8160) );
  NAND U10315 ( .A(n8161), .B(n8160), .Z(n9013) );
  OR U10316 ( .A(n8163), .B(n8162), .Z(n8167) );
  NAND U10317 ( .A(n8165), .B(n8164), .Z(n8166) );
  NAND U10318 ( .A(n8167), .B(n8166), .Z(n9010) );
  NANDN U10319 ( .A(n8169), .B(n8168), .Z(n8173) );
  NANDN U10320 ( .A(n8171), .B(n8170), .Z(n8172) );
  NAND U10321 ( .A(n8173), .B(n8172), .Z(n9011) );
  XNOR U10322 ( .A(n9010), .B(n9011), .Z(n9012) );
  XOR U10323 ( .A(n9013), .B(n9012), .Z(n9019) );
  NANDN U10324 ( .A(n8179), .B(n8178), .Z(n8183) );
  NANDN U10325 ( .A(n8181), .B(n8180), .Z(n8182) );
  NAND U10326 ( .A(n8183), .B(n8182), .Z(n9017) );
  XNOR U10327 ( .A(n9016), .B(n9017), .Z(n9018) );
  XNOR U10328 ( .A(n9019), .B(n9018), .Z(n8774) );
  NANDN U10329 ( .A(n8185), .B(n8184), .Z(n8189) );
  OR U10330 ( .A(n8187), .B(n8186), .Z(n8188) );
  NAND U10331 ( .A(n8189), .B(n8188), .Z(n8749) );
  NANDN U10332 ( .A(n8191), .B(n8190), .Z(n8195) );
  NANDN U10333 ( .A(n8193), .B(n8192), .Z(n8194) );
  NAND U10334 ( .A(n8195), .B(n8194), .Z(n8587) );
  NANDN U10335 ( .A(n8197), .B(n8196), .Z(n8201) );
  NAND U10336 ( .A(n8199), .B(n8198), .Z(n8200) );
  NAND U10337 ( .A(n8201), .B(n8200), .Z(n8585) );
  OR U10338 ( .A(n8203), .B(n8202), .Z(n8207) );
  NAND U10339 ( .A(n8205), .B(n8204), .Z(n8206) );
  AND U10340 ( .A(n8207), .B(n8206), .Z(n8584) );
  XNOR U10341 ( .A(n8585), .B(n8584), .Z(n8586) );
  XNOR U10342 ( .A(n8587), .B(n8586), .Z(n8747) );
  NANDN U10343 ( .A(n8209), .B(n8208), .Z(n8213) );
  NAND U10344 ( .A(n8211), .B(n8210), .Z(n8212) );
  AND U10345 ( .A(n8213), .B(n8212), .Z(n8746) );
  XNOR U10346 ( .A(n8747), .B(n8746), .Z(n8748) );
  XOR U10347 ( .A(n8749), .B(n8748), .Z(n8775) );
  XNOR U10348 ( .A(n8774), .B(n8775), .Z(n8776) );
  XNOR U10349 ( .A(n8777), .B(n8776), .Z(n8895) );
  XOR U10350 ( .A(n8894), .B(n8895), .Z(n8896) );
  NAND U10351 ( .A(n8215), .B(n8214), .Z(n8219) );
  OR U10352 ( .A(n8217), .B(n8216), .Z(n8218) );
  NAND U10353 ( .A(n8219), .B(n8218), .Z(n8652) );
  NANDN U10354 ( .A(n8221), .B(n8220), .Z(n8225) );
  NAND U10355 ( .A(n8223), .B(n8222), .Z(n8224) );
  NAND U10356 ( .A(n8225), .B(n8224), .Z(n8650) );
  NANDN U10357 ( .A(n8227), .B(n8226), .Z(n8231) );
  OR U10358 ( .A(n8229), .B(n8228), .Z(n8230) );
  NAND U10359 ( .A(n8231), .B(n8230), .Z(n8962) );
  NANDN U10360 ( .A(n8233), .B(n8232), .Z(n8237) );
  NAND U10361 ( .A(n8235), .B(n8234), .Z(n8236) );
  NAND U10362 ( .A(n8237), .B(n8236), .Z(n8961) );
  NANDN U10363 ( .A(n8239), .B(n8238), .Z(n8243) );
  NAND U10364 ( .A(n8241), .B(n8240), .Z(n8242) );
  NAND U10365 ( .A(n8243), .B(n8242), .Z(n8960) );
  XOR U10366 ( .A(n8962), .B(n8963), .Z(n8537) );
  NANDN U10367 ( .A(n8245), .B(n8244), .Z(n8249) );
  OR U10368 ( .A(n8247), .B(n8246), .Z(n8248) );
  NAND U10369 ( .A(n8249), .B(n8248), .Z(n8944) );
  NANDN U10370 ( .A(n8251), .B(n8250), .Z(n8255) );
  NAND U10371 ( .A(n8253), .B(n8252), .Z(n8254) );
  NAND U10372 ( .A(n8255), .B(n8254), .Z(n8501) );
  NANDN U10373 ( .A(n8257), .B(n8256), .Z(n8261) );
  NANDN U10374 ( .A(n8259), .B(n8258), .Z(n8260) );
  NAND U10375 ( .A(n8261), .B(n8260), .Z(n8499) );
  NANDN U10376 ( .A(n8263), .B(n8262), .Z(n8267) );
  NAND U10377 ( .A(n8265), .B(n8264), .Z(n8266) );
  NAND U10378 ( .A(n8267), .B(n8266), .Z(n8498) );
  XNOR U10379 ( .A(n8501), .B(n8500), .Z(n8942) );
  XOR U10380 ( .A(n8944), .B(n8945), .Z(n8534) );
  NANDN U10381 ( .A(n8273), .B(n8272), .Z(n8277) );
  NAND U10382 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U10383 ( .A(n8277), .B(n8276), .Z(n8519) );
  NANDN U10384 ( .A(n8279), .B(n8278), .Z(n8283) );
  NAND U10385 ( .A(n8281), .B(n8280), .Z(n8282) );
  NAND U10386 ( .A(n8283), .B(n8282), .Z(n8517) );
  NANDN U10387 ( .A(n8285), .B(n8284), .Z(n8289) );
  NAND U10388 ( .A(n8287), .B(n8286), .Z(n8288) );
  NAND U10389 ( .A(n8289), .B(n8288), .Z(n8516) );
  XNOR U10390 ( .A(n8519), .B(n8518), .Z(n8535) );
  XNOR U10391 ( .A(n8534), .B(n8535), .Z(n8536) );
  XOR U10392 ( .A(n8537), .B(n8536), .Z(n8649) );
  XNOR U10393 ( .A(n8650), .B(n8649), .Z(n8651) );
  XNOR U10394 ( .A(n8652), .B(n8651), .Z(n8897) );
  XNOR U10395 ( .A(n8896), .B(n8897), .Z(n8463) );
  XOR U10396 ( .A(n8462), .B(n8463), .Z(n8465) );
  XNOR U10397 ( .A(n8464), .B(n8465), .Z(n8471) );
  NANDN U10398 ( .A(n8295), .B(n8294), .Z(n8299) );
  NANDN U10399 ( .A(n8297), .B(n8296), .Z(n8298) );
  AND U10400 ( .A(n8299), .B(n8298), .Z(n8468) );
  XNOR U10401 ( .A(n8469), .B(n8468), .Z(n8470) );
  XOR U10402 ( .A(n8471), .B(n8470), .Z(n8878) );
  OR U10403 ( .A(n8301), .B(n8300), .Z(n8305) );
  NANDN U10404 ( .A(n8303), .B(n8302), .Z(n8304) );
  AND U10405 ( .A(n8305), .B(n8304), .Z(n8876) );
  NANDN U10406 ( .A(n8307), .B(n8306), .Z(n8311) );
  NAND U10407 ( .A(n8309), .B(n8308), .Z(n8310) );
  NAND U10408 ( .A(n8311), .B(n8310), .Z(n8733) );
  NANDN U10409 ( .A(n8313), .B(n8312), .Z(n8317) );
  NAND U10410 ( .A(n8315), .B(n8314), .Z(n8316) );
  NAND U10411 ( .A(n8317), .B(n8316), .Z(n8730) );
  NANDN U10412 ( .A(n8323), .B(n8322), .Z(n8327) );
  NAND U10413 ( .A(n8325), .B(n8324), .Z(n8326) );
  AND U10414 ( .A(n8327), .B(n8326), .Z(n9004) );
  NANDN U10415 ( .A(n8329), .B(n8328), .Z(n8333) );
  NANDN U10416 ( .A(n8331), .B(n8330), .Z(n8332) );
  NAND U10417 ( .A(n8333), .B(n8332), .Z(n9005) );
  NANDN U10418 ( .A(n8335), .B(n8334), .Z(n8339) );
  NAND U10419 ( .A(n8337), .B(n8336), .Z(n8338) );
  NAND U10420 ( .A(n8339), .B(n8338), .Z(n8630) );
  NANDN U10421 ( .A(n8341), .B(n8340), .Z(n8345) );
  NAND U10422 ( .A(n8343), .B(n8342), .Z(n8344) );
  NAND U10423 ( .A(n8345), .B(n8344), .Z(n8628) );
  NANDN U10424 ( .A(n8347), .B(n8346), .Z(n8351) );
  NAND U10425 ( .A(n8349), .B(n8348), .Z(n8350) );
  NAND U10426 ( .A(n8351), .B(n8350), .Z(n8627) );
  XNOR U10427 ( .A(n8630), .B(n8629), .Z(n9006) );
  NANDN U10428 ( .A(n8353), .B(n8352), .Z(n8357) );
  NAND U10429 ( .A(n8355), .B(n8354), .Z(n8356) );
  NAND U10430 ( .A(n8357), .B(n8356), .Z(n8681) );
  NANDN U10431 ( .A(n8359), .B(n8358), .Z(n8363) );
  NAND U10432 ( .A(n8361), .B(n8360), .Z(n8362) );
  AND U10433 ( .A(n8363), .B(n8362), .Z(n8989) );
  OR U10434 ( .A(n8365), .B(n8364), .Z(n8985) );
  NANDN U10435 ( .A(n8367), .B(n8366), .Z(n8371) );
  NANDN U10436 ( .A(n8369), .B(n8368), .Z(n8370) );
  NAND U10437 ( .A(n8371), .B(n8370), .Z(n8984) );
  XNOR U10438 ( .A(n8985), .B(n8984), .Z(n8986) );
  NANDN U10439 ( .A(n8373), .B(n8372), .Z(n8377) );
  NAND U10440 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U10441 ( .A(n8377), .B(n8376), .Z(n8987) );
  XNOR U10442 ( .A(n8986), .B(n8987), .Z(n8988) );
  IV U10443 ( .A(n8596), .Z(n8598) );
  NAND U10444 ( .A(n8379), .B(n8378), .Z(n8383) );
  NAND U10445 ( .A(n8381), .B(n8380), .Z(n8382) );
  NAND U10446 ( .A(n8383), .B(n8382), .Z(n8597) );
  NANDN U10447 ( .A(n8385), .B(n8384), .Z(n8389) );
  NAND U10448 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U10449 ( .A(n8389), .B(n8388), .Z(n8979) );
  NANDN U10450 ( .A(n8391), .B(n8390), .Z(n8395) );
  NAND U10451 ( .A(n8393), .B(n8392), .Z(n8394) );
  NAND U10452 ( .A(n8395), .B(n8394), .Z(n8978) );
  NANDN U10453 ( .A(n8397), .B(n8396), .Z(n8401) );
  NAND U10454 ( .A(n8399), .B(n8398), .Z(n8400) );
  NAND U10455 ( .A(n8401), .B(n8400), .Z(n8981) );
  XOR U10456 ( .A(n8980), .B(n8981), .Z(n8837) );
  NANDN U10457 ( .A(n8403), .B(n8402), .Z(n8407) );
  NAND U10458 ( .A(n8405), .B(n8404), .Z(n8406) );
  AND U10459 ( .A(n8407), .B(n8406), .Z(n8834) );
  XOR U10460 ( .A(n8837), .B(n8836), .Z(n8600) );
  XNOR U10461 ( .A(n8597), .B(n8600), .Z(n8412) );
  XOR U10462 ( .A(n8598), .B(n8412), .Z(n8682) );
  XNOR U10463 ( .A(n8681), .B(n8682), .Z(n8413) );
  XOR U10464 ( .A(n8683), .B(n8413), .Z(n8656) );
  NANDN U10465 ( .A(n8415), .B(n8414), .Z(n8419) );
  NANDN U10466 ( .A(n8417), .B(n8416), .Z(n8418) );
  NAND U10467 ( .A(n8419), .B(n8418), .Z(n8687) );
  NANDN U10468 ( .A(n8421), .B(n8420), .Z(n8425) );
  NANDN U10469 ( .A(n8423), .B(n8422), .Z(n8424) );
  NAND U10470 ( .A(n8425), .B(n8424), .Z(n8684) );
  NAND U10471 ( .A(n8427), .B(n8426), .Z(n8431) );
  OR U10472 ( .A(n8429), .B(n8428), .Z(n8430) );
  NAND U10473 ( .A(n8431), .B(n8430), .Z(n8685) );
  XNOR U10474 ( .A(n8684), .B(n8685), .Z(n8686) );
  XOR U10475 ( .A(n8687), .B(n8686), .Z(n8655) );
  XNOR U10476 ( .A(n8656), .B(n8655), .Z(n8657) );
  XNOR U10477 ( .A(n8658), .B(n8657), .Z(n8731) );
  XOR U10478 ( .A(n8730), .B(n8731), .Z(n8732) );
  XNOR U10479 ( .A(n8733), .B(n8732), .Z(n8645) );
  NAND U10480 ( .A(n8433), .B(n8432), .Z(n8437) );
  NANDN U10481 ( .A(n8435), .B(n8434), .Z(n8436) );
  NAND U10482 ( .A(n8437), .B(n8436), .Z(n8721) );
  OR U10483 ( .A(n8439), .B(n8438), .Z(n8443) );
  NAND U10484 ( .A(n8441), .B(n8440), .Z(n8442) );
  NAND U10485 ( .A(n8443), .B(n8442), .Z(n8718) );
  NANDN U10486 ( .A(n8445), .B(n8444), .Z(n8449) );
  OR U10487 ( .A(n8447), .B(n8446), .Z(n8448) );
  AND U10488 ( .A(n8449), .B(n8448), .Z(n8719) );
  XNOR U10489 ( .A(n8718), .B(n8719), .Z(n8720) );
  XNOR U10490 ( .A(n8721), .B(n8720), .Z(n8643) );
  NAND U10491 ( .A(n8451), .B(n8450), .Z(n8455) );
  NAND U10492 ( .A(n8453), .B(n8452), .Z(n8454) );
  AND U10493 ( .A(n8455), .B(n8454), .Z(n8644) );
  XOR U10494 ( .A(n8643), .B(n8644), .Z(n8646) );
  XOR U10495 ( .A(n8645), .B(n8646), .Z(n8877) );
  XNOR U10496 ( .A(n8876), .B(n8877), .Z(n8879) );
  XNOR U10497 ( .A(n8878), .B(n8879), .Z(n8459) );
  XNOR U10498 ( .A(n8458), .B(n8459), .Z(o[3]) );
  NANDN U10499 ( .A(n8457), .B(n8456), .Z(n8461) );
  NANDN U10500 ( .A(n8459), .B(n8458), .Z(n8460) );
  NAND U10501 ( .A(n8461), .B(n8460), .Z(n9292) );
  NANDN U10502 ( .A(n8463), .B(n8462), .Z(n8467) );
  NANDN U10503 ( .A(n8465), .B(n8464), .Z(n8466) );
  NAND U10504 ( .A(n8467), .B(n8466), .Z(n9281) );
  NANDN U10505 ( .A(n8469), .B(n8468), .Z(n8473) );
  NANDN U10506 ( .A(n8471), .B(n8470), .Z(n8472) );
  NAND U10507 ( .A(n8473), .B(n8472), .Z(n9300) );
  NANDN U10508 ( .A(n8475), .B(n8474), .Z(n8479) );
  NANDN U10509 ( .A(n8477), .B(n8476), .Z(n8478) );
  NAND U10510 ( .A(n8479), .B(n8478), .Z(n9149) );
  NANDN U10511 ( .A(n8481), .B(n8480), .Z(n8485) );
  NANDN U10512 ( .A(n8483), .B(n8482), .Z(n8484) );
  NAND U10513 ( .A(n8485), .B(n8484), .Z(n9147) );
  NANDN U10514 ( .A(n8487), .B(n8486), .Z(n8491) );
  NANDN U10515 ( .A(n8489), .B(n8488), .Z(n8490) );
  NAND U10516 ( .A(n8491), .B(n8490), .Z(n9255) );
  NANDN U10517 ( .A(n8493), .B(n8492), .Z(n8497) );
  NANDN U10518 ( .A(n8495), .B(n8494), .Z(n8496) );
  NAND U10519 ( .A(n8497), .B(n8496), .Z(n9252) );
  OR U10520 ( .A(n8499), .B(n8498), .Z(n8503) );
  NANDN U10521 ( .A(n8501), .B(n8500), .Z(n8502) );
  AND U10522 ( .A(n8503), .B(n8502), .Z(n9253) );
  XNOR U10523 ( .A(n9252), .B(n9253), .Z(n9254) );
  XOR U10524 ( .A(n9255), .B(n9254), .Z(n9146) );
  XNOR U10525 ( .A(n9147), .B(n9146), .Z(n9148) );
  XNOR U10526 ( .A(n9149), .B(n9148), .Z(n9150) );
  NANDN U10527 ( .A(n8505), .B(n8504), .Z(n8509) );
  NANDN U10528 ( .A(n8507), .B(n8506), .Z(n8508) );
  AND U10529 ( .A(n8509), .B(n8508), .Z(n9151) );
  XOR U10530 ( .A(n9150), .B(n9151), .Z(n9153) );
  OR U10531 ( .A(n8511), .B(n8510), .Z(n8515) );
  NANDN U10532 ( .A(n8513), .B(n8512), .Z(n8514) );
  NAND U10533 ( .A(n8515), .B(n8514), .Z(n9137) );
  OR U10534 ( .A(n8517), .B(n8516), .Z(n8521) );
  NANDN U10535 ( .A(n8519), .B(n8518), .Z(n8520) );
  NAND U10536 ( .A(n8521), .B(n8520), .Z(n9134) );
  OR U10537 ( .A(n8523), .B(n8522), .Z(n8527) );
  NANDN U10538 ( .A(n8525), .B(n8524), .Z(n8526) );
  AND U10539 ( .A(n8527), .B(n8526), .Z(n9135) );
  XNOR U10540 ( .A(n9134), .B(n9135), .Z(n9136) );
  XNOR U10541 ( .A(n9137), .B(n9136), .Z(n9152) );
  XNOR U10542 ( .A(n9153), .B(n9152), .Z(n9097) );
  NANDN U10543 ( .A(n8529), .B(n8528), .Z(n8533) );
  NAND U10544 ( .A(n8531), .B(n8530), .Z(n8532) );
  NAND U10545 ( .A(n8533), .B(n8532), .Z(n9095) );
  OR U10546 ( .A(n8543), .B(n8542), .Z(n8547) );
  NANDN U10547 ( .A(n8545), .B(n8544), .Z(n8546) );
  NAND U10548 ( .A(n8547), .B(n8546), .Z(n9043) );
  XNOR U10549 ( .A(n9042), .B(n9043), .Z(n9044) );
  XOR U10550 ( .A(n9045), .B(n9044), .Z(n9094) );
  XNOR U10551 ( .A(n9095), .B(n9094), .Z(n9096) );
  XNOR U10552 ( .A(n9097), .B(n9096), .Z(n9279) );
  NANDN U10553 ( .A(n8549), .B(n8548), .Z(n8553) );
  NAND U10554 ( .A(n8551), .B(n8550), .Z(n8552) );
  NAND U10555 ( .A(n8553), .B(n8552), .Z(n9063) );
  NANDN U10556 ( .A(n8555), .B(n8554), .Z(n8559) );
  NANDN U10557 ( .A(n8557), .B(n8556), .Z(n8558) );
  NAND U10558 ( .A(n8559), .B(n8558), .Z(n9061) );
  NANDN U10559 ( .A(n8561), .B(n8560), .Z(n8565) );
  NANDN U10560 ( .A(n8563), .B(n8562), .Z(n8564) );
  NAND U10561 ( .A(n8565), .B(n8564), .Z(n9182) );
  OR U10562 ( .A(n8567), .B(n8566), .Z(n8571) );
  NAND U10563 ( .A(n8569), .B(n8568), .Z(n8570) );
  NAND U10564 ( .A(n8571), .B(n8570), .Z(n9181) );
  OR U10565 ( .A(n8573), .B(n8572), .Z(n8577) );
  NANDN U10566 ( .A(n8575), .B(n8574), .Z(n8576) );
  NAND U10567 ( .A(n8577), .B(n8576), .Z(n9180) );
  XOR U10568 ( .A(n9182), .B(n9183), .Z(n9211) );
  OR U10569 ( .A(n8579), .B(n8578), .Z(n8583) );
  NAND U10570 ( .A(n8581), .B(n8580), .Z(n8582) );
  NAND U10571 ( .A(n8583), .B(n8582), .Z(n9208) );
  NANDN U10572 ( .A(n8585), .B(n8584), .Z(n8589) );
  NAND U10573 ( .A(n8587), .B(n8586), .Z(n8588) );
  AND U10574 ( .A(n8589), .B(n8588), .Z(n9209) );
  XNOR U10575 ( .A(n9208), .B(n9209), .Z(n9210) );
  XOR U10576 ( .A(n9211), .B(n9210), .Z(n9194) );
  OR U10577 ( .A(n8591), .B(n8590), .Z(n8595) );
  NAND U10578 ( .A(n8593), .B(n8592), .Z(n8594) );
  NAND U10579 ( .A(n8595), .B(n8594), .Z(n9207) );
  NANDN U10580 ( .A(n8596), .B(n8597), .Z(n8602) );
  NOR U10581 ( .A(n8598), .B(n8597), .Z(n8599) );
  OR U10582 ( .A(n8600), .B(n8599), .Z(n8601) );
  NAND U10583 ( .A(n8602), .B(n8601), .Z(n9205) );
  NANDN U10584 ( .A(n8604), .B(n8603), .Z(n8608) );
  NANDN U10585 ( .A(n8606), .B(n8605), .Z(n8607) );
  NAND U10586 ( .A(n8608), .B(n8607), .Z(n9229) );
  OR U10587 ( .A(n8610), .B(n8609), .Z(n8614) );
  NANDN U10588 ( .A(n8612), .B(n8611), .Z(n8613) );
  NAND U10589 ( .A(n8614), .B(n8613), .Z(n9226) );
  NAND U10590 ( .A(n8616), .B(n8615), .Z(n8620) );
  NANDN U10591 ( .A(n8618), .B(n8617), .Z(n8619) );
  AND U10592 ( .A(n8620), .B(n8619), .Z(n9227) );
  XNOR U10593 ( .A(n9226), .B(n9227), .Z(n9228) );
  XNOR U10594 ( .A(n9229), .B(n9228), .Z(n9235) );
  OR U10595 ( .A(n8622), .B(n8621), .Z(n8626) );
  NANDN U10596 ( .A(n8624), .B(n8623), .Z(n8625) );
  NAND U10597 ( .A(n8626), .B(n8625), .Z(n9233) );
  OR U10598 ( .A(n8628), .B(n8627), .Z(n8632) );
  NANDN U10599 ( .A(n8630), .B(n8629), .Z(n8631) );
  AND U10600 ( .A(n8632), .B(n8631), .Z(n9232) );
  XNOR U10601 ( .A(n9233), .B(n9232), .Z(n9234) );
  XOR U10602 ( .A(n9235), .B(n9234), .Z(n9204) );
  XNOR U10603 ( .A(n9205), .B(n9204), .Z(n9206) );
  XNOR U10604 ( .A(n9207), .B(n9206), .Z(n9192) );
  XOR U10605 ( .A(n9192), .B(n9193), .Z(n9195) );
  XOR U10606 ( .A(n9194), .B(n9195), .Z(n9060) );
  XOR U10607 ( .A(n9061), .B(n9060), .Z(n9062) );
  XNOR U10608 ( .A(n9063), .B(n9062), .Z(n9276) );
  NANDN U10609 ( .A(n8638), .B(n8637), .Z(n8642) );
  NANDN U10610 ( .A(n8640), .B(n8639), .Z(n8641) );
  NAND U10611 ( .A(n8642), .B(n8641), .Z(n9277) );
  XNOR U10612 ( .A(n9276), .B(n9277), .Z(n9278) );
  XOR U10613 ( .A(n9279), .B(n9278), .Z(n9299) );
  NANDN U10614 ( .A(n8644), .B(n8643), .Z(n8648) );
  OR U10615 ( .A(n8646), .B(n8645), .Z(n8647) );
  NAND U10616 ( .A(n8648), .B(n8647), .Z(n9298) );
  XNOR U10617 ( .A(n9299), .B(n9298), .Z(n9301) );
  XNOR U10618 ( .A(n9300), .B(n9301), .Z(n9280) );
  XNOR U10619 ( .A(n9281), .B(n9280), .Z(n9283) );
  NANDN U10620 ( .A(n8650), .B(n8649), .Z(n8654) );
  NAND U10621 ( .A(n8652), .B(n8651), .Z(n8653) );
  NAND U10622 ( .A(n8654), .B(n8653), .Z(n9101) );
  NANDN U10623 ( .A(n8660), .B(n8659), .Z(n8664) );
  NAND U10624 ( .A(n8662), .B(n8661), .Z(n8663) );
  NAND U10625 ( .A(n8664), .B(n8663), .Z(n9039) );
  NANDN U10626 ( .A(n8666), .B(n8665), .Z(n8670) );
  NAND U10627 ( .A(n8668), .B(n8667), .Z(n8669) );
  NAND U10628 ( .A(n8670), .B(n8669), .Z(n9037) );
  NANDN U10629 ( .A(n8672), .B(n8671), .Z(n8676) );
  NAND U10630 ( .A(n8674), .B(n8673), .Z(n8675) );
  AND U10631 ( .A(n8676), .B(n8675), .Z(n9036) );
  XNOR U10632 ( .A(n9037), .B(n9036), .Z(n9038) );
  XNOR U10633 ( .A(n9039), .B(n9038), .Z(n9099) );
  XNOR U10634 ( .A(n9098), .B(n9099), .Z(n9100) );
  XNOR U10635 ( .A(n9101), .B(n9100), .Z(n9266) );
  NANDN U10636 ( .A(n8685), .B(n8684), .Z(n8689) );
  NAND U10637 ( .A(n8687), .B(n8686), .Z(n8688) );
  AND U10638 ( .A(n8689), .B(n8688), .Z(n9049) );
  XOR U10639 ( .A(n9048), .B(n9049), .Z(n9051) );
  OR U10640 ( .A(n8691), .B(n8690), .Z(n8695) );
  NANDN U10641 ( .A(n8693), .B(n8692), .Z(n8694) );
  NAND U10642 ( .A(n8695), .B(n8694), .Z(n9050) );
  XNOR U10643 ( .A(n9051), .B(n9050), .Z(n9131) );
  NANDN U10644 ( .A(n8697), .B(n8696), .Z(n8701) );
  NAND U10645 ( .A(n8699), .B(n8698), .Z(n8700) );
  NAND U10646 ( .A(n8701), .B(n8700), .Z(n9128) );
  NAND U10647 ( .A(n8703), .B(n8702), .Z(n8707) );
  NANDN U10648 ( .A(n8705), .B(n8704), .Z(n8706) );
  NAND U10649 ( .A(n8707), .B(n8706), .Z(n9129) );
  XNOR U10650 ( .A(n9128), .B(n9129), .Z(n9130) );
  XOR U10651 ( .A(n9131), .B(n9130), .Z(n9123) );
  NANDN U10652 ( .A(n8709), .B(n8708), .Z(n8713) );
  NANDN U10653 ( .A(n8711), .B(n8710), .Z(n8712) );
  AND U10654 ( .A(n8713), .B(n8712), .Z(n9122) );
  XOR U10655 ( .A(n9123), .B(n9122), .Z(n9124) );
  XNOR U10656 ( .A(n9125), .B(n9124), .Z(n9264) );
  XNOR U10657 ( .A(n9264), .B(n9265), .Z(n9267) );
  XOR U10658 ( .A(n9266), .B(n9267), .Z(n9079) );
  NANDN U10659 ( .A(n8719), .B(n8718), .Z(n8723) );
  NAND U10660 ( .A(n8721), .B(n8720), .Z(n8722) );
  NAND U10661 ( .A(n8723), .B(n8722), .Z(n9077) );
  NANDN U10662 ( .A(n8725), .B(n8724), .Z(n8729) );
  NAND U10663 ( .A(n8727), .B(n8726), .Z(n8728) );
  AND U10664 ( .A(n8729), .B(n8728), .Z(n9076) );
  XNOR U10665 ( .A(n9077), .B(n9076), .Z(n9078) );
  XNOR U10666 ( .A(n9079), .B(n9078), .Z(n9307) );
  OR U10667 ( .A(n8731), .B(n8730), .Z(n8735) );
  NAND U10668 ( .A(n8733), .B(n8732), .Z(n8734) );
  NAND U10669 ( .A(n8735), .B(n8734), .Z(n9270) );
  NANDN U10670 ( .A(n8741), .B(n8740), .Z(n8745) );
  NANDN U10671 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U10672 ( .A(n8745), .B(n8744), .Z(n9189) );
  NANDN U10673 ( .A(n8747), .B(n8746), .Z(n8751) );
  NAND U10674 ( .A(n8749), .B(n8748), .Z(n8750) );
  NAND U10675 ( .A(n8751), .B(n8750), .Z(n9186) );
  NANDN U10676 ( .A(n8753), .B(n8752), .Z(n8757) );
  NANDN U10677 ( .A(n8755), .B(n8754), .Z(n8756) );
  NAND U10678 ( .A(n8757), .B(n8756), .Z(n9187) );
  XNOR U10679 ( .A(n9186), .B(n9187), .Z(n9188) );
  XNOR U10680 ( .A(n9189), .B(n9188), .Z(n9054) );
  XNOR U10681 ( .A(n9054), .B(n9055), .Z(n9056) );
  XNOR U10682 ( .A(n9057), .B(n9056), .Z(n9271) );
  XNOR U10683 ( .A(n9270), .B(n9271), .Z(n9272) );
  OR U10684 ( .A(n8763), .B(n8762), .Z(n8767) );
  NAND U10685 ( .A(n8765), .B(n8764), .Z(n8766) );
  NAND U10686 ( .A(n8767), .B(n8766), .Z(n9069) );
  NANDN U10687 ( .A(n8769), .B(n8768), .Z(n8773) );
  OR U10688 ( .A(n8771), .B(n8770), .Z(n8772) );
  NAND U10689 ( .A(n8773), .B(n8772), .Z(n9066) );
  NANDN U10690 ( .A(n8775), .B(n8774), .Z(n8779) );
  NAND U10691 ( .A(n8777), .B(n8776), .Z(n8778) );
  AND U10692 ( .A(n8779), .B(n8778), .Z(n9067) );
  XNOR U10693 ( .A(n9066), .B(n9067), .Z(n9068) );
  XOR U10694 ( .A(n9069), .B(n9068), .Z(n9273) );
  XOR U10695 ( .A(n9272), .B(n9273), .Z(n9304) );
  NANDN U10696 ( .A(n8781), .B(n8780), .Z(n8785) );
  NANDN U10697 ( .A(n8783), .B(n8782), .Z(n8784) );
  NAND U10698 ( .A(n8785), .B(n8784), .Z(n9091) );
  NAND U10699 ( .A(n8787), .B(n8786), .Z(n8791) );
  NAND U10700 ( .A(n8789), .B(n8788), .Z(n8790) );
  NAND U10701 ( .A(n8791), .B(n8790), .Z(n9075) );
  NANDN U10702 ( .A(n8793), .B(n8792), .Z(n8797) );
  NANDN U10703 ( .A(n8795), .B(n8794), .Z(n8796) );
  NAND U10704 ( .A(n8797), .B(n8796), .Z(n9110) );
  NANDN U10705 ( .A(n8799), .B(n8798), .Z(n8803) );
  NANDN U10706 ( .A(n8801), .B(n8800), .Z(n8802) );
  NAND U10707 ( .A(n8803), .B(n8802), .Z(n9159) );
  OR U10708 ( .A(n8805), .B(n8804), .Z(n8809) );
  NANDN U10709 ( .A(n8807), .B(n8806), .Z(n8808) );
  NAND U10710 ( .A(n8809), .B(n8808), .Z(n9156) );
  NANDN U10711 ( .A(n8811), .B(n8810), .Z(n8815) );
  NAND U10712 ( .A(n8813), .B(n8812), .Z(n8814) );
  AND U10713 ( .A(n8815), .B(n8814), .Z(n9157) );
  XNOR U10714 ( .A(n9156), .B(n9157), .Z(n9158) );
  XNOR U10715 ( .A(n9159), .B(n9158), .Z(n9111) );
  XNOR U10716 ( .A(n9110), .B(n9111), .Z(n9112) );
  OR U10717 ( .A(n8817), .B(n8816), .Z(n8821) );
  NANDN U10718 ( .A(n8819), .B(n8818), .Z(n8820) );
  NAND U10719 ( .A(n8821), .B(n8820), .Z(n9241) );
  OR U10720 ( .A(n8823), .B(n8822), .Z(n8827) );
  NANDN U10721 ( .A(n8825), .B(n8824), .Z(n8826) );
  NAND U10722 ( .A(n8827), .B(n8826), .Z(n9238) );
  OR U10723 ( .A(n8829), .B(n8828), .Z(n8833) );
  NANDN U10724 ( .A(n8831), .B(n8830), .Z(n8832) );
  AND U10725 ( .A(n8833), .B(n8832), .Z(n9239) );
  XNOR U10726 ( .A(n9238), .B(n9239), .Z(n9240) );
  XNOR U10727 ( .A(n9241), .B(n9240), .Z(n9201) );
  OR U10728 ( .A(n8835), .B(n8834), .Z(n8839) );
  NAND U10729 ( .A(n8837), .B(n8836), .Z(n8838) );
  NAND U10730 ( .A(n8839), .B(n8838), .Z(n9261) );
  OR U10731 ( .A(n8841), .B(n8840), .Z(n8845) );
  NANDN U10732 ( .A(n8843), .B(n8842), .Z(n8844) );
  NAND U10733 ( .A(n8845), .B(n8844), .Z(n9258) );
  OR U10734 ( .A(n8847), .B(n8846), .Z(n8851) );
  NANDN U10735 ( .A(n8849), .B(n8848), .Z(n8850) );
  AND U10736 ( .A(n8851), .B(n8850), .Z(n9259) );
  XNOR U10737 ( .A(n9258), .B(n9259), .Z(n9260) );
  XOR U10738 ( .A(n9261), .B(n9260), .Z(n9198) );
  OR U10739 ( .A(n8853), .B(n8852), .Z(n8857) );
  NANDN U10740 ( .A(n8855), .B(n8854), .Z(n8856) );
  NAND U10741 ( .A(n8857), .B(n8856), .Z(n9199) );
  XNOR U10742 ( .A(n9198), .B(n9199), .Z(n9200) );
  XOR U10743 ( .A(n9201), .B(n9200), .Z(n9113) );
  XNOR U10744 ( .A(n9112), .B(n9113), .Z(n9072) );
  OR U10745 ( .A(n8859), .B(n8858), .Z(n8863) );
  NAND U10746 ( .A(n8861), .B(n8860), .Z(n8862) );
  AND U10747 ( .A(n8863), .B(n8862), .Z(n9073) );
  XNOR U10748 ( .A(n9072), .B(n9073), .Z(n9074) );
  XOR U10749 ( .A(n9075), .B(n9074), .Z(n9088) );
  NANDN U10750 ( .A(n8865), .B(n8864), .Z(n8869) );
  NAND U10751 ( .A(n8867), .B(n8866), .Z(n8868) );
  AND U10752 ( .A(n8869), .B(n8868), .Z(n9089) );
  XNOR U10753 ( .A(n9088), .B(n9089), .Z(n9090) );
  XNOR U10754 ( .A(n9091), .B(n9090), .Z(n9305) );
  XNOR U10755 ( .A(n9304), .B(n9305), .Z(n9306) );
  XOR U10756 ( .A(n9307), .B(n9306), .Z(n9282) );
  XNOR U10757 ( .A(n9283), .B(n9282), .Z(n9293) );
  XNOR U10758 ( .A(n9292), .B(n9293), .Z(n9294) );
  OR U10759 ( .A(n8871), .B(n8870), .Z(n8875) );
  NANDN U10760 ( .A(n8873), .B(n8872), .Z(n8874) );
  AND U10761 ( .A(n8875), .B(n8874), .Z(n9286) );
  OR U10762 ( .A(n8877), .B(n8876), .Z(n8881) );
  NANDN U10763 ( .A(n8879), .B(n8878), .Z(n8880) );
  AND U10764 ( .A(n8881), .B(n8880), .Z(n9287) );
  XOR U10765 ( .A(n9286), .B(n9287), .Z(n9289) );
  NANDN U10766 ( .A(n8883), .B(n8882), .Z(n8887) );
  NAND U10767 ( .A(n8885), .B(n8884), .Z(n8886) );
  NAND U10768 ( .A(n8887), .B(n8886), .Z(n9313) );
  NAND U10769 ( .A(n8889), .B(n8888), .Z(n8893) );
  NANDN U10770 ( .A(n8891), .B(n8890), .Z(n8892) );
  NAND U10771 ( .A(n8893), .B(n8892), .Z(n9310) );
  OR U10772 ( .A(n8895), .B(n8894), .Z(n8899) );
  NANDN U10773 ( .A(n8897), .B(n8896), .Z(n8898) );
  NAND U10774 ( .A(n8899), .B(n8898), .Z(n9083) );
  NANDN U10775 ( .A(n8901), .B(n8900), .Z(n8905) );
  NANDN U10776 ( .A(n8903), .B(n8902), .Z(n8904) );
  NAND U10777 ( .A(n8905), .B(n8904), .Z(n9140) );
  NANDN U10778 ( .A(n8907), .B(n8906), .Z(n8911) );
  NAND U10779 ( .A(n8909), .B(n8908), .Z(n8910) );
  NAND U10780 ( .A(n8911), .B(n8910), .Z(n9223) );
  OR U10781 ( .A(n8913), .B(n8912), .Z(n8917) );
  NANDN U10782 ( .A(n8915), .B(n8914), .Z(n8916) );
  NAND U10783 ( .A(n8917), .B(n8916), .Z(n9221) );
  OR U10784 ( .A(n8919), .B(n8918), .Z(n8923) );
  NAND U10785 ( .A(n8921), .B(n8920), .Z(n8922) );
  AND U10786 ( .A(n8923), .B(n8922), .Z(n9220) );
  XNOR U10787 ( .A(n9221), .B(n9220), .Z(n9222) );
  XOR U10788 ( .A(n9223), .B(n9222), .Z(n9141) );
  XOR U10789 ( .A(n9140), .B(n9141), .Z(n9143) );
  NANDN U10790 ( .A(n8925), .B(n8924), .Z(n8929) );
  NAND U10791 ( .A(n8927), .B(n8926), .Z(n8928) );
  NAND U10792 ( .A(n8929), .B(n8928), .Z(n9142) );
  XNOR U10793 ( .A(n9143), .B(n9142), .Z(n9107) );
  NANDN U10794 ( .A(n8931), .B(n8930), .Z(n8935) );
  OR U10795 ( .A(n8933), .B(n8932), .Z(n8934) );
  NAND U10796 ( .A(n8935), .B(n8934), .Z(n9104) );
  NANDN U10797 ( .A(n8937), .B(n8936), .Z(n8941) );
  NAND U10798 ( .A(n8939), .B(n8938), .Z(n8940) );
  NAND U10799 ( .A(n8941), .B(n8940), .Z(n9165) );
  OR U10800 ( .A(n8943), .B(n8942), .Z(n8947) );
  NANDN U10801 ( .A(n8945), .B(n8944), .Z(n8946) );
  NAND U10802 ( .A(n8947), .B(n8946), .Z(n9162) );
  OR U10803 ( .A(n8949), .B(n8948), .Z(n8953) );
  NANDN U10804 ( .A(n8951), .B(n8950), .Z(n8952) );
  AND U10805 ( .A(n8953), .B(n8952), .Z(n9163) );
  XNOR U10806 ( .A(n9162), .B(n9163), .Z(n9164) );
  XNOR U10807 ( .A(n9165), .B(n9164), .Z(n9105) );
  XNOR U10808 ( .A(n9104), .B(n9105), .Z(n9106) );
  XNOR U10809 ( .A(n9107), .B(n9106), .Z(n9035) );
  NAND U10810 ( .A(n8955), .B(n8954), .Z(n8959) );
  OR U10811 ( .A(n8957), .B(n8956), .Z(n8958) );
  NAND U10812 ( .A(n8959), .B(n8958), .Z(n9217) );
  OR U10813 ( .A(n8961), .B(n8960), .Z(n8965) );
  NANDN U10814 ( .A(n8963), .B(n8962), .Z(n8964) );
  NAND U10815 ( .A(n8965), .B(n8964), .Z(n9170) );
  NAND U10816 ( .A(n8967), .B(n8966), .Z(n8971) );
  NAND U10817 ( .A(n8969), .B(n8968), .Z(n8970) );
  AND U10818 ( .A(n8971), .B(n8970), .Z(n9168) );
  OR U10819 ( .A(n8973), .B(n8972), .Z(n8977) );
  NANDN U10820 ( .A(n8975), .B(n8974), .Z(n8976) );
  NAND U10821 ( .A(n8977), .B(n8976), .Z(n9244) );
  OR U10822 ( .A(n8979), .B(n8978), .Z(n8983) );
  NANDN U10823 ( .A(n8981), .B(n8980), .Z(n8982) );
  AND U10824 ( .A(n8983), .B(n8982), .Z(n9245) );
  XNOR U10825 ( .A(n9244), .B(n9245), .Z(n9246) );
  OR U10826 ( .A(n8985), .B(n8984), .Z(n9251) );
  NANDN U10827 ( .A(n8987), .B(n8986), .Z(n8991) );
  NANDN U10828 ( .A(n8989), .B(n8988), .Z(n8990) );
  NAND U10829 ( .A(n8991), .B(n8990), .Z(n9250) );
  XOR U10830 ( .A(n9246), .B(n9247), .Z(n9169) );
  XOR U10831 ( .A(n9170), .B(n9171), .Z(n9214) );
  OR U10832 ( .A(n8993), .B(n8992), .Z(n8997) );
  NANDN U10833 ( .A(n8995), .B(n8994), .Z(n8996) );
  NAND U10834 ( .A(n8997), .B(n8996), .Z(n9215) );
  XNOR U10835 ( .A(n9214), .B(n9215), .Z(n9216) );
  XNOR U10836 ( .A(n9217), .B(n9216), .Z(n9033) );
  OR U10837 ( .A(n8999), .B(n8998), .Z(n9003) );
  NANDN U10838 ( .A(n9001), .B(n9000), .Z(n9002) );
  NAND U10839 ( .A(n9003), .B(n9002), .Z(n9177) );
  OR U10840 ( .A(n9005), .B(n9004), .Z(n9009) );
  NANDN U10841 ( .A(n9007), .B(n9006), .Z(n9008) );
  NAND U10842 ( .A(n9009), .B(n9008), .Z(n9174) );
  NANDN U10843 ( .A(n9011), .B(n9010), .Z(n9015) );
  NANDN U10844 ( .A(n9013), .B(n9012), .Z(n9014) );
  AND U10845 ( .A(n9015), .B(n9014), .Z(n9175) );
  XNOR U10846 ( .A(n9174), .B(n9175), .Z(n9176) );
  XNOR U10847 ( .A(n9177), .B(n9176), .Z(n9116) );
  NANDN U10848 ( .A(n9017), .B(n9016), .Z(n9021) );
  NAND U10849 ( .A(n9019), .B(n9018), .Z(n9020) );
  AND U10850 ( .A(n9021), .B(n9020), .Z(n9117) );
  XNOR U10851 ( .A(n9116), .B(n9117), .Z(n9119) );
  XNOR U10852 ( .A(n9119), .B(n9118), .Z(n9032) );
  XNOR U10853 ( .A(n9033), .B(n9032), .Z(n9034) );
  XOR U10854 ( .A(n9035), .B(n9034), .Z(n9082) );
  XNOR U10855 ( .A(n9083), .B(n9082), .Z(n9085) );
  NANDN U10856 ( .A(n9027), .B(n9026), .Z(n9031) );
  NANDN U10857 ( .A(n9029), .B(n9028), .Z(n9030) );
  NAND U10858 ( .A(n9031), .B(n9030), .Z(n9084) );
  XOR U10859 ( .A(n9085), .B(n9084), .Z(n9311) );
  XNOR U10860 ( .A(n9310), .B(n9311), .Z(n9312) );
  XOR U10861 ( .A(n9313), .B(n9312), .Z(n9288) );
  XOR U10862 ( .A(n9289), .B(n9288), .Z(n9295) );
  XNOR U10863 ( .A(n9294), .B(n9295), .Z(o[4]) );
  NANDN U10864 ( .A(n9037), .B(n9036), .Z(n9041) );
  NAND U10865 ( .A(n9039), .B(n9038), .Z(n9040) );
  NAND U10866 ( .A(n9041), .B(n9040), .Z(n9324) );
  NANDN U10867 ( .A(n9043), .B(n9042), .Z(n9047) );
  NAND U10868 ( .A(n9045), .B(n9044), .Z(n9046) );
  NAND U10869 ( .A(n9047), .B(n9046), .Z(n9322) );
  NANDN U10870 ( .A(n9049), .B(n9048), .Z(n9053) );
  OR U10871 ( .A(n9051), .B(n9050), .Z(n9052) );
  AND U10872 ( .A(n9053), .B(n9052), .Z(n9321) );
  XNOR U10873 ( .A(n9322), .B(n9321), .Z(n9323) );
  XOR U10874 ( .A(n9324), .B(n9323), .Z(n9401) );
  NANDN U10875 ( .A(n9055), .B(n9054), .Z(n9059) );
  NAND U10876 ( .A(n9057), .B(n9056), .Z(n9058) );
  AND U10877 ( .A(n9059), .B(n9058), .Z(n9402) );
  XNOR U10878 ( .A(n9401), .B(n9402), .Z(n9403) );
  XOR U10879 ( .A(n9404), .B(n9403), .Z(n9417) );
  NAND U10880 ( .A(n9061), .B(n9060), .Z(n9065) );
  NAND U10881 ( .A(n9063), .B(n9062), .Z(n9064) );
  NAND U10882 ( .A(n9065), .B(n9064), .Z(n9414) );
  NANDN U10883 ( .A(n9067), .B(n9066), .Z(n9071) );
  NANDN U10884 ( .A(n9069), .B(n9068), .Z(n9070) );
  NAND U10885 ( .A(n9071), .B(n9070), .Z(n9411) );
  XNOR U10886 ( .A(n9411), .B(n9412), .Z(n9413) );
  XOR U10887 ( .A(n9414), .B(n9413), .Z(n9418) );
  NANDN U10888 ( .A(n9077), .B(n9076), .Z(n9081) );
  NAND U10889 ( .A(n9079), .B(n9078), .Z(n9080) );
  NAND U10890 ( .A(n9081), .B(n9080), .Z(n9420) );
  XOR U10891 ( .A(n9419), .B(n9420), .Z(n9435) );
  NAND U10892 ( .A(n9083), .B(n9082), .Z(n9087) );
  OR U10893 ( .A(n9085), .B(n9084), .Z(n9086) );
  AND U10894 ( .A(n9087), .B(n9086), .Z(n9432) );
  NANDN U10895 ( .A(n9089), .B(n9088), .Z(n9093) );
  NAND U10896 ( .A(n9091), .B(n9090), .Z(n9092) );
  NAND U10897 ( .A(n9093), .B(n9092), .Z(n9433) );
  XOR U10898 ( .A(n9432), .B(n9433), .Z(n9434) );
  XOR U10899 ( .A(n9435), .B(n9434), .Z(n9318) );
  NANDN U10900 ( .A(n9099), .B(n9098), .Z(n9103) );
  NAND U10901 ( .A(n9101), .B(n9100), .Z(n9102) );
  NAND U10902 ( .A(n9103), .B(n9102), .Z(n9398) );
  NANDN U10903 ( .A(n9105), .B(n9104), .Z(n9109) );
  NAND U10904 ( .A(n9107), .B(n9106), .Z(n9108) );
  NAND U10905 ( .A(n9109), .B(n9108), .Z(n9362) );
  NANDN U10906 ( .A(n9111), .B(n9110), .Z(n9115) );
  NAND U10907 ( .A(n9113), .B(n9112), .Z(n9114) );
  NAND U10908 ( .A(n9115), .B(n9114), .Z(n9359) );
  NAND U10909 ( .A(n9117), .B(n9116), .Z(n9121) );
  NANDN U10910 ( .A(n9119), .B(n9118), .Z(n9120) );
  NAND U10911 ( .A(n9121), .B(n9120), .Z(n9360) );
  XNOR U10912 ( .A(n9359), .B(n9360), .Z(n9361) );
  XNOR U10913 ( .A(n9362), .B(n9361), .Z(n9395) );
  OR U10914 ( .A(n9123), .B(n9122), .Z(n9127) );
  NANDN U10915 ( .A(n9125), .B(n9124), .Z(n9126) );
  AND U10916 ( .A(n9127), .B(n9126), .Z(n9396) );
  XNOR U10917 ( .A(n9395), .B(n9396), .Z(n9397) );
  XNOR U10918 ( .A(n9398), .B(n9397), .Z(n9437) );
  XNOR U10919 ( .A(n9436), .B(n9437), .Z(n9439) );
  NANDN U10920 ( .A(n9129), .B(n9128), .Z(n9133) );
  NAND U10921 ( .A(n9131), .B(n9130), .Z(n9132) );
  NAND U10922 ( .A(n9133), .B(n9132), .Z(n9368) );
  NANDN U10923 ( .A(n9135), .B(n9134), .Z(n9139) );
  NAND U10924 ( .A(n9137), .B(n9136), .Z(n9138) );
  NAND U10925 ( .A(n9139), .B(n9138), .Z(n9386) );
  NANDN U10926 ( .A(n9141), .B(n9140), .Z(n9145) );
  OR U10927 ( .A(n9143), .B(n9142), .Z(n9144) );
  AND U10928 ( .A(n9145), .B(n9144), .Z(n9383) );
  XOR U10929 ( .A(n9386), .B(n9385), .Z(n9365) );
  NANDN U10930 ( .A(n9151), .B(n9150), .Z(n9155) );
  OR U10931 ( .A(n9153), .B(n9152), .Z(n9154) );
  AND U10932 ( .A(n9155), .B(n9154), .Z(n9366) );
  XNOR U10933 ( .A(n9365), .B(n9366), .Z(n9367) );
  XNOR U10934 ( .A(n9368), .B(n9367), .Z(n9410) );
  NANDN U10935 ( .A(n9157), .B(n9156), .Z(n9161) );
  NAND U10936 ( .A(n9159), .B(n9158), .Z(n9160) );
  NAND U10937 ( .A(n9161), .B(n9160), .Z(n9340) );
  NANDN U10938 ( .A(n9163), .B(n9162), .Z(n9167) );
  NAND U10939 ( .A(n9165), .B(n9164), .Z(n9166) );
  NAND U10940 ( .A(n9167), .B(n9166), .Z(n9339) );
  OR U10941 ( .A(n9169), .B(n9168), .Z(n9173) );
  NANDN U10942 ( .A(n9171), .B(n9170), .Z(n9172) );
  AND U10943 ( .A(n9173), .B(n9172), .Z(n9342) );
  XNOR U10944 ( .A(n9341), .B(n9342), .Z(n9336) );
  NANDN U10945 ( .A(n9175), .B(n9174), .Z(n9179) );
  NANDN U10946 ( .A(n9177), .B(n9176), .Z(n9178) );
  NAND U10947 ( .A(n9179), .B(n9178), .Z(n9333) );
  OR U10948 ( .A(n9181), .B(n9180), .Z(n9185) );
  NANDN U10949 ( .A(n9183), .B(n9182), .Z(n9184) );
  AND U10950 ( .A(n9185), .B(n9184), .Z(n9334) );
  XNOR U10951 ( .A(n9333), .B(n9334), .Z(n9335) );
  XOR U10952 ( .A(n9336), .B(n9335), .Z(n9374) );
  NANDN U10953 ( .A(n9187), .B(n9186), .Z(n9191) );
  NAND U10954 ( .A(n9189), .B(n9188), .Z(n9190) );
  NAND U10955 ( .A(n9191), .B(n9190), .Z(n9371) );
  NANDN U10956 ( .A(n9193), .B(n9192), .Z(n9197) );
  OR U10957 ( .A(n9195), .B(n9194), .Z(n9196) );
  NAND U10958 ( .A(n9197), .B(n9196), .Z(n9372) );
  XNOR U10959 ( .A(n9371), .B(n9372), .Z(n9373) );
  XNOR U10960 ( .A(n9374), .B(n9373), .Z(n9407) );
  NANDN U10961 ( .A(n9199), .B(n9198), .Z(n9203) );
  NAND U10962 ( .A(n9201), .B(n9200), .Z(n9202) );
  NAND U10963 ( .A(n9203), .B(n9202), .Z(n9380) );
  NANDN U10964 ( .A(n9209), .B(n9208), .Z(n9213) );
  NAND U10965 ( .A(n9211), .B(n9210), .Z(n9212) );
  NAND U10966 ( .A(n9213), .B(n9212), .Z(n9377) );
  XOR U10967 ( .A(n9380), .B(n9379), .Z(n9330) );
  NANDN U10968 ( .A(n9215), .B(n9214), .Z(n9219) );
  NAND U10969 ( .A(n9217), .B(n9216), .Z(n9218) );
  NAND U10970 ( .A(n9219), .B(n9218), .Z(n9327) );
  NANDN U10971 ( .A(n9221), .B(n9220), .Z(n9225) );
  NANDN U10972 ( .A(n9223), .B(n9222), .Z(n9224) );
  AND U10973 ( .A(n9225), .B(n9224), .Z(n9347) );
  NANDN U10974 ( .A(n9227), .B(n9226), .Z(n9231) );
  NAND U10975 ( .A(n9229), .B(n9228), .Z(n9230) );
  AND U10976 ( .A(n9231), .B(n9230), .Z(n9348) );
  NANDN U10977 ( .A(n9233), .B(n9232), .Z(n9237) );
  NAND U10978 ( .A(n9235), .B(n9234), .Z(n9236) );
  NAND U10979 ( .A(n9237), .B(n9236), .Z(n9350) );
  XOR U10980 ( .A(n9349), .B(n9350), .Z(n9391) );
  NANDN U10981 ( .A(n9239), .B(n9238), .Z(n9243) );
  NAND U10982 ( .A(n9241), .B(n9240), .Z(n9242) );
  AND U10983 ( .A(n9243), .B(n9242), .Z(n9353) );
  NANDN U10984 ( .A(n9245), .B(n9244), .Z(n9249) );
  NAND U10985 ( .A(n9247), .B(n9246), .Z(n9248) );
  AND U10986 ( .A(n9249), .B(n9248), .Z(n9354) );
  OR U10987 ( .A(n9251), .B(n9250), .Z(n9346) );
  NANDN U10988 ( .A(n9253), .B(n9252), .Z(n9257) );
  NAND U10989 ( .A(n9255), .B(n9254), .Z(n9256) );
  AND U10990 ( .A(n9257), .B(n9256), .Z(n9345) );
  NANDN U10991 ( .A(n9259), .B(n9258), .Z(n9263) );
  NANDN U10992 ( .A(n9261), .B(n9260), .Z(n9262) );
  NAND U10993 ( .A(n9263), .B(n9262), .Z(n9389) );
  XNOR U10994 ( .A(n9390), .B(n9389), .Z(n9392) );
  XOR U10995 ( .A(n9391), .B(n9392), .Z(n9328) );
  XOR U10996 ( .A(n9327), .B(n9328), .Z(n9329) );
  XOR U10997 ( .A(n9330), .B(n9329), .Z(n9408) );
  XNOR U10998 ( .A(n9407), .B(n9408), .Z(n9409) );
  XOR U10999 ( .A(n9410), .B(n9409), .Z(n9438) );
  XNOR U11000 ( .A(n9439), .B(n9438), .Z(n9316) );
  OR U11001 ( .A(n9265), .B(n9264), .Z(n9269) );
  NANDN U11002 ( .A(n9267), .B(n9266), .Z(n9268) );
  NAND U11003 ( .A(n9269), .B(n9268), .Z(n9445) );
  NANDN U11004 ( .A(n9271), .B(n9270), .Z(n9275) );
  NANDN U11005 ( .A(n9273), .B(n9272), .Z(n9274) );
  AND U11006 ( .A(n9275), .B(n9274), .Z(n9442) );
  XNOR U11007 ( .A(n9442), .B(n9443), .Z(n9444) );
  XOR U11008 ( .A(n9445), .B(n9444), .Z(n9315) );
  XOR U11009 ( .A(n9316), .B(n9315), .Z(n9317) );
  XNOR U11010 ( .A(n9318), .B(n9317), .Z(n9429) );
  OR U11011 ( .A(n9281), .B(n9280), .Z(n9285) );
  OR U11012 ( .A(n9283), .B(n9282), .Z(n9284) );
  AND U11013 ( .A(n9285), .B(n9284), .Z(n9426) );
  OR U11014 ( .A(n9287), .B(n9286), .Z(n9291) );
  NAND U11015 ( .A(n9289), .B(n9288), .Z(n9290) );
  NAND U11016 ( .A(n9291), .B(n9290), .Z(n9427) );
  XNOR U11017 ( .A(n9426), .B(n9427), .Z(n9428) );
  XNOR U11018 ( .A(n9429), .B(n9428), .Z(n9425) );
  NANDN U11019 ( .A(n9293), .B(n9292), .Z(n9297) );
  NANDN U11020 ( .A(n9295), .B(n9294), .Z(n9296) );
  NAND U11021 ( .A(n9297), .B(n9296), .Z(n9423) );
  NANDN U11022 ( .A(n9299), .B(n9298), .Z(n9303) );
  NAND U11023 ( .A(n9301), .B(n9300), .Z(n9302) );
  AND U11024 ( .A(n9303), .B(n9302), .Z(n9451) );
  NANDN U11025 ( .A(n9305), .B(n9304), .Z(n9309) );
  NAND U11026 ( .A(n9307), .B(n9306), .Z(n9308) );
  NAND U11027 ( .A(n9309), .B(n9308), .Z(n9449) );
  XOR U11028 ( .A(n9449), .B(n9448), .Z(n9450) );
  XOR U11029 ( .A(n9451), .B(n9450), .Z(n9424) );
  XNOR U11030 ( .A(n9423), .B(n9424), .Z(n9314) );
  XNOR U11031 ( .A(n9425), .B(n9314), .Z(o[5]) );
  OR U11032 ( .A(n9316), .B(n9315), .Z(n9320) );
  NANDN U11033 ( .A(n9318), .B(n9317), .Z(n9319) );
  NAND U11034 ( .A(n9320), .B(n9319), .Z(n9469) );
  NANDN U11035 ( .A(n9322), .B(n9321), .Z(n9326) );
  NANDN U11036 ( .A(n9324), .B(n9323), .Z(n9325) );
  NAND U11037 ( .A(n9326), .B(n9325), .Z(n9485) );
  OR U11038 ( .A(n9328), .B(n9327), .Z(n9332) );
  NAND U11039 ( .A(n9330), .B(n9329), .Z(n9331) );
  AND U11040 ( .A(n9332), .B(n9331), .Z(n9484) );
  XNOR U11041 ( .A(n9485), .B(n9484), .Z(n9487) );
  NANDN U11042 ( .A(n9334), .B(n9333), .Z(n9338) );
  NANDN U11043 ( .A(n9336), .B(n9335), .Z(n9337) );
  AND U11044 ( .A(n9338), .B(n9337), .Z(n9502) );
  OR U11045 ( .A(n9340), .B(n9339), .Z(n9344) );
  NAND U11046 ( .A(n9342), .B(n9341), .Z(n9343) );
  NAND U11047 ( .A(n9344), .B(n9343), .Z(n9500) );
  OR U11048 ( .A(n9346), .B(n9345), .Z(n9507) );
  OR U11049 ( .A(n9348), .B(n9347), .Z(n9352) );
  NANDN U11050 ( .A(n9350), .B(n9349), .Z(n9351) );
  AND U11051 ( .A(n9352), .B(n9351), .Z(n9506) );
  XNOR U11052 ( .A(n9507), .B(n9506), .Z(n9508) );
  OR U11053 ( .A(n9354), .B(n9353), .Z(n9358) );
  NANDN U11054 ( .A(n9356), .B(n9355), .Z(n9357) );
  AND U11055 ( .A(n9358), .B(n9357), .Z(n9509) );
  XOR U11056 ( .A(n9500), .B(n9501), .Z(n9503) );
  XOR U11057 ( .A(n9487), .B(n9486), .Z(n9481) );
  NANDN U11058 ( .A(n9360), .B(n9359), .Z(n9364) );
  NAND U11059 ( .A(n9362), .B(n9361), .Z(n9363) );
  NAND U11060 ( .A(n9364), .B(n9363), .Z(n9478) );
  NANDN U11061 ( .A(n9366), .B(n9365), .Z(n9370) );
  NAND U11062 ( .A(n9368), .B(n9367), .Z(n9369) );
  NAND U11063 ( .A(n9370), .B(n9369), .Z(n9489) );
  NANDN U11064 ( .A(n9372), .B(n9371), .Z(n9376) );
  NAND U11065 ( .A(n9374), .B(n9373), .Z(n9375) );
  NAND U11066 ( .A(n9376), .B(n9375), .Z(n9488) );
  OR U11067 ( .A(n9378), .B(n9377), .Z(n9382) );
  NANDN U11068 ( .A(n9380), .B(n9379), .Z(n9381) );
  NAND U11069 ( .A(n9382), .B(n9381), .Z(n9497) );
  OR U11070 ( .A(n9384), .B(n9383), .Z(n9388) );
  NANDN U11071 ( .A(n9386), .B(n9385), .Z(n9387) );
  AND U11072 ( .A(n9388), .B(n9387), .Z(n9494) );
  OR U11073 ( .A(n9390), .B(n9389), .Z(n9394) );
  NANDN U11074 ( .A(n9392), .B(n9391), .Z(n9393) );
  NAND U11075 ( .A(n9394), .B(n9393), .Z(n9495) );
  XNOR U11076 ( .A(n9497), .B(n9496), .Z(n9491) );
  XNOR U11077 ( .A(n9490), .B(n9491), .Z(n9479) );
  XNOR U11078 ( .A(n9478), .B(n9479), .Z(n9480) );
  XNOR U11079 ( .A(n9481), .B(n9480), .Z(n9519) );
  NANDN U11080 ( .A(n9396), .B(n9395), .Z(n9400) );
  NAND U11081 ( .A(n9398), .B(n9397), .Z(n9399) );
  AND U11082 ( .A(n9400), .B(n9399), .Z(n9518) );
  XOR U11083 ( .A(n9519), .B(n9518), .Z(n9520) );
  NANDN U11084 ( .A(n9402), .B(n9401), .Z(n9406) );
  NAND U11085 ( .A(n9404), .B(n9403), .Z(n9405) );
  NAND U11086 ( .A(n9406), .B(n9405), .Z(n9515) );
  NANDN U11087 ( .A(n9412), .B(n9411), .Z(n9416) );
  NAND U11088 ( .A(n9414), .B(n9413), .Z(n9415) );
  AND U11089 ( .A(n9416), .B(n9415), .Z(n9513) );
  XNOR U11090 ( .A(n9515), .B(n9514), .Z(n9521) );
  XOR U11091 ( .A(n9520), .B(n9521), .Z(n9466) );
  OR U11092 ( .A(n9418), .B(n9417), .Z(n9422) );
  NANDN U11093 ( .A(n9420), .B(n9419), .Z(n9421) );
  AND U11094 ( .A(n9422), .B(n9421), .Z(n9467) );
  XNOR U11095 ( .A(n9466), .B(n9467), .Z(n9468) );
  XOR U11096 ( .A(n9469), .B(n9468), .Z(n9455) );
  XOR U11097 ( .A(n9455), .B(n9454), .Z(n9457) );
  OR U11098 ( .A(n9427), .B(n9426), .Z(n9431) );
  OR U11099 ( .A(n9429), .B(n9428), .Z(n9430) );
  NAND U11100 ( .A(n9431), .B(n9430), .Z(n9463) );
  OR U11101 ( .A(n9437), .B(n9436), .Z(n9441) );
  NANDN U11102 ( .A(n9439), .B(n9438), .Z(n9440) );
  NAND U11103 ( .A(n9441), .B(n9440), .Z(n9472) );
  OR U11104 ( .A(n9443), .B(n9442), .Z(n9447) );
  OR U11105 ( .A(n9445), .B(n9444), .Z(n9446) );
  AND U11106 ( .A(n9447), .B(n9446), .Z(n9473) );
  XNOR U11107 ( .A(n9472), .B(n9473), .Z(n9474) );
  XOR U11108 ( .A(n9475), .B(n9474), .Z(n9460) );
  OR U11109 ( .A(n9449), .B(n9448), .Z(n9453) );
  NANDN U11110 ( .A(n9451), .B(n9450), .Z(n9452) );
  NAND U11111 ( .A(n9453), .B(n9452), .Z(n9461) );
  XNOR U11112 ( .A(n9460), .B(n9461), .Z(n9462) );
  XOR U11113 ( .A(n9463), .B(n9462), .Z(n9456) );
  XOR U11114 ( .A(n9457), .B(n9456), .Z(o[6]) );
  NANDN U11115 ( .A(n9455), .B(n9454), .Z(n9459) );
  OR U11116 ( .A(n9457), .B(n9456), .Z(n9458) );
  AND U11117 ( .A(n9459), .B(n9458), .Z(n9525) );
  OR U11118 ( .A(n9461), .B(n9460), .Z(n9465) );
  OR U11119 ( .A(n9463), .B(n9462), .Z(n9464) );
  NAND U11120 ( .A(n9465), .B(n9464), .Z(n9528) );
  NANDN U11121 ( .A(n9467), .B(n9466), .Z(n9471) );
  NAND U11122 ( .A(n9469), .B(n9468), .Z(n9470) );
  AND U11123 ( .A(n9471), .B(n9470), .Z(n9534) );
  NANDN U11124 ( .A(n9473), .B(n9472), .Z(n9477) );
  NAND U11125 ( .A(n9475), .B(n9474), .Z(n9476) );
  NAND U11126 ( .A(n9477), .B(n9476), .Z(n9532) );
  NANDN U11127 ( .A(n9479), .B(n9478), .Z(n9483) );
  NANDN U11128 ( .A(n9481), .B(n9480), .Z(n9482) );
  NAND U11129 ( .A(n9483), .B(n9482), .Z(n9549) );
  XNOR U11130 ( .A(n9549), .B(n9548), .Z(n9550) );
  OR U11131 ( .A(n9489), .B(n9488), .Z(n9493) );
  NANDN U11132 ( .A(n9491), .B(n9490), .Z(n9492) );
  AND U11133 ( .A(n9493), .B(n9492), .Z(n9542) );
  OR U11134 ( .A(n9495), .B(n9494), .Z(n9499) );
  NAND U11135 ( .A(n9497), .B(n9496), .Z(n9498) );
  AND U11136 ( .A(n9499), .B(n9498), .Z(n9544) );
  NANDN U11137 ( .A(n9501), .B(n9500), .Z(n9505) );
  OR U11138 ( .A(n9503), .B(n9502), .Z(n9504) );
  NAND U11139 ( .A(n9505), .B(n9504), .Z(n9539) );
  OR U11140 ( .A(n9507), .B(n9506), .Z(n9511) );
  OR U11141 ( .A(n9509), .B(n9508), .Z(n9510) );
  AND U11142 ( .A(n9511), .B(n9510), .Z(n9540) );
  XOR U11143 ( .A(n9539), .B(n9540), .Z(n9543) );
  XNOR U11144 ( .A(n9544), .B(n9543), .Z(n9541) );
  XNOR U11145 ( .A(n9550), .B(n9551), .Z(n9537) );
  OR U11146 ( .A(n9513), .B(n9512), .Z(n9517) );
  NAND U11147 ( .A(n9515), .B(n9514), .Z(n9516) );
  NAND U11148 ( .A(n9517), .B(n9516), .Z(n9536) );
  OR U11149 ( .A(n9519), .B(n9518), .Z(n9523) );
  NANDN U11150 ( .A(n9521), .B(n9520), .Z(n9522) );
  AND U11151 ( .A(n9523), .B(n9522), .Z(n9535) );
  XNOR U11152 ( .A(n9536), .B(n9535), .Z(n9538) );
  XOR U11153 ( .A(n9537), .B(n9538), .Z(n9531) );
  XNOR U11154 ( .A(n9532), .B(n9531), .Z(n9533) );
  XOR U11155 ( .A(n9534), .B(n9533), .Z(n9526) );
  XOR U11156 ( .A(n9528), .B(n9526), .Z(n9524) );
  XOR U11157 ( .A(n9525), .B(n9524), .Z(o[7]) );
  NANDN U11158 ( .A(n9525), .B(n9526), .Z(n9530) );
  XNOR U11159 ( .A(n9526), .B(n9525), .Z(n9527) );
  NANDN U11160 ( .A(n9528), .B(n9527), .Z(n9529) );
  NAND U11161 ( .A(n9530), .B(n9529), .Z(n9562) );
  NANDN U11162 ( .A(n9540), .B(n9539), .Z(n9565) );
  NOR U11163 ( .A(n9542), .B(n9541), .Z(n9564) );
  XOR U11164 ( .A(n9565), .B(n9564), .Z(n9547) );
  NOR U11165 ( .A(n9544), .B(n9543), .Z(n9545) );
  NAND U11166 ( .A(n9545), .B(n9565), .Z(n9546) );
  AND U11167 ( .A(n9547), .B(n9546), .Z(n9556) );
  NANDN U11168 ( .A(n9549), .B(n9548), .Z(n9553) );
  NAND U11169 ( .A(n9551), .B(n9550), .Z(n9552) );
  NAND U11170 ( .A(n9553), .B(n9552), .Z(n9555) );
  XNOR U11171 ( .A(n9556), .B(n9555), .Z(n9557) );
  XNOR U11172 ( .A(n9558), .B(n9557), .Z(n9563) );
  XNOR U11173 ( .A(n9561), .B(n9563), .Z(n9554) );
  XNOR U11174 ( .A(n9562), .B(n9554), .Z(o[8]) );
  NANDN U11175 ( .A(n9556), .B(n9555), .Z(n9560) );
  NANDN U11176 ( .A(n9558), .B(n9557), .Z(n9559) );
  NAND U11177 ( .A(n9560), .B(n9559), .Z(n9569) );
  NANDN U11178 ( .A(n9565), .B(n9564), .Z(n9567) );
  XOR U11179 ( .A(n9568), .B(n9567), .Z(n9566) );
  XOR U11180 ( .A(n9569), .B(n9566), .Z(o[9]) );
endmodule

