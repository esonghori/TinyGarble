
module FA_4093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module FA_4094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module COMP_N4096 ( A, B, O );
  input [4095:0] A;
  input [4095:0] B;
  output O;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096;
  wire   [4095:1] C;

  FA_4093 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n4096), .CI(1'b1), 
        .CO(C[1]) );
  FA_8188 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n4095), .CI(C[1]), 
        .CO(C[2]) );
  FA_8187 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n4094), .CI(C[2]), 
        .CO(C[3]) );
  FA_8186 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n4093), .CI(C[3]), 
        .CO(C[4]) );
  FA_8185 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n4092), .CI(C[4]), 
        .CO(C[5]) );
  FA_8184 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n4091), .CI(C[5]), 
        .CO(C[6]) );
  FA_8183 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n4090), .CI(C[6]), 
        .CO(C[7]) );
  FA_8182 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n4089), .CI(C[7]), 
        .CO(C[8]) );
  FA_8181 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n4088), .CI(C[8]), 
        .CO(C[9]) );
  FA_8180 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n4087), .CI(C[9]), 
        .CO(C[10]) );
  FA_8179 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n4086), .CI(C[10]), 
        .CO(C[11]) );
  FA_8178 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n4085), .CI(C[11]), 
        .CO(C[12]) );
  FA_8177 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n4084), .CI(C[12]), 
        .CO(C[13]) );
  FA_8176 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n4083), .CI(C[13]), 
        .CO(C[14]) );
  FA_8175 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n4082), .CI(C[14]), 
        .CO(C[15]) );
  FA_8174 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n4081), .CI(C[15]), 
        .CO(C[16]) );
  FA_8173 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n4080), .CI(C[16]), 
        .CO(C[17]) );
  FA_8172 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n4079), .CI(C[17]), 
        .CO(C[18]) );
  FA_8171 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n4078), .CI(C[18]), 
        .CO(C[19]) );
  FA_8170 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n4077), .CI(C[19]), 
        .CO(C[20]) );
  FA_8169 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n4076), .CI(C[20]), 
        .CO(C[21]) );
  FA_8168 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n4075), .CI(C[21]), 
        .CO(C[22]) );
  FA_8167 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n4074), .CI(C[22]), 
        .CO(C[23]) );
  FA_8166 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n4073), .CI(C[23]), 
        .CO(C[24]) );
  FA_8165 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n4072), .CI(C[24]), 
        .CO(C[25]) );
  FA_8164 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n4071), .CI(C[25]), 
        .CO(C[26]) );
  FA_8163 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n4070), .CI(C[26]), 
        .CO(C[27]) );
  FA_8162 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n4069), .CI(C[27]), 
        .CO(C[28]) );
  FA_8161 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n4068), .CI(C[28]), 
        .CO(C[29]) );
  FA_8160 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n4067), .CI(C[29]), 
        .CO(C[30]) );
  FA_8159 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n4066), .CI(C[30]), 
        .CO(C[31]) );
  FA_8158 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n4065), .CI(C[31]), 
        .CO(C[32]) );
  FA_8157 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n4064), .CI(C[32]), 
        .CO(C[33]) );
  FA_8156 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n4063), .CI(C[33]), 
        .CO(C[34]) );
  FA_8155 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n4062), .CI(C[34]), 
        .CO(C[35]) );
  FA_8154 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n4061), .CI(C[35]), 
        .CO(C[36]) );
  FA_8153 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n4060), .CI(C[36]), 
        .CO(C[37]) );
  FA_8152 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n4059), .CI(C[37]), 
        .CO(C[38]) );
  FA_8151 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n4058), .CI(C[38]), 
        .CO(C[39]) );
  FA_8150 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n4057), .CI(C[39]), 
        .CO(C[40]) );
  FA_8149 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n4056), .CI(C[40]), 
        .CO(C[41]) );
  FA_8148 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n4055), .CI(C[41]), 
        .CO(C[42]) );
  FA_8147 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n4054), .CI(C[42]), 
        .CO(C[43]) );
  FA_8146 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n4053), .CI(C[43]), 
        .CO(C[44]) );
  FA_8145 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n4052), .CI(C[44]), 
        .CO(C[45]) );
  FA_8144 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n4051), .CI(C[45]), 
        .CO(C[46]) );
  FA_8143 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n4050), .CI(C[46]), 
        .CO(C[47]) );
  FA_8142 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n4049), .CI(C[47]), 
        .CO(C[48]) );
  FA_8141 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n4048), .CI(C[48]), 
        .CO(C[49]) );
  FA_8140 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n4047), .CI(C[49]), 
        .CO(C[50]) );
  FA_8139 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n4046), .CI(C[50]), 
        .CO(C[51]) );
  FA_8138 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n4045), .CI(C[51]), 
        .CO(C[52]) );
  FA_8137 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n4044), .CI(C[52]), 
        .CO(C[53]) );
  FA_8136 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n4043), .CI(C[53]), 
        .CO(C[54]) );
  FA_8135 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n4042), .CI(C[54]), 
        .CO(C[55]) );
  FA_8134 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n4041), .CI(C[55]), 
        .CO(C[56]) );
  FA_8133 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n4040), .CI(C[56]), 
        .CO(C[57]) );
  FA_8132 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n4039), .CI(C[57]), 
        .CO(C[58]) );
  FA_8131 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n4038), .CI(C[58]), 
        .CO(C[59]) );
  FA_8130 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n4037), .CI(C[59]), 
        .CO(C[60]) );
  FA_8129 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n4036), .CI(C[60]), 
        .CO(C[61]) );
  FA_8128 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n4035), .CI(C[61]), 
        .CO(C[62]) );
  FA_8127 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n4034), .CI(C[62]), 
        .CO(C[63]) );
  FA_8126 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n4033), .CI(C[63]), 
        .CO(C[64]) );
  FA_8125 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n4032), .CI(C[64]), 
        .CO(C[65]) );
  FA_8124 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n4031), .CI(C[65]), 
        .CO(C[66]) );
  FA_8123 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n4030), .CI(C[66]), 
        .CO(C[67]) );
  FA_8122 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n4029), .CI(C[67]), 
        .CO(C[68]) );
  FA_8121 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n4028), .CI(C[68]), 
        .CO(C[69]) );
  FA_8120 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n4027), .CI(C[69]), 
        .CO(C[70]) );
  FA_8119 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n4026), .CI(C[70]), 
        .CO(C[71]) );
  FA_8118 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n4025), .CI(C[71]), 
        .CO(C[72]) );
  FA_8117 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n4024), .CI(C[72]), 
        .CO(C[73]) );
  FA_8116 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n4023), .CI(C[73]), 
        .CO(C[74]) );
  FA_8115 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n4022), .CI(C[74]), 
        .CO(C[75]) );
  FA_8114 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n4021), .CI(C[75]), 
        .CO(C[76]) );
  FA_8113 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n4020), .CI(C[76]), 
        .CO(C[77]) );
  FA_8112 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n4019), .CI(C[77]), 
        .CO(C[78]) );
  FA_8111 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n4018), .CI(C[78]), 
        .CO(C[79]) );
  FA_8110 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n4017), .CI(C[79]), 
        .CO(C[80]) );
  FA_8109 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n4016), .CI(C[80]), 
        .CO(C[81]) );
  FA_8108 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n4015), .CI(C[81]), 
        .CO(C[82]) );
  FA_8107 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n4014), .CI(C[82]), 
        .CO(C[83]) );
  FA_8106 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n4013), .CI(C[83]), 
        .CO(C[84]) );
  FA_8105 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n4012), .CI(C[84]), 
        .CO(C[85]) );
  FA_8104 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n4011), .CI(C[85]), 
        .CO(C[86]) );
  FA_8103 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n4010), .CI(C[86]), 
        .CO(C[87]) );
  FA_8102 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n4009), .CI(C[87]), 
        .CO(C[88]) );
  FA_8101 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n4008), .CI(C[88]), 
        .CO(C[89]) );
  FA_8100 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n4007), .CI(C[89]), 
        .CO(C[90]) );
  FA_8099 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n4006), .CI(C[90]), 
        .CO(C[91]) );
  FA_8098 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n4005), .CI(C[91]), 
        .CO(C[92]) );
  FA_8097 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n4004), .CI(C[92]), 
        .CO(C[93]) );
  FA_8096 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n4003), .CI(C[93]), 
        .CO(C[94]) );
  FA_8095 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n4002), .CI(C[94]), 
        .CO(C[95]) );
  FA_8094 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n4001), .CI(C[95]), 
        .CO(C[96]) );
  FA_8093 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n4000), .CI(C[96]), 
        .CO(C[97]) );
  FA_8092 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n3999), .CI(C[97]), 
        .CO(C[98]) );
  FA_8091 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n3998), .CI(C[98]), 
        .CO(C[99]) );
  FA_8090 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n3997), .CI(C[99]), 
        .CO(C[100]) );
  FA_8089 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n3996), .CI(
        C[100]), .CO(C[101]) );
  FA_8088 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n3995), .CI(
        C[101]), .CO(C[102]) );
  FA_8087 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n3994), .CI(
        C[102]), .CO(C[103]) );
  FA_8086 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n3993), .CI(
        C[103]), .CO(C[104]) );
  FA_8085 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n3992), .CI(
        C[104]), .CO(C[105]) );
  FA_8084 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n3991), .CI(
        C[105]), .CO(C[106]) );
  FA_8083 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n3990), .CI(
        C[106]), .CO(C[107]) );
  FA_8082 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n3989), .CI(
        C[107]), .CO(C[108]) );
  FA_8081 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n3988), .CI(
        C[108]), .CO(C[109]) );
  FA_8080 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n3987), .CI(
        C[109]), .CO(C[110]) );
  FA_8079 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n3986), .CI(
        C[110]), .CO(C[111]) );
  FA_8078 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n3985), .CI(
        C[111]), .CO(C[112]) );
  FA_8077 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n3984), .CI(
        C[112]), .CO(C[113]) );
  FA_8076 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n3983), .CI(
        C[113]), .CO(C[114]) );
  FA_8075 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n3982), .CI(
        C[114]), .CO(C[115]) );
  FA_8074 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n3981), .CI(
        C[115]), .CO(C[116]) );
  FA_8073 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n3980), .CI(
        C[116]), .CO(C[117]) );
  FA_8072 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n3979), .CI(
        C[117]), .CO(C[118]) );
  FA_8071 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n3978), .CI(
        C[118]), .CO(C[119]) );
  FA_8070 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n3977), .CI(
        C[119]), .CO(C[120]) );
  FA_8069 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n3976), .CI(
        C[120]), .CO(C[121]) );
  FA_8068 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n3975), .CI(
        C[121]), .CO(C[122]) );
  FA_8067 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n3974), .CI(
        C[122]), .CO(C[123]) );
  FA_8066 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n3973), .CI(
        C[123]), .CO(C[124]) );
  FA_8065 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n3972), .CI(
        C[124]), .CO(C[125]) );
  FA_8064 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n3971), .CI(
        C[125]), .CO(C[126]) );
  FA_8063 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n3970), .CI(
        C[126]), .CO(C[127]) );
  FA_8062 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n3969), .CI(
        C[127]), .CO(C[128]) );
  FA_8061 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n3968), .CI(
        C[128]), .CO(C[129]) );
  FA_8060 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n3967), .CI(
        C[129]), .CO(C[130]) );
  FA_8059 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n3966), .CI(
        C[130]), .CO(C[131]) );
  FA_8058 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n3965), .CI(
        C[131]), .CO(C[132]) );
  FA_8057 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n3964), .CI(
        C[132]), .CO(C[133]) );
  FA_8056 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n3963), .CI(
        C[133]), .CO(C[134]) );
  FA_8055 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n3962), .CI(
        C[134]), .CO(C[135]) );
  FA_8054 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n3961), .CI(
        C[135]), .CO(C[136]) );
  FA_8053 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n3960), .CI(
        C[136]), .CO(C[137]) );
  FA_8052 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n3959), .CI(
        C[137]), .CO(C[138]) );
  FA_8051 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n3958), .CI(
        C[138]), .CO(C[139]) );
  FA_8050 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n3957), .CI(
        C[139]), .CO(C[140]) );
  FA_8049 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n3956), .CI(
        C[140]), .CO(C[141]) );
  FA_8048 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n3955), .CI(
        C[141]), .CO(C[142]) );
  FA_8047 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n3954), .CI(
        C[142]), .CO(C[143]) );
  FA_8046 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n3953), .CI(
        C[143]), .CO(C[144]) );
  FA_8045 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n3952), .CI(
        C[144]), .CO(C[145]) );
  FA_8044 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n3951), .CI(
        C[145]), .CO(C[146]) );
  FA_8043 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n3950), .CI(
        C[146]), .CO(C[147]) );
  FA_8042 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n3949), .CI(
        C[147]), .CO(C[148]) );
  FA_8041 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n3948), .CI(
        C[148]), .CO(C[149]) );
  FA_8040 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n3947), .CI(
        C[149]), .CO(C[150]) );
  FA_8039 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n3946), .CI(
        C[150]), .CO(C[151]) );
  FA_8038 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n3945), .CI(
        C[151]), .CO(C[152]) );
  FA_8037 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n3944), .CI(
        C[152]), .CO(C[153]) );
  FA_8036 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n3943), .CI(
        C[153]), .CO(C[154]) );
  FA_8035 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n3942), .CI(
        C[154]), .CO(C[155]) );
  FA_8034 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n3941), .CI(
        C[155]), .CO(C[156]) );
  FA_8033 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n3940), .CI(
        C[156]), .CO(C[157]) );
  FA_8032 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n3939), .CI(
        C[157]), .CO(C[158]) );
  FA_8031 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n3938), .CI(
        C[158]), .CO(C[159]) );
  FA_8030 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n3937), .CI(
        C[159]), .CO(C[160]) );
  FA_8029 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n3936), .CI(
        C[160]), .CO(C[161]) );
  FA_8028 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n3935), .CI(
        C[161]), .CO(C[162]) );
  FA_8027 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n3934), .CI(
        C[162]), .CO(C[163]) );
  FA_8026 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n3933), .CI(
        C[163]), .CO(C[164]) );
  FA_8025 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n3932), .CI(
        C[164]), .CO(C[165]) );
  FA_8024 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n3931), .CI(
        C[165]), .CO(C[166]) );
  FA_8023 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n3930), .CI(
        C[166]), .CO(C[167]) );
  FA_8022 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n3929), .CI(
        C[167]), .CO(C[168]) );
  FA_8021 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n3928), .CI(
        C[168]), .CO(C[169]) );
  FA_8020 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n3927), .CI(
        C[169]), .CO(C[170]) );
  FA_8019 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n3926), .CI(
        C[170]), .CO(C[171]) );
  FA_8018 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n3925), .CI(
        C[171]), .CO(C[172]) );
  FA_8017 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n3924), .CI(
        C[172]), .CO(C[173]) );
  FA_8016 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n3923), .CI(
        C[173]), .CO(C[174]) );
  FA_8015 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n3922), .CI(
        C[174]), .CO(C[175]) );
  FA_8014 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n3921), .CI(
        C[175]), .CO(C[176]) );
  FA_8013 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n3920), .CI(
        C[176]), .CO(C[177]) );
  FA_8012 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n3919), .CI(
        C[177]), .CO(C[178]) );
  FA_8011 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n3918), .CI(
        C[178]), .CO(C[179]) );
  FA_8010 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n3917), .CI(
        C[179]), .CO(C[180]) );
  FA_8009 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n3916), .CI(
        C[180]), .CO(C[181]) );
  FA_8008 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n3915), .CI(
        C[181]), .CO(C[182]) );
  FA_8007 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n3914), .CI(
        C[182]), .CO(C[183]) );
  FA_8006 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n3913), .CI(
        C[183]), .CO(C[184]) );
  FA_8005 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n3912), .CI(
        C[184]), .CO(C[185]) );
  FA_8004 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n3911), .CI(
        C[185]), .CO(C[186]) );
  FA_8003 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n3910), .CI(
        C[186]), .CO(C[187]) );
  FA_8002 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n3909), .CI(
        C[187]), .CO(C[188]) );
  FA_8001 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n3908), .CI(
        C[188]), .CO(C[189]) );
  FA_8000 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n3907), .CI(
        C[189]), .CO(C[190]) );
  FA_7999 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n3906), .CI(
        C[190]), .CO(C[191]) );
  FA_7998 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n3905), .CI(
        C[191]), .CO(C[192]) );
  FA_7997 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n3904), .CI(
        C[192]), .CO(C[193]) );
  FA_7996 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n3903), .CI(
        C[193]), .CO(C[194]) );
  FA_7995 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n3902), .CI(
        C[194]), .CO(C[195]) );
  FA_7994 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n3901), .CI(
        C[195]), .CO(C[196]) );
  FA_7993 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n3900), .CI(
        C[196]), .CO(C[197]) );
  FA_7992 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n3899), .CI(
        C[197]), .CO(C[198]) );
  FA_7991 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n3898), .CI(
        C[198]), .CO(C[199]) );
  FA_7990 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n3897), .CI(
        C[199]), .CO(C[200]) );
  FA_7989 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n3896), .CI(
        C[200]), .CO(C[201]) );
  FA_7988 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n3895), .CI(
        C[201]), .CO(C[202]) );
  FA_7987 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n3894), .CI(
        C[202]), .CO(C[203]) );
  FA_7986 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n3893), .CI(
        C[203]), .CO(C[204]) );
  FA_7985 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n3892), .CI(
        C[204]), .CO(C[205]) );
  FA_7984 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n3891), .CI(
        C[205]), .CO(C[206]) );
  FA_7983 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n3890), .CI(
        C[206]), .CO(C[207]) );
  FA_7982 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n3889), .CI(
        C[207]), .CO(C[208]) );
  FA_7981 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n3888), .CI(
        C[208]), .CO(C[209]) );
  FA_7980 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n3887), .CI(
        C[209]), .CO(C[210]) );
  FA_7979 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n3886), .CI(
        C[210]), .CO(C[211]) );
  FA_7978 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n3885), .CI(
        C[211]), .CO(C[212]) );
  FA_7977 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n3884), .CI(
        C[212]), .CO(C[213]) );
  FA_7976 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n3883), .CI(
        C[213]), .CO(C[214]) );
  FA_7975 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n3882), .CI(
        C[214]), .CO(C[215]) );
  FA_7974 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n3881), .CI(
        C[215]), .CO(C[216]) );
  FA_7973 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n3880), .CI(
        C[216]), .CO(C[217]) );
  FA_7972 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n3879), .CI(
        C[217]), .CO(C[218]) );
  FA_7971 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n3878), .CI(
        C[218]), .CO(C[219]) );
  FA_7970 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n3877), .CI(
        C[219]), .CO(C[220]) );
  FA_7969 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n3876), .CI(
        C[220]), .CO(C[221]) );
  FA_7968 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n3875), .CI(
        C[221]), .CO(C[222]) );
  FA_7967 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n3874), .CI(
        C[222]), .CO(C[223]) );
  FA_7966 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n3873), .CI(
        C[223]), .CO(C[224]) );
  FA_7965 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n3872), .CI(
        C[224]), .CO(C[225]) );
  FA_7964 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n3871), .CI(
        C[225]), .CO(C[226]) );
  FA_7963 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n3870), .CI(
        C[226]), .CO(C[227]) );
  FA_7962 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n3869), .CI(
        C[227]), .CO(C[228]) );
  FA_7961 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n3868), .CI(
        C[228]), .CO(C[229]) );
  FA_7960 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n3867), .CI(
        C[229]), .CO(C[230]) );
  FA_7959 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n3866), .CI(
        C[230]), .CO(C[231]) );
  FA_7958 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n3865), .CI(
        C[231]), .CO(C[232]) );
  FA_7957 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n3864), .CI(
        C[232]), .CO(C[233]) );
  FA_7956 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n3863), .CI(
        C[233]), .CO(C[234]) );
  FA_7955 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n3862), .CI(
        C[234]), .CO(C[235]) );
  FA_7954 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n3861), .CI(
        C[235]), .CO(C[236]) );
  FA_7953 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n3860), .CI(
        C[236]), .CO(C[237]) );
  FA_7952 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n3859), .CI(
        C[237]), .CO(C[238]) );
  FA_7951 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n3858), .CI(
        C[238]), .CO(C[239]) );
  FA_7950 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n3857), .CI(
        C[239]), .CO(C[240]) );
  FA_7949 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n3856), .CI(
        C[240]), .CO(C[241]) );
  FA_7948 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n3855), .CI(
        C[241]), .CO(C[242]) );
  FA_7947 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n3854), .CI(
        C[242]), .CO(C[243]) );
  FA_7946 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n3853), .CI(
        C[243]), .CO(C[244]) );
  FA_7945 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n3852), .CI(
        C[244]), .CO(C[245]) );
  FA_7944 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n3851), .CI(
        C[245]), .CO(C[246]) );
  FA_7943 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n3850), .CI(
        C[246]), .CO(C[247]) );
  FA_7942 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n3849), .CI(
        C[247]), .CO(C[248]) );
  FA_7941 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n3848), .CI(
        C[248]), .CO(C[249]) );
  FA_7940 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n3847), .CI(
        C[249]), .CO(C[250]) );
  FA_7939 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n3846), .CI(
        C[250]), .CO(C[251]) );
  FA_7938 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n3845), .CI(
        C[251]), .CO(C[252]) );
  FA_7937 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n3844), .CI(
        C[252]), .CO(C[253]) );
  FA_7936 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n3843), .CI(
        C[253]), .CO(C[254]) );
  FA_7935 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n3842), .CI(
        C[254]), .CO(C[255]) );
  FA_7934 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n3841), .CI(
        C[255]), .CO(C[256]) );
  FA_7933 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n3840), .CI(
        C[256]), .CO(C[257]) );
  FA_7932 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n3839), .CI(
        C[257]), .CO(C[258]) );
  FA_7931 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n3838), .CI(
        C[258]), .CO(C[259]) );
  FA_7930 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n3837), .CI(
        C[259]), .CO(C[260]) );
  FA_7929 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n3836), .CI(
        C[260]), .CO(C[261]) );
  FA_7928 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n3835), .CI(
        C[261]), .CO(C[262]) );
  FA_7927 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n3834), .CI(
        C[262]), .CO(C[263]) );
  FA_7926 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n3833), .CI(
        C[263]), .CO(C[264]) );
  FA_7925 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n3832), .CI(
        C[264]), .CO(C[265]) );
  FA_7924 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n3831), .CI(
        C[265]), .CO(C[266]) );
  FA_7923 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n3830), .CI(
        C[266]), .CO(C[267]) );
  FA_7922 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n3829), .CI(
        C[267]), .CO(C[268]) );
  FA_7921 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n3828), .CI(
        C[268]), .CO(C[269]) );
  FA_7920 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n3827), .CI(
        C[269]), .CO(C[270]) );
  FA_7919 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n3826), .CI(
        C[270]), .CO(C[271]) );
  FA_7918 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n3825), .CI(
        C[271]), .CO(C[272]) );
  FA_7917 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n3824), .CI(
        C[272]), .CO(C[273]) );
  FA_7916 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n3823), .CI(
        C[273]), .CO(C[274]) );
  FA_7915 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n3822), .CI(
        C[274]), .CO(C[275]) );
  FA_7914 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n3821), .CI(
        C[275]), .CO(C[276]) );
  FA_7913 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n3820), .CI(
        C[276]), .CO(C[277]) );
  FA_7912 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n3819), .CI(
        C[277]), .CO(C[278]) );
  FA_7911 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n3818), .CI(
        C[278]), .CO(C[279]) );
  FA_7910 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n3817), .CI(
        C[279]), .CO(C[280]) );
  FA_7909 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n3816), .CI(
        C[280]), .CO(C[281]) );
  FA_7908 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n3815), .CI(
        C[281]), .CO(C[282]) );
  FA_7907 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n3814), .CI(
        C[282]), .CO(C[283]) );
  FA_7906 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n3813), .CI(
        C[283]), .CO(C[284]) );
  FA_7905 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n3812), .CI(
        C[284]), .CO(C[285]) );
  FA_7904 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n3811), .CI(
        C[285]), .CO(C[286]) );
  FA_7903 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n3810), .CI(
        C[286]), .CO(C[287]) );
  FA_7902 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n3809), .CI(
        C[287]), .CO(C[288]) );
  FA_7901 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n3808), .CI(
        C[288]), .CO(C[289]) );
  FA_7900 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n3807), .CI(
        C[289]), .CO(C[290]) );
  FA_7899 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n3806), .CI(
        C[290]), .CO(C[291]) );
  FA_7898 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n3805), .CI(
        C[291]), .CO(C[292]) );
  FA_7897 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n3804), .CI(
        C[292]), .CO(C[293]) );
  FA_7896 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n3803), .CI(
        C[293]), .CO(C[294]) );
  FA_7895 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n3802), .CI(
        C[294]), .CO(C[295]) );
  FA_7894 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n3801), .CI(
        C[295]), .CO(C[296]) );
  FA_7893 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n3800), .CI(
        C[296]), .CO(C[297]) );
  FA_7892 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n3799), .CI(
        C[297]), .CO(C[298]) );
  FA_7891 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n3798), .CI(
        C[298]), .CO(C[299]) );
  FA_7890 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n3797), .CI(
        C[299]), .CO(C[300]) );
  FA_7889 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n3796), .CI(
        C[300]), .CO(C[301]) );
  FA_7888 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n3795), .CI(
        C[301]), .CO(C[302]) );
  FA_7887 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n3794), .CI(
        C[302]), .CO(C[303]) );
  FA_7886 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n3793), .CI(
        C[303]), .CO(C[304]) );
  FA_7885 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n3792), .CI(
        C[304]), .CO(C[305]) );
  FA_7884 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n3791), .CI(
        C[305]), .CO(C[306]) );
  FA_7883 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n3790), .CI(
        C[306]), .CO(C[307]) );
  FA_7882 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n3789), .CI(
        C[307]), .CO(C[308]) );
  FA_7881 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n3788), .CI(
        C[308]), .CO(C[309]) );
  FA_7880 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n3787), .CI(
        C[309]), .CO(C[310]) );
  FA_7879 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n3786), .CI(
        C[310]), .CO(C[311]) );
  FA_7878 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n3785), .CI(
        C[311]), .CO(C[312]) );
  FA_7877 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n3784), .CI(
        C[312]), .CO(C[313]) );
  FA_7876 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n3783), .CI(
        C[313]), .CO(C[314]) );
  FA_7875 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n3782), .CI(
        C[314]), .CO(C[315]) );
  FA_7874 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n3781), .CI(
        C[315]), .CO(C[316]) );
  FA_7873 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n3780), .CI(
        C[316]), .CO(C[317]) );
  FA_7872 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n3779), .CI(
        C[317]), .CO(C[318]) );
  FA_7871 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n3778), .CI(
        C[318]), .CO(C[319]) );
  FA_7870 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n3777), .CI(
        C[319]), .CO(C[320]) );
  FA_7869 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n3776), .CI(
        C[320]), .CO(C[321]) );
  FA_7868 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n3775), .CI(
        C[321]), .CO(C[322]) );
  FA_7867 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n3774), .CI(
        C[322]), .CO(C[323]) );
  FA_7866 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n3773), .CI(
        C[323]), .CO(C[324]) );
  FA_7865 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n3772), .CI(
        C[324]), .CO(C[325]) );
  FA_7864 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n3771), .CI(
        C[325]), .CO(C[326]) );
  FA_7863 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n3770), .CI(
        C[326]), .CO(C[327]) );
  FA_7862 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n3769), .CI(
        C[327]), .CO(C[328]) );
  FA_7861 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n3768), .CI(
        C[328]), .CO(C[329]) );
  FA_7860 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n3767), .CI(
        C[329]), .CO(C[330]) );
  FA_7859 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n3766), .CI(
        C[330]), .CO(C[331]) );
  FA_7858 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n3765), .CI(
        C[331]), .CO(C[332]) );
  FA_7857 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n3764), .CI(
        C[332]), .CO(C[333]) );
  FA_7856 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n3763), .CI(
        C[333]), .CO(C[334]) );
  FA_7855 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n3762), .CI(
        C[334]), .CO(C[335]) );
  FA_7854 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n3761), .CI(
        C[335]), .CO(C[336]) );
  FA_7853 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n3760), .CI(
        C[336]), .CO(C[337]) );
  FA_7852 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n3759), .CI(
        C[337]), .CO(C[338]) );
  FA_7851 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n3758), .CI(
        C[338]), .CO(C[339]) );
  FA_7850 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n3757), .CI(
        C[339]), .CO(C[340]) );
  FA_7849 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n3756), .CI(
        C[340]), .CO(C[341]) );
  FA_7848 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n3755), .CI(
        C[341]), .CO(C[342]) );
  FA_7847 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n3754), .CI(
        C[342]), .CO(C[343]) );
  FA_7846 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n3753), .CI(
        C[343]), .CO(C[344]) );
  FA_7845 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n3752), .CI(
        C[344]), .CO(C[345]) );
  FA_7844 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n3751), .CI(
        C[345]), .CO(C[346]) );
  FA_7843 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n3750), .CI(
        C[346]), .CO(C[347]) );
  FA_7842 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n3749), .CI(
        C[347]), .CO(C[348]) );
  FA_7841 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n3748), .CI(
        C[348]), .CO(C[349]) );
  FA_7840 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n3747), .CI(
        C[349]), .CO(C[350]) );
  FA_7839 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n3746), .CI(
        C[350]), .CO(C[351]) );
  FA_7838 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n3745), .CI(
        C[351]), .CO(C[352]) );
  FA_7837 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n3744), .CI(
        C[352]), .CO(C[353]) );
  FA_7836 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n3743), .CI(
        C[353]), .CO(C[354]) );
  FA_7835 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n3742), .CI(
        C[354]), .CO(C[355]) );
  FA_7834 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n3741), .CI(
        C[355]), .CO(C[356]) );
  FA_7833 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n3740), .CI(
        C[356]), .CO(C[357]) );
  FA_7832 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n3739), .CI(
        C[357]), .CO(C[358]) );
  FA_7831 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n3738), .CI(
        C[358]), .CO(C[359]) );
  FA_7830 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n3737), .CI(
        C[359]), .CO(C[360]) );
  FA_7829 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n3736), .CI(
        C[360]), .CO(C[361]) );
  FA_7828 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n3735), .CI(
        C[361]), .CO(C[362]) );
  FA_7827 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n3734), .CI(
        C[362]), .CO(C[363]) );
  FA_7826 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n3733), .CI(
        C[363]), .CO(C[364]) );
  FA_7825 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n3732), .CI(
        C[364]), .CO(C[365]) );
  FA_7824 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n3731), .CI(
        C[365]), .CO(C[366]) );
  FA_7823 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n3730), .CI(
        C[366]), .CO(C[367]) );
  FA_7822 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n3729), .CI(
        C[367]), .CO(C[368]) );
  FA_7821 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n3728), .CI(
        C[368]), .CO(C[369]) );
  FA_7820 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n3727), .CI(
        C[369]), .CO(C[370]) );
  FA_7819 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n3726), .CI(
        C[370]), .CO(C[371]) );
  FA_7818 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n3725), .CI(
        C[371]), .CO(C[372]) );
  FA_7817 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n3724), .CI(
        C[372]), .CO(C[373]) );
  FA_7816 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n3723), .CI(
        C[373]), .CO(C[374]) );
  FA_7815 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n3722), .CI(
        C[374]), .CO(C[375]) );
  FA_7814 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n3721), .CI(
        C[375]), .CO(C[376]) );
  FA_7813 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n3720), .CI(
        C[376]), .CO(C[377]) );
  FA_7812 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n3719), .CI(
        C[377]), .CO(C[378]) );
  FA_7811 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n3718), .CI(
        C[378]), .CO(C[379]) );
  FA_7810 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n3717), .CI(
        C[379]), .CO(C[380]) );
  FA_7809 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n3716), .CI(
        C[380]), .CO(C[381]) );
  FA_7808 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n3715), .CI(
        C[381]), .CO(C[382]) );
  FA_7807 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n3714), .CI(
        C[382]), .CO(C[383]) );
  FA_7806 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n3713), .CI(
        C[383]), .CO(C[384]) );
  FA_7805 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n3712), .CI(
        C[384]), .CO(C[385]) );
  FA_7804 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n3711), .CI(
        C[385]), .CO(C[386]) );
  FA_7803 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n3710), .CI(
        C[386]), .CO(C[387]) );
  FA_7802 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n3709), .CI(
        C[387]), .CO(C[388]) );
  FA_7801 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n3708), .CI(
        C[388]), .CO(C[389]) );
  FA_7800 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n3707), .CI(
        C[389]), .CO(C[390]) );
  FA_7799 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n3706), .CI(
        C[390]), .CO(C[391]) );
  FA_7798 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n3705), .CI(
        C[391]), .CO(C[392]) );
  FA_7797 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n3704), .CI(
        C[392]), .CO(C[393]) );
  FA_7796 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n3703), .CI(
        C[393]), .CO(C[394]) );
  FA_7795 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n3702), .CI(
        C[394]), .CO(C[395]) );
  FA_7794 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n3701), .CI(
        C[395]), .CO(C[396]) );
  FA_7793 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n3700), .CI(
        C[396]), .CO(C[397]) );
  FA_7792 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n3699), .CI(
        C[397]), .CO(C[398]) );
  FA_7791 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n3698), .CI(
        C[398]), .CO(C[399]) );
  FA_7790 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n3697), .CI(
        C[399]), .CO(C[400]) );
  FA_7789 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n3696), .CI(
        C[400]), .CO(C[401]) );
  FA_7788 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n3695), .CI(
        C[401]), .CO(C[402]) );
  FA_7787 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n3694), .CI(
        C[402]), .CO(C[403]) );
  FA_7786 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n3693), .CI(
        C[403]), .CO(C[404]) );
  FA_7785 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n3692), .CI(
        C[404]), .CO(C[405]) );
  FA_7784 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n3691), .CI(
        C[405]), .CO(C[406]) );
  FA_7783 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n3690), .CI(
        C[406]), .CO(C[407]) );
  FA_7782 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n3689), .CI(
        C[407]), .CO(C[408]) );
  FA_7781 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n3688), .CI(
        C[408]), .CO(C[409]) );
  FA_7780 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n3687), .CI(
        C[409]), .CO(C[410]) );
  FA_7779 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n3686), .CI(
        C[410]), .CO(C[411]) );
  FA_7778 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n3685), .CI(
        C[411]), .CO(C[412]) );
  FA_7777 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n3684), .CI(
        C[412]), .CO(C[413]) );
  FA_7776 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n3683), .CI(
        C[413]), .CO(C[414]) );
  FA_7775 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n3682), .CI(
        C[414]), .CO(C[415]) );
  FA_7774 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n3681), .CI(
        C[415]), .CO(C[416]) );
  FA_7773 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n3680), .CI(
        C[416]), .CO(C[417]) );
  FA_7772 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n3679), .CI(
        C[417]), .CO(C[418]) );
  FA_7771 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n3678), .CI(
        C[418]), .CO(C[419]) );
  FA_7770 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n3677), .CI(
        C[419]), .CO(C[420]) );
  FA_7769 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n3676), .CI(
        C[420]), .CO(C[421]) );
  FA_7768 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n3675), .CI(
        C[421]), .CO(C[422]) );
  FA_7767 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n3674), .CI(
        C[422]), .CO(C[423]) );
  FA_7766 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n3673), .CI(
        C[423]), .CO(C[424]) );
  FA_7765 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n3672), .CI(
        C[424]), .CO(C[425]) );
  FA_7764 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n3671), .CI(
        C[425]), .CO(C[426]) );
  FA_7763 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n3670), .CI(
        C[426]), .CO(C[427]) );
  FA_7762 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n3669), .CI(
        C[427]), .CO(C[428]) );
  FA_7761 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n3668), .CI(
        C[428]), .CO(C[429]) );
  FA_7760 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n3667), .CI(
        C[429]), .CO(C[430]) );
  FA_7759 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n3666), .CI(
        C[430]), .CO(C[431]) );
  FA_7758 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n3665), .CI(
        C[431]), .CO(C[432]) );
  FA_7757 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n3664), .CI(
        C[432]), .CO(C[433]) );
  FA_7756 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n3663), .CI(
        C[433]), .CO(C[434]) );
  FA_7755 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n3662), .CI(
        C[434]), .CO(C[435]) );
  FA_7754 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n3661), .CI(
        C[435]), .CO(C[436]) );
  FA_7753 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n3660), .CI(
        C[436]), .CO(C[437]) );
  FA_7752 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n3659), .CI(
        C[437]), .CO(C[438]) );
  FA_7751 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n3658), .CI(
        C[438]), .CO(C[439]) );
  FA_7750 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n3657), .CI(
        C[439]), .CO(C[440]) );
  FA_7749 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n3656), .CI(
        C[440]), .CO(C[441]) );
  FA_7748 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n3655), .CI(
        C[441]), .CO(C[442]) );
  FA_7747 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n3654), .CI(
        C[442]), .CO(C[443]) );
  FA_7746 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n3653), .CI(
        C[443]), .CO(C[444]) );
  FA_7745 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n3652), .CI(
        C[444]), .CO(C[445]) );
  FA_7744 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n3651), .CI(
        C[445]), .CO(C[446]) );
  FA_7743 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n3650), .CI(
        C[446]), .CO(C[447]) );
  FA_7742 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n3649), .CI(
        C[447]), .CO(C[448]) );
  FA_7741 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n3648), .CI(
        C[448]), .CO(C[449]) );
  FA_7740 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n3647), .CI(
        C[449]), .CO(C[450]) );
  FA_7739 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n3646), .CI(
        C[450]), .CO(C[451]) );
  FA_7738 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n3645), .CI(
        C[451]), .CO(C[452]) );
  FA_7737 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n3644), .CI(
        C[452]), .CO(C[453]) );
  FA_7736 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n3643), .CI(
        C[453]), .CO(C[454]) );
  FA_7735 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n3642), .CI(
        C[454]), .CO(C[455]) );
  FA_7734 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n3641), .CI(
        C[455]), .CO(C[456]) );
  FA_7733 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n3640), .CI(
        C[456]), .CO(C[457]) );
  FA_7732 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n3639), .CI(
        C[457]), .CO(C[458]) );
  FA_7731 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n3638), .CI(
        C[458]), .CO(C[459]) );
  FA_7730 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n3637), .CI(
        C[459]), .CO(C[460]) );
  FA_7729 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n3636), .CI(
        C[460]), .CO(C[461]) );
  FA_7728 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n3635), .CI(
        C[461]), .CO(C[462]) );
  FA_7727 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n3634), .CI(
        C[462]), .CO(C[463]) );
  FA_7726 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n3633), .CI(
        C[463]), .CO(C[464]) );
  FA_7725 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n3632), .CI(
        C[464]), .CO(C[465]) );
  FA_7724 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n3631), .CI(
        C[465]), .CO(C[466]) );
  FA_7723 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n3630), .CI(
        C[466]), .CO(C[467]) );
  FA_7722 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n3629), .CI(
        C[467]), .CO(C[468]) );
  FA_7721 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n3628), .CI(
        C[468]), .CO(C[469]) );
  FA_7720 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n3627), .CI(
        C[469]), .CO(C[470]) );
  FA_7719 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n3626), .CI(
        C[470]), .CO(C[471]) );
  FA_7718 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n3625), .CI(
        C[471]), .CO(C[472]) );
  FA_7717 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n3624), .CI(
        C[472]), .CO(C[473]) );
  FA_7716 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n3623), .CI(
        C[473]), .CO(C[474]) );
  FA_7715 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n3622), .CI(
        C[474]), .CO(C[475]) );
  FA_7714 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n3621), .CI(
        C[475]), .CO(C[476]) );
  FA_7713 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n3620), .CI(
        C[476]), .CO(C[477]) );
  FA_7712 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n3619), .CI(
        C[477]), .CO(C[478]) );
  FA_7711 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n3618), .CI(
        C[478]), .CO(C[479]) );
  FA_7710 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n3617), .CI(
        C[479]), .CO(C[480]) );
  FA_7709 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n3616), .CI(
        C[480]), .CO(C[481]) );
  FA_7708 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n3615), .CI(
        C[481]), .CO(C[482]) );
  FA_7707 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n3614), .CI(
        C[482]), .CO(C[483]) );
  FA_7706 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n3613), .CI(
        C[483]), .CO(C[484]) );
  FA_7705 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n3612), .CI(
        C[484]), .CO(C[485]) );
  FA_7704 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n3611), .CI(
        C[485]), .CO(C[486]) );
  FA_7703 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n3610), .CI(
        C[486]), .CO(C[487]) );
  FA_7702 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n3609), .CI(
        C[487]), .CO(C[488]) );
  FA_7701 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n3608), .CI(
        C[488]), .CO(C[489]) );
  FA_7700 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n3607), .CI(
        C[489]), .CO(C[490]) );
  FA_7699 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n3606), .CI(
        C[490]), .CO(C[491]) );
  FA_7698 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n3605), .CI(
        C[491]), .CO(C[492]) );
  FA_7697 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n3604), .CI(
        C[492]), .CO(C[493]) );
  FA_7696 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n3603), .CI(
        C[493]), .CO(C[494]) );
  FA_7695 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n3602), .CI(
        C[494]), .CO(C[495]) );
  FA_7694 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n3601), .CI(
        C[495]), .CO(C[496]) );
  FA_7693 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n3600), .CI(
        C[496]), .CO(C[497]) );
  FA_7692 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n3599), .CI(
        C[497]), .CO(C[498]) );
  FA_7691 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n3598), .CI(
        C[498]), .CO(C[499]) );
  FA_7690 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n3597), .CI(
        C[499]), .CO(C[500]) );
  FA_7689 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n3596), .CI(
        C[500]), .CO(C[501]) );
  FA_7688 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n3595), .CI(
        C[501]), .CO(C[502]) );
  FA_7687 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n3594), .CI(
        C[502]), .CO(C[503]) );
  FA_7686 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n3593), .CI(
        C[503]), .CO(C[504]) );
  FA_7685 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n3592), .CI(
        C[504]), .CO(C[505]) );
  FA_7684 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n3591), .CI(
        C[505]), .CO(C[506]) );
  FA_7683 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n3590), .CI(
        C[506]), .CO(C[507]) );
  FA_7682 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n3589), .CI(
        C[507]), .CO(C[508]) );
  FA_7681 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n3588), .CI(
        C[508]), .CO(C[509]) );
  FA_7680 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n3587), .CI(
        C[509]), .CO(C[510]) );
  FA_7679 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n3586), .CI(
        C[510]), .CO(C[511]) );
  FA_7678 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n3585), .CI(
        C[511]), .CO(C[512]) );
  FA_7677 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(n3584), .CI(C[512]), 
        .CO(C[513]) );
  FA_7676 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(n3583), .CI(C[513]), 
        .CO(C[514]) );
  FA_7675 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(n3582), .CI(C[514]), 
        .CO(C[515]) );
  FA_7674 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(n3581), .CI(C[515]), 
        .CO(C[516]) );
  FA_7673 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(n3580), .CI(C[516]), 
        .CO(C[517]) );
  FA_7672 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(n3579), .CI(C[517]), 
        .CO(C[518]) );
  FA_7671 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(n3578), .CI(C[518]), 
        .CO(C[519]) );
  FA_7670 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(n3577), .CI(C[519]), 
        .CO(C[520]) );
  FA_7669 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(n3576), .CI(C[520]), 
        .CO(C[521]) );
  FA_7668 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(n3575), .CI(C[521]), 
        .CO(C[522]) );
  FA_7667 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(n3574), .CI(C[522]), .CO(C[523]) );
  FA_7666 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(n3573), .CI(C[523]), .CO(C[524]) );
  FA_7665 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(n3572), .CI(C[524]), .CO(C[525]) );
  FA_7664 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(n3571), .CI(C[525]), .CO(C[526]) );
  FA_7663 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(n3570), .CI(C[526]), .CO(C[527]) );
  FA_7662 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(n3569), .CI(C[527]), .CO(C[528]) );
  FA_7661 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(n3568), .CI(C[528]), .CO(C[529]) );
  FA_7660 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(n3567), .CI(C[529]), .CO(C[530]) );
  FA_7659 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(n3566), .CI(C[530]), .CO(C[531]) );
  FA_7658 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(n3565), .CI(C[531]), .CO(C[532]) );
  FA_7657 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(n3564), .CI(C[532]), .CO(C[533]) );
  FA_7656 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(n3563), .CI(C[533]), .CO(C[534]) );
  FA_7655 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(n3562), .CI(C[534]), .CO(C[535]) );
  FA_7654 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(n3561), .CI(C[535]), .CO(C[536]) );
  FA_7653 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(n3560), .CI(C[536]), .CO(C[537]) );
  FA_7652 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(n3559), .CI(C[537]), .CO(C[538]) );
  FA_7651 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(n3558), .CI(C[538]), .CO(C[539]) );
  FA_7650 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(n3557), .CI(C[539]), .CO(C[540]) );
  FA_7649 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(n3556), .CI(C[540]), .CO(C[541]) );
  FA_7648 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(n3555), .CI(C[541]), .CO(C[542]) );
  FA_7647 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(n3554), .CI(C[542]), .CO(C[543]) );
  FA_7646 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(n3553), .CI(C[543]), .CO(C[544]) );
  FA_7645 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(n3552), .CI(C[544]), .CO(C[545]) );
  FA_7644 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(n3551), .CI(C[545]), .CO(C[546]) );
  FA_7643 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(n3550), .CI(C[546]), .CO(C[547]) );
  FA_7642 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(n3549), .CI(C[547]), .CO(C[548]) );
  FA_7641 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(n3548), .CI(C[548]), .CO(C[549]) );
  FA_7640 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(n3547), .CI(C[549]), .CO(C[550]) );
  FA_7639 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(n3546), .CI(C[550]), .CO(C[551]) );
  FA_7638 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(n3545), .CI(C[551]), .CO(C[552]) );
  FA_7637 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(n3544), .CI(C[552]), .CO(C[553]) );
  FA_7636 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(n3543), .CI(C[553]), .CO(C[554]) );
  FA_7635 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(n3542), .CI(C[554]), .CO(C[555]) );
  FA_7634 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(n3541), .CI(C[555]), .CO(C[556]) );
  FA_7633 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(n3540), .CI(C[556]), .CO(C[557]) );
  FA_7632 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(n3539), .CI(C[557]), .CO(C[558]) );
  FA_7631 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(n3538), .CI(C[558]), .CO(C[559]) );
  FA_7630 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(n3537), .CI(C[559]), .CO(C[560]) );
  FA_7629 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(n3536), .CI(C[560]), .CO(C[561]) );
  FA_7628 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(n3535), .CI(C[561]), .CO(C[562]) );
  FA_7627 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(n3534), .CI(C[562]), .CO(C[563]) );
  FA_7626 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(n3533), .CI(C[563]), .CO(C[564]) );
  FA_7625 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(n3532), .CI(C[564]), .CO(C[565]) );
  FA_7624 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(n3531), .CI(C[565]), .CO(C[566]) );
  FA_7623 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(n3530), .CI(C[566]), .CO(C[567]) );
  FA_7622 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(n3529), .CI(C[567]), .CO(C[568]) );
  FA_7621 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(n3528), .CI(C[568]), .CO(C[569]) );
  FA_7620 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(n3527), .CI(C[569]), .CO(C[570]) );
  FA_7619 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(n3526), .CI(C[570]), .CO(C[571]) );
  FA_7618 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(n3525), .CI(C[571]), .CO(C[572]) );
  FA_7617 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(n3524), .CI(C[572]), .CO(C[573]) );
  FA_7616 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(n3523), .CI(C[573]), .CO(C[574]) );
  FA_7615 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(n3522), .CI(C[574]), .CO(C[575]) );
  FA_7614 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(n3521), .CI(C[575]), .CO(C[576]) );
  FA_7613 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(n3520), .CI(C[576]), .CO(C[577]) );
  FA_7612 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(n3519), .CI(C[577]), .CO(C[578]) );
  FA_7611 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(n3518), .CI(C[578]), .CO(C[579]) );
  FA_7610 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(n3517), .CI(C[579]), .CO(C[580]) );
  FA_7609 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(n3516), .CI(C[580]), .CO(C[581]) );
  FA_7608 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(n3515), .CI(C[581]), .CO(C[582]) );
  FA_7607 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(n3514), .CI(C[582]), .CO(C[583]) );
  FA_7606 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(n3513), .CI(C[583]), .CO(C[584]) );
  FA_7605 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(n3512), .CI(C[584]), .CO(C[585]) );
  FA_7604 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(n3511), .CI(C[585]), .CO(C[586]) );
  FA_7603 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(n3510), .CI(C[586]), .CO(C[587]) );
  FA_7602 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(n3509), .CI(C[587]), .CO(C[588]) );
  FA_7601 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(n3508), .CI(C[588]), .CO(C[589]) );
  FA_7600 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(n3507), .CI(C[589]), .CO(C[590]) );
  FA_7599 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(n3506), .CI(C[590]), .CO(C[591]) );
  FA_7598 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(n3505), .CI(C[591]), .CO(C[592]) );
  FA_7597 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(n3504), .CI(C[592]), .CO(C[593]) );
  FA_7596 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(n3503), .CI(C[593]), .CO(C[594]) );
  FA_7595 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(n3502), .CI(C[594]), .CO(C[595]) );
  FA_7594 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(n3501), .CI(C[595]), .CO(C[596]) );
  FA_7593 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(n3500), .CI(C[596]), .CO(C[597]) );
  FA_7592 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(n3499), .CI(C[597]), .CO(C[598]) );
  FA_7591 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(n3498), .CI(C[598]), .CO(C[599]) );
  FA_7590 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(n3497), .CI(C[599]), .CO(C[600]) );
  FA_7589 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(n3496), .CI(C[600]), .CO(C[601]) );
  FA_7588 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(n3495), .CI(C[601]), .CO(C[602]) );
  FA_7587 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(n3494), .CI(C[602]), .CO(C[603]) );
  FA_7586 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(n3493), .CI(C[603]), .CO(C[604]) );
  FA_7585 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(n3492), .CI(C[604]), .CO(C[605]) );
  FA_7584 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(n3491), .CI(C[605]), .CO(C[606]) );
  FA_7583 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(n3490), .CI(C[606]), .CO(C[607]) );
  FA_7582 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(n3489), .CI(C[607]), .CO(C[608]) );
  FA_7581 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(n3488), .CI(C[608]), .CO(C[609]) );
  FA_7580 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(n3487), .CI(C[609]), .CO(C[610]) );
  FA_7579 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(n3486), .CI(C[610]), .CO(C[611]) );
  FA_7578 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(n3485), .CI(C[611]), .CO(C[612]) );
  FA_7577 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(n3484), .CI(
        C[612]), .CO(C[613]) );
  FA_7576 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(n3483), .CI(
        C[613]), .CO(C[614]) );
  FA_7575 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(n3482), .CI(
        C[614]), .CO(C[615]) );
  FA_7574 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(n3481), .CI(
        C[615]), .CO(C[616]) );
  FA_7573 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(n3480), .CI(
        C[616]), .CO(C[617]) );
  FA_7572 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(n3479), .CI(
        C[617]), .CO(C[618]) );
  FA_7571 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(n3478), .CI(
        C[618]), .CO(C[619]) );
  FA_7570 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(n3477), .CI(
        C[619]), .CO(C[620]) );
  FA_7569 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(n3476), .CI(
        C[620]), .CO(C[621]) );
  FA_7568 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(n3475), .CI(
        C[621]), .CO(C[622]) );
  FA_7567 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(n3474), .CI(
        C[622]), .CO(C[623]) );
  FA_7566 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(n3473), .CI(
        C[623]), .CO(C[624]) );
  FA_7565 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(n3472), .CI(
        C[624]), .CO(C[625]) );
  FA_7564 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(n3471), .CI(
        C[625]), .CO(C[626]) );
  FA_7563 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(n3470), .CI(
        C[626]), .CO(C[627]) );
  FA_7562 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(n3469), .CI(
        C[627]), .CO(C[628]) );
  FA_7561 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(n3468), .CI(
        C[628]), .CO(C[629]) );
  FA_7560 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(n3467), .CI(
        C[629]), .CO(C[630]) );
  FA_7559 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(n3466), .CI(
        C[630]), .CO(C[631]) );
  FA_7558 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(n3465), .CI(
        C[631]), .CO(C[632]) );
  FA_7557 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(n3464), .CI(
        C[632]), .CO(C[633]) );
  FA_7556 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(n3463), .CI(
        C[633]), .CO(C[634]) );
  FA_7555 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(n3462), .CI(
        C[634]), .CO(C[635]) );
  FA_7554 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(n3461), .CI(
        C[635]), .CO(C[636]) );
  FA_7553 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(n3460), .CI(
        C[636]), .CO(C[637]) );
  FA_7552 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(n3459), .CI(
        C[637]), .CO(C[638]) );
  FA_7551 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(n3458), .CI(
        C[638]), .CO(C[639]) );
  FA_7550 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(n3457), .CI(
        C[639]), .CO(C[640]) );
  FA_7549 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(n3456), .CI(
        C[640]), .CO(C[641]) );
  FA_7548 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(n3455), .CI(
        C[641]), .CO(C[642]) );
  FA_7547 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(n3454), .CI(
        C[642]), .CO(C[643]) );
  FA_7546 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(n3453), .CI(
        C[643]), .CO(C[644]) );
  FA_7545 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(n3452), .CI(
        C[644]), .CO(C[645]) );
  FA_7544 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(n3451), .CI(
        C[645]), .CO(C[646]) );
  FA_7543 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(n3450), .CI(
        C[646]), .CO(C[647]) );
  FA_7542 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(n3449), .CI(
        C[647]), .CO(C[648]) );
  FA_7541 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(n3448), .CI(
        C[648]), .CO(C[649]) );
  FA_7540 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(n3447), .CI(
        C[649]), .CO(C[650]) );
  FA_7539 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(n3446), .CI(
        C[650]), .CO(C[651]) );
  FA_7538 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(n3445), .CI(
        C[651]), .CO(C[652]) );
  FA_7537 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(n3444), .CI(
        C[652]), .CO(C[653]) );
  FA_7536 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(n3443), .CI(
        C[653]), .CO(C[654]) );
  FA_7535 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(n3442), .CI(
        C[654]), .CO(C[655]) );
  FA_7534 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(n3441), .CI(
        C[655]), .CO(C[656]) );
  FA_7533 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(n3440), .CI(
        C[656]), .CO(C[657]) );
  FA_7532 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(n3439), .CI(
        C[657]), .CO(C[658]) );
  FA_7531 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(n3438), .CI(
        C[658]), .CO(C[659]) );
  FA_7530 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(n3437), .CI(
        C[659]), .CO(C[660]) );
  FA_7529 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(n3436), .CI(
        C[660]), .CO(C[661]) );
  FA_7528 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(n3435), .CI(
        C[661]), .CO(C[662]) );
  FA_7527 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(n3434), .CI(
        C[662]), .CO(C[663]) );
  FA_7526 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(n3433), .CI(
        C[663]), .CO(C[664]) );
  FA_7525 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(n3432), .CI(
        C[664]), .CO(C[665]) );
  FA_7524 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(n3431), .CI(
        C[665]), .CO(C[666]) );
  FA_7523 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(n3430), .CI(
        C[666]), .CO(C[667]) );
  FA_7522 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(n3429), .CI(
        C[667]), .CO(C[668]) );
  FA_7521 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(n3428), .CI(
        C[668]), .CO(C[669]) );
  FA_7520 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(n3427), .CI(
        C[669]), .CO(C[670]) );
  FA_7519 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(n3426), .CI(
        C[670]), .CO(C[671]) );
  FA_7518 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(n3425), .CI(
        C[671]), .CO(C[672]) );
  FA_7517 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(n3424), .CI(
        C[672]), .CO(C[673]) );
  FA_7516 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(n3423), .CI(
        C[673]), .CO(C[674]) );
  FA_7515 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(n3422), .CI(
        C[674]), .CO(C[675]) );
  FA_7514 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(n3421), .CI(
        C[675]), .CO(C[676]) );
  FA_7513 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(n3420), .CI(
        C[676]), .CO(C[677]) );
  FA_7512 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(n3419), .CI(
        C[677]), .CO(C[678]) );
  FA_7511 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(n3418), .CI(
        C[678]), .CO(C[679]) );
  FA_7510 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(n3417), .CI(
        C[679]), .CO(C[680]) );
  FA_7509 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(n3416), .CI(
        C[680]), .CO(C[681]) );
  FA_7508 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(n3415), .CI(
        C[681]), .CO(C[682]) );
  FA_7507 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(n3414), .CI(
        C[682]), .CO(C[683]) );
  FA_7506 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(n3413), .CI(
        C[683]), .CO(C[684]) );
  FA_7505 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(n3412), .CI(
        C[684]), .CO(C[685]) );
  FA_7504 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(n3411), .CI(
        C[685]), .CO(C[686]) );
  FA_7503 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(n3410), .CI(
        C[686]), .CO(C[687]) );
  FA_7502 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(n3409), .CI(
        C[687]), .CO(C[688]) );
  FA_7501 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(n3408), .CI(
        C[688]), .CO(C[689]) );
  FA_7500 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(n3407), .CI(
        C[689]), .CO(C[690]) );
  FA_7499 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(n3406), .CI(
        C[690]), .CO(C[691]) );
  FA_7498 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(n3405), .CI(
        C[691]), .CO(C[692]) );
  FA_7497 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(n3404), .CI(
        C[692]), .CO(C[693]) );
  FA_7496 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(n3403), .CI(
        C[693]), .CO(C[694]) );
  FA_7495 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(n3402), .CI(
        C[694]), .CO(C[695]) );
  FA_7494 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(n3401), .CI(
        C[695]), .CO(C[696]) );
  FA_7493 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(n3400), .CI(
        C[696]), .CO(C[697]) );
  FA_7492 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(n3399), .CI(
        C[697]), .CO(C[698]) );
  FA_7491 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(n3398), .CI(
        C[698]), .CO(C[699]) );
  FA_7490 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(n3397), .CI(
        C[699]), .CO(C[700]) );
  FA_7489 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(n3396), .CI(
        C[700]), .CO(C[701]) );
  FA_7488 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(n3395), .CI(
        C[701]), .CO(C[702]) );
  FA_7487 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(n3394), .CI(
        C[702]), .CO(C[703]) );
  FA_7486 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(n3393), .CI(
        C[703]), .CO(C[704]) );
  FA_7485 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(n3392), .CI(
        C[704]), .CO(C[705]) );
  FA_7484 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(n3391), .CI(
        C[705]), .CO(C[706]) );
  FA_7483 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(n3390), .CI(
        C[706]), .CO(C[707]) );
  FA_7482 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(n3389), .CI(
        C[707]), .CO(C[708]) );
  FA_7481 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(n3388), .CI(
        C[708]), .CO(C[709]) );
  FA_7480 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(n3387), .CI(
        C[709]), .CO(C[710]) );
  FA_7479 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(n3386), .CI(
        C[710]), .CO(C[711]) );
  FA_7478 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(n3385), .CI(
        C[711]), .CO(C[712]) );
  FA_7477 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(n3384), .CI(
        C[712]), .CO(C[713]) );
  FA_7476 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(n3383), .CI(
        C[713]), .CO(C[714]) );
  FA_7475 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(n3382), .CI(
        C[714]), .CO(C[715]) );
  FA_7474 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(n3381), .CI(
        C[715]), .CO(C[716]) );
  FA_7473 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(n3380), .CI(
        C[716]), .CO(C[717]) );
  FA_7472 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(n3379), .CI(
        C[717]), .CO(C[718]) );
  FA_7471 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(n3378), .CI(
        C[718]), .CO(C[719]) );
  FA_7470 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(n3377), .CI(
        C[719]), .CO(C[720]) );
  FA_7469 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(n3376), .CI(
        C[720]), .CO(C[721]) );
  FA_7468 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(n3375), .CI(
        C[721]), .CO(C[722]) );
  FA_7467 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(n3374), .CI(
        C[722]), .CO(C[723]) );
  FA_7466 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(n3373), .CI(
        C[723]), .CO(C[724]) );
  FA_7465 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(n3372), .CI(
        C[724]), .CO(C[725]) );
  FA_7464 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(n3371), .CI(
        C[725]), .CO(C[726]) );
  FA_7463 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(n3370), .CI(
        C[726]), .CO(C[727]) );
  FA_7462 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(n3369), .CI(
        C[727]), .CO(C[728]) );
  FA_7461 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(n3368), .CI(
        C[728]), .CO(C[729]) );
  FA_7460 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(n3367), .CI(
        C[729]), .CO(C[730]) );
  FA_7459 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(n3366), .CI(
        C[730]), .CO(C[731]) );
  FA_7458 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(n3365), .CI(
        C[731]), .CO(C[732]) );
  FA_7457 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(n3364), .CI(
        C[732]), .CO(C[733]) );
  FA_7456 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(n3363), .CI(
        C[733]), .CO(C[734]) );
  FA_7455 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(n3362), .CI(
        C[734]), .CO(C[735]) );
  FA_7454 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(n3361), .CI(
        C[735]), .CO(C[736]) );
  FA_7453 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(n3360), .CI(
        C[736]), .CO(C[737]) );
  FA_7452 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(n3359), .CI(
        C[737]), .CO(C[738]) );
  FA_7451 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(n3358), .CI(
        C[738]), .CO(C[739]) );
  FA_7450 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(n3357), .CI(
        C[739]), .CO(C[740]) );
  FA_7449 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(n3356), .CI(
        C[740]), .CO(C[741]) );
  FA_7448 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(n3355), .CI(
        C[741]), .CO(C[742]) );
  FA_7447 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(n3354), .CI(
        C[742]), .CO(C[743]) );
  FA_7446 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(n3353), .CI(
        C[743]), .CO(C[744]) );
  FA_7445 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(n3352), .CI(
        C[744]), .CO(C[745]) );
  FA_7444 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(n3351), .CI(
        C[745]), .CO(C[746]) );
  FA_7443 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(n3350), .CI(
        C[746]), .CO(C[747]) );
  FA_7442 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(n3349), .CI(
        C[747]), .CO(C[748]) );
  FA_7441 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(n3348), .CI(
        C[748]), .CO(C[749]) );
  FA_7440 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(n3347), .CI(
        C[749]), .CO(C[750]) );
  FA_7439 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(n3346), .CI(
        C[750]), .CO(C[751]) );
  FA_7438 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(n3345), .CI(
        C[751]), .CO(C[752]) );
  FA_7437 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(n3344), .CI(
        C[752]), .CO(C[753]) );
  FA_7436 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(n3343), .CI(
        C[753]), .CO(C[754]) );
  FA_7435 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(n3342), .CI(
        C[754]), .CO(C[755]) );
  FA_7434 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(n3341), .CI(
        C[755]), .CO(C[756]) );
  FA_7433 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(n3340), .CI(
        C[756]), .CO(C[757]) );
  FA_7432 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(n3339), .CI(
        C[757]), .CO(C[758]) );
  FA_7431 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(n3338), .CI(
        C[758]), .CO(C[759]) );
  FA_7430 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(n3337), .CI(
        C[759]), .CO(C[760]) );
  FA_7429 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(n3336), .CI(
        C[760]), .CO(C[761]) );
  FA_7428 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(n3335), .CI(
        C[761]), .CO(C[762]) );
  FA_7427 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(n3334), .CI(
        C[762]), .CO(C[763]) );
  FA_7426 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(n3333), .CI(
        C[763]), .CO(C[764]) );
  FA_7425 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(n3332), .CI(
        C[764]), .CO(C[765]) );
  FA_7424 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(n3331), .CI(
        C[765]), .CO(C[766]) );
  FA_7423 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(n3330), .CI(
        C[766]), .CO(C[767]) );
  FA_7422 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(n3329), .CI(
        C[767]), .CO(C[768]) );
  FA_7421 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(n3328), .CI(
        C[768]), .CO(C[769]) );
  FA_7420 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(n3327), .CI(
        C[769]), .CO(C[770]) );
  FA_7419 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(n3326), .CI(
        C[770]), .CO(C[771]) );
  FA_7418 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(n3325), .CI(
        C[771]), .CO(C[772]) );
  FA_7417 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(n3324), .CI(
        C[772]), .CO(C[773]) );
  FA_7416 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(n3323), .CI(
        C[773]), .CO(C[774]) );
  FA_7415 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(n3322), .CI(
        C[774]), .CO(C[775]) );
  FA_7414 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(n3321), .CI(
        C[775]), .CO(C[776]) );
  FA_7413 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(n3320), .CI(
        C[776]), .CO(C[777]) );
  FA_7412 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(n3319), .CI(
        C[777]), .CO(C[778]) );
  FA_7411 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(n3318), .CI(
        C[778]), .CO(C[779]) );
  FA_7410 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(n3317), .CI(
        C[779]), .CO(C[780]) );
  FA_7409 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(n3316), .CI(
        C[780]), .CO(C[781]) );
  FA_7408 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(n3315), .CI(
        C[781]), .CO(C[782]) );
  FA_7407 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(n3314), .CI(
        C[782]), .CO(C[783]) );
  FA_7406 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(n3313), .CI(
        C[783]), .CO(C[784]) );
  FA_7405 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(n3312), .CI(
        C[784]), .CO(C[785]) );
  FA_7404 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(n3311), .CI(
        C[785]), .CO(C[786]) );
  FA_7403 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(n3310), .CI(
        C[786]), .CO(C[787]) );
  FA_7402 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(n3309), .CI(
        C[787]), .CO(C[788]) );
  FA_7401 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(n3308), .CI(
        C[788]), .CO(C[789]) );
  FA_7400 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(n3307), .CI(
        C[789]), .CO(C[790]) );
  FA_7399 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(n3306), .CI(
        C[790]), .CO(C[791]) );
  FA_7398 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(n3305), .CI(
        C[791]), .CO(C[792]) );
  FA_7397 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(n3304), .CI(
        C[792]), .CO(C[793]) );
  FA_7396 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(n3303), .CI(
        C[793]), .CO(C[794]) );
  FA_7395 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(n3302), .CI(
        C[794]), .CO(C[795]) );
  FA_7394 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(n3301), .CI(
        C[795]), .CO(C[796]) );
  FA_7393 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(n3300), .CI(
        C[796]), .CO(C[797]) );
  FA_7392 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(n3299), .CI(
        C[797]), .CO(C[798]) );
  FA_7391 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(n3298), .CI(
        C[798]), .CO(C[799]) );
  FA_7390 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(n3297), .CI(
        C[799]), .CO(C[800]) );
  FA_7389 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(n3296), .CI(
        C[800]), .CO(C[801]) );
  FA_7388 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(n3295), .CI(
        C[801]), .CO(C[802]) );
  FA_7387 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(n3294), .CI(
        C[802]), .CO(C[803]) );
  FA_7386 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(n3293), .CI(
        C[803]), .CO(C[804]) );
  FA_7385 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(n3292), .CI(
        C[804]), .CO(C[805]) );
  FA_7384 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(n3291), .CI(
        C[805]), .CO(C[806]) );
  FA_7383 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(n3290), .CI(
        C[806]), .CO(C[807]) );
  FA_7382 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(n3289), .CI(
        C[807]), .CO(C[808]) );
  FA_7381 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(n3288), .CI(
        C[808]), .CO(C[809]) );
  FA_7380 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(n3287), .CI(
        C[809]), .CO(C[810]) );
  FA_7379 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(n3286), .CI(
        C[810]), .CO(C[811]) );
  FA_7378 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(n3285), .CI(
        C[811]), .CO(C[812]) );
  FA_7377 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(n3284), .CI(
        C[812]), .CO(C[813]) );
  FA_7376 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(n3283), .CI(
        C[813]), .CO(C[814]) );
  FA_7375 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(n3282), .CI(
        C[814]), .CO(C[815]) );
  FA_7374 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(n3281), .CI(
        C[815]), .CO(C[816]) );
  FA_7373 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(n3280), .CI(
        C[816]), .CO(C[817]) );
  FA_7372 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(n3279), .CI(
        C[817]), .CO(C[818]) );
  FA_7371 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(n3278), .CI(
        C[818]), .CO(C[819]) );
  FA_7370 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(n3277), .CI(
        C[819]), .CO(C[820]) );
  FA_7369 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(n3276), .CI(
        C[820]), .CO(C[821]) );
  FA_7368 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(n3275), .CI(
        C[821]), .CO(C[822]) );
  FA_7367 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(n3274), .CI(
        C[822]), .CO(C[823]) );
  FA_7366 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(n3273), .CI(
        C[823]), .CO(C[824]) );
  FA_7365 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(n3272), .CI(
        C[824]), .CO(C[825]) );
  FA_7364 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(n3271), .CI(
        C[825]), .CO(C[826]) );
  FA_7363 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(n3270), .CI(
        C[826]), .CO(C[827]) );
  FA_7362 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(n3269), .CI(
        C[827]), .CO(C[828]) );
  FA_7361 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(n3268), .CI(
        C[828]), .CO(C[829]) );
  FA_7360 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(n3267), .CI(
        C[829]), .CO(C[830]) );
  FA_7359 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(n3266), .CI(
        C[830]), .CO(C[831]) );
  FA_7358 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(n3265), .CI(
        C[831]), .CO(C[832]) );
  FA_7357 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(n3264), .CI(
        C[832]), .CO(C[833]) );
  FA_7356 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(n3263), .CI(
        C[833]), .CO(C[834]) );
  FA_7355 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(n3262), .CI(
        C[834]), .CO(C[835]) );
  FA_7354 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(n3261), .CI(
        C[835]), .CO(C[836]) );
  FA_7353 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(n3260), .CI(
        C[836]), .CO(C[837]) );
  FA_7352 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(n3259), .CI(
        C[837]), .CO(C[838]) );
  FA_7351 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(n3258), .CI(
        C[838]), .CO(C[839]) );
  FA_7350 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(n3257), .CI(
        C[839]), .CO(C[840]) );
  FA_7349 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(n3256), .CI(
        C[840]), .CO(C[841]) );
  FA_7348 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(n3255), .CI(
        C[841]), .CO(C[842]) );
  FA_7347 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(n3254), .CI(
        C[842]), .CO(C[843]) );
  FA_7346 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(n3253), .CI(
        C[843]), .CO(C[844]) );
  FA_7345 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(n3252), .CI(
        C[844]), .CO(C[845]) );
  FA_7344 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(n3251), .CI(
        C[845]), .CO(C[846]) );
  FA_7343 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(n3250), .CI(
        C[846]), .CO(C[847]) );
  FA_7342 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(n3249), .CI(
        C[847]), .CO(C[848]) );
  FA_7341 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(n3248), .CI(
        C[848]), .CO(C[849]) );
  FA_7340 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(n3247), .CI(
        C[849]), .CO(C[850]) );
  FA_7339 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(n3246), .CI(
        C[850]), .CO(C[851]) );
  FA_7338 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(n3245), .CI(
        C[851]), .CO(C[852]) );
  FA_7337 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(n3244), .CI(
        C[852]), .CO(C[853]) );
  FA_7336 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(n3243), .CI(
        C[853]), .CO(C[854]) );
  FA_7335 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(n3242), .CI(
        C[854]), .CO(C[855]) );
  FA_7334 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(n3241), .CI(
        C[855]), .CO(C[856]) );
  FA_7333 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(n3240), .CI(
        C[856]), .CO(C[857]) );
  FA_7332 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(n3239), .CI(
        C[857]), .CO(C[858]) );
  FA_7331 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(n3238), .CI(
        C[858]), .CO(C[859]) );
  FA_7330 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(n3237), .CI(
        C[859]), .CO(C[860]) );
  FA_7329 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(n3236), .CI(
        C[860]), .CO(C[861]) );
  FA_7328 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(n3235), .CI(
        C[861]), .CO(C[862]) );
  FA_7327 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(n3234), .CI(
        C[862]), .CO(C[863]) );
  FA_7326 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(n3233), .CI(
        C[863]), .CO(C[864]) );
  FA_7325 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(n3232), .CI(
        C[864]), .CO(C[865]) );
  FA_7324 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(n3231), .CI(
        C[865]), .CO(C[866]) );
  FA_7323 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(n3230), .CI(
        C[866]), .CO(C[867]) );
  FA_7322 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(n3229), .CI(
        C[867]), .CO(C[868]) );
  FA_7321 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(n3228), .CI(
        C[868]), .CO(C[869]) );
  FA_7320 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(n3227), .CI(
        C[869]), .CO(C[870]) );
  FA_7319 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(n3226), .CI(
        C[870]), .CO(C[871]) );
  FA_7318 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(n3225), .CI(
        C[871]), .CO(C[872]) );
  FA_7317 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(n3224), .CI(
        C[872]), .CO(C[873]) );
  FA_7316 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(n3223), .CI(
        C[873]), .CO(C[874]) );
  FA_7315 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(n3222), .CI(
        C[874]), .CO(C[875]) );
  FA_7314 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(n3221), .CI(
        C[875]), .CO(C[876]) );
  FA_7313 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(n3220), .CI(
        C[876]), .CO(C[877]) );
  FA_7312 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(n3219), .CI(
        C[877]), .CO(C[878]) );
  FA_7311 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(n3218), .CI(
        C[878]), .CO(C[879]) );
  FA_7310 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(n3217), .CI(
        C[879]), .CO(C[880]) );
  FA_7309 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(n3216), .CI(
        C[880]), .CO(C[881]) );
  FA_7308 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(n3215), .CI(
        C[881]), .CO(C[882]) );
  FA_7307 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(n3214), .CI(
        C[882]), .CO(C[883]) );
  FA_7306 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(n3213), .CI(
        C[883]), .CO(C[884]) );
  FA_7305 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(n3212), .CI(
        C[884]), .CO(C[885]) );
  FA_7304 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(n3211), .CI(
        C[885]), .CO(C[886]) );
  FA_7303 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(n3210), .CI(
        C[886]), .CO(C[887]) );
  FA_7302 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(n3209), .CI(
        C[887]), .CO(C[888]) );
  FA_7301 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(n3208), .CI(
        C[888]), .CO(C[889]) );
  FA_7300 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(n3207), .CI(
        C[889]), .CO(C[890]) );
  FA_7299 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(n3206), .CI(
        C[890]), .CO(C[891]) );
  FA_7298 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(n3205), .CI(
        C[891]), .CO(C[892]) );
  FA_7297 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(n3204), .CI(
        C[892]), .CO(C[893]) );
  FA_7296 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(n3203), .CI(
        C[893]), .CO(C[894]) );
  FA_7295 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(n3202), .CI(
        C[894]), .CO(C[895]) );
  FA_7294 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(n3201), .CI(
        C[895]), .CO(C[896]) );
  FA_7293 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(n3200), .CI(
        C[896]), .CO(C[897]) );
  FA_7292 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(n3199), .CI(
        C[897]), .CO(C[898]) );
  FA_7291 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(n3198), .CI(
        C[898]), .CO(C[899]) );
  FA_7290 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(n3197), .CI(
        C[899]), .CO(C[900]) );
  FA_7289 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(n3196), .CI(
        C[900]), .CO(C[901]) );
  FA_7288 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(n3195), .CI(
        C[901]), .CO(C[902]) );
  FA_7287 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(n3194), .CI(
        C[902]), .CO(C[903]) );
  FA_7286 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(n3193), .CI(
        C[903]), .CO(C[904]) );
  FA_7285 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(n3192), .CI(
        C[904]), .CO(C[905]) );
  FA_7284 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(n3191), .CI(
        C[905]), .CO(C[906]) );
  FA_7283 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(n3190), .CI(
        C[906]), .CO(C[907]) );
  FA_7282 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(n3189), .CI(
        C[907]), .CO(C[908]) );
  FA_7281 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(n3188), .CI(
        C[908]), .CO(C[909]) );
  FA_7280 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(n3187), .CI(
        C[909]), .CO(C[910]) );
  FA_7279 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(n3186), .CI(
        C[910]), .CO(C[911]) );
  FA_7278 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(n3185), .CI(
        C[911]), .CO(C[912]) );
  FA_7277 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(n3184), .CI(
        C[912]), .CO(C[913]) );
  FA_7276 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(n3183), .CI(
        C[913]), .CO(C[914]) );
  FA_7275 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(n3182), .CI(
        C[914]), .CO(C[915]) );
  FA_7274 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(n3181), .CI(
        C[915]), .CO(C[916]) );
  FA_7273 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(n3180), .CI(
        C[916]), .CO(C[917]) );
  FA_7272 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(n3179), .CI(
        C[917]), .CO(C[918]) );
  FA_7271 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(n3178), .CI(
        C[918]), .CO(C[919]) );
  FA_7270 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(n3177), .CI(
        C[919]), .CO(C[920]) );
  FA_7269 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(n3176), .CI(
        C[920]), .CO(C[921]) );
  FA_7268 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(n3175), .CI(
        C[921]), .CO(C[922]) );
  FA_7267 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(n3174), .CI(
        C[922]), .CO(C[923]) );
  FA_7266 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(n3173), .CI(
        C[923]), .CO(C[924]) );
  FA_7265 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(n3172), .CI(
        C[924]), .CO(C[925]) );
  FA_7264 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(n3171), .CI(
        C[925]), .CO(C[926]) );
  FA_7263 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(n3170), .CI(
        C[926]), .CO(C[927]) );
  FA_7262 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(n3169), .CI(
        C[927]), .CO(C[928]) );
  FA_7261 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(n3168), .CI(
        C[928]), .CO(C[929]) );
  FA_7260 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(n3167), .CI(
        C[929]), .CO(C[930]) );
  FA_7259 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(n3166), .CI(
        C[930]), .CO(C[931]) );
  FA_7258 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(n3165), .CI(
        C[931]), .CO(C[932]) );
  FA_7257 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(n3164), .CI(
        C[932]), .CO(C[933]) );
  FA_7256 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(n3163), .CI(
        C[933]), .CO(C[934]) );
  FA_7255 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(n3162), .CI(
        C[934]), .CO(C[935]) );
  FA_7254 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(n3161), .CI(
        C[935]), .CO(C[936]) );
  FA_7253 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(n3160), .CI(
        C[936]), .CO(C[937]) );
  FA_7252 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(n3159), .CI(
        C[937]), .CO(C[938]) );
  FA_7251 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(n3158), .CI(
        C[938]), .CO(C[939]) );
  FA_7250 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(n3157), .CI(
        C[939]), .CO(C[940]) );
  FA_7249 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(n3156), .CI(
        C[940]), .CO(C[941]) );
  FA_7248 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(n3155), .CI(
        C[941]), .CO(C[942]) );
  FA_7247 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(n3154), .CI(
        C[942]), .CO(C[943]) );
  FA_7246 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(n3153), .CI(
        C[943]), .CO(C[944]) );
  FA_7245 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(n3152), .CI(
        C[944]), .CO(C[945]) );
  FA_7244 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(n3151), .CI(
        C[945]), .CO(C[946]) );
  FA_7243 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(n3150), .CI(
        C[946]), .CO(C[947]) );
  FA_7242 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(n3149), .CI(
        C[947]), .CO(C[948]) );
  FA_7241 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(n3148), .CI(
        C[948]), .CO(C[949]) );
  FA_7240 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(n3147), .CI(
        C[949]), .CO(C[950]) );
  FA_7239 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(n3146), .CI(
        C[950]), .CO(C[951]) );
  FA_7238 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(n3145), .CI(
        C[951]), .CO(C[952]) );
  FA_7237 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(n3144), .CI(
        C[952]), .CO(C[953]) );
  FA_7236 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(n3143), .CI(
        C[953]), .CO(C[954]) );
  FA_7235 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(n3142), .CI(
        C[954]), .CO(C[955]) );
  FA_7234 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(n3141), .CI(
        C[955]), .CO(C[956]) );
  FA_7233 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(n3140), .CI(
        C[956]), .CO(C[957]) );
  FA_7232 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(n3139), .CI(
        C[957]), .CO(C[958]) );
  FA_7231 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(n3138), .CI(
        C[958]), .CO(C[959]) );
  FA_7230 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(n3137), .CI(
        C[959]), .CO(C[960]) );
  FA_7229 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(n3136), .CI(
        C[960]), .CO(C[961]) );
  FA_7228 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(n3135), .CI(
        C[961]), .CO(C[962]) );
  FA_7227 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(n3134), .CI(
        C[962]), .CO(C[963]) );
  FA_7226 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(n3133), .CI(
        C[963]), .CO(C[964]) );
  FA_7225 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(n3132), .CI(
        C[964]), .CO(C[965]) );
  FA_7224 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(n3131), .CI(
        C[965]), .CO(C[966]) );
  FA_7223 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(n3130), .CI(
        C[966]), .CO(C[967]) );
  FA_7222 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(n3129), .CI(
        C[967]), .CO(C[968]) );
  FA_7221 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(n3128), .CI(
        C[968]), .CO(C[969]) );
  FA_7220 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(n3127), .CI(
        C[969]), .CO(C[970]) );
  FA_7219 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(n3126), .CI(
        C[970]), .CO(C[971]) );
  FA_7218 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(n3125), .CI(
        C[971]), .CO(C[972]) );
  FA_7217 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(n3124), .CI(
        C[972]), .CO(C[973]) );
  FA_7216 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(n3123), .CI(
        C[973]), .CO(C[974]) );
  FA_7215 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(n3122), .CI(
        C[974]), .CO(C[975]) );
  FA_7214 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(n3121), .CI(
        C[975]), .CO(C[976]) );
  FA_7213 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(n3120), .CI(
        C[976]), .CO(C[977]) );
  FA_7212 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(n3119), .CI(
        C[977]), .CO(C[978]) );
  FA_7211 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(n3118), .CI(
        C[978]), .CO(C[979]) );
  FA_7210 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(n3117), .CI(
        C[979]), .CO(C[980]) );
  FA_7209 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(n3116), .CI(
        C[980]), .CO(C[981]) );
  FA_7208 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(n3115), .CI(
        C[981]), .CO(C[982]) );
  FA_7207 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(n3114), .CI(
        C[982]), .CO(C[983]) );
  FA_7206 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(n3113), .CI(
        C[983]), .CO(C[984]) );
  FA_7205 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(n3112), .CI(
        C[984]), .CO(C[985]) );
  FA_7204 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(n3111), .CI(
        C[985]), .CO(C[986]) );
  FA_7203 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(n3110), .CI(
        C[986]), .CO(C[987]) );
  FA_7202 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(n3109), .CI(
        C[987]), .CO(C[988]) );
  FA_7201 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(n3108), .CI(
        C[988]), .CO(C[989]) );
  FA_7200 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(n3107), .CI(
        C[989]), .CO(C[990]) );
  FA_7199 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(n3106), .CI(
        C[990]), .CO(C[991]) );
  FA_7198 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(n3105), .CI(
        C[991]), .CO(C[992]) );
  FA_7197 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(n3104), .CI(
        C[992]), .CO(C[993]) );
  FA_7196 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(n3103), .CI(
        C[993]), .CO(C[994]) );
  FA_7195 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(n3102), .CI(
        C[994]), .CO(C[995]) );
  FA_7194 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(n3101), .CI(
        C[995]), .CO(C[996]) );
  FA_7193 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(n3100), .CI(
        C[996]), .CO(C[997]) );
  FA_7192 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(n3099), .CI(
        C[997]), .CO(C[998]) );
  FA_7191 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(n3098), .CI(
        C[998]), .CO(C[999]) );
  FA_7190 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(n3097), .CI(
        C[999]), .CO(C[1000]) );
  FA_7189 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(n3096), .CI(
        C[1000]), .CO(C[1001]) );
  FA_7188 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(n3095), .CI(
        C[1001]), .CO(C[1002]) );
  FA_7187 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(n3094), .CI(
        C[1002]), .CO(C[1003]) );
  FA_7186 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(n3093), .CI(
        C[1003]), .CO(C[1004]) );
  FA_7185 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(n3092), .CI(
        C[1004]), .CO(C[1005]) );
  FA_7184 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(n3091), .CI(
        C[1005]), .CO(C[1006]) );
  FA_7183 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(n3090), .CI(
        C[1006]), .CO(C[1007]) );
  FA_7182 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(n3089), .CI(
        C[1007]), .CO(C[1008]) );
  FA_7181 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(n3088), .CI(
        C[1008]), .CO(C[1009]) );
  FA_7180 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(n3087), .CI(
        C[1009]), .CO(C[1010]) );
  FA_7179 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(n3086), .CI(
        C[1010]), .CO(C[1011]) );
  FA_7178 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(n3085), .CI(
        C[1011]), .CO(C[1012]) );
  FA_7177 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(n3084), .CI(
        C[1012]), .CO(C[1013]) );
  FA_7176 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(n3083), .CI(
        C[1013]), .CO(C[1014]) );
  FA_7175 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(n3082), .CI(
        C[1014]), .CO(C[1015]) );
  FA_7174 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(n3081), .CI(
        C[1015]), .CO(C[1016]) );
  FA_7173 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(n3080), .CI(
        C[1016]), .CO(C[1017]) );
  FA_7172 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(n3079), .CI(
        C[1017]), .CO(C[1018]) );
  FA_7171 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(n3078), .CI(
        C[1018]), .CO(C[1019]) );
  FA_7170 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(n3077), .CI(
        C[1019]), .CO(C[1020]) );
  FA_7169 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(A[1020]), .B(n3076), .CI(
        C[1020]), .CO(C[1021]) );
  FA_7168 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(A[1021]), .B(n3075), .CI(
        C[1021]), .CO(C[1022]) );
  FA_7167 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(A[1022]), .B(n3074), .CI(
        C[1022]), .CO(C[1023]) );
  FA_7166 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(A[1023]), .B(n3073), .CI(
        C[1023]), .CO(C[1024]) );
  FA_7165 \FA_INST_0[2].FA_INST_1[0].FA_  ( .A(A[1024]), .B(n3072), .CI(
        C[1024]), .CO(C[1025]) );
  FA_7164 \FA_INST_0[2].FA_INST_1[1].FA_  ( .A(A[1025]), .B(n3071), .CI(
        C[1025]), .CO(C[1026]) );
  FA_7163 \FA_INST_0[2].FA_INST_1[2].FA_  ( .A(A[1026]), .B(n3070), .CI(
        C[1026]), .CO(C[1027]) );
  FA_7162 \FA_INST_0[2].FA_INST_1[3].FA_  ( .A(A[1027]), .B(n3069), .CI(
        C[1027]), .CO(C[1028]) );
  FA_7161 \FA_INST_0[2].FA_INST_1[4].FA_  ( .A(A[1028]), .B(n3068), .CI(
        C[1028]), .CO(C[1029]) );
  FA_7160 \FA_INST_0[2].FA_INST_1[5].FA_  ( .A(A[1029]), .B(n3067), .CI(
        C[1029]), .CO(C[1030]) );
  FA_7159 \FA_INST_0[2].FA_INST_1[6].FA_  ( .A(A[1030]), .B(n3066), .CI(
        C[1030]), .CO(C[1031]) );
  FA_7158 \FA_INST_0[2].FA_INST_1[7].FA_  ( .A(A[1031]), .B(n3065), .CI(
        C[1031]), .CO(C[1032]) );
  FA_7157 \FA_INST_0[2].FA_INST_1[8].FA_  ( .A(A[1032]), .B(n3064), .CI(
        C[1032]), .CO(C[1033]) );
  FA_7156 \FA_INST_0[2].FA_INST_1[9].FA_  ( .A(A[1033]), .B(n3063), .CI(
        C[1033]), .CO(C[1034]) );
  FA_7155 \FA_INST_0[2].FA_INST_1[10].FA_  ( .A(A[1034]), .B(n3062), .CI(
        C[1034]), .CO(C[1035]) );
  FA_7154 \FA_INST_0[2].FA_INST_1[11].FA_  ( .A(A[1035]), .B(n3061), .CI(
        C[1035]), .CO(C[1036]) );
  FA_7153 \FA_INST_0[2].FA_INST_1[12].FA_  ( .A(A[1036]), .B(n3060), .CI(
        C[1036]), .CO(C[1037]) );
  FA_7152 \FA_INST_0[2].FA_INST_1[13].FA_  ( .A(A[1037]), .B(n3059), .CI(
        C[1037]), .CO(C[1038]) );
  FA_7151 \FA_INST_0[2].FA_INST_1[14].FA_  ( .A(A[1038]), .B(n3058), .CI(
        C[1038]), .CO(C[1039]) );
  FA_7150 \FA_INST_0[2].FA_INST_1[15].FA_  ( .A(A[1039]), .B(n3057), .CI(
        C[1039]), .CO(C[1040]) );
  FA_7149 \FA_INST_0[2].FA_INST_1[16].FA_  ( .A(A[1040]), .B(n3056), .CI(
        C[1040]), .CO(C[1041]) );
  FA_7148 \FA_INST_0[2].FA_INST_1[17].FA_  ( .A(A[1041]), .B(n3055), .CI(
        C[1041]), .CO(C[1042]) );
  FA_7147 \FA_INST_0[2].FA_INST_1[18].FA_  ( .A(A[1042]), .B(n3054), .CI(
        C[1042]), .CO(C[1043]) );
  FA_7146 \FA_INST_0[2].FA_INST_1[19].FA_  ( .A(A[1043]), .B(n3053), .CI(
        C[1043]), .CO(C[1044]) );
  FA_7145 \FA_INST_0[2].FA_INST_1[20].FA_  ( .A(A[1044]), .B(n3052), .CI(
        C[1044]), .CO(C[1045]) );
  FA_7144 \FA_INST_0[2].FA_INST_1[21].FA_  ( .A(A[1045]), .B(n3051), .CI(
        C[1045]), .CO(C[1046]) );
  FA_7143 \FA_INST_0[2].FA_INST_1[22].FA_  ( .A(A[1046]), .B(n3050), .CI(
        C[1046]), .CO(C[1047]) );
  FA_7142 \FA_INST_0[2].FA_INST_1[23].FA_  ( .A(A[1047]), .B(n3049), .CI(
        C[1047]), .CO(C[1048]) );
  FA_7141 \FA_INST_0[2].FA_INST_1[24].FA_  ( .A(A[1048]), .B(n3048), .CI(
        C[1048]), .CO(C[1049]) );
  FA_7140 \FA_INST_0[2].FA_INST_1[25].FA_  ( .A(A[1049]), .B(n3047), .CI(
        C[1049]), .CO(C[1050]) );
  FA_7139 \FA_INST_0[2].FA_INST_1[26].FA_  ( .A(A[1050]), .B(n3046), .CI(
        C[1050]), .CO(C[1051]) );
  FA_7138 \FA_INST_0[2].FA_INST_1[27].FA_  ( .A(A[1051]), .B(n3045), .CI(
        C[1051]), .CO(C[1052]) );
  FA_7137 \FA_INST_0[2].FA_INST_1[28].FA_  ( .A(A[1052]), .B(n3044), .CI(
        C[1052]), .CO(C[1053]) );
  FA_7136 \FA_INST_0[2].FA_INST_1[29].FA_  ( .A(A[1053]), .B(n3043), .CI(
        C[1053]), .CO(C[1054]) );
  FA_7135 \FA_INST_0[2].FA_INST_1[30].FA_  ( .A(A[1054]), .B(n3042), .CI(
        C[1054]), .CO(C[1055]) );
  FA_7134 \FA_INST_0[2].FA_INST_1[31].FA_  ( .A(A[1055]), .B(n3041), .CI(
        C[1055]), .CO(C[1056]) );
  FA_7133 \FA_INST_0[2].FA_INST_1[32].FA_  ( .A(A[1056]), .B(n3040), .CI(
        C[1056]), .CO(C[1057]) );
  FA_7132 \FA_INST_0[2].FA_INST_1[33].FA_  ( .A(A[1057]), .B(n3039), .CI(
        C[1057]), .CO(C[1058]) );
  FA_7131 \FA_INST_0[2].FA_INST_1[34].FA_  ( .A(A[1058]), .B(n3038), .CI(
        C[1058]), .CO(C[1059]) );
  FA_7130 \FA_INST_0[2].FA_INST_1[35].FA_  ( .A(A[1059]), .B(n3037), .CI(
        C[1059]), .CO(C[1060]) );
  FA_7129 \FA_INST_0[2].FA_INST_1[36].FA_  ( .A(A[1060]), .B(n3036), .CI(
        C[1060]), .CO(C[1061]) );
  FA_7128 \FA_INST_0[2].FA_INST_1[37].FA_  ( .A(A[1061]), .B(n3035), .CI(
        C[1061]), .CO(C[1062]) );
  FA_7127 \FA_INST_0[2].FA_INST_1[38].FA_  ( .A(A[1062]), .B(n3034), .CI(
        C[1062]), .CO(C[1063]) );
  FA_7126 \FA_INST_0[2].FA_INST_1[39].FA_  ( .A(A[1063]), .B(n3033), .CI(
        C[1063]), .CO(C[1064]) );
  FA_7125 \FA_INST_0[2].FA_INST_1[40].FA_  ( .A(A[1064]), .B(n3032), .CI(
        C[1064]), .CO(C[1065]) );
  FA_7124 \FA_INST_0[2].FA_INST_1[41].FA_  ( .A(A[1065]), .B(n3031), .CI(
        C[1065]), .CO(C[1066]) );
  FA_7123 \FA_INST_0[2].FA_INST_1[42].FA_  ( .A(A[1066]), .B(n3030), .CI(
        C[1066]), .CO(C[1067]) );
  FA_7122 \FA_INST_0[2].FA_INST_1[43].FA_  ( .A(A[1067]), .B(n3029), .CI(
        C[1067]), .CO(C[1068]) );
  FA_7121 \FA_INST_0[2].FA_INST_1[44].FA_  ( .A(A[1068]), .B(n3028), .CI(
        C[1068]), .CO(C[1069]) );
  FA_7120 \FA_INST_0[2].FA_INST_1[45].FA_  ( .A(A[1069]), .B(n3027), .CI(
        C[1069]), .CO(C[1070]) );
  FA_7119 \FA_INST_0[2].FA_INST_1[46].FA_  ( .A(A[1070]), .B(n3026), .CI(
        C[1070]), .CO(C[1071]) );
  FA_7118 \FA_INST_0[2].FA_INST_1[47].FA_  ( .A(A[1071]), .B(n3025), .CI(
        C[1071]), .CO(C[1072]) );
  FA_7117 \FA_INST_0[2].FA_INST_1[48].FA_  ( .A(A[1072]), .B(n3024), .CI(
        C[1072]), .CO(C[1073]) );
  FA_7116 \FA_INST_0[2].FA_INST_1[49].FA_  ( .A(A[1073]), .B(n3023), .CI(
        C[1073]), .CO(C[1074]) );
  FA_7115 \FA_INST_0[2].FA_INST_1[50].FA_  ( .A(A[1074]), .B(n3022), .CI(
        C[1074]), .CO(C[1075]) );
  FA_7114 \FA_INST_0[2].FA_INST_1[51].FA_  ( .A(A[1075]), .B(n3021), .CI(
        C[1075]), .CO(C[1076]) );
  FA_7113 \FA_INST_0[2].FA_INST_1[52].FA_  ( .A(A[1076]), .B(n3020), .CI(
        C[1076]), .CO(C[1077]) );
  FA_7112 \FA_INST_0[2].FA_INST_1[53].FA_  ( .A(A[1077]), .B(n3019), .CI(
        C[1077]), .CO(C[1078]) );
  FA_7111 \FA_INST_0[2].FA_INST_1[54].FA_  ( .A(A[1078]), .B(n3018), .CI(
        C[1078]), .CO(C[1079]) );
  FA_7110 \FA_INST_0[2].FA_INST_1[55].FA_  ( .A(A[1079]), .B(n3017), .CI(
        C[1079]), .CO(C[1080]) );
  FA_7109 \FA_INST_0[2].FA_INST_1[56].FA_  ( .A(A[1080]), .B(n3016), .CI(
        C[1080]), .CO(C[1081]) );
  FA_7108 \FA_INST_0[2].FA_INST_1[57].FA_  ( .A(A[1081]), .B(n3015), .CI(
        C[1081]), .CO(C[1082]) );
  FA_7107 \FA_INST_0[2].FA_INST_1[58].FA_  ( .A(A[1082]), .B(n3014), .CI(
        C[1082]), .CO(C[1083]) );
  FA_7106 \FA_INST_0[2].FA_INST_1[59].FA_  ( .A(A[1083]), .B(n3013), .CI(
        C[1083]), .CO(C[1084]) );
  FA_7105 \FA_INST_0[2].FA_INST_1[60].FA_  ( .A(A[1084]), .B(n3012), .CI(
        C[1084]), .CO(C[1085]) );
  FA_7104 \FA_INST_0[2].FA_INST_1[61].FA_  ( .A(A[1085]), .B(n3011), .CI(
        C[1085]), .CO(C[1086]) );
  FA_7103 \FA_INST_0[2].FA_INST_1[62].FA_  ( .A(A[1086]), .B(n3010), .CI(
        C[1086]), .CO(C[1087]) );
  FA_7102 \FA_INST_0[2].FA_INST_1[63].FA_  ( .A(A[1087]), .B(n3009), .CI(
        C[1087]), .CO(C[1088]) );
  FA_7101 \FA_INST_0[2].FA_INST_1[64].FA_  ( .A(A[1088]), .B(n3008), .CI(
        C[1088]), .CO(C[1089]) );
  FA_7100 \FA_INST_0[2].FA_INST_1[65].FA_  ( .A(A[1089]), .B(n3007), .CI(
        C[1089]), .CO(C[1090]) );
  FA_7099 \FA_INST_0[2].FA_INST_1[66].FA_  ( .A(A[1090]), .B(n3006), .CI(
        C[1090]), .CO(C[1091]) );
  FA_7098 \FA_INST_0[2].FA_INST_1[67].FA_  ( .A(A[1091]), .B(n3005), .CI(
        C[1091]), .CO(C[1092]) );
  FA_7097 \FA_INST_0[2].FA_INST_1[68].FA_  ( .A(A[1092]), .B(n3004), .CI(
        C[1092]), .CO(C[1093]) );
  FA_7096 \FA_INST_0[2].FA_INST_1[69].FA_  ( .A(A[1093]), .B(n3003), .CI(
        C[1093]), .CO(C[1094]) );
  FA_7095 \FA_INST_0[2].FA_INST_1[70].FA_  ( .A(A[1094]), .B(n3002), .CI(
        C[1094]), .CO(C[1095]) );
  FA_7094 \FA_INST_0[2].FA_INST_1[71].FA_  ( .A(A[1095]), .B(n3001), .CI(
        C[1095]), .CO(C[1096]) );
  FA_7093 \FA_INST_0[2].FA_INST_1[72].FA_  ( .A(A[1096]), .B(n3000), .CI(
        C[1096]), .CO(C[1097]) );
  FA_7092 \FA_INST_0[2].FA_INST_1[73].FA_  ( .A(A[1097]), .B(n2999), .CI(
        C[1097]), .CO(C[1098]) );
  FA_7091 \FA_INST_0[2].FA_INST_1[74].FA_  ( .A(A[1098]), .B(n2998), .CI(
        C[1098]), .CO(C[1099]) );
  FA_7090 \FA_INST_0[2].FA_INST_1[75].FA_  ( .A(A[1099]), .B(n2997), .CI(
        C[1099]), .CO(C[1100]) );
  FA_7089 \FA_INST_0[2].FA_INST_1[76].FA_  ( .A(A[1100]), .B(n2996), .CI(
        C[1100]), .CO(C[1101]) );
  FA_7088 \FA_INST_0[2].FA_INST_1[77].FA_  ( .A(A[1101]), .B(n2995), .CI(
        C[1101]), .CO(C[1102]) );
  FA_7087 \FA_INST_0[2].FA_INST_1[78].FA_  ( .A(A[1102]), .B(n2994), .CI(
        C[1102]), .CO(C[1103]) );
  FA_7086 \FA_INST_0[2].FA_INST_1[79].FA_  ( .A(A[1103]), .B(n2993), .CI(
        C[1103]), .CO(C[1104]) );
  FA_7085 \FA_INST_0[2].FA_INST_1[80].FA_  ( .A(A[1104]), .B(n2992), .CI(
        C[1104]), .CO(C[1105]) );
  FA_7084 \FA_INST_0[2].FA_INST_1[81].FA_  ( .A(A[1105]), .B(n2991), .CI(
        C[1105]), .CO(C[1106]) );
  FA_7083 \FA_INST_0[2].FA_INST_1[82].FA_  ( .A(A[1106]), .B(n2990), .CI(
        C[1106]), .CO(C[1107]) );
  FA_7082 \FA_INST_0[2].FA_INST_1[83].FA_  ( .A(A[1107]), .B(n2989), .CI(
        C[1107]), .CO(C[1108]) );
  FA_7081 \FA_INST_0[2].FA_INST_1[84].FA_  ( .A(A[1108]), .B(n2988), .CI(
        C[1108]), .CO(C[1109]) );
  FA_7080 \FA_INST_0[2].FA_INST_1[85].FA_  ( .A(A[1109]), .B(n2987), .CI(
        C[1109]), .CO(C[1110]) );
  FA_7079 \FA_INST_0[2].FA_INST_1[86].FA_  ( .A(A[1110]), .B(n2986), .CI(
        C[1110]), .CO(C[1111]) );
  FA_7078 \FA_INST_0[2].FA_INST_1[87].FA_  ( .A(A[1111]), .B(n2985), .CI(
        C[1111]), .CO(C[1112]) );
  FA_7077 \FA_INST_0[2].FA_INST_1[88].FA_  ( .A(A[1112]), .B(n2984), .CI(
        C[1112]), .CO(C[1113]) );
  FA_7076 \FA_INST_0[2].FA_INST_1[89].FA_  ( .A(A[1113]), .B(n2983), .CI(
        C[1113]), .CO(C[1114]) );
  FA_7075 \FA_INST_0[2].FA_INST_1[90].FA_  ( .A(A[1114]), .B(n2982), .CI(
        C[1114]), .CO(C[1115]) );
  FA_7074 \FA_INST_0[2].FA_INST_1[91].FA_  ( .A(A[1115]), .B(n2981), .CI(
        C[1115]), .CO(C[1116]) );
  FA_7073 \FA_INST_0[2].FA_INST_1[92].FA_  ( .A(A[1116]), .B(n2980), .CI(
        C[1116]), .CO(C[1117]) );
  FA_7072 \FA_INST_0[2].FA_INST_1[93].FA_  ( .A(A[1117]), .B(n2979), .CI(
        C[1117]), .CO(C[1118]) );
  FA_7071 \FA_INST_0[2].FA_INST_1[94].FA_  ( .A(A[1118]), .B(n2978), .CI(
        C[1118]), .CO(C[1119]) );
  FA_7070 \FA_INST_0[2].FA_INST_1[95].FA_  ( .A(A[1119]), .B(n2977), .CI(
        C[1119]), .CO(C[1120]) );
  FA_7069 \FA_INST_0[2].FA_INST_1[96].FA_  ( .A(A[1120]), .B(n2976), .CI(
        C[1120]), .CO(C[1121]) );
  FA_7068 \FA_INST_0[2].FA_INST_1[97].FA_  ( .A(A[1121]), .B(n2975), .CI(
        C[1121]), .CO(C[1122]) );
  FA_7067 \FA_INST_0[2].FA_INST_1[98].FA_  ( .A(A[1122]), .B(n2974), .CI(
        C[1122]), .CO(C[1123]) );
  FA_7066 \FA_INST_0[2].FA_INST_1[99].FA_  ( .A(A[1123]), .B(n2973), .CI(
        C[1123]), .CO(C[1124]) );
  FA_7065 \FA_INST_0[2].FA_INST_1[100].FA_  ( .A(A[1124]), .B(n2972), .CI(
        C[1124]), .CO(C[1125]) );
  FA_7064 \FA_INST_0[2].FA_INST_1[101].FA_  ( .A(A[1125]), .B(n2971), .CI(
        C[1125]), .CO(C[1126]) );
  FA_7063 \FA_INST_0[2].FA_INST_1[102].FA_  ( .A(A[1126]), .B(n2970), .CI(
        C[1126]), .CO(C[1127]) );
  FA_7062 \FA_INST_0[2].FA_INST_1[103].FA_  ( .A(A[1127]), .B(n2969), .CI(
        C[1127]), .CO(C[1128]) );
  FA_7061 \FA_INST_0[2].FA_INST_1[104].FA_  ( .A(A[1128]), .B(n2968), .CI(
        C[1128]), .CO(C[1129]) );
  FA_7060 \FA_INST_0[2].FA_INST_1[105].FA_  ( .A(A[1129]), .B(n2967), .CI(
        C[1129]), .CO(C[1130]) );
  FA_7059 \FA_INST_0[2].FA_INST_1[106].FA_  ( .A(A[1130]), .B(n2966), .CI(
        C[1130]), .CO(C[1131]) );
  FA_7058 \FA_INST_0[2].FA_INST_1[107].FA_  ( .A(A[1131]), .B(n2965), .CI(
        C[1131]), .CO(C[1132]) );
  FA_7057 \FA_INST_0[2].FA_INST_1[108].FA_  ( .A(A[1132]), .B(n2964), .CI(
        C[1132]), .CO(C[1133]) );
  FA_7056 \FA_INST_0[2].FA_INST_1[109].FA_  ( .A(A[1133]), .B(n2963), .CI(
        C[1133]), .CO(C[1134]) );
  FA_7055 \FA_INST_0[2].FA_INST_1[110].FA_  ( .A(A[1134]), .B(n2962), .CI(
        C[1134]), .CO(C[1135]) );
  FA_7054 \FA_INST_0[2].FA_INST_1[111].FA_  ( .A(A[1135]), .B(n2961), .CI(
        C[1135]), .CO(C[1136]) );
  FA_7053 \FA_INST_0[2].FA_INST_1[112].FA_  ( .A(A[1136]), .B(n2960), .CI(
        C[1136]), .CO(C[1137]) );
  FA_7052 \FA_INST_0[2].FA_INST_1[113].FA_  ( .A(A[1137]), .B(n2959), .CI(
        C[1137]), .CO(C[1138]) );
  FA_7051 \FA_INST_0[2].FA_INST_1[114].FA_  ( .A(A[1138]), .B(n2958), .CI(
        C[1138]), .CO(C[1139]) );
  FA_7050 \FA_INST_0[2].FA_INST_1[115].FA_  ( .A(A[1139]), .B(n2957), .CI(
        C[1139]), .CO(C[1140]) );
  FA_7049 \FA_INST_0[2].FA_INST_1[116].FA_  ( .A(A[1140]), .B(n2956), .CI(
        C[1140]), .CO(C[1141]) );
  FA_7048 \FA_INST_0[2].FA_INST_1[117].FA_  ( .A(A[1141]), .B(n2955), .CI(
        C[1141]), .CO(C[1142]) );
  FA_7047 \FA_INST_0[2].FA_INST_1[118].FA_  ( .A(A[1142]), .B(n2954), .CI(
        C[1142]), .CO(C[1143]) );
  FA_7046 \FA_INST_0[2].FA_INST_1[119].FA_  ( .A(A[1143]), .B(n2953), .CI(
        C[1143]), .CO(C[1144]) );
  FA_7045 \FA_INST_0[2].FA_INST_1[120].FA_  ( .A(A[1144]), .B(n2952), .CI(
        C[1144]), .CO(C[1145]) );
  FA_7044 \FA_INST_0[2].FA_INST_1[121].FA_  ( .A(A[1145]), .B(n2951), .CI(
        C[1145]), .CO(C[1146]) );
  FA_7043 \FA_INST_0[2].FA_INST_1[122].FA_  ( .A(A[1146]), .B(n2950), .CI(
        C[1146]), .CO(C[1147]) );
  FA_7042 \FA_INST_0[2].FA_INST_1[123].FA_  ( .A(A[1147]), .B(n2949), .CI(
        C[1147]), .CO(C[1148]) );
  FA_7041 \FA_INST_0[2].FA_INST_1[124].FA_  ( .A(A[1148]), .B(n2948), .CI(
        C[1148]), .CO(C[1149]) );
  FA_7040 \FA_INST_0[2].FA_INST_1[125].FA_  ( .A(A[1149]), .B(n2947), .CI(
        C[1149]), .CO(C[1150]) );
  FA_7039 \FA_INST_0[2].FA_INST_1[126].FA_  ( .A(A[1150]), .B(n2946), .CI(
        C[1150]), .CO(C[1151]) );
  FA_7038 \FA_INST_0[2].FA_INST_1[127].FA_  ( .A(A[1151]), .B(n2945), .CI(
        C[1151]), .CO(C[1152]) );
  FA_7037 \FA_INST_0[2].FA_INST_1[128].FA_  ( .A(A[1152]), .B(n2944), .CI(
        C[1152]), .CO(C[1153]) );
  FA_7036 \FA_INST_0[2].FA_INST_1[129].FA_  ( .A(A[1153]), .B(n2943), .CI(
        C[1153]), .CO(C[1154]) );
  FA_7035 \FA_INST_0[2].FA_INST_1[130].FA_  ( .A(A[1154]), .B(n2942), .CI(
        C[1154]), .CO(C[1155]) );
  FA_7034 \FA_INST_0[2].FA_INST_1[131].FA_  ( .A(A[1155]), .B(n2941), .CI(
        C[1155]), .CO(C[1156]) );
  FA_7033 \FA_INST_0[2].FA_INST_1[132].FA_  ( .A(A[1156]), .B(n2940), .CI(
        C[1156]), .CO(C[1157]) );
  FA_7032 \FA_INST_0[2].FA_INST_1[133].FA_  ( .A(A[1157]), .B(n2939), .CI(
        C[1157]), .CO(C[1158]) );
  FA_7031 \FA_INST_0[2].FA_INST_1[134].FA_  ( .A(A[1158]), .B(n2938), .CI(
        C[1158]), .CO(C[1159]) );
  FA_7030 \FA_INST_0[2].FA_INST_1[135].FA_  ( .A(A[1159]), .B(n2937), .CI(
        C[1159]), .CO(C[1160]) );
  FA_7029 \FA_INST_0[2].FA_INST_1[136].FA_  ( .A(A[1160]), .B(n2936), .CI(
        C[1160]), .CO(C[1161]) );
  FA_7028 \FA_INST_0[2].FA_INST_1[137].FA_  ( .A(A[1161]), .B(n2935), .CI(
        C[1161]), .CO(C[1162]) );
  FA_7027 \FA_INST_0[2].FA_INST_1[138].FA_  ( .A(A[1162]), .B(n2934), .CI(
        C[1162]), .CO(C[1163]) );
  FA_7026 \FA_INST_0[2].FA_INST_1[139].FA_  ( .A(A[1163]), .B(n2933), .CI(
        C[1163]), .CO(C[1164]) );
  FA_7025 \FA_INST_0[2].FA_INST_1[140].FA_  ( .A(A[1164]), .B(n2932), .CI(
        C[1164]), .CO(C[1165]) );
  FA_7024 \FA_INST_0[2].FA_INST_1[141].FA_  ( .A(A[1165]), .B(n2931), .CI(
        C[1165]), .CO(C[1166]) );
  FA_7023 \FA_INST_0[2].FA_INST_1[142].FA_  ( .A(A[1166]), .B(n2930), .CI(
        C[1166]), .CO(C[1167]) );
  FA_7022 \FA_INST_0[2].FA_INST_1[143].FA_  ( .A(A[1167]), .B(n2929), .CI(
        C[1167]), .CO(C[1168]) );
  FA_7021 \FA_INST_0[2].FA_INST_1[144].FA_  ( .A(A[1168]), .B(n2928), .CI(
        C[1168]), .CO(C[1169]) );
  FA_7020 \FA_INST_0[2].FA_INST_1[145].FA_  ( .A(A[1169]), .B(n2927), .CI(
        C[1169]), .CO(C[1170]) );
  FA_7019 \FA_INST_0[2].FA_INST_1[146].FA_  ( .A(A[1170]), .B(n2926), .CI(
        C[1170]), .CO(C[1171]) );
  FA_7018 \FA_INST_0[2].FA_INST_1[147].FA_  ( .A(A[1171]), .B(n2925), .CI(
        C[1171]), .CO(C[1172]) );
  FA_7017 \FA_INST_0[2].FA_INST_1[148].FA_  ( .A(A[1172]), .B(n2924), .CI(
        C[1172]), .CO(C[1173]) );
  FA_7016 \FA_INST_0[2].FA_INST_1[149].FA_  ( .A(A[1173]), .B(n2923), .CI(
        C[1173]), .CO(C[1174]) );
  FA_7015 \FA_INST_0[2].FA_INST_1[150].FA_  ( .A(A[1174]), .B(n2922), .CI(
        C[1174]), .CO(C[1175]) );
  FA_7014 \FA_INST_0[2].FA_INST_1[151].FA_  ( .A(A[1175]), .B(n2921), .CI(
        C[1175]), .CO(C[1176]) );
  FA_7013 \FA_INST_0[2].FA_INST_1[152].FA_  ( .A(A[1176]), .B(n2920), .CI(
        C[1176]), .CO(C[1177]) );
  FA_7012 \FA_INST_0[2].FA_INST_1[153].FA_  ( .A(A[1177]), .B(n2919), .CI(
        C[1177]), .CO(C[1178]) );
  FA_7011 \FA_INST_0[2].FA_INST_1[154].FA_  ( .A(A[1178]), .B(n2918), .CI(
        C[1178]), .CO(C[1179]) );
  FA_7010 \FA_INST_0[2].FA_INST_1[155].FA_  ( .A(A[1179]), .B(n2917), .CI(
        C[1179]), .CO(C[1180]) );
  FA_7009 \FA_INST_0[2].FA_INST_1[156].FA_  ( .A(A[1180]), .B(n2916), .CI(
        C[1180]), .CO(C[1181]) );
  FA_7008 \FA_INST_0[2].FA_INST_1[157].FA_  ( .A(A[1181]), .B(n2915), .CI(
        C[1181]), .CO(C[1182]) );
  FA_7007 \FA_INST_0[2].FA_INST_1[158].FA_  ( .A(A[1182]), .B(n2914), .CI(
        C[1182]), .CO(C[1183]) );
  FA_7006 \FA_INST_0[2].FA_INST_1[159].FA_  ( .A(A[1183]), .B(n2913), .CI(
        C[1183]), .CO(C[1184]) );
  FA_7005 \FA_INST_0[2].FA_INST_1[160].FA_  ( .A(A[1184]), .B(n2912), .CI(
        C[1184]), .CO(C[1185]) );
  FA_7004 \FA_INST_0[2].FA_INST_1[161].FA_  ( .A(A[1185]), .B(n2911), .CI(
        C[1185]), .CO(C[1186]) );
  FA_7003 \FA_INST_0[2].FA_INST_1[162].FA_  ( .A(A[1186]), .B(n2910), .CI(
        C[1186]), .CO(C[1187]) );
  FA_7002 \FA_INST_0[2].FA_INST_1[163].FA_  ( .A(A[1187]), .B(n2909), .CI(
        C[1187]), .CO(C[1188]) );
  FA_7001 \FA_INST_0[2].FA_INST_1[164].FA_  ( .A(A[1188]), .B(n2908), .CI(
        C[1188]), .CO(C[1189]) );
  FA_7000 \FA_INST_0[2].FA_INST_1[165].FA_  ( .A(A[1189]), .B(n2907), .CI(
        C[1189]), .CO(C[1190]) );
  FA_6999 \FA_INST_0[2].FA_INST_1[166].FA_  ( .A(A[1190]), .B(n2906), .CI(
        C[1190]), .CO(C[1191]) );
  FA_6998 \FA_INST_0[2].FA_INST_1[167].FA_  ( .A(A[1191]), .B(n2905), .CI(
        C[1191]), .CO(C[1192]) );
  FA_6997 \FA_INST_0[2].FA_INST_1[168].FA_  ( .A(A[1192]), .B(n2904), .CI(
        C[1192]), .CO(C[1193]) );
  FA_6996 \FA_INST_0[2].FA_INST_1[169].FA_  ( .A(A[1193]), .B(n2903), .CI(
        C[1193]), .CO(C[1194]) );
  FA_6995 \FA_INST_0[2].FA_INST_1[170].FA_  ( .A(A[1194]), .B(n2902), .CI(
        C[1194]), .CO(C[1195]) );
  FA_6994 \FA_INST_0[2].FA_INST_1[171].FA_  ( .A(A[1195]), .B(n2901), .CI(
        C[1195]), .CO(C[1196]) );
  FA_6993 \FA_INST_0[2].FA_INST_1[172].FA_  ( .A(A[1196]), .B(n2900), .CI(
        C[1196]), .CO(C[1197]) );
  FA_6992 \FA_INST_0[2].FA_INST_1[173].FA_  ( .A(A[1197]), .B(n2899), .CI(
        C[1197]), .CO(C[1198]) );
  FA_6991 \FA_INST_0[2].FA_INST_1[174].FA_  ( .A(A[1198]), .B(n2898), .CI(
        C[1198]), .CO(C[1199]) );
  FA_6990 \FA_INST_0[2].FA_INST_1[175].FA_  ( .A(A[1199]), .B(n2897), .CI(
        C[1199]), .CO(C[1200]) );
  FA_6989 \FA_INST_0[2].FA_INST_1[176].FA_  ( .A(A[1200]), .B(n2896), .CI(
        C[1200]), .CO(C[1201]) );
  FA_6988 \FA_INST_0[2].FA_INST_1[177].FA_  ( .A(A[1201]), .B(n2895), .CI(
        C[1201]), .CO(C[1202]) );
  FA_6987 \FA_INST_0[2].FA_INST_1[178].FA_  ( .A(A[1202]), .B(n2894), .CI(
        C[1202]), .CO(C[1203]) );
  FA_6986 \FA_INST_0[2].FA_INST_1[179].FA_  ( .A(A[1203]), .B(n2893), .CI(
        C[1203]), .CO(C[1204]) );
  FA_6985 \FA_INST_0[2].FA_INST_1[180].FA_  ( .A(A[1204]), .B(n2892), .CI(
        C[1204]), .CO(C[1205]) );
  FA_6984 \FA_INST_0[2].FA_INST_1[181].FA_  ( .A(A[1205]), .B(n2891), .CI(
        C[1205]), .CO(C[1206]) );
  FA_6983 \FA_INST_0[2].FA_INST_1[182].FA_  ( .A(A[1206]), .B(n2890), .CI(
        C[1206]), .CO(C[1207]) );
  FA_6982 \FA_INST_0[2].FA_INST_1[183].FA_  ( .A(A[1207]), .B(n2889), .CI(
        C[1207]), .CO(C[1208]) );
  FA_6981 \FA_INST_0[2].FA_INST_1[184].FA_  ( .A(A[1208]), .B(n2888), .CI(
        C[1208]), .CO(C[1209]) );
  FA_6980 \FA_INST_0[2].FA_INST_1[185].FA_  ( .A(A[1209]), .B(n2887), .CI(
        C[1209]), .CO(C[1210]) );
  FA_6979 \FA_INST_0[2].FA_INST_1[186].FA_  ( .A(A[1210]), .B(n2886), .CI(
        C[1210]), .CO(C[1211]) );
  FA_6978 \FA_INST_0[2].FA_INST_1[187].FA_  ( .A(A[1211]), .B(n2885), .CI(
        C[1211]), .CO(C[1212]) );
  FA_6977 \FA_INST_0[2].FA_INST_1[188].FA_  ( .A(A[1212]), .B(n2884), .CI(
        C[1212]), .CO(C[1213]) );
  FA_6976 \FA_INST_0[2].FA_INST_1[189].FA_  ( .A(A[1213]), .B(n2883), .CI(
        C[1213]), .CO(C[1214]) );
  FA_6975 \FA_INST_0[2].FA_INST_1[190].FA_  ( .A(A[1214]), .B(n2882), .CI(
        C[1214]), .CO(C[1215]) );
  FA_6974 \FA_INST_0[2].FA_INST_1[191].FA_  ( .A(A[1215]), .B(n2881), .CI(
        C[1215]), .CO(C[1216]) );
  FA_6973 \FA_INST_0[2].FA_INST_1[192].FA_  ( .A(A[1216]), .B(n2880), .CI(
        C[1216]), .CO(C[1217]) );
  FA_6972 \FA_INST_0[2].FA_INST_1[193].FA_  ( .A(A[1217]), .B(n2879), .CI(
        C[1217]), .CO(C[1218]) );
  FA_6971 \FA_INST_0[2].FA_INST_1[194].FA_  ( .A(A[1218]), .B(n2878), .CI(
        C[1218]), .CO(C[1219]) );
  FA_6970 \FA_INST_0[2].FA_INST_1[195].FA_  ( .A(A[1219]), .B(n2877), .CI(
        C[1219]), .CO(C[1220]) );
  FA_6969 \FA_INST_0[2].FA_INST_1[196].FA_  ( .A(A[1220]), .B(n2876), .CI(
        C[1220]), .CO(C[1221]) );
  FA_6968 \FA_INST_0[2].FA_INST_1[197].FA_  ( .A(A[1221]), .B(n2875), .CI(
        C[1221]), .CO(C[1222]) );
  FA_6967 \FA_INST_0[2].FA_INST_1[198].FA_  ( .A(A[1222]), .B(n2874), .CI(
        C[1222]), .CO(C[1223]) );
  FA_6966 \FA_INST_0[2].FA_INST_1[199].FA_  ( .A(A[1223]), .B(n2873), .CI(
        C[1223]), .CO(C[1224]) );
  FA_6965 \FA_INST_0[2].FA_INST_1[200].FA_  ( .A(A[1224]), .B(n2872), .CI(
        C[1224]), .CO(C[1225]) );
  FA_6964 \FA_INST_0[2].FA_INST_1[201].FA_  ( .A(A[1225]), .B(n2871), .CI(
        C[1225]), .CO(C[1226]) );
  FA_6963 \FA_INST_0[2].FA_INST_1[202].FA_  ( .A(A[1226]), .B(n2870), .CI(
        C[1226]), .CO(C[1227]) );
  FA_6962 \FA_INST_0[2].FA_INST_1[203].FA_  ( .A(A[1227]), .B(n2869), .CI(
        C[1227]), .CO(C[1228]) );
  FA_6961 \FA_INST_0[2].FA_INST_1[204].FA_  ( .A(A[1228]), .B(n2868), .CI(
        C[1228]), .CO(C[1229]) );
  FA_6960 \FA_INST_0[2].FA_INST_1[205].FA_  ( .A(A[1229]), .B(n2867), .CI(
        C[1229]), .CO(C[1230]) );
  FA_6959 \FA_INST_0[2].FA_INST_1[206].FA_  ( .A(A[1230]), .B(n2866), .CI(
        C[1230]), .CO(C[1231]) );
  FA_6958 \FA_INST_0[2].FA_INST_1[207].FA_  ( .A(A[1231]), .B(n2865), .CI(
        C[1231]), .CO(C[1232]) );
  FA_6957 \FA_INST_0[2].FA_INST_1[208].FA_  ( .A(A[1232]), .B(n2864), .CI(
        C[1232]), .CO(C[1233]) );
  FA_6956 \FA_INST_0[2].FA_INST_1[209].FA_  ( .A(A[1233]), .B(n2863), .CI(
        C[1233]), .CO(C[1234]) );
  FA_6955 \FA_INST_0[2].FA_INST_1[210].FA_  ( .A(A[1234]), .B(n2862), .CI(
        C[1234]), .CO(C[1235]) );
  FA_6954 \FA_INST_0[2].FA_INST_1[211].FA_  ( .A(A[1235]), .B(n2861), .CI(
        C[1235]), .CO(C[1236]) );
  FA_6953 \FA_INST_0[2].FA_INST_1[212].FA_  ( .A(A[1236]), .B(n2860), .CI(
        C[1236]), .CO(C[1237]) );
  FA_6952 \FA_INST_0[2].FA_INST_1[213].FA_  ( .A(A[1237]), .B(n2859), .CI(
        C[1237]), .CO(C[1238]) );
  FA_6951 \FA_INST_0[2].FA_INST_1[214].FA_  ( .A(A[1238]), .B(n2858), .CI(
        C[1238]), .CO(C[1239]) );
  FA_6950 \FA_INST_0[2].FA_INST_1[215].FA_  ( .A(A[1239]), .B(n2857), .CI(
        C[1239]), .CO(C[1240]) );
  FA_6949 \FA_INST_0[2].FA_INST_1[216].FA_  ( .A(A[1240]), .B(n2856), .CI(
        C[1240]), .CO(C[1241]) );
  FA_6948 \FA_INST_0[2].FA_INST_1[217].FA_  ( .A(A[1241]), .B(n2855), .CI(
        C[1241]), .CO(C[1242]) );
  FA_6947 \FA_INST_0[2].FA_INST_1[218].FA_  ( .A(A[1242]), .B(n2854), .CI(
        C[1242]), .CO(C[1243]) );
  FA_6946 \FA_INST_0[2].FA_INST_1[219].FA_  ( .A(A[1243]), .B(n2853), .CI(
        C[1243]), .CO(C[1244]) );
  FA_6945 \FA_INST_0[2].FA_INST_1[220].FA_  ( .A(A[1244]), .B(n2852), .CI(
        C[1244]), .CO(C[1245]) );
  FA_6944 \FA_INST_0[2].FA_INST_1[221].FA_  ( .A(A[1245]), .B(n2851), .CI(
        C[1245]), .CO(C[1246]) );
  FA_6943 \FA_INST_0[2].FA_INST_1[222].FA_  ( .A(A[1246]), .B(n2850), .CI(
        C[1246]), .CO(C[1247]) );
  FA_6942 \FA_INST_0[2].FA_INST_1[223].FA_  ( .A(A[1247]), .B(n2849), .CI(
        C[1247]), .CO(C[1248]) );
  FA_6941 \FA_INST_0[2].FA_INST_1[224].FA_  ( .A(A[1248]), .B(n2848), .CI(
        C[1248]), .CO(C[1249]) );
  FA_6940 \FA_INST_0[2].FA_INST_1[225].FA_  ( .A(A[1249]), .B(n2847), .CI(
        C[1249]), .CO(C[1250]) );
  FA_6939 \FA_INST_0[2].FA_INST_1[226].FA_  ( .A(A[1250]), .B(n2846), .CI(
        C[1250]), .CO(C[1251]) );
  FA_6938 \FA_INST_0[2].FA_INST_1[227].FA_  ( .A(A[1251]), .B(n2845), .CI(
        C[1251]), .CO(C[1252]) );
  FA_6937 \FA_INST_0[2].FA_INST_1[228].FA_  ( .A(A[1252]), .B(n2844), .CI(
        C[1252]), .CO(C[1253]) );
  FA_6936 \FA_INST_0[2].FA_INST_1[229].FA_  ( .A(A[1253]), .B(n2843), .CI(
        C[1253]), .CO(C[1254]) );
  FA_6935 \FA_INST_0[2].FA_INST_1[230].FA_  ( .A(A[1254]), .B(n2842), .CI(
        C[1254]), .CO(C[1255]) );
  FA_6934 \FA_INST_0[2].FA_INST_1[231].FA_  ( .A(A[1255]), .B(n2841), .CI(
        C[1255]), .CO(C[1256]) );
  FA_6933 \FA_INST_0[2].FA_INST_1[232].FA_  ( .A(A[1256]), .B(n2840), .CI(
        C[1256]), .CO(C[1257]) );
  FA_6932 \FA_INST_0[2].FA_INST_1[233].FA_  ( .A(A[1257]), .B(n2839), .CI(
        C[1257]), .CO(C[1258]) );
  FA_6931 \FA_INST_0[2].FA_INST_1[234].FA_  ( .A(A[1258]), .B(n2838), .CI(
        C[1258]), .CO(C[1259]) );
  FA_6930 \FA_INST_0[2].FA_INST_1[235].FA_  ( .A(A[1259]), .B(n2837), .CI(
        C[1259]), .CO(C[1260]) );
  FA_6929 \FA_INST_0[2].FA_INST_1[236].FA_  ( .A(A[1260]), .B(n2836), .CI(
        C[1260]), .CO(C[1261]) );
  FA_6928 \FA_INST_0[2].FA_INST_1[237].FA_  ( .A(A[1261]), .B(n2835), .CI(
        C[1261]), .CO(C[1262]) );
  FA_6927 \FA_INST_0[2].FA_INST_1[238].FA_  ( .A(A[1262]), .B(n2834), .CI(
        C[1262]), .CO(C[1263]) );
  FA_6926 \FA_INST_0[2].FA_INST_1[239].FA_  ( .A(A[1263]), .B(n2833), .CI(
        C[1263]), .CO(C[1264]) );
  FA_6925 \FA_INST_0[2].FA_INST_1[240].FA_  ( .A(A[1264]), .B(n2832), .CI(
        C[1264]), .CO(C[1265]) );
  FA_6924 \FA_INST_0[2].FA_INST_1[241].FA_  ( .A(A[1265]), .B(n2831), .CI(
        C[1265]), .CO(C[1266]) );
  FA_6923 \FA_INST_0[2].FA_INST_1[242].FA_  ( .A(A[1266]), .B(n2830), .CI(
        C[1266]), .CO(C[1267]) );
  FA_6922 \FA_INST_0[2].FA_INST_1[243].FA_  ( .A(A[1267]), .B(n2829), .CI(
        C[1267]), .CO(C[1268]) );
  FA_6921 \FA_INST_0[2].FA_INST_1[244].FA_  ( .A(A[1268]), .B(n2828), .CI(
        C[1268]), .CO(C[1269]) );
  FA_6920 \FA_INST_0[2].FA_INST_1[245].FA_  ( .A(A[1269]), .B(n2827), .CI(
        C[1269]), .CO(C[1270]) );
  FA_6919 \FA_INST_0[2].FA_INST_1[246].FA_  ( .A(A[1270]), .B(n2826), .CI(
        C[1270]), .CO(C[1271]) );
  FA_6918 \FA_INST_0[2].FA_INST_1[247].FA_  ( .A(A[1271]), .B(n2825), .CI(
        C[1271]), .CO(C[1272]) );
  FA_6917 \FA_INST_0[2].FA_INST_1[248].FA_  ( .A(A[1272]), .B(n2824), .CI(
        C[1272]), .CO(C[1273]) );
  FA_6916 \FA_INST_0[2].FA_INST_1[249].FA_  ( .A(A[1273]), .B(n2823), .CI(
        C[1273]), .CO(C[1274]) );
  FA_6915 \FA_INST_0[2].FA_INST_1[250].FA_  ( .A(A[1274]), .B(n2822), .CI(
        C[1274]), .CO(C[1275]) );
  FA_6914 \FA_INST_0[2].FA_INST_1[251].FA_  ( .A(A[1275]), .B(n2821), .CI(
        C[1275]), .CO(C[1276]) );
  FA_6913 \FA_INST_0[2].FA_INST_1[252].FA_  ( .A(A[1276]), .B(n2820), .CI(
        C[1276]), .CO(C[1277]) );
  FA_6912 \FA_INST_0[2].FA_INST_1[253].FA_  ( .A(A[1277]), .B(n2819), .CI(
        C[1277]), .CO(C[1278]) );
  FA_6911 \FA_INST_0[2].FA_INST_1[254].FA_  ( .A(A[1278]), .B(n2818), .CI(
        C[1278]), .CO(C[1279]) );
  FA_6910 \FA_INST_0[2].FA_INST_1[255].FA_  ( .A(A[1279]), .B(n2817), .CI(
        C[1279]), .CO(C[1280]) );
  FA_6909 \FA_INST_0[2].FA_INST_1[256].FA_  ( .A(A[1280]), .B(n2816), .CI(
        C[1280]), .CO(C[1281]) );
  FA_6908 \FA_INST_0[2].FA_INST_1[257].FA_  ( .A(A[1281]), .B(n2815), .CI(
        C[1281]), .CO(C[1282]) );
  FA_6907 \FA_INST_0[2].FA_INST_1[258].FA_  ( .A(A[1282]), .B(n2814), .CI(
        C[1282]), .CO(C[1283]) );
  FA_6906 \FA_INST_0[2].FA_INST_1[259].FA_  ( .A(A[1283]), .B(n2813), .CI(
        C[1283]), .CO(C[1284]) );
  FA_6905 \FA_INST_0[2].FA_INST_1[260].FA_  ( .A(A[1284]), .B(n2812), .CI(
        C[1284]), .CO(C[1285]) );
  FA_6904 \FA_INST_0[2].FA_INST_1[261].FA_  ( .A(A[1285]), .B(n2811), .CI(
        C[1285]), .CO(C[1286]) );
  FA_6903 \FA_INST_0[2].FA_INST_1[262].FA_  ( .A(A[1286]), .B(n2810), .CI(
        C[1286]), .CO(C[1287]) );
  FA_6902 \FA_INST_0[2].FA_INST_1[263].FA_  ( .A(A[1287]), .B(n2809), .CI(
        C[1287]), .CO(C[1288]) );
  FA_6901 \FA_INST_0[2].FA_INST_1[264].FA_  ( .A(A[1288]), .B(n2808), .CI(
        C[1288]), .CO(C[1289]) );
  FA_6900 \FA_INST_0[2].FA_INST_1[265].FA_  ( .A(A[1289]), .B(n2807), .CI(
        C[1289]), .CO(C[1290]) );
  FA_6899 \FA_INST_0[2].FA_INST_1[266].FA_  ( .A(A[1290]), .B(n2806), .CI(
        C[1290]), .CO(C[1291]) );
  FA_6898 \FA_INST_0[2].FA_INST_1[267].FA_  ( .A(A[1291]), .B(n2805), .CI(
        C[1291]), .CO(C[1292]) );
  FA_6897 \FA_INST_0[2].FA_INST_1[268].FA_  ( .A(A[1292]), .B(n2804), .CI(
        C[1292]), .CO(C[1293]) );
  FA_6896 \FA_INST_0[2].FA_INST_1[269].FA_  ( .A(A[1293]), .B(n2803), .CI(
        C[1293]), .CO(C[1294]) );
  FA_6895 \FA_INST_0[2].FA_INST_1[270].FA_  ( .A(A[1294]), .B(n2802), .CI(
        C[1294]), .CO(C[1295]) );
  FA_6894 \FA_INST_0[2].FA_INST_1[271].FA_  ( .A(A[1295]), .B(n2801), .CI(
        C[1295]), .CO(C[1296]) );
  FA_6893 \FA_INST_0[2].FA_INST_1[272].FA_  ( .A(A[1296]), .B(n2800), .CI(
        C[1296]), .CO(C[1297]) );
  FA_6892 \FA_INST_0[2].FA_INST_1[273].FA_  ( .A(A[1297]), .B(n2799), .CI(
        C[1297]), .CO(C[1298]) );
  FA_6891 \FA_INST_0[2].FA_INST_1[274].FA_  ( .A(A[1298]), .B(n2798), .CI(
        C[1298]), .CO(C[1299]) );
  FA_6890 \FA_INST_0[2].FA_INST_1[275].FA_  ( .A(A[1299]), .B(n2797), .CI(
        C[1299]), .CO(C[1300]) );
  FA_6889 \FA_INST_0[2].FA_INST_1[276].FA_  ( .A(A[1300]), .B(n2796), .CI(
        C[1300]), .CO(C[1301]) );
  FA_6888 \FA_INST_0[2].FA_INST_1[277].FA_  ( .A(A[1301]), .B(n2795), .CI(
        C[1301]), .CO(C[1302]) );
  FA_6887 \FA_INST_0[2].FA_INST_1[278].FA_  ( .A(A[1302]), .B(n2794), .CI(
        C[1302]), .CO(C[1303]) );
  FA_6886 \FA_INST_0[2].FA_INST_1[279].FA_  ( .A(A[1303]), .B(n2793), .CI(
        C[1303]), .CO(C[1304]) );
  FA_6885 \FA_INST_0[2].FA_INST_1[280].FA_  ( .A(A[1304]), .B(n2792), .CI(
        C[1304]), .CO(C[1305]) );
  FA_6884 \FA_INST_0[2].FA_INST_1[281].FA_  ( .A(A[1305]), .B(n2791), .CI(
        C[1305]), .CO(C[1306]) );
  FA_6883 \FA_INST_0[2].FA_INST_1[282].FA_  ( .A(A[1306]), .B(n2790), .CI(
        C[1306]), .CO(C[1307]) );
  FA_6882 \FA_INST_0[2].FA_INST_1[283].FA_  ( .A(A[1307]), .B(n2789), .CI(
        C[1307]), .CO(C[1308]) );
  FA_6881 \FA_INST_0[2].FA_INST_1[284].FA_  ( .A(A[1308]), .B(n2788), .CI(
        C[1308]), .CO(C[1309]) );
  FA_6880 \FA_INST_0[2].FA_INST_1[285].FA_  ( .A(A[1309]), .B(n2787), .CI(
        C[1309]), .CO(C[1310]) );
  FA_6879 \FA_INST_0[2].FA_INST_1[286].FA_  ( .A(A[1310]), .B(n2786), .CI(
        C[1310]), .CO(C[1311]) );
  FA_6878 \FA_INST_0[2].FA_INST_1[287].FA_  ( .A(A[1311]), .B(n2785), .CI(
        C[1311]), .CO(C[1312]) );
  FA_6877 \FA_INST_0[2].FA_INST_1[288].FA_  ( .A(A[1312]), .B(n2784), .CI(
        C[1312]), .CO(C[1313]) );
  FA_6876 \FA_INST_0[2].FA_INST_1[289].FA_  ( .A(A[1313]), .B(n2783), .CI(
        C[1313]), .CO(C[1314]) );
  FA_6875 \FA_INST_0[2].FA_INST_1[290].FA_  ( .A(A[1314]), .B(n2782), .CI(
        C[1314]), .CO(C[1315]) );
  FA_6874 \FA_INST_0[2].FA_INST_1[291].FA_  ( .A(A[1315]), .B(n2781), .CI(
        C[1315]), .CO(C[1316]) );
  FA_6873 \FA_INST_0[2].FA_INST_1[292].FA_  ( .A(A[1316]), .B(n2780), .CI(
        C[1316]), .CO(C[1317]) );
  FA_6872 \FA_INST_0[2].FA_INST_1[293].FA_  ( .A(A[1317]), .B(n2779), .CI(
        C[1317]), .CO(C[1318]) );
  FA_6871 \FA_INST_0[2].FA_INST_1[294].FA_  ( .A(A[1318]), .B(n2778), .CI(
        C[1318]), .CO(C[1319]) );
  FA_6870 \FA_INST_0[2].FA_INST_1[295].FA_  ( .A(A[1319]), .B(n2777), .CI(
        C[1319]), .CO(C[1320]) );
  FA_6869 \FA_INST_0[2].FA_INST_1[296].FA_  ( .A(A[1320]), .B(n2776), .CI(
        C[1320]), .CO(C[1321]) );
  FA_6868 \FA_INST_0[2].FA_INST_1[297].FA_  ( .A(A[1321]), .B(n2775), .CI(
        C[1321]), .CO(C[1322]) );
  FA_6867 \FA_INST_0[2].FA_INST_1[298].FA_  ( .A(A[1322]), .B(n2774), .CI(
        C[1322]), .CO(C[1323]) );
  FA_6866 \FA_INST_0[2].FA_INST_1[299].FA_  ( .A(A[1323]), .B(n2773), .CI(
        C[1323]), .CO(C[1324]) );
  FA_6865 \FA_INST_0[2].FA_INST_1[300].FA_  ( .A(A[1324]), .B(n2772), .CI(
        C[1324]), .CO(C[1325]) );
  FA_6864 \FA_INST_0[2].FA_INST_1[301].FA_  ( .A(A[1325]), .B(n2771), .CI(
        C[1325]), .CO(C[1326]) );
  FA_6863 \FA_INST_0[2].FA_INST_1[302].FA_  ( .A(A[1326]), .B(n2770), .CI(
        C[1326]), .CO(C[1327]) );
  FA_6862 \FA_INST_0[2].FA_INST_1[303].FA_  ( .A(A[1327]), .B(n2769), .CI(
        C[1327]), .CO(C[1328]) );
  FA_6861 \FA_INST_0[2].FA_INST_1[304].FA_  ( .A(A[1328]), .B(n2768), .CI(
        C[1328]), .CO(C[1329]) );
  FA_6860 \FA_INST_0[2].FA_INST_1[305].FA_  ( .A(A[1329]), .B(n2767), .CI(
        C[1329]), .CO(C[1330]) );
  FA_6859 \FA_INST_0[2].FA_INST_1[306].FA_  ( .A(A[1330]), .B(n2766), .CI(
        C[1330]), .CO(C[1331]) );
  FA_6858 \FA_INST_0[2].FA_INST_1[307].FA_  ( .A(A[1331]), .B(n2765), .CI(
        C[1331]), .CO(C[1332]) );
  FA_6857 \FA_INST_0[2].FA_INST_1[308].FA_  ( .A(A[1332]), .B(n2764), .CI(
        C[1332]), .CO(C[1333]) );
  FA_6856 \FA_INST_0[2].FA_INST_1[309].FA_  ( .A(A[1333]), .B(n2763), .CI(
        C[1333]), .CO(C[1334]) );
  FA_6855 \FA_INST_0[2].FA_INST_1[310].FA_  ( .A(A[1334]), .B(n2762), .CI(
        C[1334]), .CO(C[1335]) );
  FA_6854 \FA_INST_0[2].FA_INST_1[311].FA_  ( .A(A[1335]), .B(n2761), .CI(
        C[1335]), .CO(C[1336]) );
  FA_6853 \FA_INST_0[2].FA_INST_1[312].FA_  ( .A(A[1336]), .B(n2760), .CI(
        C[1336]), .CO(C[1337]) );
  FA_6852 \FA_INST_0[2].FA_INST_1[313].FA_  ( .A(A[1337]), .B(n2759), .CI(
        C[1337]), .CO(C[1338]) );
  FA_6851 \FA_INST_0[2].FA_INST_1[314].FA_  ( .A(A[1338]), .B(n2758), .CI(
        C[1338]), .CO(C[1339]) );
  FA_6850 \FA_INST_0[2].FA_INST_1[315].FA_  ( .A(A[1339]), .B(n2757), .CI(
        C[1339]), .CO(C[1340]) );
  FA_6849 \FA_INST_0[2].FA_INST_1[316].FA_  ( .A(A[1340]), .B(n2756), .CI(
        C[1340]), .CO(C[1341]) );
  FA_6848 \FA_INST_0[2].FA_INST_1[317].FA_  ( .A(A[1341]), .B(n2755), .CI(
        C[1341]), .CO(C[1342]) );
  FA_6847 \FA_INST_0[2].FA_INST_1[318].FA_  ( .A(A[1342]), .B(n2754), .CI(
        C[1342]), .CO(C[1343]) );
  FA_6846 \FA_INST_0[2].FA_INST_1[319].FA_  ( .A(A[1343]), .B(n2753), .CI(
        C[1343]), .CO(C[1344]) );
  FA_6845 \FA_INST_0[2].FA_INST_1[320].FA_  ( .A(A[1344]), .B(n2752), .CI(
        C[1344]), .CO(C[1345]) );
  FA_6844 \FA_INST_0[2].FA_INST_1[321].FA_  ( .A(A[1345]), .B(n2751), .CI(
        C[1345]), .CO(C[1346]) );
  FA_6843 \FA_INST_0[2].FA_INST_1[322].FA_  ( .A(A[1346]), .B(n2750), .CI(
        C[1346]), .CO(C[1347]) );
  FA_6842 \FA_INST_0[2].FA_INST_1[323].FA_  ( .A(A[1347]), .B(n2749), .CI(
        C[1347]), .CO(C[1348]) );
  FA_6841 \FA_INST_0[2].FA_INST_1[324].FA_  ( .A(A[1348]), .B(n2748), .CI(
        C[1348]), .CO(C[1349]) );
  FA_6840 \FA_INST_0[2].FA_INST_1[325].FA_  ( .A(A[1349]), .B(n2747), .CI(
        C[1349]), .CO(C[1350]) );
  FA_6839 \FA_INST_0[2].FA_INST_1[326].FA_  ( .A(A[1350]), .B(n2746), .CI(
        C[1350]), .CO(C[1351]) );
  FA_6838 \FA_INST_0[2].FA_INST_1[327].FA_  ( .A(A[1351]), .B(n2745), .CI(
        C[1351]), .CO(C[1352]) );
  FA_6837 \FA_INST_0[2].FA_INST_1[328].FA_  ( .A(A[1352]), .B(n2744), .CI(
        C[1352]), .CO(C[1353]) );
  FA_6836 \FA_INST_0[2].FA_INST_1[329].FA_  ( .A(A[1353]), .B(n2743), .CI(
        C[1353]), .CO(C[1354]) );
  FA_6835 \FA_INST_0[2].FA_INST_1[330].FA_  ( .A(A[1354]), .B(n2742), .CI(
        C[1354]), .CO(C[1355]) );
  FA_6834 \FA_INST_0[2].FA_INST_1[331].FA_  ( .A(A[1355]), .B(n2741), .CI(
        C[1355]), .CO(C[1356]) );
  FA_6833 \FA_INST_0[2].FA_INST_1[332].FA_  ( .A(A[1356]), .B(n2740), .CI(
        C[1356]), .CO(C[1357]) );
  FA_6832 \FA_INST_0[2].FA_INST_1[333].FA_  ( .A(A[1357]), .B(n2739), .CI(
        C[1357]), .CO(C[1358]) );
  FA_6831 \FA_INST_0[2].FA_INST_1[334].FA_  ( .A(A[1358]), .B(n2738), .CI(
        C[1358]), .CO(C[1359]) );
  FA_6830 \FA_INST_0[2].FA_INST_1[335].FA_  ( .A(A[1359]), .B(n2737), .CI(
        C[1359]), .CO(C[1360]) );
  FA_6829 \FA_INST_0[2].FA_INST_1[336].FA_  ( .A(A[1360]), .B(n2736), .CI(
        C[1360]), .CO(C[1361]) );
  FA_6828 \FA_INST_0[2].FA_INST_1[337].FA_  ( .A(A[1361]), .B(n2735), .CI(
        C[1361]), .CO(C[1362]) );
  FA_6827 \FA_INST_0[2].FA_INST_1[338].FA_  ( .A(A[1362]), .B(n2734), .CI(
        C[1362]), .CO(C[1363]) );
  FA_6826 \FA_INST_0[2].FA_INST_1[339].FA_  ( .A(A[1363]), .B(n2733), .CI(
        C[1363]), .CO(C[1364]) );
  FA_6825 \FA_INST_0[2].FA_INST_1[340].FA_  ( .A(A[1364]), .B(n2732), .CI(
        C[1364]), .CO(C[1365]) );
  FA_6824 \FA_INST_0[2].FA_INST_1[341].FA_  ( .A(A[1365]), .B(n2731), .CI(
        C[1365]), .CO(C[1366]) );
  FA_6823 \FA_INST_0[2].FA_INST_1[342].FA_  ( .A(A[1366]), .B(n2730), .CI(
        C[1366]), .CO(C[1367]) );
  FA_6822 \FA_INST_0[2].FA_INST_1[343].FA_  ( .A(A[1367]), .B(n2729), .CI(
        C[1367]), .CO(C[1368]) );
  FA_6821 \FA_INST_0[2].FA_INST_1[344].FA_  ( .A(A[1368]), .B(n2728), .CI(
        C[1368]), .CO(C[1369]) );
  FA_6820 \FA_INST_0[2].FA_INST_1[345].FA_  ( .A(A[1369]), .B(n2727), .CI(
        C[1369]), .CO(C[1370]) );
  FA_6819 \FA_INST_0[2].FA_INST_1[346].FA_  ( .A(A[1370]), .B(n2726), .CI(
        C[1370]), .CO(C[1371]) );
  FA_6818 \FA_INST_0[2].FA_INST_1[347].FA_  ( .A(A[1371]), .B(n2725), .CI(
        C[1371]), .CO(C[1372]) );
  FA_6817 \FA_INST_0[2].FA_INST_1[348].FA_  ( .A(A[1372]), .B(n2724), .CI(
        C[1372]), .CO(C[1373]) );
  FA_6816 \FA_INST_0[2].FA_INST_1[349].FA_  ( .A(A[1373]), .B(n2723), .CI(
        C[1373]), .CO(C[1374]) );
  FA_6815 \FA_INST_0[2].FA_INST_1[350].FA_  ( .A(A[1374]), .B(n2722), .CI(
        C[1374]), .CO(C[1375]) );
  FA_6814 \FA_INST_0[2].FA_INST_1[351].FA_  ( .A(A[1375]), .B(n2721), .CI(
        C[1375]), .CO(C[1376]) );
  FA_6813 \FA_INST_0[2].FA_INST_1[352].FA_  ( .A(A[1376]), .B(n2720), .CI(
        C[1376]), .CO(C[1377]) );
  FA_6812 \FA_INST_0[2].FA_INST_1[353].FA_  ( .A(A[1377]), .B(n2719), .CI(
        C[1377]), .CO(C[1378]) );
  FA_6811 \FA_INST_0[2].FA_INST_1[354].FA_  ( .A(A[1378]), .B(n2718), .CI(
        C[1378]), .CO(C[1379]) );
  FA_6810 \FA_INST_0[2].FA_INST_1[355].FA_  ( .A(A[1379]), .B(n2717), .CI(
        C[1379]), .CO(C[1380]) );
  FA_6809 \FA_INST_0[2].FA_INST_1[356].FA_  ( .A(A[1380]), .B(n2716), .CI(
        C[1380]), .CO(C[1381]) );
  FA_6808 \FA_INST_0[2].FA_INST_1[357].FA_  ( .A(A[1381]), .B(n2715), .CI(
        C[1381]), .CO(C[1382]) );
  FA_6807 \FA_INST_0[2].FA_INST_1[358].FA_  ( .A(A[1382]), .B(n2714), .CI(
        C[1382]), .CO(C[1383]) );
  FA_6806 \FA_INST_0[2].FA_INST_1[359].FA_  ( .A(A[1383]), .B(n2713), .CI(
        C[1383]), .CO(C[1384]) );
  FA_6805 \FA_INST_0[2].FA_INST_1[360].FA_  ( .A(A[1384]), .B(n2712), .CI(
        C[1384]), .CO(C[1385]) );
  FA_6804 \FA_INST_0[2].FA_INST_1[361].FA_  ( .A(A[1385]), .B(n2711), .CI(
        C[1385]), .CO(C[1386]) );
  FA_6803 \FA_INST_0[2].FA_INST_1[362].FA_  ( .A(A[1386]), .B(n2710), .CI(
        C[1386]), .CO(C[1387]) );
  FA_6802 \FA_INST_0[2].FA_INST_1[363].FA_  ( .A(A[1387]), .B(n2709), .CI(
        C[1387]), .CO(C[1388]) );
  FA_6801 \FA_INST_0[2].FA_INST_1[364].FA_  ( .A(A[1388]), .B(n2708), .CI(
        C[1388]), .CO(C[1389]) );
  FA_6800 \FA_INST_0[2].FA_INST_1[365].FA_  ( .A(A[1389]), .B(n2707), .CI(
        C[1389]), .CO(C[1390]) );
  FA_6799 \FA_INST_0[2].FA_INST_1[366].FA_  ( .A(A[1390]), .B(n2706), .CI(
        C[1390]), .CO(C[1391]) );
  FA_6798 \FA_INST_0[2].FA_INST_1[367].FA_  ( .A(A[1391]), .B(n2705), .CI(
        C[1391]), .CO(C[1392]) );
  FA_6797 \FA_INST_0[2].FA_INST_1[368].FA_  ( .A(A[1392]), .B(n2704), .CI(
        C[1392]), .CO(C[1393]) );
  FA_6796 \FA_INST_0[2].FA_INST_1[369].FA_  ( .A(A[1393]), .B(n2703), .CI(
        C[1393]), .CO(C[1394]) );
  FA_6795 \FA_INST_0[2].FA_INST_1[370].FA_  ( .A(A[1394]), .B(n2702), .CI(
        C[1394]), .CO(C[1395]) );
  FA_6794 \FA_INST_0[2].FA_INST_1[371].FA_  ( .A(A[1395]), .B(n2701), .CI(
        C[1395]), .CO(C[1396]) );
  FA_6793 \FA_INST_0[2].FA_INST_1[372].FA_  ( .A(A[1396]), .B(n2700), .CI(
        C[1396]), .CO(C[1397]) );
  FA_6792 \FA_INST_0[2].FA_INST_1[373].FA_  ( .A(A[1397]), .B(n2699), .CI(
        C[1397]), .CO(C[1398]) );
  FA_6791 \FA_INST_0[2].FA_INST_1[374].FA_  ( .A(A[1398]), .B(n2698), .CI(
        C[1398]), .CO(C[1399]) );
  FA_6790 \FA_INST_0[2].FA_INST_1[375].FA_  ( .A(A[1399]), .B(n2697), .CI(
        C[1399]), .CO(C[1400]) );
  FA_6789 \FA_INST_0[2].FA_INST_1[376].FA_  ( .A(A[1400]), .B(n2696), .CI(
        C[1400]), .CO(C[1401]) );
  FA_6788 \FA_INST_0[2].FA_INST_1[377].FA_  ( .A(A[1401]), .B(n2695), .CI(
        C[1401]), .CO(C[1402]) );
  FA_6787 \FA_INST_0[2].FA_INST_1[378].FA_  ( .A(A[1402]), .B(n2694), .CI(
        C[1402]), .CO(C[1403]) );
  FA_6786 \FA_INST_0[2].FA_INST_1[379].FA_  ( .A(A[1403]), .B(n2693), .CI(
        C[1403]), .CO(C[1404]) );
  FA_6785 \FA_INST_0[2].FA_INST_1[380].FA_  ( .A(A[1404]), .B(n2692), .CI(
        C[1404]), .CO(C[1405]) );
  FA_6784 \FA_INST_0[2].FA_INST_1[381].FA_  ( .A(A[1405]), .B(n2691), .CI(
        C[1405]), .CO(C[1406]) );
  FA_6783 \FA_INST_0[2].FA_INST_1[382].FA_  ( .A(A[1406]), .B(n2690), .CI(
        C[1406]), .CO(C[1407]) );
  FA_6782 \FA_INST_0[2].FA_INST_1[383].FA_  ( .A(A[1407]), .B(n2689), .CI(
        C[1407]), .CO(C[1408]) );
  FA_6781 \FA_INST_0[2].FA_INST_1[384].FA_  ( .A(A[1408]), .B(n2688), .CI(
        C[1408]), .CO(C[1409]) );
  FA_6780 \FA_INST_0[2].FA_INST_1[385].FA_  ( .A(A[1409]), .B(n2687), .CI(
        C[1409]), .CO(C[1410]) );
  FA_6779 \FA_INST_0[2].FA_INST_1[386].FA_  ( .A(A[1410]), .B(n2686), .CI(
        C[1410]), .CO(C[1411]) );
  FA_6778 \FA_INST_0[2].FA_INST_1[387].FA_  ( .A(A[1411]), .B(n2685), .CI(
        C[1411]), .CO(C[1412]) );
  FA_6777 \FA_INST_0[2].FA_INST_1[388].FA_  ( .A(A[1412]), .B(n2684), .CI(
        C[1412]), .CO(C[1413]) );
  FA_6776 \FA_INST_0[2].FA_INST_1[389].FA_  ( .A(A[1413]), .B(n2683), .CI(
        C[1413]), .CO(C[1414]) );
  FA_6775 \FA_INST_0[2].FA_INST_1[390].FA_  ( .A(A[1414]), .B(n2682), .CI(
        C[1414]), .CO(C[1415]) );
  FA_6774 \FA_INST_0[2].FA_INST_1[391].FA_  ( .A(A[1415]), .B(n2681), .CI(
        C[1415]), .CO(C[1416]) );
  FA_6773 \FA_INST_0[2].FA_INST_1[392].FA_  ( .A(A[1416]), .B(n2680), .CI(
        C[1416]), .CO(C[1417]) );
  FA_6772 \FA_INST_0[2].FA_INST_1[393].FA_  ( .A(A[1417]), .B(n2679), .CI(
        C[1417]), .CO(C[1418]) );
  FA_6771 \FA_INST_0[2].FA_INST_1[394].FA_  ( .A(A[1418]), .B(n2678), .CI(
        C[1418]), .CO(C[1419]) );
  FA_6770 \FA_INST_0[2].FA_INST_1[395].FA_  ( .A(A[1419]), .B(n2677), .CI(
        C[1419]), .CO(C[1420]) );
  FA_6769 \FA_INST_0[2].FA_INST_1[396].FA_  ( .A(A[1420]), .B(n2676), .CI(
        C[1420]), .CO(C[1421]) );
  FA_6768 \FA_INST_0[2].FA_INST_1[397].FA_  ( .A(A[1421]), .B(n2675), .CI(
        C[1421]), .CO(C[1422]) );
  FA_6767 \FA_INST_0[2].FA_INST_1[398].FA_  ( .A(A[1422]), .B(n2674), .CI(
        C[1422]), .CO(C[1423]) );
  FA_6766 \FA_INST_0[2].FA_INST_1[399].FA_  ( .A(A[1423]), .B(n2673), .CI(
        C[1423]), .CO(C[1424]) );
  FA_6765 \FA_INST_0[2].FA_INST_1[400].FA_  ( .A(A[1424]), .B(n2672), .CI(
        C[1424]), .CO(C[1425]) );
  FA_6764 \FA_INST_0[2].FA_INST_1[401].FA_  ( .A(A[1425]), .B(n2671), .CI(
        C[1425]), .CO(C[1426]) );
  FA_6763 \FA_INST_0[2].FA_INST_1[402].FA_  ( .A(A[1426]), .B(n2670), .CI(
        C[1426]), .CO(C[1427]) );
  FA_6762 \FA_INST_0[2].FA_INST_1[403].FA_  ( .A(A[1427]), .B(n2669), .CI(
        C[1427]), .CO(C[1428]) );
  FA_6761 \FA_INST_0[2].FA_INST_1[404].FA_  ( .A(A[1428]), .B(n2668), .CI(
        C[1428]), .CO(C[1429]) );
  FA_6760 \FA_INST_0[2].FA_INST_1[405].FA_  ( .A(A[1429]), .B(n2667), .CI(
        C[1429]), .CO(C[1430]) );
  FA_6759 \FA_INST_0[2].FA_INST_1[406].FA_  ( .A(A[1430]), .B(n2666), .CI(
        C[1430]), .CO(C[1431]) );
  FA_6758 \FA_INST_0[2].FA_INST_1[407].FA_  ( .A(A[1431]), .B(n2665), .CI(
        C[1431]), .CO(C[1432]) );
  FA_6757 \FA_INST_0[2].FA_INST_1[408].FA_  ( .A(A[1432]), .B(n2664), .CI(
        C[1432]), .CO(C[1433]) );
  FA_6756 \FA_INST_0[2].FA_INST_1[409].FA_  ( .A(A[1433]), .B(n2663), .CI(
        C[1433]), .CO(C[1434]) );
  FA_6755 \FA_INST_0[2].FA_INST_1[410].FA_  ( .A(A[1434]), .B(n2662), .CI(
        C[1434]), .CO(C[1435]) );
  FA_6754 \FA_INST_0[2].FA_INST_1[411].FA_  ( .A(A[1435]), .B(n2661), .CI(
        C[1435]), .CO(C[1436]) );
  FA_6753 \FA_INST_0[2].FA_INST_1[412].FA_  ( .A(A[1436]), .B(n2660), .CI(
        C[1436]), .CO(C[1437]) );
  FA_6752 \FA_INST_0[2].FA_INST_1[413].FA_  ( .A(A[1437]), .B(n2659), .CI(
        C[1437]), .CO(C[1438]) );
  FA_6751 \FA_INST_0[2].FA_INST_1[414].FA_  ( .A(A[1438]), .B(n2658), .CI(
        C[1438]), .CO(C[1439]) );
  FA_6750 \FA_INST_0[2].FA_INST_1[415].FA_  ( .A(A[1439]), .B(n2657), .CI(
        C[1439]), .CO(C[1440]) );
  FA_6749 \FA_INST_0[2].FA_INST_1[416].FA_  ( .A(A[1440]), .B(n2656), .CI(
        C[1440]), .CO(C[1441]) );
  FA_6748 \FA_INST_0[2].FA_INST_1[417].FA_  ( .A(A[1441]), .B(n2655), .CI(
        C[1441]), .CO(C[1442]) );
  FA_6747 \FA_INST_0[2].FA_INST_1[418].FA_  ( .A(A[1442]), .B(n2654), .CI(
        C[1442]), .CO(C[1443]) );
  FA_6746 \FA_INST_0[2].FA_INST_1[419].FA_  ( .A(A[1443]), .B(n2653), .CI(
        C[1443]), .CO(C[1444]) );
  FA_6745 \FA_INST_0[2].FA_INST_1[420].FA_  ( .A(A[1444]), .B(n2652), .CI(
        C[1444]), .CO(C[1445]) );
  FA_6744 \FA_INST_0[2].FA_INST_1[421].FA_  ( .A(A[1445]), .B(n2651), .CI(
        C[1445]), .CO(C[1446]) );
  FA_6743 \FA_INST_0[2].FA_INST_1[422].FA_  ( .A(A[1446]), .B(n2650), .CI(
        C[1446]), .CO(C[1447]) );
  FA_6742 \FA_INST_0[2].FA_INST_1[423].FA_  ( .A(A[1447]), .B(n2649), .CI(
        C[1447]), .CO(C[1448]) );
  FA_6741 \FA_INST_0[2].FA_INST_1[424].FA_  ( .A(A[1448]), .B(n2648), .CI(
        C[1448]), .CO(C[1449]) );
  FA_6740 \FA_INST_0[2].FA_INST_1[425].FA_  ( .A(A[1449]), .B(n2647), .CI(
        C[1449]), .CO(C[1450]) );
  FA_6739 \FA_INST_0[2].FA_INST_1[426].FA_  ( .A(A[1450]), .B(n2646), .CI(
        C[1450]), .CO(C[1451]) );
  FA_6738 \FA_INST_0[2].FA_INST_1[427].FA_  ( .A(A[1451]), .B(n2645), .CI(
        C[1451]), .CO(C[1452]) );
  FA_6737 \FA_INST_0[2].FA_INST_1[428].FA_  ( .A(A[1452]), .B(n2644), .CI(
        C[1452]), .CO(C[1453]) );
  FA_6736 \FA_INST_0[2].FA_INST_1[429].FA_  ( .A(A[1453]), .B(n2643), .CI(
        C[1453]), .CO(C[1454]) );
  FA_6735 \FA_INST_0[2].FA_INST_1[430].FA_  ( .A(A[1454]), .B(n2642), .CI(
        C[1454]), .CO(C[1455]) );
  FA_6734 \FA_INST_0[2].FA_INST_1[431].FA_  ( .A(A[1455]), .B(n2641), .CI(
        C[1455]), .CO(C[1456]) );
  FA_6733 \FA_INST_0[2].FA_INST_1[432].FA_  ( .A(A[1456]), .B(n2640), .CI(
        C[1456]), .CO(C[1457]) );
  FA_6732 \FA_INST_0[2].FA_INST_1[433].FA_  ( .A(A[1457]), .B(n2639), .CI(
        C[1457]), .CO(C[1458]) );
  FA_6731 \FA_INST_0[2].FA_INST_1[434].FA_  ( .A(A[1458]), .B(n2638), .CI(
        C[1458]), .CO(C[1459]) );
  FA_6730 \FA_INST_0[2].FA_INST_1[435].FA_  ( .A(A[1459]), .B(n2637), .CI(
        C[1459]), .CO(C[1460]) );
  FA_6729 \FA_INST_0[2].FA_INST_1[436].FA_  ( .A(A[1460]), .B(n2636), .CI(
        C[1460]), .CO(C[1461]) );
  FA_6728 \FA_INST_0[2].FA_INST_1[437].FA_  ( .A(A[1461]), .B(n2635), .CI(
        C[1461]), .CO(C[1462]) );
  FA_6727 \FA_INST_0[2].FA_INST_1[438].FA_  ( .A(A[1462]), .B(n2634), .CI(
        C[1462]), .CO(C[1463]) );
  FA_6726 \FA_INST_0[2].FA_INST_1[439].FA_  ( .A(A[1463]), .B(n2633), .CI(
        C[1463]), .CO(C[1464]) );
  FA_6725 \FA_INST_0[2].FA_INST_1[440].FA_  ( .A(A[1464]), .B(n2632), .CI(
        C[1464]), .CO(C[1465]) );
  FA_6724 \FA_INST_0[2].FA_INST_1[441].FA_  ( .A(A[1465]), .B(n2631), .CI(
        C[1465]), .CO(C[1466]) );
  FA_6723 \FA_INST_0[2].FA_INST_1[442].FA_  ( .A(A[1466]), .B(n2630), .CI(
        C[1466]), .CO(C[1467]) );
  FA_6722 \FA_INST_0[2].FA_INST_1[443].FA_  ( .A(A[1467]), .B(n2629), .CI(
        C[1467]), .CO(C[1468]) );
  FA_6721 \FA_INST_0[2].FA_INST_1[444].FA_  ( .A(A[1468]), .B(n2628), .CI(
        C[1468]), .CO(C[1469]) );
  FA_6720 \FA_INST_0[2].FA_INST_1[445].FA_  ( .A(A[1469]), .B(n2627), .CI(
        C[1469]), .CO(C[1470]) );
  FA_6719 \FA_INST_0[2].FA_INST_1[446].FA_  ( .A(A[1470]), .B(n2626), .CI(
        C[1470]), .CO(C[1471]) );
  FA_6718 \FA_INST_0[2].FA_INST_1[447].FA_  ( .A(A[1471]), .B(n2625), .CI(
        C[1471]), .CO(C[1472]) );
  FA_6717 \FA_INST_0[2].FA_INST_1[448].FA_  ( .A(A[1472]), .B(n2624), .CI(
        C[1472]), .CO(C[1473]) );
  FA_6716 \FA_INST_0[2].FA_INST_1[449].FA_  ( .A(A[1473]), .B(n2623), .CI(
        C[1473]), .CO(C[1474]) );
  FA_6715 \FA_INST_0[2].FA_INST_1[450].FA_  ( .A(A[1474]), .B(n2622), .CI(
        C[1474]), .CO(C[1475]) );
  FA_6714 \FA_INST_0[2].FA_INST_1[451].FA_  ( .A(A[1475]), .B(n2621), .CI(
        C[1475]), .CO(C[1476]) );
  FA_6713 \FA_INST_0[2].FA_INST_1[452].FA_  ( .A(A[1476]), .B(n2620), .CI(
        C[1476]), .CO(C[1477]) );
  FA_6712 \FA_INST_0[2].FA_INST_1[453].FA_  ( .A(A[1477]), .B(n2619), .CI(
        C[1477]), .CO(C[1478]) );
  FA_6711 \FA_INST_0[2].FA_INST_1[454].FA_  ( .A(A[1478]), .B(n2618), .CI(
        C[1478]), .CO(C[1479]) );
  FA_6710 \FA_INST_0[2].FA_INST_1[455].FA_  ( .A(A[1479]), .B(n2617), .CI(
        C[1479]), .CO(C[1480]) );
  FA_6709 \FA_INST_0[2].FA_INST_1[456].FA_  ( .A(A[1480]), .B(n2616), .CI(
        C[1480]), .CO(C[1481]) );
  FA_6708 \FA_INST_0[2].FA_INST_1[457].FA_  ( .A(A[1481]), .B(n2615), .CI(
        C[1481]), .CO(C[1482]) );
  FA_6707 \FA_INST_0[2].FA_INST_1[458].FA_  ( .A(A[1482]), .B(n2614), .CI(
        C[1482]), .CO(C[1483]) );
  FA_6706 \FA_INST_0[2].FA_INST_1[459].FA_  ( .A(A[1483]), .B(n2613), .CI(
        C[1483]), .CO(C[1484]) );
  FA_6705 \FA_INST_0[2].FA_INST_1[460].FA_  ( .A(A[1484]), .B(n2612), .CI(
        C[1484]), .CO(C[1485]) );
  FA_6704 \FA_INST_0[2].FA_INST_1[461].FA_  ( .A(A[1485]), .B(n2611), .CI(
        C[1485]), .CO(C[1486]) );
  FA_6703 \FA_INST_0[2].FA_INST_1[462].FA_  ( .A(A[1486]), .B(n2610), .CI(
        C[1486]), .CO(C[1487]) );
  FA_6702 \FA_INST_0[2].FA_INST_1[463].FA_  ( .A(A[1487]), .B(n2609), .CI(
        C[1487]), .CO(C[1488]) );
  FA_6701 \FA_INST_0[2].FA_INST_1[464].FA_  ( .A(A[1488]), .B(n2608), .CI(
        C[1488]), .CO(C[1489]) );
  FA_6700 \FA_INST_0[2].FA_INST_1[465].FA_  ( .A(A[1489]), .B(n2607), .CI(
        C[1489]), .CO(C[1490]) );
  FA_6699 \FA_INST_0[2].FA_INST_1[466].FA_  ( .A(A[1490]), .B(n2606), .CI(
        C[1490]), .CO(C[1491]) );
  FA_6698 \FA_INST_0[2].FA_INST_1[467].FA_  ( .A(A[1491]), .B(n2605), .CI(
        C[1491]), .CO(C[1492]) );
  FA_6697 \FA_INST_0[2].FA_INST_1[468].FA_  ( .A(A[1492]), .B(n2604), .CI(
        C[1492]), .CO(C[1493]) );
  FA_6696 \FA_INST_0[2].FA_INST_1[469].FA_  ( .A(A[1493]), .B(n2603), .CI(
        C[1493]), .CO(C[1494]) );
  FA_6695 \FA_INST_0[2].FA_INST_1[470].FA_  ( .A(A[1494]), .B(n2602), .CI(
        C[1494]), .CO(C[1495]) );
  FA_6694 \FA_INST_0[2].FA_INST_1[471].FA_  ( .A(A[1495]), .B(n2601), .CI(
        C[1495]), .CO(C[1496]) );
  FA_6693 \FA_INST_0[2].FA_INST_1[472].FA_  ( .A(A[1496]), .B(n2600), .CI(
        C[1496]), .CO(C[1497]) );
  FA_6692 \FA_INST_0[2].FA_INST_1[473].FA_  ( .A(A[1497]), .B(n2599), .CI(
        C[1497]), .CO(C[1498]) );
  FA_6691 \FA_INST_0[2].FA_INST_1[474].FA_  ( .A(A[1498]), .B(n2598), .CI(
        C[1498]), .CO(C[1499]) );
  FA_6690 \FA_INST_0[2].FA_INST_1[475].FA_  ( .A(A[1499]), .B(n2597), .CI(
        C[1499]), .CO(C[1500]) );
  FA_6689 \FA_INST_0[2].FA_INST_1[476].FA_  ( .A(A[1500]), .B(n2596), .CI(
        C[1500]), .CO(C[1501]) );
  FA_6688 \FA_INST_0[2].FA_INST_1[477].FA_  ( .A(A[1501]), .B(n2595), .CI(
        C[1501]), .CO(C[1502]) );
  FA_6687 \FA_INST_0[2].FA_INST_1[478].FA_  ( .A(A[1502]), .B(n2594), .CI(
        C[1502]), .CO(C[1503]) );
  FA_6686 \FA_INST_0[2].FA_INST_1[479].FA_  ( .A(A[1503]), .B(n2593), .CI(
        C[1503]), .CO(C[1504]) );
  FA_6685 \FA_INST_0[2].FA_INST_1[480].FA_  ( .A(A[1504]), .B(n2592), .CI(
        C[1504]), .CO(C[1505]) );
  FA_6684 \FA_INST_0[2].FA_INST_1[481].FA_  ( .A(A[1505]), .B(n2591), .CI(
        C[1505]), .CO(C[1506]) );
  FA_6683 \FA_INST_0[2].FA_INST_1[482].FA_  ( .A(A[1506]), .B(n2590), .CI(
        C[1506]), .CO(C[1507]) );
  FA_6682 \FA_INST_0[2].FA_INST_1[483].FA_  ( .A(A[1507]), .B(n2589), .CI(
        C[1507]), .CO(C[1508]) );
  FA_6681 \FA_INST_0[2].FA_INST_1[484].FA_  ( .A(A[1508]), .B(n2588), .CI(
        C[1508]), .CO(C[1509]) );
  FA_6680 \FA_INST_0[2].FA_INST_1[485].FA_  ( .A(A[1509]), .B(n2587), .CI(
        C[1509]), .CO(C[1510]) );
  FA_6679 \FA_INST_0[2].FA_INST_1[486].FA_  ( .A(A[1510]), .B(n2586), .CI(
        C[1510]), .CO(C[1511]) );
  FA_6678 \FA_INST_0[2].FA_INST_1[487].FA_  ( .A(A[1511]), .B(n2585), .CI(
        C[1511]), .CO(C[1512]) );
  FA_6677 \FA_INST_0[2].FA_INST_1[488].FA_  ( .A(A[1512]), .B(n2584), .CI(
        C[1512]), .CO(C[1513]) );
  FA_6676 \FA_INST_0[2].FA_INST_1[489].FA_  ( .A(A[1513]), .B(n2583), .CI(
        C[1513]), .CO(C[1514]) );
  FA_6675 \FA_INST_0[2].FA_INST_1[490].FA_  ( .A(A[1514]), .B(n2582), .CI(
        C[1514]), .CO(C[1515]) );
  FA_6674 \FA_INST_0[2].FA_INST_1[491].FA_  ( .A(A[1515]), .B(n2581), .CI(
        C[1515]), .CO(C[1516]) );
  FA_6673 \FA_INST_0[2].FA_INST_1[492].FA_  ( .A(A[1516]), .B(n2580), .CI(
        C[1516]), .CO(C[1517]) );
  FA_6672 \FA_INST_0[2].FA_INST_1[493].FA_  ( .A(A[1517]), .B(n2579), .CI(
        C[1517]), .CO(C[1518]) );
  FA_6671 \FA_INST_0[2].FA_INST_1[494].FA_  ( .A(A[1518]), .B(n2578), .CI(
        C[1518]), .CO(C[1519]) );
  FA_6670 \FA_INST_0[2].FA_INST_1[495].FA_  ( .A(A[1519]), .B(n2577), .CI(
        C[1519]), .CO(C[1520]) );
  FA_6669 \FA_INST_0[2].FA_INST_1[496].FA_  ( .A(A[1520]), .B(n2576), .CI(
        C[1520]), .CO(C[1521]) );
  FA_6668 \FA_INST_0[2].FA_INST_1[497].FA_  ( .A(A[1521]), .B(n2575), .CI(
        C[1521]), .CO(C[1522]) );
  FA_6667 \FA_INST_0[2].FA_INST_1[498].FA_  ( .A(A[1522]), .B(n2574), .CI(
        C[1522]), .CO(C[1523]) );
  FA_6666 \FA_INST_0[2].FA_INST_1[499].FA_  ( .A(A[1523]), .B(n2573), .CI(
        C[1523]), .CO(C[1524]) );
  FA_6665 \FA_INST_0[2].FA_INST_1[500].FA_  ( .A(A[1524]), .B(n2572), .CI(
        C[1524]), .CO(C[1525]) );
  FA_6664 \FA_INST_0[2].FA_INST_1[501].FA_  ( .A(A[1525]), .B(n2571), .CI(
        C[1525]), .CO(C[1526]) );
  FA_6663 \FA_INST_0[2].FA_INST_1[502].FA_  ( .A(A[1526]), .B(n2570), .CI(
        C[1526]), .CO(C[1527]) );
  FA_6662 \FA_INST_0[2].FA_INST_1[503].FA_  ( .A(A[1527]), .B(n2569), .CI(
        C[1527]), .CO(C[1528]) );
  FA_6661 \FA_INST_0[2].FA_INST_1[504].FA_  ( .A(A[1528]), .B(n2568), .CI(
        C[1528]), .CO(C[1529]) );
  FA_6660 \FA_INST_0[2].FA_INST_1[505].FA_  ( .A(A[1529]), .B(n2567), .CI(
        C[1529]), .CO(C[1530]) );
  FA_6659 \FA_INST_0[2].FA_INST_1[506].FA_  ( .A(A[1530]), .B(n2566), .CI(
        C[1530]), .CO(C[1531]) );
  FA_6658 \FA_INST_0[2].FA_INST_1[507].FA_  ( .A(A[1531]), .B(n2565), .CI(
        C[1531]), .CO(C[1532]) );
  FA_6657 \FA_INST_0[2].FA_INST_1[508].FA_  ( .A(A[1532]), .B(n2564), .CI(
        C[1532]), .CO(C[1533]) );
  FA_6656 \FA_INST_0[2].FA_INST_1[509].FA_  ( .A(A[1533]), .B(n2563), .CI(
        C[1533]), .CO(C[1534]) );
  FA_6655 \FA_INST_0[2].FA_INST_1[510].FA_  ( .A(A[1534]), .B(n2562), .CI(
        C[1534]), .CO(C[1535]) );
  FA_6654 \FA_INST_0[2].FA_INST_1[511].FA_  ( .A(A[1535]), .B(n2561), .CI(
        C[1535]), .CO(C[1536]) );
  FA_6653 \FA_INST_0[3].FA_INST_1[0].FA_  ( .A(A[1536]), .B(n2560), .CI(
        C[1536]), .CO(C[1537]) );
  FA_6652 \FA_INST_0[3].FA_INST_1[1].FA_  ( .A(A[1537]), .B(n2559), .CI(
        C[1537]), .CO(C[1538]) );
  FA_6651 \FA_INST_0[3].FA_INST_1[2].FA_  ( .A(A[1538]), .B(n2558), .CI(
        C[1538]), .CO(C[1539]) );
  FA_6650 \FA_INST_0[3].FA_INST_1[3].FA_  ( .A(A[1539]), .B(n2557), .CI(
        C[1539]), .CO(C[1540]) );
  FA_6649 \FA_INST_0[3].FA_INST_1[4].FA_  ( .A(A[1540]), .B(n2556), .CI(
        C[1540]), .CO(C[1541]) );
  FA_6648 \FA_INST_0[3].FA_INST_1[5].FA_  ( .A(A[1541]), .B(n2555), .CI(
        C[1541]), .CO(C[1542]) );
  FA_6647 \FA_INST_0[3].FA_INST_1[6].FA_  ( .A(A[1542]), .B(n2554), .CI(
        C[1542]), .CO(C[1543]) );
  FA_6646 \FA_INST_0[3].FA_INST_1[7].FA_  ( .A(A[1543]), .B(n2553), .CI(
        C[1543]), .CO(C[1544]) );
  FA_6645 \FA_INST_0[3].FA_INST_1[8].FA_  ( .A(A[1544]), .B(n2552), .CI(
        C[1544]), .CO(C[1545]) );
  FA_6644 \FA_INST_0[3].FA_INST_1[9].FA_  ( .A(A[1545]), .B(n2551), .CI(
        C[1545]), .CO(C[1546]) );
  FA_6643 \FA_INST_0[3].FA_INST_1[10].FA_  ( .A(A[1546]), .B(n2550), .CI(
        C[1546]), .CO(C[1547]) );
  FA_6642 \FA_INST_0[3].FA_INST_1[11].FA_  ( .A(A[1547]), .B(n2549), .CI(
        C[1547]), .CO(C[1548]) );
  FA_6641 \FA_INST_0[3].FA_INST_1[12].FA_  ( .A(A[1548]), .B(n2548), .CI(
        C[1548]), .CO(C[1549]) );
  FA_6640 \FA_INST_0[3].FA_INST_1[13].FA_  ( .A(A[1549]), .B(n2547), .CI(
        C[1549]), .CO(C[1550]) );
  FA_6639 \FA_INST_0[3].FA_INST_1[14].FA_  ( .A(A[1550]), .B(n2546), .CI(
        C[1550]), .CO(C[1551]) );
  FA_6638 \FA_INST_0[3].FA_INST_1[15].FA_  ( .A(A[1551]), .B(n2545), .CI(
        C[1551]), .CO(C[1552]) );
  FA_6637 \FA_INST_0[3].FA_INST_1[16].FA_  ( .A(A[1552]), .B(n2544), .CI(
        C[1552]), .CO(C[1553]) );
  FA_6636 \FA_INST_0[3].FA_INST_1[17].FA_  ( .A(A[1553]), .B(n2543), .CI(
        C[1553]), .CO(C[1554]) );
  FA_6635 \FA_INST_0[3].FA_INST_1[18].FA_  ( .A(A[1554]), .B(n2542), .CI(
        C[1554]), .CO(C[1555]) );
  FA_6634 \FA_INST_0[3].FA_INST_1[19].FA_  ( .A(A[1555]), .B(n2541), .CI(
        C[1555]), .CO(C[1556]) );
  FA_6633 \FA_INST_0[3].FA_INST_1[20].FA_  ( .A(A[1556]), .B(n2540), .CI(
        C[1556]), .CO(C[1557]) );
  FA_6632 \FA_INST_0[3].FA_INST_1[21].FA_  ( .A(A[1557]), .B(n2539), .CI(
        C[1557]), .CO(C[1558]) );
  FA_6631 \FA_INST_0[3].FA_INST_1[22].FA_  ( .A(A[1558]), .B(n2538), .CI(
        C[1558]), .CO(C[1559]) );
  FA_6630 \FA_INST_0[3].FA_INST_1[23].FA_  ( .A(A[1559]), .B(n2537), .CI(
        C[1559]), .CO(C[1560]) );
  FA_6629 \FA_INST_0[3].FA_INST_1[24].FA_  ( .A(A[1560]), .B(n2536), .CI(
        C[1560]), .CO(C[1561]) );
  FA_6628 \FA_INST_0[3].FA_INST_1[25].FA_  ( .A(A[1561]), .B(n2535), .CI(
        C[1561]), .CO(C[1562]) );
  FA_6627 \FA_INST_0[3].FA_INST_1[26].FA_  ( .A(A[1562]), .B(n2534), .CI(
        C[1562]), .CO(C[1563]) );
  FA_6626 \FA_INST_0[3].FA_INST_1[27].FA_  ( .A(A[1563]), .B(n2533), .CI(
        C[1563]), .CO(C[1564]) );
  FA_6625 \FA_INST_0[3].FA_INST_1[28].FA_  ( .A(A[1564]), .B(n2532), .CI(
        C[1564]), .CO(C[1565]) );
  FA_6624 \FA_INST_0[3].FA_INST_1[29].FA_  ( .A(A[1565]), .B(n2531), .CI(
        C[1565]), .CO(C[1566]) );
  FA_6623 \FA_INST_0[3].FA_INST_1[30].FA_  ( .A(A[1566]), .B(n2530), .CI(
        C[1566]), .CO(C[1567]) );
  FA_6622 \FA_INST_0[3].FA_INST_1[31].FA_  ( .A(A[1567]), .B(n2529), .CI(
        C[1567]), .CO(C[1568]) );
  FA_6621 \FA_INST_0[3].FA_INST_1[32].FA_  ( .A(A[1568]), .B(n2528), .CI(
        C[1568]), .CO(C[1569]) );
  FA_6620 \FA_INST_0[3].FA_INST_1[33].FA_  ( .A(A[1569]), .B(n2527), .CI(
        C[1569]), .CO(C[1570]) );
  FA_6619 \FA_INST_0[3].FA_INST_1[34].FA_  ( .A(A[1570]), .B(n2526), .CI(
        C[1570]), .CO(C[1571]) );
  FA_6618 \FA_INST_0[3].FA_INST_1[35].FA_  ( .A(A[1571]), .B(n2525), .CI(
        C[1571]), .CO(C[1572]) );
  FA_6617 \FA_INST_0[3].FA_INST_1[36].FA_  ( .A(A[1572]), .B(n2524), .CI(
        C[1572]), .CO(C[1573]) );
  FA_6616 \FA_INST_0[3].FA_INST_1[37].FA_  ( .A(A[1573]), .B(n2523), .CI(
        C[1573]), .CO(C[1574]) );
  FA_6615 \FA_INST_0[3].FA_INST_1[38].FA_  ( .A(A[1574]), .B(n2522), .CI(
        C[1574]), .CO(C[1575]) );
  FA_6614 \FA_INST_0[3].FA_INST_1[39].FA_  ( .A(A[1575]), .B(n2521), .CI(
        C[1575]), .CO(C[1576]) );
  FA_6613 \FA_INST_0[3].FA_INST_1[40].FA_  ( .A(A[1576]), .B(n2520), .CI(
        C[1576]), .CO(C[1577]) );
  FA_6612 \FA_INST_0[3].FA_INST_1[41].FA_  ( .A(A[1577]), .B(n2519), .CI(
        C[1577]), .CO(C[1578]) );
  FA_6611 \FA_INST_0[3].FA_INST_1[42].FA_  ( .A(A[1578]), .B(n2518), .CI(
        C[1578]), .CO(C[1579]) );
  FA_6610 \FA_INST_0[3].FA_INST_1[43].FA_  ( .A(A[1579]), .B(n2517), .CI(
        C[1579]), .CO(C[1580]) );
  FA_6609 \FA_INST_0[3].FA_INST_1[44].FA_  ( .A(A[1580]), .B(n2516), .CI(
        C[1580]), .CO(C[1581]) );
  FA_6608 \FA_INST_0[3].FA_INST_1[45].FA_  ( .A(A[1581]), .B(n2515), .CI(
        C[1581]), .CO(C[1582]) );
  FA_6607 \FA_INST_0[3].FA_INST_1[46].FA_  ( .A(A[1582]), .B(n2514), .CI(
        C[1582]), .CO(C[1583]) );
  FA_6606 \FA_INST_0[3].FA_INST_1[47].FA_  ( .A(A[1583]), .B(n2513), .CI(
        C[1583]), .CO(C[1584]) );
  FA_6605 \FA_INST_0[3].FA_INST_1[48].FA_  ( .A(A[1584]), .B(n2512), .CI(
        C[1584]), .CO(C[1585]) );
  FA_6604 \FA_INST_0[3].FA_INST_1[49].FA_  ( .A(A[1585]), .B(n2511), .CI(
        C[1585]), .CO(C[1586]) );
  FA_6603 \FA_INST_0[3].FA_INST_1[50].FA_  ( .A(A[1586]), .B(n2510), .CI(
        C[1586]), .CO(C[1587]) );
  FA_6602 \FA_INST_0[3].FA_INST_1[51].FA_  ( .A(A[1587]), .B(n2509), .CI(
        C[1587]), .CO(C[1588]) );
  FA_6601 \FA_INST_0[3].FA_INST_1[52].FA_  ( .A(A[1588]), .B(n2508), .CI(
        C[1588]), .CO(C[1589]) );
  FA_6600 \FA_INST_0[3].FA_INST_1[53].FA_  ( .A(A[1589]), .B(n2507), .CI(
        C[1589]), .CO(C[1590]) );
  FA_6599 \FA_INST_0[3].FA_INST_1[54].FA_  ( .A(A[1590]), .B(n2506), .CI(
        C[1590]), .CO(C[1591]) );
  FA_6598 \FA_INST_0[3].FA_INST_1[55].FA_  ( .A(A[1591]), .B(n2505), .CI(
        C[1591]), .CO(C[1592]) );
  FA_6597 \FA_INST_0[3].FA_INST_1[56].FA_  ( .A(A[1592]), .B(n2504), .CI(
        C[1592]), .CO(C[1593]) );
  FA_6596 \FA_INST_0[3].FA_INST_1[57].FA_  ( .A(A[1593]), .B(n2503), .CI(
        C[1593]), .CO(C[1594]) );
  FA_6595 \FA_INST_0[3].FA_INST_1[58].FA_  ( .A(A[1594]), .B(n2502), .CI(
        C[1594]), .CO(C[1595]) );
  FA_6594 \FA_INST_0[3].FA_INST_1[59].FA_  ( .A(A[1595]), .B(n2501), .CI(
        C[1595]), .CO(C[1596]) );
  FA_6593 \FA_INST_0[3].FA_INST_1[60].FA_  ( .A(A[1596]), .B(n2500), .CI(
        C[1596]), .CO(C[1597]) );
  FA_6592 \FA_INST_0[3].FA_INST_1[61].FA_  ( .A(A[1597]), .B(n2499), .CI(
        C[1597]), .CO(C[1598]) );
  FA_6591 \FA_INST_0[3].FA_INST_1[62].FA_  ( .A(A[1598]), .B(n2498), .CI(
        C[1598]), .CO(C[1599]) );
  FA_6590 \FA_INST_0[3].FA_INST_1[63].FA_  ( .A(A[1599]), .B(n2497), .CI(
        C[1599]), .CO(C[1600]) );
  FA_6589 \FA_INST_0[3].FA_INST_1[64].FA_  ( .A(A[1600]), .B(n2496), .CI(
        C[1600]), .CO(C[1601]) );
  FA_6588 \FA_INST_0[3].FA_INST_1[65].FA_  ( .A(A[1601]), .B(n2495), .CI(
        C[1601]), .CO(C[1602]) );
  FA_6587 \FA_INST_0[3].FA_INST_1[66].FA_  ( .A(A[1602]), .B(n2494), .CI(
        C[1602]), .CO(C[1603]) );
  FA_6586 \FA_INST_0[3].FA_INST_1[67].FA_  ( .A(A[1603]), .B(n2493), .CI(
        C[1603]), .CO(C[1604]) );
  FA_6585 \FA_INST_0[3].FA_INST_1[68].FA_  ( .A(A[1604]), .B(n2492), .CI(
        C[1604]), .CO(C[1605]) );
  FA_6584 \FA_INST_0[3].FA_INST_1[69].FA_  ( .A(A[1605]), .B(n2491), .CI(
        C[1605]), .CO(C[1606]) );
  FA_6583 \FA_INST_0[3].FA_INST_1[70].FA_  ( .A(A[1606]), .B(n2490), .CI(
        C[1606]), .CO(C[1607]) );
  FA_6582 \FA_INST_0[3].FA_INST_1[71].FA_  ( .A(A[1607]), .B(n2489), .CI(
        C[1607]), .CO(C[1608]) );
  FA_6581 \FA_INST_0[3].FA_INST_1[72].FA_  ( .A(A[1608]), .B(n2488), .CI(
        C[1608]), .CO(C[1609]) );
  FA_6580 \FA_INST_0[3].FA_INST_1[73].FA_  ( .A(A[1609]), .B(n2487), .CI(
        C[1609]), .CO(C[1610]) );
  FA_6579 \FA_INST_0[3].FA_INST_1[74].FA_  ( .A(A[1610]), .B(n2486), .CI(
        C[1610]), .CO(C[1611]) );
  FA_6578 \FA_INST_0[3].FA_INST_1[75].FA_  ( .A(A[1611]), .B(n2485), .CI(
        C[1611]), .CO(C[1612]) );
  FA_6577 \FA_INST_0[3].FA_INST_1[76].FA_  ( .A(A[1612]), .B(n2484), .CI(
        C[1612]), .CO(C[1613]) );
  FA_6576 \FA_INST_0[3].FA_INST_1[77].FA_  ( .A(A[1613]), .B(n2483), .CI(
        C[1613]), .CO(C[1614]) );
  FA_6575 \FA_INST_0[3].FA_INST_1[78].FA_  ( .A(A[1614]), .B(n2482), .CI(
        C[1614]), .CO(C[1615]) );
  FA_6574 \FA_INST_0[3].FA_INST_1[79].FA_  ( .A(A[1615]), .B(n2481), .CI(
        C[1615]), .CO(C[1616]) );
  FA_6573 \FA_INST_0[3].FA_INST_1[80].FA_  ( .A(A[1616]), .B(n2480), .CI(
        C[1616]), .CO(C[1617]) );
  FA_6572 \FA_INST_0[3].FA_INST_1[81].FA_  ( .A(A[1617]), .B(n2479), .CI(
        C[1617]), .CO(C[1618]) );
  FA_6571 \FA_INST_0[3].FA_INST_1[82].FA_  ( .A(A[1618]), .B(n2478), .CI(
        C[1618]), .CO(C[1619]) );
  FA_6570 \FA_INST_0[3].FA_INST_1[83].FA_  ( .A(A[1619]), .B(n2477), .CI(
        C[1619]), .CO(C[1620]) );
  FA_6569 \FA_INST_0[3].FA_INST_1[84].FA_  ( .A(A[1620]), .B(n2476), .CI(
        C[1620]), .CO(C[1621]) );
  FA_6568 \FA_INST_0[3].FA_INST_1[85].FA_  ( .A(A[1621]), .B(n2475), .CI(
        C[1621]), .CO(C[1622]) );
  FA_6567 \FA_INST_0[3].FA_INST_1[86].FA_  ( .A(A[1622]), .B(n2474), .CI(
        C[1622]), .CO(C[1623]) );
  FA_6566 \FA_INST_0[3].FA_INST_1[87].FA_  ( .A(A[1623]), .B(n2473), .CI(
        C[1623]), .CO(C[1624]) );
  FA_6565 \FA_INST_0[3].FA_INST_1[88].FA_  ( .A(A[1624]), .B(n2472), .CI(
        C[1624]), .CO(C[1625]) );
  FA_6564 \FA_INST_0[3].FA_INST_1[89].FA_  ( .A(A[1625]), .B(n2471), .CI(
        C[1625]), .CO(C[1626]) );
  FA_6563 \FA_INST_0[3].FA_INST_1[90].FA_  ( .A(A[1626]), .B(n2470), .CI(
        C[1626]), .CO(C[1627]) );
  FA_6562 \FA_INST_0[3].FA_INST_1[91].FA_  ( .A(A[1627]), .B(n2469), .CI(
        C[1627]), .CO(C[1628]) );
  FA_6561 \FA_INST_0[3].FA_INST_1[92].FA_  ( .A(A[1628]), .B(n2468), .CI(
        C[1628]), .CO(C[1629]) );
  FA_6560 \FA_INST_0[3].FA_INST_1[93].FA_  ( .A(A[1629]), .B(n2467), .CI(
        C[1629]), .CO(C[1630]) );
  FA_6559 \FA_INST_0[3].FA_INST_1[94].FA_  ( .A(A[1630]), .B(n2466), .CI(
        C[1630]), .CO(C[1631]) );
  FA_6558 \FA_INST_0[3].FA_INST_1[95].FA_  ( .A(A[1631]), .B(n2465), .CI(
        C[1631]), .CO(C[1632]) );
  FA_6557 \FA_INST_0[3].FA_INST_1[96].FA_  ( .A(A[1632]), .B(n2464), .CI(
        C[1632]), .CO(C[1633]) );
  FA_6556 \FA_INST_0[3].FA_INST_1[97].FA_  ( .A(A[1633]), .B(n2463), .CI(
        C[1633]), .CO(C[1634]) );
  FA_6555 \FA_INST_0[3].FA_INST_1[98].FA_  ( .A(A[1634]), .B(n2462), .CI(
        C[1634]), .CO(C[1635]) );
  FA_6554 \FA_INST_0[3].FA_INST_1[99].FA_  ( .A(A[1635]), .B(n2461), .CI(
        C[1635]), .CO(C[1636]) );
  FA_6553 \FA_INST_0[3].FA_INST_1[100].FA_  ( .A(A[1636]), .B(n2460), .CI(
        C[1636]), .CO(C[1637]) );
  FA_6552 \FA_INST_0[3].FA_INST_1[101].FA_  ( .A(A[1637]), .B(n2459), .CI(
        C[1637]), .CO(C[1638]) );
  FA_6551 \FA_INST_0[3].FA_INST_1[102].FA_  ( .A(A[1638]), .B(n2458), .CI(
        C[1638]), .CO(C[1639]) );
  FA_6550 \FA_INST_0[3].FA_INST_1[103].FA_  ( .A(A[1639]), .B(n2457), .CI(
        C[1639]), .CO(C[1640]) );
  FA_6549 \FA_INST_0[3].FA_INST_1[104].FA_  ( .A(A[1640]), .B(n2456), .CI(
        C[1640]), .CO(C[1641]) );
  FA_6548 \FA_INST_0[3].FA_INST_1[105].FA_  ( .A(A[1641]), .B(n2455), .CI(
        C[1641]), .CO(C[1642]) );
  FA_6547 \FA_INST_0[3].FA_INST_1[106].FA_  ( .A(A[1642]), .B(n2454), .CI(
        C[1642]), .CO(C[1643]) );
  FA_6546 \FA_INST_0[3].FA_INST_1[107].FA_  ( .A(A[1643]), .B(n2453), .CI(
        C[1643]), .CO(C[1644]) );
  FA_6545 \FA_INST_0[3].FA_INST_1[108].FA_  ( .A(A[1644]), .B(n2452), .CI(
        C[1644]), .CO(C[1645]) );
  FA_6544 \FA_INST_0[3].FA_INST_1[109].FA_  ( .A(A[1645]), .B(n2451), .CI(
        C[1645]), .CO(C[1646]) );
  FA_6543 \FA_INST_0[3].FA_INST_1[110].FA_  ( .A(A[1646]), .B(n2450), .CI(
        C[1646]), .CO(C[1647]) );
  FA_6542 \FA_INST_0[3].FA_INST_1[111].FA_  ( .A(A[1647]), .B(n2449), .CI(
        C[1647]), .CO(C[1648]) );
  FA_6541 \FA_INST_0[3].FA_INST_1[112].FA_  ( .A(A[1648]), .B(n2448), .CI(
        C[1648]), .CO(C[1649]) );
  FA_6540 \FA_INST_0[3].FA_INST_1[113].FA_  ( .A(A[1649]), .B(n2447), .CI(
        C[1649]), .CO(C[1650]) );
  FA_6539 \FA_INST_0[3].FA_INST_1[114].FA_  ( .A(A[1650]), .B(n2446), .CI(
        C[1650]), .CO(C[1651]) );
  FA_6538 \FA_INST_0[3].FA_INST_1[115].FA_  ( .A(A[1651]), .B(n2445), .CI(
        C[1651]), .CO(C[1652]) );
  FA_6537 \FA_INST_0[3].FA_INST_1[116].FA_  ( .A(A[1652]), .B(n2444), .CI(
        C[1652]), .CO(C[1653]) );
  FA_6536 \FA_INST_0[3].FA_INST_1[117].FA_  ( .A(A[1653]), .B(n2443), .CI(
        C[1653]), .CO(C[1654]) );
  FA_6535 \FA_INST_0[3].FA_INST_1[118].FA_  ( .A(A[1654]), .B(n2442), .CI(
        C[1654]), .CO(C[1655]) );
  FA_6534 \FA_INST_0[3].FA_INST_1[119].FA_  ( .A(A[1655]), .B(n2441), .CI(
        C[1655]), .CO(C[1656]) );
  FA_6533 \FA_INST_0[3].FA_INST_1[120].FA_  ( .A(A[1656]), .B(n2440), .CI(
        C[1656]), .CO(C[1657]) );
  FA_6532 \FA_INST_0[3].FA_INST_1[121].FA_  ( .A(A[1657]), .B(n2439), .CI(
        C[1657]), .CO(C[1658]) );
  FA_6531 \FA_INST_0[3].FA_INST_1[122].FA_  ( .A(A[1658]), .B(n2438), .CI(
        C[1658]), .CO(C[1659]) );
  FA_6530 \FA_INST_0[3].FA_INST_1[123].FA_  ( .A(A[1659]), .B(n2437), .CI(
        C[1659]), .CO(C[1660]) );
  FA_6529 \FA_INST_0[3].FA_INST_1[124].FA_  ( .A(A[1660]), .B(n2436), .CI(
        C[1660]), .CO(C[1661]) );
  FA_6528 \FA_INST_0[3].FA_INST_1[125].FA_  ( .A(A[1661]), .B(n2435), .CI(
        C[1661]), .CO(C[1662]) );
  FA_6527 \FA_INST_0[3].FA_INST_1[126].FA_  ( .A(A[1662]), .B(n2434), .CI(
        C[1662]), .CO(C[1663]) );
  FA_6526 \FA_INST_0[3].FA_INST_1[127].FA_  ( .A(A[1663]), .B(n2433), .CI(
        C[1663]), .CO(C[1664]) );
  FA_6525 \FA_INST_0[3].FA_INST_1[128].FA_  ( .A(A[1664]), .B(n2432), .CI(
        C[1664]), .CO(C[1665]) );
  FA_6524 \FA_INST_0[3].FA_INST_1[129].FA_  ( .A(A[1665]), .B(n2431), .CI(
        C[1665]), .CO(C[1666]) );
  FA_6523 \FA_INST_0[3].FA_INST_1[130].FA_  ( .A(A[1666]), .B(n2430), .CI(
        C[1666]), .CO(C[1667]) );
  FA_6522 \FA_INST_0[3].FA_INST_1[131].FA_  ( .A(A[1667]), .B(n2429), .CI(
        C[1667]), .CO(C[1668]) );
  FA_6521 \FA_INST_0[3].FA_INST_1[132].FA_  ( .A(A[1668]), .B(n2428), .CI(
        C[1668]), .CO(C[1669]) );
  FA_6520 \FA_INST_0[3].FA_INST_1[133].FA_  ( .A(A[1669]), .B(n2427), .CI(
        C[1669]), .CO(C[1670]) );
  FA_6519 \FA_INST_0[3].FA_INST_1[134].FA_  ( .A(A[1670]), .B(n2426), .CI(
        C[1670]), .CO(C[1671]) );
  FA_6518 \FA_INST_0[3].FA_INST_1[135].FA_  ( .A(A[1671]), .B(n2425), .CI(
        C[1671]), .CO(C[1672]) );
  FA_6517 \FA_INST_0[3].FA_INST_1[136].FA_  ( .A(A[1672]), .B(n2424), .CI(
        C[1672]), .CO(C[1673]) );
  FA_6516 \FA_INST_0[3].FA_INST_1[137].FA_  ( .A(A[1673]), .B(n2423), .CI(
        C[1673]), .CO(C[1674]) );
  FA_6515 \FA_INST_0[3].FA_INST_1[138].FA_  ( .A(A[1674]), .B(n2422), .CI(
        C[1674]), .CO(C[1675]) );
  FA_6514 \FA_INST_0[3].FA_INST_1[139].FA_  ( .A(A[1675]), .B(n2421), .CI(
        C[1675]), .CO(C[1676]) );
  FA_6513 \FA_INST_0[3].FA_INST_1[140].FA_  ( .A(A[1676]), .B(n2420), .CI(
        C[1676]), .CO(C[1677]) );
  FA_6512 \FA_INST_0[3].FA_INST_1[141].FA_  ( .A(A[1677]), .B(n2419), .CI(
        C[1677]), .CO(C[1678]) );
  FA_6511 \FA_INST_0[3].FA_INST_1[142].FA_  ( .A(A[1678]), .B(n2418), .CI(
        C[1678]), .CO(C[1679]) );
  FA_6510 \FA_INST_0[3].FA_INST_1[143].FA_  ( .A(A[1679]), .B(n2417), .CI(
        C[1679]), .CO(C[1680]) );
  FA_6509 \FA_INST_0[3].FA_INST_1[144].FA_  ( .A(A[1680]), .B(n2416), .CI(
        C[1680]), .CO(C[1681]) );
  FA_6508 \FA_INST_0[3].FA_INST_1[145].FA_  ( .A(A[1681]), .B(n2415), .CI(
        C[1681]), .CO(C[1682]) );
  FA_6507 \FA_INST_0[3].FA_INST_1[146].FA_  ( .A(A[1682]), .B(n2414), .CI(
        C[1682]), .CO(C[1683]) );
  FA_6506 \FA_INST_0[3].FA_INST_1[147].FA_  ( .A(A[1683]), .B(n2413), .CI(
        C[1683]), .CO(C[1684]) );
  FA_6505 \FA_INST_0[3].FA_INST_1[148].FA_  ( .A(A[1684]), .B(n2412), .CI(
        C[1684]), .CO(C[1685]) );
  FA_6504 \FA_INST_0[3].FA_INST_1[149].FA_  ( .A(A[1685]), .B(n2411), .CI(
        C[1685]), .CO(C[1686]) );
  FA_6503 \FA_INST_0[3].FA_INST_1[150].FA_  ( .A(A[1686]), .B(n2410), .CI(
        C[1686]), .CO(C[1687]) );
  FA_6502 \FA_INST_0[3].FA_INST_1[151].FA_  ( .A(A[1687]), .B(n2409), .CI(
        C[1687]), .CO(C[1688]) );
  FA_6501 \FA_INST_0[3].FA_INST_1[152].FA_  ( .A(A[1688]), .B(n2408), .CI(
        C[1688]), .CO(C[1689]) );
  FA_6500 \FA_INST_0[3].FA_INST_1[153].FA_  ( .A(A[1689]), .B(n2407), .CI(
        C[1689]), .CO(C[1690]) );
  FA_6499 \FA_INST_0[3].FA_INST_1[154].FA_  ( .A(A[1690]), .B(n2406), .CI(
        C[1690]), .CO(C[1691]) );
  FA_6498 \FA_INST_0[3].FA_INST_1[155].FA_  ( .A(A[1691]), .B(n2405), .CI(
        C[1691]), .CO(C[1692]) );
  FA_6497 \FA_INST_0[3].FA_INST_1[156].FA_  ( .A(A[1692]), .B(n2404), .CI(
        C[1692]), .CO(C[1693]) );
  FA_6496 \FA_INST_0[3].FA_INST_1[157].FA_  ( .A(A[1693]), .B(n2403), .CI(
        C[1693]), .CO(C[1694]) );
  FA_6495 \FA_INST_0[3].FA_INST_1[158].FA_  ( .A(A[1694]), .B(n2402), .CI(
        C[1694]), .CO(C[1695]) );
  FA_6494 \FA_INST_0[3].FA_INST_1[159].FA_  ( .A(A[1695]), .B(n2401), .CI(
        C[1695]), .CO(C[1696]) );
  FA_6493 \FA_INST_0[3].FA_INST_1[160].FA_  ( .A(A[1696]), .B(n2400), .CI(
        C[1696]), .CO(C[1697]) );
  FA_6492 \FA_INST_0[3].FA_INST_1[161].FA_  ( .A(A[1697]), .B(n2399), .CI(
        C[1697]), .CO(C[1698]) );
  FA_6491 \FA_INST_0[3].FA_INST_1[162].FA_  ( .A(A[1698]), .B(n2398), .CI(
        C[1698]), .CO(C[1699]) );
  FA_6490 \FA_INST_0[3].FA_INST_1[163].FA_  ( .A(A[1699]), .B(n2397), .CI(
        C[1699]), .CO(C[1700]) );
  FA_6489 \FA_INST_0[3].FA_INST_1[164].FA_  ( .A(A[1700]), .B(n2396), .CI(
        C[1700]), .CO(C[1701]) );
  FA_6488 \FA_INST_0[3].FA_INST_1[165].FA_  ( .A(A[1701]), .B(n2395), .CI(
        C[1701]), .CO(C[1702]) );
  FA_6487 \FA_INST_0[3].FA_INST_1[166].FA_  ( .A(A[1702]), .B(n2394), .CI(
        C[1702]), .CO(C[1703]) );
  FA_6486 \FA_INST_0[3].FA_INST_1[167].FA_  ( .A(A[1703]), .B(n2393), .CI(
        C[1703]), .CO(C[1704]) );
  FA_6485 \FA_INST_0[3].FA_INST_1[168].FA_  ( .A(A[1704]), .B(n2392), .CI(
        C[1704]), .CO(C[1705]) );
  FA_6484 \FA_INST_0[3].FA_INST_1[169].FA_  ( .A(A[1705]), .B(n2391), .CI(
        C[1705]), .CO(C[1706]) );
  FA_6483 \FA_INST_0[3].FA_INST_1[170].FA_  ( .A(A[1706]), .B(n2390), .CI(
        C[1706]), .CO(C[1707]) );
  FA_6482 \FA_INST_0[3].FA_INST_1[171].FA_  ( .A(A[1707]), .B(n2389), .CI(
        C[1707]), .CO(C[1708]) );
  FA_6481 \FA_INST_0[3].FA_INST_1[172].FA_  ( .A(A[1708]), .B(n2388), .CI(
        C[1708]), .CO(C[1709]) );
  FA_6480 \FA_INST_0[3].FA_INST_1[173].FA_  ( .A(A[1709]), .B(n2387), .CI(
        C[1709]), .CO(C[1710]) );
  FA_6479 \FA_INST_0[3].FA_INST_1[174].FA_  ( .A(A[1710]), .B(n2386), .CI(
        C[1710]), .CO(C[1711]) );
  FA_6478 \FA_INST_0[3].FA_INST_1[175].FA_  ( .A(A[1711]), .B(n2385), .CI(
        C[1711]), .CO(C[1712]) );
  FA_6477 \FA_INST_0[3].FA_INST_1[176].FA_  ( .A(A[1712]), .B(n2384), .CI(
        C[1712]), .CO(C[1713]) );
  FA_6476 \FA_INST_0[3].FA_INST_1[177].FA_  ( .A(A[1713]), .B(n2383), .CI(
        C[1713]), .CO(C[1714]) );
  FA_6475 \FA_INST_0[3].FA_INST_1[178].FA_  ( .A(A[1714]), .B(n2382), .CI(
        C[1714]), .CO(C[1715]) );
  FA_6474 \FA_INST_0[3].FA_INST_1[179].FA_  ( .A(A[1715]), .B(n2381), .CI(
        C[1715]), .CO(C[1716]) );
  FA_6473 \FA_INST_0[3].FA_INST_1[180].FA_  ( .A(A[1716]), .B(n2380), .CI(
        C[1716]), .CO(C[1717]) );
  FA_6472 \FA_INST_0[3].FA_INST_1[181].FA_  ( .A(A[1717]), .B(n2379), .CI(
        C[1717]), .CO(C[1718]) );
  FA_6471 \FA_INST_0[3].FA_INST_1[182].FA_  ( .A(A[1718]), .B(n2378), .CI(
        C[1718]), .CO(C[1719]) );
  FA_6470 \FA_INST_0[3].FA_INST_1[183].FA_  ( .A(A[1719]), .B(n2377), .CI(
        C[1719]), .CO(C[1720]) );
  FA_6469 \FA_INST_0[3].FA_INST_1[184].FA_  ( .A(A[1720]), .B(n2376), .CI(
        C[1720]), .CO(C[1721]) );
  FA_6468 \FA_INST_0[3].FA_INST_1[185].FA_  ( .A(A[1721]), .B(n2375), .CI(
        C[1721]), .CO(C[1722]) );
  FA_6467 \FA_INST_0[3].FA_INST_1[186].FA_  ( .A(A[1722]), .B(n2374), .CI(
        C[1722]), .CO(C[1723]) );
  FA_6466 \FA_INST_0[3].FA_INST_1[187].FA_  ( .A(A[1723]), .B(n2373), .CI(
        C[1723]), .CO(C[1724]) );
  FA_6465 \FA_INST_0[3].FA_INST_1[188].FA_  ( .A(A[1724]), .B(n2372), .CI(
        C[1724]), .CO(C[1725]) );
  FA_6464 \FA_INST_0[3].FA_INST_1[189].FA_  ( .A(A[1725]), .B(n2371), .CI(
        C[1725]), .CO(C[1726]) );
  FA_6463 \FA_INST_0[3].FA_INST_1[190].FA_  ( .A(A[1726]), .B(n2370), .CI(
        C[1726]), .CO(C[1727]) );
  FA_6462 \FA_INST_0[3].FA_INST_1[191].FA_  ( .A(A[1727]), .B(n2369), .CI(
        C[1727]), .CO(C[1728]) );
  FA_6461 \FA_INST_0[3].FA_INST_1[192].FA_  ( .A(A[1728]), .B(n2368), .CI(
        C[1728]), .CO(C[1729]) );
  FA_6460 \FA_INST_0[3].FA_INST_1[193].FA_  ( .A(A[1729]), .B(n2367), .CI(
        C[1729]), .CO(C[1730]) );
  FA_6459 \FA_INST_0[3].FA_INST_1[194].FA_  ( .A(A[1730]), .B(n2366), .CI(
        C[1730]), .CO(C[1731]) );
  FA_6458 \FA_INST_0[3].FA_INST_1[195].FA_  ( .A(A[1731]), .B(n2365), .CI(
        C[1731]), .CO(C[1732]) );
  FA_6457 \FA_INST_0[3].FA_INST_1[196].FA_  ( .A(A[1732]), .B(n2364), .CI(
        C[1732]), .CO(C[1733]) );
  FA_6456 \FA_INST_0[3].FA_INST_1[197].FA_  ( .A(A[1733]), .B(n2363), .CI(
        C[1733]), .CO(C[1734]) );
  FA_6455 \FA_INST_0[3].FA_INST_1[198].FA_  ( .A(A[1734]), .B(n2362), .CI(
        C[1734]), .CO(C[1735]) );
  FA_6454 \FA_INST_0[3].FA_INST_1[199].FA_  ( .A(A[1735]), .B(n2361), .CI(
        C[1735]), .CO(C[1736]) );
  FA_6453 \FA_INST_0[3].FA_INST_1[200].FA_  ( .A(A[1736]), .B(n2360), .CI(
        C[1736]), .CO(C[1737]) );
  FA_6452 \FA_INST_0[3].FA_INST_1[201].FA_  ( .A(A[1737]), .B(n2359), .CI(
        C[1737]), .CO(C[1738]) );
  FA_6451 \FA_INST_0[3].FA_INST_1[202].FA_  ( .A(A[1738]), .B(n2358), .CI(
        C[1738]), .CO(C[1739]) );
  FA_6450 \FA_INST_0[3].FA_INST_1[203].FA_  ( .A(A[1739]), .B(n2357), .CI(
        C[1739]), .CO(C[1740]) );
  FA_6449 \FA_INST_0[3].FA_INST_1[204].FA_  ( .A(A[1740]), .B(n2356), .CI(
        C[1740]), .CO(C[1741]) );
  FA_6448 \FA_INST_0[3].FA_INST_1[205].FA_  ( .A(A[1741]), .B(n2355), .CI(
        C[1741]), .CO(C[1742]) );
  FA_6447 \FA_INST_0[3].FA_INST_1[206].FA_  ( .A(A[1742]), .B(n2354), .CI(
        C[1742]), .CO(C[1743]) );
  FA_6446 \FA_INST_0[3].FA_INST_1[207].FA_  ( .A(A[1743]), .B(n2353), .CI(
        C[1743]), .CO(C[1744]) );
  FA_6445 \FA_INST_0[3].FA_INST_1[208].FA_  ( .A(A[1744]), .B(n2352), .CI(
        C[1744]), .CO(C[1745]) );
  FA_6444 \FA_INST_0[3].FA_INST_1[209].FA_  ( .A(A[1745]), .B(n2351), .CI(
        C[1745]), .CO(C[1746]) );
  FA_6443 \FA_INST_0[3].FA_INST_1[210].FA_  ( .A(A[1746]), .B(n2350), .CI(
        C[1746]), .CO(C[1747]) );
  FA_6442 \FA_INST_0[3].FA_INST_1[211].FA_  ( .A(A[1747]), .B(n2349), .CI(
        C[1747]), .CO(C[1748]) );
  FA_6441 \FA_INST_0[3].FA_INST_1[212].FA_  ( .A(A[1748]), .B(n2348), .CI(
        C[1748]), .CO(C[1749]) );
  FA_6440 \FA_INST_0[3].FA_INST_1[213].FA_  ( .A(A[1749]), .B(n2347), .CI(
        C[1749]), .CO(C[1750]) );
  FA_6439 \FA_INST_0[3].FA_INST_1[214].FA_  ( .A(A[1750]), .B(n2346), .CI(
        C[1750]), .CO(C[1751]) );
  FA_6438 \FA_INST_0[3].FA_INST_1[215].FA_  ( .A(A[1751]), .B(n2345), .CI(
        C[1751]), .CO(C[1752]) );
  FA_6437 \FA_INST_0[3].FA_INST_1[216].FA_  ( .A(A[1752]), .B(n2344), .CI(
        C[1752]), .CO(C[1753]) );
  FA_6436 \FA_INST_0[3].FA_INST_1[217].FA_  ( .A(A[1753]), .B(n2343), .CI(
        C[1753]), .CO(C[1754]) );
  FA_6435 \FA_INST_0[3].FA_INST_1[218].FA_  ( .A(A[1754]), .B(n2342), .CI(
        C[1754]), .CO(C[1755]) );
  FA_6434 \FA_INST_0[3].FA_INST_1[219].FA_  ( .A(A[1755]), .B(n2341), .CI(
        C[1755]), .CO(C[1756]) );
  FA_6433 \FA_INST_0[3].FA_INST_1[220].FA_  ( .A(A[1756]), .B(n2340), .CI(
        C[1756]), .CO(C[1757]) );
  FA_6432 \FA_INST_0[3].FA_INST_1[221].FA_  ( .A(A[1757]), .B(n2339), .CI(
        C[1757]), .CO(C[1758]) );
  FA_6431 \FA_INST_0[3].FA_INST_1[222].FA_  ( .A(A[1758]), .B(n2338), .CI(
        C[1758]), .CO(C[1759]) );
  FA_6430 \FA_INST_0[3].FA_INST_1[223].FA_  ( .A(A[1759]), .B(n2337), .CI(
        C[1759]), .CO(C[1760]) );
  FA_6429 \FA_INST_0[3].FA_INST_1[224].FA_  ( .A(A[1760]), .B(n2336), .CI(
        C[1760]), .CO(C[1761]) );
  FA_6428 \FA_INST_0[3].FA_INST_1[225].FA_  ( .A(A[1761]), .B(n2335), .CI(
        C[1761]), .CO(C[1762]) );
  FA_6427 \FA_INST_0[3].FA_INST_1[226].FA_  ( .A(A[1762]), .B(n2334), .CI(
        C[1762]), .CO(C[1763]) );
  FA_6426 \FA_INST_0[3].FA_INST_1[227].FA_  ( .A(A[1763]), .B(n2333), .CI(
        C[1763]), .CO(C[1764]) );
  FA_6425 \FA_INST_0[3].FA_INST_1[228].FA_  ( .A(A[1764]), .B(n2332), .CI(
        C[1764]), .CO(C[1765]) );
  FA_6424 \FA_INST_0[3].FA_INST_1[229].FA_  ( .A(A[1765]), .B(n2331), .CI(
        C[1765]), .CO(C[1766]) );
  FA_6423 \FA_INST_0[3].FA_INST_1[230].FA_  ( .A(A[1766]), .B(n2330), .CI(
        C[1766]), .CO(C[1767]) );
  FA_6422 \FA_INST_0[3].FA_INST_1[231].FA_  ( .A(A[1767]), .B(n2329), .CI(
        C[1767]), .CO(C[1768]) );
  FA_6421 \FA_INST_0[3].FA_INST_1[232].FA_  ( .A(A[1768]), .B(n2328), .CI(
        C[1768]), .CO(C[1769]) );
  FA_6420 \FA_INST_0[3].FA_INST_1[233].FA_  ( .A(A[1769]), .B(n2327), .CI(
        C[1769]), .CO(C[1770]) );
  FA_6419 \FA_INST_0[3].FA_INST_1[234].FA_  ( .A(A[1770]), .B(n2326), .CI(
        C[1770]), .CO(C[1771]) );
  FA_6418 \FA_INST_0[3].FA_INST_1[235].FA_  ( .A(A[1771]), .B(n2325), .CI(
        C[1771]), .CO(C[1772]) );
  FA_6417 \FA_INST_0[3].FA_INST_1[236].FA_  ( .A(A[1772]), .B(n2324), .CI(
        C[1772]), .CO(C[1773]) );
  FA_6416 \FA_INST_0[3].FA_INST_1[237].FA_  ( .A(A[1773]), .B(n2323), .CI(
        C[1773]), .CO(C[1774]) );
  FA_6415 \FA_INST_0[3].FA_INST_1[238].FA_  ( .A(A[1774]), .B(n2322), .CI(
        C[1774]), .CO(C[1775]) );
  FA_6414 \FA_INST_0[3].FA_INST_1[239].FA_  ( .A(A[1775]), .B(n2321), .CI(
        C[1775]), .CO(C[1776]) );
  FA_6413 \FA_INST_0[3].FA_INST_1[240].FA_  ( .A(A[1776]), .B(n2320), .CI(
        C[1776]), .CO(C[1777]) );
  FA_6412 \FA_INST_0[3].FA_INST_1[241].FA_  ( .A(A[1777]), .B(n2319), .CI(
        C[1777]), .CO(C[1778]) );
  FA_6411 \FA_INST_0[3].FA_INST_1[242].FA_  ( .A(A[1778]), .B(n2318), .CI(
        C[1778]), .CO(C[1779]) );
  FA_6410 \FA_INST_0[3].FA_INST_1[243].FA_  ( .A(A[1779]), .B(n2317), .CI(
        C[1779]), .CO(C[1780]) );
  FA_6409 \FA_INST_0[3].FA_INST_1[244].FA_  ( .A(A[1780]), .B(n2316), .CI(
        C[1780]), .CO(C[1781]) );
  FA_6408 \FA_INST_0[3].FA_INST_1[245].FA_  ( .A(A[1781]), .B(n2315), .CI(
        C[1781]), .CO(C[1782]) );
  FA_6407 \FA_INST_0[3].FA_INST_1[246].FA_  ( .A(A[1782]), .B(n2314), .CI(
        C[1782]), .CO(C[1783]) );
  FA_6406 \FA_INST_0[3].FA_INST_1[247].FA_  ( .A(A[1783]), .B(n2313), .CI(
        C[1783]), .CO(C[1784]) );
  FA_6405 \FA_INST_0[3].FA_INST_1[248].FA_  ( .A(A[1784]), .B(n2312), .CI(
        C[1784]), .CO(C[1785]) );
  FA_6404 \FA_INST_0[3].FA_INST_1[249].FA_  ( .A(A[1785]), .B(n2311), .CI(
        C[1785]), .CO(C[1786]) );
  FA_6403 \FA_INST_0[3].FA_INST_1[250].FA_  ( .A(A[1786]), .B(n2310), .CI(
        C[1786]), .CO(C[1787]) );
  FA_6402 \FA_INST_0[3].FA_INST_1[251].FA_  ( .A(A[1787]), .B(n2309), .CI(
        C[1787]), .CO(C[1788]) );
  FA_6401 \FA_INST_0[3].FA_INST_1[252].FA_  ( .A(A[1788]), .B(n2308), .CI(
        C[1788]), .CO(C[1789]) );
  FA_6400 \FA_INST_0[3].FA_INST_1[253].FA_  ( .A(A[1789]), .B(n2307), .CI(
        C[1789]), .CO(C[1790]) );
  FA_6399 \FA_INST_0[3].FA_INST_1[254].FA_  ( .A(A[1790]), .B(n2306), .CI(
        C[1790]), .CO(C[1791]) );
  FA_6398 \FA_INST_0[3].FA_INST_1[255].FA_  ( .A(A[1791]), .B(n2305), .CI(
        C[1791]), .CO(C[1792]) );
  FA_6397 \FA_INST_0[3].FA_INST_1[256].FA_  ( .A(A[1792]), .B(n2304), .CI(
        C[1792]), .CO(C[1793]) );
  FA_6396 \FA_INST_0[3].FA_INST_1[257].FA_  ( .A(A[1793]), .B(n2303), .CI(
        C[1793]), .CO(C[1794]) );
  FA_6395 \FA_INST_0[3].FA_INST_1[258].FA_  ( .A(A[1794]), .B(n2302), .CI(
        C[1794]), .CO(C[1795]) );
  FA_6394 \FA_INST_0[3].FA_INST_1[259].FA_  ( .A(A[1795]), .B(n2301), .CI(
        C[1795]), .CO(C[1796]) );
  FA_6393 \FA_INST_0[3].FA_INST_1[260].FA_  ( .A(A[1796]), .B(n2300), .CI(
        C[1796]), .CO(C[1797]) );
  FA_6392 \FA_INST_0[3].FA_INST_1[261].FA_  ( .A(A[1797]), .B(n2299), .CI(
        C[1797]), .CO(C[1798]) );
  FA_6391 \FA_INST_0[3].FA_INST_1[262].FA_  ( .A(A[1798]), .B(n2298), .CI(
        C[1798]), .CO(C[1799]) );
  FA_6390 \FA_INST_0[3].FA_INST_1[263].FA_  ( .A(A[1799]), .B(n2297), .CI(
        C[1799]), .CO(C[1800]) );
  FA_6389 \FA_INST_0[3].FA_INST_1[264].FA_  ( .A(A[1800]), .B(n2296), .CI(
        C[1800]), .CO(C[1801]) );
  FA_6388 \FA_INST_0[3].FA_INST_1[265].FA_  ( .A(A[1801]), .B(n2295), .CI(
        C[1801]), .CO(C[1802]) );
  FA_6387 \FA_INST_0[3].FA_INST_1[266].FA_  ( .A(A[1802]), .B(n2294), .CI(
        C[1802]), .CO(C[1803]) );
  FA_6386 \FA_INST_0[3].FA_INST_1[267].FA_  ( .A(A[1803]), .B(n2293), .CI(
        C[1803]), .CO(C[1804]) );
  FA_6385 \FA_INST_0[3].FA_INST_1[268].FA_  ( .A(A[1804]), .B(n2292), .CI(
        C[1804]), .CO(C[1805]) );
  FA_6384 \FA_INST_0[3].FA_INST_1[269].FA_  ( .A(A[1805]), .B(n2291), .CI(
        C[1805]), .CO(C[1806]) );
  FA_6383 \FA_INST_0[3].FA_INST_1[270].FA_  ( .A(A[1806]), .B(n2290), .CI(
        C[1806]), .CO(C[1807]) );
  FA_6382 \FA_INST_0[3].FA_INST_1[271].FA_  ( .A(A[1807]), .B(n2289), .CI(
        C[1807]), .CO(C[1808]) );
  FA_6381 \FA_INST_0[3].FA_INST_1[272].FA_  ( .A(A[1808]), .B(n2288), .CI(
        C[1808]), .CO(C[1809]) );
  FA_6380 \FA_INST_0[3].FA_INST_1[273].FA_  ( .A(A[1809]), .B(n2287), .CI(
        C[1809]), .CO(C[1810]) );
  FA_6379 \FA_INST_0[3].FA_INST_1[274].FA_  ( .A(A[1810]), .B(n2286), .CI(
        C[1810]), .CO(C[1811]) );
  FA_6378 \FA_INST_0[3].FA_INST_1[275].FA_  ( .A(A[1811]), .B(n2285), .CI(
        C[1811]), .CO(C[1812]) );
  FA_6377 \FA_INST_0[3].FA_INST_1[276].FA_  ( .A(A[1812]), .B(n2284), .CI(
        C[1812]), .CO(C[1813]) );
  FA_6376 \FA_INST_0[3].FA_INST_1[277].FA_  ( .A(A[1813]), .B(n2283), .CI(
        C[1813]), .CO(C[1814]) );
  FA_6375 \FA_INST_0[3].FA_INST_1[278].FA_  ( .A(A[1814]), .B(n2282), .CI(
        C[1814]), .CO(C[1815]) );
  FA_6374 \FA_INST_0[3].FA_INST_1[279].FA_  ( .A(A[1815]), .B(n2281), .CI(
        C[1815]), .CO(C[1816]) );
  FA_6373 \FA_INST_0[3].FA_INST_1[280].FA_  ( .A(A[1816]), .B(n2280), .CI(
        C[1816]), .CO(C[1817]) );
  FA_6372 \FA_INST_0[3].FA_INST_1[281].FA_  ( .A(A[1817]), .B(n2279), .CI(
        C[1817]), .CO(C[1818]) );
  FA_6371 \FA_INST_0[3].FA_INST_1[282].FA_  ( .A(A[1818]), .B(n2278), .CI(
        C[1818]), .CO(C[1819]) );
  FA_6370 \FA_INST_0[3].FA_INST_1[283].FA_  ( .A(A[1819]), .B(n2277), .CI(
        C[1819]), .CO(C[1820]) );
  FA_6369 \FA_INST_0[3].FA_INST_1[284].FA_  ( .A(A[1820]), .B(n2276), .CI(
        C[1820]), .CO(C[1821]) );
  FA_6368 \FA_INST_0[3].FA_INST_1[285].FA_  ( .A(A[1821]), .B(n2275), .CI(
        C[1821]), .CO(C[1822]) );
  FA_6367 \FA_INST_0[3].FA_INST_1[286].FA_  ( .A(A[1822]), .B(n2274), .CI(
        C[1822]), .CO(C[1823]) );
  FA_6366 \FA_INST_0[3].FA_INST_1[287].FA_  ( .A(A[1823]), .B(n2273), .CI(
        C[1823]), .CO(C[1824]) );
  FA_6365 \FA_INST_0[3].FA_INST_1[288].FA_  ( .A(A[1824]), .B(n2272), .CI(
        C[1824]), .CO(C[1825]) );
  FA_6364 \FA_INST_0[3].FA_INST_1[289].FA_  ( .A(A[1825]), .B(n2271), .CI(
        C[1825]), .CO(C[1826]) );
  FA_6363 \FA_INST_0[3].FA_INST_1[290].FA_  ( .A(A[1826]), .B(n2270), .CI(
        C[1826]), .CO(C[1827]) );
  FA_6362 \FA_INST_0[3].FA_INST_1[291].FA_  ( .A(A[1827]), .B(n2269), .CI(
        C[1827]), .CO(C[1828]) );
  FA_6361 \FA_INST_0[3].FA_INST_1[292].FA_  ( .A(A[1828]), .B(n2268), .CI(
        C[1828]), .CO(C[1829]) );
  FA_6360 \FA_INST_0[3].FA_INST_1[293].FA_  ( .A(A[1829]), .B(n2267), .CI(
        C[1829]), .CO(C[1830]) );
  FA_6359 \FA_INST_0[3].FA_INST_1[294].FA_  ( .A(A[1830]), .B(n2266), .CI(
        C[1830]), .CO(C[1831]) );
  FA_6358 \FA_INST_0[3].FA_INST_1[295].FA_  ( .A(A[1831]), .B(n2265), .CI(
        C[1831]), .CO(C[1832]) );
  FA_6357 \FA_INST_0[3].FA_INST_1[296].FA_  ( .A(A[1832]), .B(n2264), .CI(
        C[1832]), .CO(C[1833]) );
  FA_6356 \FA_INST_0[3].FA_INST_1[297].FA_  ( .A(A[1833]), .B(n2263), .CI(
        C[1833]), .CO(C[1834]) );
  FA_6355 \FA_INST_0[3].FA_INST_1[298].FA_  ( .A(A[1834]), .B(n2262), .CI(
        C[1834]), .CO(C[1835]) );
  FA_6354 \FA_INST_0[3].FA_INST_1[299].FA_  ( .A(A[1835]), .B(n2261), .CI(
        C[1835]), .CO(C[1836]) );
  FA_6353 \FA_INST_0[3].FA_INST_1[300].FA_  ( .A(A[1836]), .B(n2260), .CI(
        C[1836]), .CO(C[1837]) );
  FA_6352 \FA_INST_0[3].FA_INST_1[301].FA_  ( .A(A[1837]), .B(n2259), .CI(
        C[1837]), .CO(C[1838]) );
  FA_6351 \FA_INST_0[3].FA_INST_1[302].FA_  ( .A(A[1838]), .B(n2258), .CI(
        C[1838]), .CO(C[1839]) );
  FA_6350 \FA_INST_0[3].FA_INST_1[303].FA_  ( .A(A[1839]), .B(n2257), .CI(
        C[1839]), .CO(C[1840]) );
  FA_6349 \FA_INST_0[3].FA_INST_1[304].FA_  ( .A(A[1840]), .B(n2256), .CI(
        C[1840]), .CO(C[1841]) );
  FA_6348 \FA_INST_0[3].FA_INST_1[305].FA_  ( .A(A[1841]), .B(n2255), .CI(
        C[1841]), .CO(C[1842]) );
  FA_6347 \FA_INST_0[3].FA_INST_1[306].FA_  ( .A(A[1842]), .B(n2254), .CI(
        C[1842]), .CO(C[1843]) );
  FA_6346 \FA_INST_0[3].FA_INST_1[307].FA_  ( .A(A[1843]), .B(n2253), .CI(
        C[1843]), .CO(C[1844]) );
  FA_6345 \FA_INST_0[3].FA_INST_1[308].FA_  ( .A(A[1844]), .B(n2252), .CI(
        C[1844]), .CO(C[1845]) );
  FA_6344 \FA_INST_0[3].FA_INST_1[309].FA_  ( .A(A[1845]), .B(n2251), .CI(
        C[1845]), .CO(C[1846]) );
  FA_6343 \FA_INST_0[3].FA_INST_1[310].FA_  ( .A(A[1846]), .B(n2250), .CI(
        C[1846]), .CO(C[1847]) );
  FA_6342 \FA_INST_0[3].FA_INST_1[311].FA_  ( .A(A[1847]), .B(n2249), .CI(
        C[1847]), .CO(C[1848]) );
  FA_6341 \FA_INST_0[3].FA_INST_1[312].FA_  ( .A(A[1848]), .B(n2248), .CI(
        C[1848]), .CO(C[1849]) );
  FA_6340 \FA_INST_0[3].FA_INST_1[313].FA_  ( .A(A[1849]), .B(n2247), .CI(
        C[1849]), .CO(C[1850]) );
  FA_6339 \FA_INST_0[3].FA_INST_1[314].FA_  ( .A(A[1850]), .B(n2246), .CI(
        C[1850]), .CO(C[1851]) );
  FA_6338 \FA_INST_0[3].FA_INST_1[315].FA_  ( .A(A[1851]), .B(n2245), .CI(
        C[1851]), .CO(C[1852]) );
  FA_6337 \FA_INST_0[3].FA_INST_1[316].FA_  ( .A(A[1852]), .B(n2244), .CI(
        C[1852]), .CO(C[1853]) );
  FA_6336 \FA_INST_0[3].FA_INST_1[317].FA_  ( .A(A[1853]), .B(n2243), .CI(
        C[1853]), .CO(C[1854]) );
  FA_6335 \FA_INST_0[3].FA_INST_1[318].FA_  ( .A(A[1854]), .B(n2242), .CI(
        C[1854]), .CO(C[1855]) );
  FA_6334 \FA_INST_0[3].FA_INST_1[319].FA_  ( .A(A[1855]), .B(n2241), .CI(
        C[1855]), .CO(C[1856]) );
  FA_6333 \FA_INST_0[3].FA_INST_1[320].FA_  ( .A(A[1856]), .B(n2240), .CI(
        C[1856]), .CO(C[1857]) );
  FA_6332 \FA_INST_0[3].FA_INST_1[321].FA_  ( .A(A[1857]), .B(n2239), .CI(
        C[1857]), .CO(C[1858]) );
  FA_6331 \FA_INST_0[3].FA_INST_1[322].FA_  ( .A(A[1858]), .B(n2238), .CI(
        C[1858]), .CO(C[1859]) );
  FA_6330 \FA_INST_0[3].FA_INST_1[323].FA_  ( .A(A[1859]), .B(n2237), .CI(
        C[1859]), .CO(C[1860]) );
  FA_6329 \FA_INST_0[3].FA_INST_1[324].FA_  ( .A(A[1860]), .B(n2236), .CI(
        C[1860]), .CO(C[1861]) );
  FA_6328 \FA_INST_0[3].FA_INST_1[325].FA_  ( .A(A[1861]), .B(n2235), .CI(
        C[1861]), .CO(C[1862]) );
  FA_6327 \FA_INST_0[3].FA_INST_1[326].FA_  ( .A(A[1862]), .B(n2234), .CI(
        C[1862]), .CO(C[1863]) );
  FA_6326 \FA_INST_0[3].FA_INST_1[327].FA_  ( .A(A[1863]), .B(n2233), .CI(
        C[1863]), .CO(C[1864]) );
  FA_6325 \FA_INST_0[3].FA_INST_1[328].FA_  ( .A(A[1864]), .B(n2232), .CI(
        C[1864]), .CO(C[1865]) );
  FA_6324 \FA_INST_0[3].FA_INST_1[329].FA_  ( .A(A[1865]), .B(n2231), .CI(
        C[1865]), .CO(C[1866]) );
  FA_6323 \FA_INST_0[3].FA_INST_1[330].FA_  ( .A(A[1866]), .B(n2230), .CI(
        C[1866]), .CO(C[1867]) );
  FA_6322 \FA_INST_0[3].FA_INST_1[331].FA_  ( .A(A[1867]), .B(n2229), .CI(
        C[1867]), .CO(C[1868]) );
  FA_6321 \FA_INST_0[3].FA_INST_1[332].FA_  ( .A(A[1868]), .B(n2228), .CI(
        C[1868]), .CO(C[1869]) );
  FA_6320 \FA_INST_0[3].FA_INST_1[333].FA_  ( .A(A[1869]), .B(n2227), .CI(
        C[1869]), .CO(C[1870]) );
  FA_6319 \FA_INST_0[3].FA_INST_1[334].FA_  ( .A(A[1870]), .B(n2226), .CI(
        C[1870]), .CO(C[1871]) );
  FA_6318 \FA_INST_0[3].FA_INST_1[335].FA_  ( .A(A[1871]), .B(n2225), .CI(
        C[1871]), .CO(C[1872]) );
  FA_6317 \FA_INST_0[3].FA_INST_1[336].FA_  ( .A(A[1872]), .B(n2224), .CI(
        C[1872]), .CO(C[1873]) );
  FA_6316 \FA_INST_0[3].FA_INST_1[337].FA_  ( .A(A[1873]), .B(n2223), .CI(
        C[1873]), .CO(C[1874]) );
  FA_6315 \FA_INST_0[3].FA_INST_1[338].FA_  ( .A(A[1874]), .B(n2222), .CI(
        C[1874]), .CO(C[1875]) );
  FA_6314 \FA_INST_0[3].FA_INST_1[339].FA_  ( .A(A[1875]), .B(n2221), .CI(
        C[1875]), .CO(C[1876]) );
  FA_6313 \FA_INST_0[3].FA_INST_1[340].FA_  ( .A(A[1876]), .B(n2220), .CI(
        C[1876]), .CO(C[1877]) );
  FA_6312 \FA_INST_0[3].FA_INST_1[341].FA_  ( .A(A[1877]), .B(n2219), .CI(
        C[1877]), .CO(C[1878]) );
  FA_6311 \FA_INST_0[3].FA_INST_1[342].FA_  ( .A(A[1878]), .B(n2218), .CI(
        C[1878]), .CO(C[1879]) );
  FA_6310 \FA_INST_0[3].FA_INST_1[343].FA_  ( .A(A[1879]), .B(n2217), .CI(
        C[1879]), .CO(C[1880]) );
  FA_6309 \FA_INST_0[3].FA_INST_1[344].FA_  ( .A(A[1880]), .B(n2216), .CI(
        C[1880]), .CO(C[1881]) );
  FA_6308 \FA_INST_0[3].FA_INST_1[345].FA_  ( .A(A[1881]), .B(n2215), .CI(
        C[1881]), .CO(C[1882]) );
  FA_6307 \FA_INST_0[3].FA_INST_1[346].FA_  ( .A(A[1882]), .B(n2214), .CI(
        C[1882]), .CO(C[1883]) );
  FA_6306 \FA_INST_0[3].FA_INST_1[347].FA_  ( .A(A[1883]), .B(n2213), .CI(
        C[1883]), .CO(C[1884]) );
  FA_6305 \FA_INST_0[3].FA_INST_1[348].FA_  ( .A(A[1884]), .B(n2212), .CI(
        C[1884]), .CO(C[1885]) );
  FA_6304 \FA_INST_0[3].FA_INST_1[349].FA_  ( .A(A[1885]), .B(n2211), .CI(
        C[1885]), .CO(C[1886]) );
  FA_6303 \FA_INST_0[3].FA_INST_1[350].FA_  ( .A(A[1886]), .B(n2210), .CI(
        C[1886]), .CO(C[1887]) );
  FA_6302 \FA_INST_0[3].FA_INST_1[351].FA_  ( .A(A[1887]), .B(n2209), .CI(
        C[1887]), .CO(C[1888]) );
  FA_6301 \FA_INST_0[3].FA_INST_1[352].FA_  ( .A(A[1888]), .B(n2208), .CI(
        C[1888]), .CO(C[1889]) );
  FA_6300 \FA_INST_0[3].FA_INST_1[353].FA_  ( .A(A[1889]), .B(n2207), .CI(
        C[1889]), .CO(C[1890]) );
  FA_6299 \FA_INST_0[3].FA_INST_1[354].FA_  ( .A(A[1890]), .B(n2206), .CI(
        C[1890]), .CO(C[1891]) );
  FA_6298 \FA_INST_0[3].FA_INST_1[355].FA_  ( .A(A[1891]), .B(n2205), .CI(
        C[1891]), .CO(C[1892]) );
  FA_6297 \FA_INST_0[3].FA_INST_1[356].FA_  ( .A(A[1892]), .B(n2204), .CI(
        C[1892]), .CO(C[1893]) );
  FA_6296 \FA_INST_0[3].FA_INST_1[357].FA_  ( .A(A[1893]), .B(n2203), .CI(
        C[1893]), .CO(C[1894]) );
  FA_6295 \FA_INST_0[3].FA_INST_1[358].FA_  ( .A(A[1894]), .B(n2202), .CI(
        C[1894]), .CO(C[1895]) );
  FA_6294 \FA_INST_0[3].FA_INST_1[359].FA_  ( .A(A[1895]), .B(n2201), .CI(
        C[1895]), .CO(C[1896]) );
  FA_6293 \FA_INST_0[3].FA_INST_1[360].FA_  ( .A(A[1896]), .B(n2200), .CI(
        C[1896]), .CO(C[1897]) );
  FA_6292 \FA_INST_0[3].FA_INST_1[361].FA_  ( .A(A[1897]), .B(n2199), .CI(
        C[1897]), .CO(C[1898]) );
  FA_6291 \FA_INST_0[3].FA_INST_1[362].FA_  ( .A(A[1898]), .B(n2198), .CI(
        C[1898]), .CO(C[1899]) );
  FA_6290 \FA_INST_0[3].FA_INST_1[363].FA_  ( .A(A[1899]), .B(n2197), .CI(
        C[1899]), .CO(C[1900]) );
  FA_6289 \FA_INST_0[3].FA_INST_1[364].FA_  ( .A(A[1900]), .B(n2196), .CI(
        C[1900]), .CO(C[1901]) );
  FA_6288 \FA_INST_0[3].FA_INST_1[365].FA_  ( .A(A[1901]), .B(n2195), .CI(
        C[1901]), .CO(C[1902]) );
  FA_6287 \FA_INST_0[3].FA_INST_1[366].FA_  ( .A(A[1902]), .B(n2194), .CI(
        C[1902]), .CO(C[1903]) );
  FA_6286 \FA_INST_0[3].FA_INST_1[367].FA_  ( .A(A[1903]), .B(n2193), .CI(
        C[1903]), .CO(C[1904]) );
  FA_6285 \FA_INST_0[3].FA_INST_1[368].FA_  ( .A(A[1904]), .B(n2192), .CI(
        C[1904]), .CO(C[1905]) );
  FA_6284 \FA_INST_0[3].FA_INST_1[369].FA_  ( .A(A[1905]), .B(n2191), .CI(
        C[1905]), .CO(C[1906]) );
  FA_6283 \FA_INST_0[3].FA_INST_1[370].FA_  ( .A(A[1906]), .B(n2190), .CI(
        C[1906]), .CO(C[1907]) );
  FA_6282 \FA_INST_0[3].FA_INST_1[371].FA_  ( .A(A[1907]), .B(n2189), .CI(
        C[1907]), .CO(C[1908]) );
  FA_6281 \FA_INST_0[3].FA_INST_1[372].FA_  ( .A(A[1908]), .B(n2188), .CI(
        C[1908]), .CO(C[1909]) );
  FA_6280 \FA_INST_0[3].FA_INST_1[373].FA_  ( .A(A[1909]), .B(n2187), .CI(
        C[1909]), .CO(C[1910]) );
  FA_6279 \FA_INST_0[3].FA_INST_1[374].FA_  ( .A(A[1910]), .B(n2186), .CI(
        C[1910]), .CO(C[1911]) );
  FA_6278 \FA_INST_0[3].FA_INST_1[375].FA_  ( .A(A[1911]), .B(n2185), .CI(
        C[1911]), .CO(C[1912]) );
  FA_6277 \FA_INST_0[3].FA_INST_1[376].FA_  ( .A(A[1912]), .B(n2184), .CI(
        C[1912]), .CO(C[1913]) );
  FA_6276 \FA_INST_0[3].FA_INST_1[377].FA_  ( .A(A[1913]), .B(n2183), .CI(
        C[1913]), .CO(C[1914]) );
  FA_6275 \FA_INST_0[3].FA_INST_1[378].FA_  ( .A(A[1914]), .B(n2182), .CI(
        C[1914]), .CO(C[1915]) );
  FA_6274 \FA_INST_0[3].FA_INST_1[379].FA_  ( .A(A[1915]), .B(n2181), .CI(
        C[1915]), .CO(C[1916]) );
  FA_6273 \FA_INST_0[3].FA_INST_1[380].FA_  ( .A(A[1916]), .B(n2180), .CI(
        C[1916]), .CO(C[1917]) );
  FA_6272 \FA_INST_0[3].FA_INST_1[381].FA_  ( .A(A[1917]), .B(n2179), .CI(
        C[1917]), .CO(C[1918]) );
  FA_6271 \FA_INST_0[3].FA_INST_1[382].FA_  ( .A(A[1918]), .B(n2178), .CI(
        C[1918]), .CO(C[1919]) );
  FA_6270 \FA_INST_0[3].FA_INST_1[383].FA_  ( .A(A[1919]), .B(n2177), .CI(
        C[1919]), .CO(C[1920]) );
  FA_6269 \FA_INST_0[3].FA_INST_1[384].FA_  ( .A(A[1920]), .B(n2176), .CI(
        C[1920]), .CO(C[1921]) );
  FA_6268 \FA_INST_0[3].FA_INST_1[385].FA_  ( .A(A[1921]), .B(n2175), .CI(
        C[1921]), .CO(C[1922]) );
  FA_6267 \FA_INST_0[3].FA_INST_1[386].FA_  ( .A(A[1922]), .B(n2174), .CI(
        C[1922]), .CO(C[1923]) );
  FA_6266 \FA_INST_0[3].FA_INST_1[387].FA_  ( .A(A[1923]), .B(n2173), .CI(
        C[1923]), .CO(C[1924]) );
  FA_6265 \FA_INST_0[3].FA_INST_1[388].FA_  ( .A(A[1924]), .B(n2172), .CI(
        C[1924]), .CO(C[1925]) );
  FA_6264 \FA_INST_0[3].FA_INST_1[389].FA_  ( .A(A[1925]), .B(n2171), .CI(
        C[1925]), .CO(C[1926]) );
  FA_6263 \FA_INST_0[3].FA_INST_1[390].FA_  ( .A(A[1926]), .B(n2170), .CI(
        C[1926]), .CO(C[1927]) );
  FA_6262 \FA_INST_0[3].FA_INST_1[391].FA_  ( .A(A[1927]), .B(n2169), .CI(
        C[1927]), .CO(C[1928]) );
  FA_6261 \FA_INST_0[3].FA_INST_1[392].FA_  ( .A(A[1928]), .B(n2168), .CI(
        C[1928]), .CO(C[1929]) );
  FA_6260 \FA_INST_0[3].FA_INST_1[393].FA_  ( .A(A[1929]), .B(n2167), .CI(
        C[1929]), .CO(C[1930]) );
  FA_6259 \FA_INST_0[3].FA_INST_1[394].FA_  ( .A(A[1930]), .B(n2166), .CI(
        C[1930]), .CO(C[1931]) );
  FA_6258 \FA_INST_0[3].FA_INST_1[395].FA_  ( .A(A[1931]), .B(n2165), .CI(
        C[1931]), .CO(C[1932]) );
  FA_6257 \FA_INST_0[3].FA_INST_1[396].FA_  ( .A(A[1932]), .B(n2164), .CI(
        C[1932]), .CO(C[1933]) );
  FA_6256 \FA_INST_0[3].FA_INST_1[397].FA_  ( .A(A[1933]), .B(n2163), .CI(
        C[1933]), .CO(C[1934]) );
  FA_6255 \FA_INST_0[3].FA_INST_1[398].FA_  ( .A(A[1934]), .B(n2162), .CI(
        C[1934]), .CO(C[1935]) );
  FA_6254 \FA_INST_0[3].FA_INST_1[399].FA_  ( .A(A[1935]), .B(n2161), .CI(
        C[1935]), .CO(C[1936]) );
  FA_6253 \FA_INST_0[3].FA_INST_1[400].FA_  ( .A(A[1936]), .B(n2160), .CI(
        C[1936]), .CO(C[1937]) );
  FA_6252 \FA_INST_0[3].FA_INST_1[401].FA_  ( .A(A[1937]), .B(n2159), .CI(
        C[1937]), .CO(C[1938]) );
  FA_6251 \FA_INST_0[3].FA_INST_1[402].FA_  ( .A(A[1938]), .B(n2158), .CI(
        C[1938]), .CO(C[1939]) );
  FA_6250 \FA_INST_0[3].FA_INST_1[403].FA_  ( .A(A[1939]), .B(n2157), .CI(
        C[1939]), .CO(C[1940]) );
  FA_6249 \FA_INST_0[3].FA_INST_1[404].FA_  ( .A(A[1940]), .B(n2156), .CI(
        C[1940]), .CO(C[1941]) );
  FA_6248 \FA_INST_0[3].FA_INST_1[405].FA_  ( .A(A[1941]), .B(n2155), .CI(
        C[1941]), .CO(C[1942]) );
  FA_6247 \FA_INST_0[3].FA_INST_1[406].FA_  ( .A(A[1942]), .B(n2154), .CI(
        C[1942]), .CO(C[1943]) );
  FA_6246 \FA_INST_0[3].FA_INST_1[407].FA_  ( .A(A[1943]), .B(n2153), .CI(
        C[1943]), .CO(C[1944]) );
  FA_6245 \FA_INST_0[3].FA_INST_1[408].FA_  ( .A(A[1944]), .B(n2152), .CI(
        C[1944]), .CO(C[1945]) );
  FA_6244 \FA_INST_0[3].FA_INST_1[409].FA_  ( .A(A[1945]), .B(n2151), .CI(
        C[1945]), .CO(C[1946]) );
  FA_6243 \FA_INST_0[3].FA_INST_1[410].FA_  ( .A(A[1946]), .B(n2150), .CI(
        C[1946]), .CO(C[1947]) );
  FA_6242 \FA_INST_0[3].FA_INST_1[411].FA_  ( .A(A[1947]), .B(n2149), .CI(
        C[1947]), .CO(C[1948]) );
  FA_6241 \FA_INST_0[3].FA_INST_1[412].FA_  ( .A(A[1948]), .B(n2148), .CI(
        C[1948]), .CO(C[1949]) );
  FA_6240 \FA_INST_0[3].FA_INST_1[413].FA_  ( .A(A[1949]), .B(n2147), .CI(
        C[1949]), .CO(C[1950]) );
  FA_6239 \FA_INST_0[3].FA_INST_1[414].FA_  ( .A(A[1950]), .B(n2146), .CI(
        C[1950]), .CO(C[1951]) );
  FA_6238 \FA_INST_0[3].FA_INST_1[415].FA_  ( .A(A[1951]), .B(n2145), .CI(
        C[1951]), .CO(C[1952]) );
  FA_6237 \FA_INST_0[3].FA_INST_1[416].FA_  ( .A(A[1952]), .B(n2144), .CI(
        C[1952]), .CO(C[1953]) );
  FA_6236 \FA_INST_0[3].FA_INST_1[417].FA_  ( .A(A[1953]), .B(n2143), .CI(
        C[1953]), .CO(C[1954]) );
  FA_6235 \FA_INST_0[3].FA_INST_1[418].FA_  ( .A(A[1954]), .B(n2142), .CI(
        C[1954]), .CO(C[1955]) );
  FA_6234 \FA_INST_0[3].FA_INST_1[419].FA_  ( .A(A[1955]), .B(n2141), .CI(
        C[1955]), .CO(C[1956]) );
  FA_6233 \FA_INST_0[3].FA_INST_1[420].FA_  ( .A(A[1956]), .B(n2140), .CI(
        C[1956]), .CO(C[1957]) );
  FA_6232 \FA_INST_0[3].FA_INST_1[421].FA_  ( .A(A[1957]), .B(n2139), .CI(
        C[1957]), .CO(C[1958]) );
  FA_6231 \FA_INST_0[3].FA_INST_1[422].FA_  ( .A(A[1958]), .B(n2138), .CI(
        C[1958]), .CO(C[1959]) );
  FA_6230 \FA_INST_0[3].FA_INST_1[423].FA_  ( .A(A[1959]), .B(n2137), .CI(
        C[1959]), .CO(C[1960]) );
  FA_6229 \FA_INST_0[3].FA_INST_1[424].FA_  ( .A(A[1960]), .B(n2136), .CI(
        C[1960]), .CO(C[1961]) );
  FA_6228 \FA_INST_0[3].FA_INST_1[425].FA_  ( .A(A[1961]), .B(n2135), .CI(
        C[1961]), .CO(C[1962]) );
  FA_6227 \FA_INST_0[3].FA_INST_1[426].FA_  ( .A(A[1962]), .B(n2134), .CI(
        C[1962]), .CO(C[1963]) );
  FA_6226 \FA_INST_0[3].FA_INST_1[427].FA_  ( .A(A[1963]), .B(n2133), .CI(
        C[1963]), .CO(C[1964]) );
  FA_6225 \FA_INST_0[3].FA_INST_1[428].FA_  ( .A(A[1964]), .B(n2132), .CI(
        C[1964]), .CO(C[1965]) );
  FA_6224 \FA_INST_0[3].FA_INST_1[429].FA_  ( .A(A[1965]), .B(n2131), .CI(
        C[1965]), .CO(C[1966]) );
  FA_6223 \FA_INST_0[3].FA_INST_1[430].FA_  ( .A(A[1966]), .B(n2130), .CI(
        C[1966]), .CO(C[1967]) );
  FA_6222 \FA_INST_0[3].FA_INST_1[431].FA_  ( .A(A[1967]), .B(n2129), .CI(
        C[1967]), .CO(C[1968]) );
  FA_6221 \FA_INST_0[3].FA_INST_1[432].FA_  ( .A(A[1968]), .B(n2128), .CI(
        C[1968]), .CO(C[1969]) );
  FA_6220 \FA_INST_0[3].FA_INST_1[433].FA_  ( .A(A[1969]), .B(n2127), .CI(
        C[1969]), .CO(C[1970]) );
  FA_6219 \FA_INST_0[3].FA_INST_1[434].FA_  ( .A(A[1970]), .B(n2126), .CI(
        C[1970]), .CO(C[1971]) );
  FA_6218 \FA_INST_0[3].FA_INST_1[435].FA_  ( .A(A[1971]), .B(n2125), .CI(
        C[1971]), .CO(C[1972]) );
  FA_6217 \FA_INST_0[3].FA_INST_1[436].FA_  ( .A(A[1972]), .B(n2124), .CI(
        C[1972]), .CO(C[1973]) );
  FA_6216 \FA_INST_0[3].FA_INST_1[437].FA_  ( .A(A[1973]), .B(n2123), .CI(
        C[1973]), .CO(C[1974]) );
  FA_6215 \FA_INST_0[3].FA_INST_1[438].FA_  ( .A(A[1974]), .B(n2122), .CI(
        C[1974]), .CO(C[1975]) );
  FA_6214 \FA_INST_0[3].FA_INST_1[439].FA_  ( .A(A[1975]), .B(n2121), .CI(
        C[1975]), .CO(C[1976]) );
  FA_6213 \FA_INST_0[3].FA_INST_1[440].FA_  ( .A(A[1976]), .B(n2120), .CI(
        C[1976]), .CO(C[1977]) );
  FA_6212 \FA_INST_0[3].FA_INST_1[441].FA_  ( .A(A[1977]), .B(n2119), .CI(
        C[1977]), .CO(C[1978]) );
  FA_6211 \FA_INST_0[3].FA_INST_1[442].FA_  ( .A(A[1978]), .B(n2118), .CI(
        C[1978]), .CO(C[1979]) );
  FA_6210 \FA_INST_0[3].FA_INST_1[443].FA_  ( .A(A[1979]), .B(n2117), .CI(
        C[1979]), .CO(C[1980]) );
  FA_6209 \FA_INST_0[3].FA_INST_1[444].FA_  ( .A(A[1980]), .B(n2116), .CI(
        C[1980]), .CO(C[1981]) );
  FA_6208 \FA_INST_0[3].FA_INST_1[445].FA_  ( .A(A[1981]), .B(n2115), .CI(
        C[1981]), .CO(C[1982]) );
  FA_6207 \FA_INST_0[3].FA_INST_1[446].FA_  ( .A(A[1982]), .B(n2114), .CI(
        C[1982]), .CO(C[1983]) );
  FA_6206 \FA_INST_0[3].FA_INST_1[447].FA_  ( .A(A[1983]), .B(n2113), .CI(
        C[1983]), .CO(C[1984]) );
  FA_6205 \FA_INST_0[3].FA_INST_1[448].FA_  ( .A(A[1984]), .B(n2112), .CI(
        C[1984]), .CO(C[1985]) );
  FA_6204 \FA_INST_0[3].FA_INST_1[449].FA_  ( .A(A[1985]), .B(n2111), .CI(
        C[1985]), .CO(C[1986]) );
  FA_6203 \FA_INST_0[3].FA_INST_1[450].FA_  ( .A(A[1986]), .B(n2110), .CI(
        C[1986]), .CO(C[1987]) );
  FA_6202 \FA_INST_0[3].FA_INST_1[451].FA_  ( .A(A[1987]), .B(n2109), .CI(
        C[1987]), .CO(C[1988]) );
  FA_6201 \FA_INST_0[3].FA_INST_1[452].FA_  ( .A(A[1988]), .B(n2108), .CI(
        C[1988]), .CO(C[1989]) );
  FA_6200 \FA_INST_0[3].FA_INST_1[453].FA_  ( .A(A[1989]), .B(n2107), .CI(
        C[1989]), .CO(C[1990]) );
  FA_6199 \FA_INST_0[3].FA_INST_1[454].FA_  ( .A(A[1990]), .B(n2106), .CI(
        C[1990]), .CO(C[1991]) );
  FA_6198 \FA_INST_0[3].FA_INST_1[455].FA_  ( .A(A[1991]), .B(n2105), .CI(
        C[1991]), .CO(C[1992]) );
  FA_6197 \FA_INST_0[3].FA_INST_1[456].FA_  ( .A(A[1992]), .B(n2104), .CI(
        C[1992]), .CO(C[1993]) );
  FA_6196 \FA_INST_0[3].FA_INST_1[457].FA_  ( .A(A[1993]), .B(n2103), .CI(
        C[1993]), .CO(C[1994]) );
  FA_6195 \FA_INST_0[3].FA_INST_1[458].FA_  ( .A(A[1994]), .B(n2102), .CI(
        C[1994]), .CO(C[1995]) );
  FA_6194 \FA_INST_0[3].FA_INST_1[459].FA_  ( .A(A[1995]), .B(n2101), .CI(
        C[1995]), .CO(C[1996]) );
  FA_6193 \FA_INST_0[3].FA_INST_1[460].FA_  ( .A(A[1996]), .B(n2100), .CI(
        C[1996]), .CO(C[1997]) );
  FA_6192 \FA_INST_0[3].FA_INST_1[461].FA_  ( .A(A[1997]), .B(n2099), .CI(
        C[1997]), .CO(C[1998]) );
  FA_6191 \FA_INST_0[3].FA_INST_1[462].FA_  ( .A(A[1998]), .B(n2098), .CI(
        C[1998]), .CO(C[1999]) );
  FA_6190 \FA_INST_0[3].FA_INST_1[463].FA_  ( .A(A[1999]), .B(n2097), .CI(
        C[1999]), .CO(C[2000]) );
  FA_6189 \FA_INST_0[3].FA_INST_1[464].FA_  ( .A(A[2000]), .B(n2096), .CI(
        C[2000]), .CO(C[2001]) );
  FA_6188 \FA_INST_0[3].FA_INST_1[465].FA_  ( .A(A[2001]), .B(n2095), .CI(
        C[2001]), .CO(C[2002]) );
  FA_6187 \FA_INST_0[3].FA_INST_1[466].FA_  ( .A(A[2002]), .B(n2094), .CI(
        C[2002]), .CO(C[2003]) );
  FA_6186 \FA_INST_0[3].FA_INST_1[467].FA_  ( .A(A[2003]), .B(n2093), .CI(
        C[2003]), .CO(C[2004]) );
  FA_6185 \FA_INST_0[3].FA_INST_1[468].FA_  ( .A(A[2004]), .B(n2092), .CI(
        C[2004]), .CO(C[2005]) );
  FA_6184 \FA_INST_0[3].FA_INST_1[469].FA_  ( .A(A[2005]), .B(n2091), .CI(
        C[2005]), .CO(C[2006]) );
  FA_6183 \FA_INST_0[3].FA_INST_1[470].FA_  ( .A(A[2006]), .B(n2090), .CI(
        C[2006]), .CO(C[2007]) );
  FA_6182 \FA_INST_0[3].FA_INST_1[471].FA_  ( .A(A[2007]), .B(n2089), .CI(
        C[2007]), .CO(C[2008]) );
  FA_6181 \FA_INST_0[3].FA_INST_1[472].FA_  ( .A(A[2008]), .B(n2088), .CI(
        C[2008]), .CO(C[2009]) );
  FA_6180 \FA_INST_0[3].FA_INST_1[473].FA_  ( .A(A[2009]), .B(n2087), .CI(
        C[2009]), .CO(C[2010]) );
  FA_6179 \FA_INST_0[3].FA_INST_1[474].FA_  ( .A(A[2010]), .B(n2086), .CI(
        C[2010]), .CO(C[2011]) );
  FA_6178 \FA_INST_0[3].FA_INST_1[475].FA_  ( .A(A[2011]), .B(n2085), .CI(
        C[2011]), .CO(C[2012]) );
  FA_6177 \FA_INST_0[3].FA_INST_1[476].FA_  ( .A(A[2012]), .B(n2084), .CI(
        C[2012]), .CO(C[2013]) );
  FA_6176 \FA_INST_0[3].FA_INST_1[477].FA_  ( .A(A[2013]), .B(n2083), .CI(
        C[2013]), .CO(C[2014]) );
  FA_6175 \FA_INST_0[3].FA_INST_1[478].FA_  ( .A(A[2014]), .B(n2082), .CI(
        C[2014]), .CO(C[2015]) );
  FA_6174 \FA_INST_0[3].FA_INST_1[479].FA_  ( .A(A[2015]), .B(n2081), .CI(
        C[2015]), .CO(C[2016]) );
  FA_6173 \FA_INST_0[3].FA_INST_1[480].FA_  ( .A(A[2016]), .B(n2080), .CI(
        C[2016]), .CO(C[2017]) );
  FA_6172 \FA_INST_0[3].FA_INST_1[481].FA_  ( .A(A[2017]), .B(n2079), .CI(
        C[2017]), .CO(C[2018]) );
  FA_6171 \FA_INST_0[3].FA_INST_1[482].FA_  ( .A(A[2018]), .B(n2078), .CI(
        C[2018]), .CO(C[2019]) );
  FA_6170 \FA_INST_0[3].FA_INST_1[483].FA_  ( .A(A[2019]), .B(n2077), .CI(
        C[2019]), .CO(C[2020]) );
  FA_6169 \FA_INST_0[3].FA_INST_1[484].FA_  ( .A(A[2020]), .B(n2076), .CI(
        C[2020]), .CO(C[2021]) );
  FA_6168 \FA_INST_0[3].FA_INST_1[485].FA_  ( .A(A[2021]), .B(n2075), .CI(
        C[2021]), .CO(C[2022]) );
  FA_6167 \FA_INST_0[3].FA_INST_1[486].FA_  ( .A(A[2022]), .B(n2074), .CI(
        C[2022]), .CO(C[2023]) );
  FA_6166 \FA_INST_0[3].FA_INST_1[487].FA_  ( .A(A[2023]), .B(n2073), .CI(
        C[2023]), .CO(C[2024]) );
  FA_6165 \FA_INST_0[3].FA_INST_1[488].FA_  ( .A(A[2024]), .B(n2072), .CI(
        C[2024]), .CO(C[2025]) );
  FA_6164 \FA_INST_0[3].FA_INST_1[489].FA_  ( .A(A[2025]), .B(n2071), .CI(
        C[2025]), .CO(C[2026]) );
  FA_6163 \FA_INST_0[3].FA_INST_1[490].FA_  ( .A(A[2026]), .B(n2070), .CI(
        C[2026]), .CO(C[2027]) );
  FA_6162 \FA_INST_0[3].FA_INST_1[491].FA_  ( .A(A[2027]), .B(n2069), .CI(
        C[2027]), .CO(C[2028]) );
  FA_6161 \FA_INST_0[3].FA_INST_1[492].FA_  ( .A(A[2028]), .B(n2068), .CI(
        C[2028]), .CO(C[2029]) );
  FA_6160 \FA_INST_0[3].FA_INST_1[493].FA_  ( .A(A[2029]), .B(n2067), .CI(
        C[2029]), .CO(C[2030]) );
  FA_6159 \FA_INST_0[3].FA_INST_1[494].FA_  ( .A(A[2030]), .B(n2066), .CI(
        C[2030]), .CO(C[2031]) );
  FA_6158 \FA_INST_0[3].FA_INST_1[495].FA_  ( .A(A[2031]), .B(n2065), .CI(
        C[2031]), .CO(C[2032]) );
  FA_6157 \FA_INST_0[3].FA_INST_1[496].FA_  ( .A(A[2032]), .B(n2064), .CI(
        C[2032]), .CO(C[2033]) );
  FA_6156 \FA_INST_0[3].FA_INST_1[497].FA_  ( .A(A[2033]), .B(n2063), .CI(
        C[2033]), .CO(C[2034]) );
  FA_6155 \FA_INST_0[3].FA_INST_1[498].FA_  ( .A(A[2034]), .B(n2062), .CI(
        C[2034]), .CO(C[2035]) );
  FA_6154 \FA_INST_0[3].FA_INST_1[499].FA_  ( .A(A[2035]), .B(n2061), .CI(
        C[2035]), .CO(C[2036]) );
  FA_6153 \FA_INST_0[3].FA_INST_1[500].FA_  ( .A(A[2036]), .B(n2060), .CI(
        C[2036]), .CO(C[2037]) );
  FA_6152 \FA_INST_0[3].FA_INST_1[501].FA_  ( .A(A[2037]), .B(n2059), .CI(
        C[2037]), .CO(C[2038]) );
  FA_6151 \FA_INST_0[3].FA_INST_1[502].FA_  ( .A(A[2038]), .B(n2058), .CI(
        C[2038]), .CO(C[2039]) );
  FA_6150 \FA_INST_0[3].FA_INST_1[503].FA_  ( .A(A[2039]), .B(n2057), .CI(
        C[2039]), .CO(C[2040]) );
  FA_6149 \FA_INST_0[3].FA_INST_1[504].FA_  ( .A(A[2040]), .B(n2056), .CI(
        C[2040]), .CO(C[2041]) );
  FA_6148 \FA_INST_0[3].FA_INST_1[505].FA_  ( .A(A[2041]), .B(n2055), .CI(
        C[2041]), .CO(C[2042]) );
  FA_6147 \FA_INST_0[3].FA_INST_1[506].FA_  ( .A(A[2042]), .B(n2054), .CI(
        C[2042]), .CO(C[2043]) );
  FA_6146 \FA_INST_0[3].FA_INST_1[507].FA_  ( .A(A[2043]), .B(n2053), .CI(
        C[2043]), .CO(C[2044]) );
  FA_6145 \FA_INST_0[3].FA_INST_1[508].FA_  ( .A(A[2044]), .B(n2052), .CI(
        C[2044]), .CO(C[2045]) );
  FA_6144 \FA_INST_0[3].FA_INST_1[509].FA_  ( .A(A[2045]), .B(n2051), .CI(
        C[2045]), .CO(C[2046]) );
  FA_6143 \FA_INST_0[3].FA_INST_1[510].FA_  ( .A(A[2046]), .B(n2050), .CI(
        C[2046]), .CO(C[2047]) );
  FA_6142 \FA_INST_0[3].FA_INST_1[511].FA_  ( .A(A[2047]), .B(n2049), .CI(
        C[2047]), .CO(C[2048]) );
  FA_6141 \FA_INST_0[4].FA_INST_1[0].FA_  ( .A(A[2048]), .B(n2048), .CI(
        C[2048]), .CO(C[2049]) );
  FA_6140 \FA_INST_0[4].FA_INST_1[1].FA_  ( .A(A[2049]), .B(n2047), .CI(
        C[2049]), .CO(C[2050]) );
  FA_6139 \FA_INST_0[4].FA_INST_1[2].FA_  ( .A(A[2050]), .B(n2046), .CI(
        C[2050]), .CO(C[2051]) );
  FA_6138 \FA_INST_0[4].FA_INST_1[3].FA_  ( .A(A[2051]), .B(n2045), .CI(
        C[2051]), .CO(C[2052]) );
  FA_6137 \FA_INST_0[4].FA_INST_1[4].FA_  ( .A(A[2052]), .B(n2044), .CI(
        C[2052]), .CO(C[2053]) );
  FA_6136 \FA_INST_0[4].FA_INST_1[5].FA_  ( .A(A[2053]), .B(n2043), .CI(
        C[2053]), .CO(C[2054]) );
  FA_6135 \FA_INST_0[4].FA_INST_1[6].FA_  ( .A(A[2054]), .B(n2042), .CI(
        C[2054]), .CO(C[2055]) );
  FA_6134 \FA_INST_0[4].FA_INST_1[7].FA_  ( .A(A[2055]), .B(n2041), .CI(
        C[2055]), .CO(C[2056]) );
  FA_6133 \FA_INST_0[4].FA_INST_1[8].FA_  ( .A(A[2056]), .B(n2040), .CI(
        C[2056]), .CO(C[2057]) );
  FA_6132 \FA_INST_0[4].FA_INST_1[9].FA_  ( .A(A[2057]), .B(n2039), .CI(
        C[2057]), .CO(C[2058]) );
  FA_6131 \FA_INST_0[4].FA_INST_1[10].FA_  ( .A(A[2058]), .B(n2038), .CI(
        C[2058]), .CO(C[2059]) );
  FA_6130 \FA_INST_0[4].FA_INST_1[11].FA_  ( .A(A[2059]), .B(n2037), .CI(
        C[2059]), .CO(C[2060]) );
  FA_6129 \FA_INST_0[4].FA_INST_1[12].FA_  ( .A(A[2060]), .B(n2036), .CI(
        C[2060]), .CO(C[2061]) );
  FA_6128 \FA_INST_0[4].FA_INST_1[13].FA_  ( .A(A[2061]), .B(n2035), .CI(
        C[2061]), .CO(C[2062]) );
  FA_6127 \FA_INST_0[4].FA_INST_1[14].FA_  ( .A(A[2062]), .B(n2034), .CI(
        C[2062]), .CO(C[2063]) );
  FA_6126 \FA_INST_0[4].FA_INST_1[15].FA_  ( .A(A[2063]), .B(n2033), .CI(
        C[2063]), .CO(C[2064]) );
  FA_6125 \FA_INST_0[4].FA_INST_1[16].FA_  ( .A(A[2064]), .B(n2032), .CI(
        C[2064]), .CO(C[2065]) );
  FA_6124 \FA_INST_0[4].FA_INST_1[17].FA_  ( .A(A[2065]), .B(n2031), .CI(
        C[2065]), .CO(C[2066]) );
  FA_6123 \FA_INST_0[4].FA_INST_1[18].FA_  ( .A(A[2066]), .B(n2030), .CI(
        C[2066]), .CO(C[2067]) );
  FA_6122 \FA_INST_0[4].FA_INST_1[19].FA_  ( .A(A[2067]), .B(n2029), .CI(
        C[2067]), .CO(C[2068]) );
  FA_6121 \FA_INST_0[4].FA_INST_1[20].FA_  ( .A(A[2068]), .B(n2028), .CI(
        C[2068]), .CO(C[2069]) );
  FA_6120 \FA_INST_0[4].FA_INST_1[21].FA_  ( .A(A[2069]), .B(n2027), .CI(
        C[2069]), .CO(C[2070]) );
  FA_6119 \FA_INST_0[4].FA_INST_1[22].FA_  ( .A(A[2070]), .B(n2026), .CI(
        C[2070]), .CO(C[2071]) );
  FA_6118 \FA_INST_0[4].FA_INST_1[23].FA_  ( .A(A[2071]), .B(n2025), .CI(
        C[2071]), .CO(C[2072]) );
  FA_6117 \FA_INST_0[4].FA_INST_1[24].FA_  ( .A(A[2072]), .B(n2024), .CI(
        C[2072]), .CO(C[2073]) );
  FA_6116 \FA_INST_0[4].FA_INST_1[25].FA_  ( .A(A[2073]), .B(n2023), .CI(
        C[2073]), .CO(C[2074]) );
  FA_6115 \FA_INST_0[4].FA_INST_1[26].FA_  ( .A(A[2074]), .B(n2022), .CI(
        C[2074]), .CO(C[2075]) );
  FA_6114 \FA_INST_0[4].FA_INST_1[27].FA_  ( .A(A[2075]), .B(n2021), .CI(
        C[2075]), .CO(C[2076]) );
  FA_6113 \FA_INST_0[4].FA_INST_1[28].FA_  ( .A(A[2076]), .B(n2020), .CI(
        C[2076]), .CO(C[2077]) );
  FA_6112 \FA_INST_0[4].FA_INST_1[29].FA_  ( .A(A[2077]), .B(n2019), .CI(
        C[2077]), .CO(C[2078]) );
  FA_6111 \FA_INST_0[4].FA_INST_1[30].FA_  ( .A(A[2078]), .B(n2018), .CI(
        C[2078]), .CO(C[2079]) );
  FA_6110 \FA_INST_0[4].FA_INST_1[31].FA_  ( .A(A[2079]), .B(n2017), .CI(
        C[2079]), .CO(C[2080]) );
  FA_6109 \FA_INST_0[4].FA_INST_1[32].FA_  ( .A(A[2080]), .B(n2016), .CI(
        C[2080]), .CO(C[2081]) );
  FA_6108 \FA_INST_0[4].FA_INST_1[33].FA_  ( .A(A[2081]), .B(n2015), .CI(
        C[2081]), .CO(C[2082]) );
  FA_6107 \FA_INST_0[4].FA_INST_1[34].FA_  ( .A(A[2082]), .B(n2014), .CI(
        C[2082]), .CO(C[2083]) );
  FA_6106 \FA_INST_0[4].FA_INST_1[35].FA_  ( .A(A[2083]), .B(n2013), .CI(
        C[2083]), .CO(C[2084]) );
  FA_6105 \FA_INST_0[4].FA_INST_1[36].FA_  ( .A(A[2084]), .B(n2012), .CI(
        C[2084]), .CO(C[2085]) );
  FA_6104 \FA_INST_0[4].FA_INST_1[37].FA_  ( .A(A[2085]), .B(n2011), .CI(
        C[2085]), .CO(C[2086]) );
  FA_6103 \FA_INST_0[4].FA_INST_1[38].FA_  ( .A(A[2086]), .B(n2010), .CI(
        C[2086]), .CO(C[2087]) );
  FA_6102 \FA_INST_0[4].FA_INST_1[39].FA_  ( .A(A[2087]), .B(n2009), .CI(
        C[2087]), .CO(C[2088]) );
  FA_6101 \FA_INST_0[4].FA_INST_1[40].FA_  ( .A(A[2088]), .B(n2008), .CI(
        C[2088]), .CO(C[2089]) );
  FA_6100 \FA_INST_0[4].FA_INST_1[41].FA_  ( .A(A[2089]), .B(n2007), .CI(
        C[2089]), .CO(C[2090]) );
  FA_6099 \FA_INST_0[4].FA_INST_1[42].FA_  ( .A(A[2090]), .B(n2006), .CI(
        C[2090]), .CO(C[2091]) );
  FA_6098 \FA_INST_0[4].FA_INST_1[43].FA_  ( .A(A[2091]), .B(n2005), .CI(
        C[2091]), .CO(C[2092]) );
  FA_6097 \FA_INST_0[4].FA_INST_1[44].FA_  ( .A(A[2092]), .B(n2004), .CI(
        C[2092]), .CO(C[2093]) );
  FA_6096 \FA_INST_0[4].FA_INST_1[45].FA_  ( .A(A[2093]), .B(n2003), .CI(
        C[2093]), .CO(C[2094]) );
  FA_6095 \FA_INST_0[4].FA_INST_1[46].FA_  ( .A(A[2094]), .B(n2002), .CI(
        C[2094]), .CO(C[2095]) );
  FA_6094 \FA_INST_0[4].FA_INST_1[47].FA_  ( .A(A[2095]), .B(n2001), .CI(
        C[2095]), .CO(C[2096]) );
  FA_6093 \FA_INST_0[4].FA_INST_1[48].FA_  ( .A(A[2096]), .B(n2000), .CI(
        C[2096]), .CO(C[2097]) );
  FA_6092 \FA_INST_0[4].FA_INST_1[49].FA_  ( .A(A[2097]), .B(n1999), .CI(
        C[2097]), .CO(C[2098]) );
  FA_6091 \FA_INST_0[4].FA_INST_1[50].FA_  ( .A(A[2098]), .B(n1998), .CI(
        C[2098]), .CO(C[2099]) );
  FA_6090 \FA_INST_0[4].FA_INST_1[51].FA_  ( .A(A[2099]), .B(n1997), .CI(
        C[2099]), .CO(C[2100]) );
  FA_6089 \FA_INST_0[4].FA_INST_1[52].FA_  ( .A(A[2100]), .B(n1996), .CI(
        C[2100]), .CO(C[2101]) );
  FA_6088 \FA_INST_0[4].FA_INST_1[53].FA_  ( .A(A[2101]), .B(n1995), .CI(
        C[2101]), .CO(C[2102]) );
  FA_6087 \FA_INST_0[4].FA_INST_1[54].FA_  ( .A(A[2102]), .B(n1994), .CI(
        C[2102]), .CO(C[2103]) );
  FA_6086 \FA_INST_0[4].FA_INST_1[55].FA_  ( .A(A[2103]), .B(n1993), .CI(
        C[2103]), .CO(C[2104]) );
  FA_6085 \FA_INST_0[4].FA_INST_1[56].FA_  ( .A(A[2104]), .B(n1992), .CI(
        C[2104]), .CO(C[2105]) );
  FA_6084 \FA_INST_0[4].FA_INST_1[57].FA_  ( .A(A[2105]), .B(n1991), .CI(
        C[2105]), .CO(C[2106]) );
  FA_6083 \FA_INST_0[4].FA_INST_1[58].FA_  ( .A(A[2106]), .B(n1990), .CI(
        C[2106]), .CO(C[2107]) );
  FA_6082 \FA_INST_0[4].FA_INST_1[59].FA_  ( .A(A[2107]), .B(n1989), .CI(
        C[2107]), .CO(C[2108]) );
  FA_6081 \FA_INST_0[4].FA_INST_1[60].FA_  ( .A(A[2108]), .B(n1988), .CI(
        C[2108]), .CO(C[2109]) );
  FA_6080 \FA_INST_0[4].FA_INST_1[61].FA_  ( .A(A[2109]), .B(n1987), .CI(
        C[2109]), .CO(C[2110]) );
  FA_6079 \FA_INST_0[4].FA_INST_1[62].FA_  ( .A(A[2110]), .B(n1986), .CI(
        C[2110]), .CO(C[2111]) );
  FA_6078 \FA_INST_0[4].FA_INST_1[63].FA_  ( .A(A[2111]), .B(n1985), .CI(
        C[2111]), .CO(C[2112]) );
  FA_6077 \FA_INST_0[4].FA_INST_1[64].FA_  ( .A(A[2112]), .B(n1984), .CI(
        C[2112]), .CO(C[2113]) );
  FA_6076 \FA_INST_0[4].FA_INST_1[65].FA_  ( .A(A[2113]), .B(n1983), .CI(
        C[2113]), .CO(C[2114]) );
  FA_6075 \FA_INST_0[4].FA_INST_1[66].FA_  ( .A(A[2114]), .B(n1982), .CI(
        C[2114]), .CO(C[2115]) );
  FA_6074 \FA_INST_0[4].FA_INST_1[67].FA_  ( .A(A[2115]), .B(n1981), .CI(
        C[2115]), .CO(C[2116]) );
  FA_6073 \FA_INST_0[4].FA_INST_1[68].FA_  ( .A(A[2116]), .B(n1980), .CI(
        C[2116]), .CO(C[2117]) );
  FA_6072 \FA_INST_0[4].FA_INST_1[69].FA_  ( .A(A[2117]), .B(n1979), .CI(
        C[2117]), .CO(C[2118]) );
  FA_6071 \FA_INST_0[4].FA_INST_1[70].FA_  ( .A(A[2118]), .B(n1978), .CI(
        C[2118]), .CO(C[2119]) );
  FA_6070 \FA_INST_0[4].FA_INST_1[71].FA_  ( .A(A[2119]), .B(n1977), .CI(
        C[2119]), .CO(C[2120]) );
  FA_6069 \FA_INST_0[4].FA_INST_1[72].FA_  ( .A(A[2120]), .B(n1976), .CI(
        C[2120]), .CO(C[2121]) );
  FA_6068 \FA_INST_0[4].FA_INST_1[73].FA_  ( .A(A[2121]), .B(n1975), .CI(
        C[2121]), .CO(C[2122]) );
  FA_6067 \FA_INST_0[4].FA_INST_1[74].FA_  ( .A(A[2122]), .B(n1974), .CI(
        C[2122]), .CO(C[2123]) );
  FA_6066 \FA_INST_0[4].FA_INST_1[75].FA_  ( .A(A[2123]), .B(n1973), .CI(
        C[2123]), .CO(C[2124]) );
  FA_6065 \FA_INST_0[4].FA_INST_1[76].FA_  ( .A(A[2124]), .B(n1972), .CI(
        C[2124]), .CO(C[2125]) );
  FA_6064 \FA_INST_0[4].FA_INST_1[77].FA_  ( .A(A[2125]), .B(n1971), .CI(
        C[2125]), .CO(C[2126]) );
  FA_6063 \FA_INST_0[4].FA_INST_1[78].FA_  ( .A(A[2126]), .B(n1970), .CI(
        C[2126]), .CO(C[2127]) );
  FA_6062 \FA_INST_0[4].FA_INST_1[79].FA_  ( .A(A[2127]), .B(n1969), .CI(
        C[2127]), .CO(C[2128]) );
  FA_6061 \FA_INST_0[4].FA_INST_1[80].FA_  ( .A(A[2128]), .B(n1968), .CI(
        C[2128]), .CO(C[2129]) );
  FA_6060 \FA_INST_0[4].FA_INST_1[81].FA_  ( .A(A[2129]), .B(n1967), .CI(
        C[2129]), .CO(C[2130]) );
  FA_6059 \FA_INST_0[4].FA_INST_1[82].FA_  ( .A(A[2130]), .B(n1966), .CI(
        C[2130]), .CO(C[2131]) );
  FA_6058 \FA_INST_0[4].FA_INST_1[83].FA_  ( .A(A[2131]), .B(n1965), .CI(
        C[2131]), .CO(C[2132]) );
  FA_6057 \FA_INST_0[4].FA_INST_1[84].FA_  ( .A(A[2132]), .B(n1964), .CI(
        C[2132]), .CO(C[2133]) );
  FA_6056 \FA_INST_0[4].FA_INST_1[85].FA_  ( .A(A[2133]), .B(n1963), .CI(
        C[2133]), .CO(C[2134]) );
  FA_6055 \FA_INST_0[4].FA_INST_1[86].FA_  ( .A(A[2134]), .B(n1962), .CI(
        C[2134]), .CO(C[2135]) );
  FA_6054 \FA_INST_0[4].FA_INST_1[87].FA_  ( .A(A[2135]), .B(n1961), .CI(
        C[2135]), .CO(C[2136]) );
  FA_6053 \FA_INST_0[4].FA_INST_1[88].FA_  ( .A(A[2136]), .B(n1960), .CI(
        C[2136]), .CO(C[2137]) );
  FA_6052 \FA_INST_0[4].FA_INST_1[89].FA_  ( .A(A[2137]), .B(n1959), .CI(
        C[2137]), .CO(C[2138]) );
  FA_6051 \FA_INST_0[4].FA_INST_1[90].FA_  ( .A(A[2138]), .B(n1958), .CI(
        C[2138]), .CO(C[2139]) );
  FA_6050 \FA_INST_0[4].FA_INST_1[91].FA_  ( .A(A[2139]), .B(n1957), .CI(
        C[2139]), .CO(C[2140]) );
  FA_6049 \FA_INST_0[4].FA_INST_1[92].FA_  ( .A(A[2140]), .B(n1956), .CI(
        C[2140]), .CO(C[2141]) );
  FA_6048 \FA_INST_0[4].FA_INST_1[93].FA_  ( .A(A[2141]), .B(n1955), .CI(
        C[2141]), .CO(C[2142]) );
  FA_6047 \FA_INST_0[4].FA_INST_1[94].FA_  ( .A(A[2142]), .B(n1954), .CI(
        C[2142]), .CO(C[2143]) );
  FA_6046 \FA_INST_0[4].FA_INST_1[95].FA_  ( .A(A[2143]), .B(n1953), .CI(
        C[2143]), .CO(C[2144]) );
  FA_6045 \FA_INST_0[4].FA_INST_1[96].FA_  ( .A(A[2144]), .B(n1952), .CI(
        C[2144]), .CO(C[2145]) );
  FA_6044 \FA_INST_0[4].FA_INST_1[97].FA_  ( .A(A[2145]), .B(n1951), .CI(
        C[2145]), .CO(C[2146]) );
  FA_6043 \FA_INST_0[4].FA_INST_1[98].FA_  ( .A(A[2146]), .B(n1950), .CI(
        C[2146]), .CO(C[2147]) );
  FA_6042 \FA_INST_0[4].FA_INST_1[99].FA_  ( .A(A[2147]), .B(n1949), .CI(
        C[2147]), .CO(C[2148]) );
  FA_6041 \FA_INST_0[4].FA_INST_1[100].FA_  ( .A(A[2148]), .B(n1948), .CI(
        C[2148]), .CO(C[2149]) );
  FA_6040 \FA_INST_0[4].FA_INST_1[101].FA_  ( .A(A[2149]), .B(n1947), .CI(
        C[2149]), .CO(C[2150]) );
  FA_6039 \FA_INST_0[4].FA_INST_1[102].FA_  ( .A(A[2150]), .B(n1946), .CI(
        C[2150]), .CO(C[2151]) );
  FA_6038 \FA_INST_0[4].FA_INST_1[103].FA_  ( .A(A[2151]), .B(n1945), .CI(
        C[2151]), .CO(C[2152]) );
  FA_6037 \FA_INST_0[4].FA_INST_1[104].FA_  ( .A(A[2152]), .B(n1944), .CI(
        C[2152]), .CO(C[2153]) );
  FA_6036 \FA_INST_0[4].FA_INST_1[105].FA_  ( .A(A[2153]), .B(n1943), .CI(
        C[2153]), .CO(C[2154]) );
  FA_6035 \FA_INST_0[4].FA_INST_1[106].FA_  ( .A(A[2154]), .B(n1942), .CI(
        C[2154]), .CO(C[2155]) );
  FA_6034 \FA_INST_0[4].FA_INST_1[107].FA_  ( .A(A[2155]), .B(n1941), .CI(
        C[2155]), .CO(C[2156]) );
  FA_6033 \FA_INST_0[4].FA_INST_1[108].FA_  ( .A(A[2156]), .B(n1940), .CI(
        C[2156]), .CO(C[2157]) );
  FA_6032 \FA_INST_0[4].FA_INST_1[109].FA_  ( .A(A[2157]), .B(n1939), .CI(
        C[2157]), .CO(C[2158]) );
  FA_6031 \FA_INST_0[4].FA_INST_1[110].FA_  ( .A(A[2158]), .B(n1938), .CI(
        C[2158]), .CO(C[2159]) );
  FA_6030 \FA_INST_0[4].FA_INST_1[111].FA_  ( .A(A[2159]), .B(n1937), .CI(
        C[2159]), .CO(C[2160]) );
  FA_6029 \FA_INST_0[4].FA_INST_1[112].FA_  ( .A(A[2160]), .B(n1936), .CI(
        C[2160]), .CO(C[2161]) );
  FA_6028 \FA_INST_0[4].FA_INST_1[113].FA_  ( .A(A[2161]), .B(n1935), .CI(
        C[2161]), .CO(C[2162]) );
  FA_6027 \FA_INST_0[4].FA_INST_1[114].FA_  ( .A(A[2162]), .B(n1934), .CI(
        C[2162]), .CO(C[2163]) );
  FA_6026 \FA_INST_0[4].FA_INST_1[115].FA_  ( .A(A[2163]), .B(n1933), .CI(
        C[2163]), .CO(C[2164]) );
  FA_6025 \FA_INST_0[4].FA_INST_1[116].FA_  ( .A(A[2164]), .B(n1932), .CI(
        C[2164]), .CO(C[2165]) );
  FA_6024 \FA_INST_0[4].FA_INST_1[117].FA_  ( .A(A[2165]), .B(n1931), .CI(
        C[2165]), .CO(C[2166]) );
  FA_6023 \FA_INST_0[4].FA_INST_1[118].FA_  ( .A(A[2166]), .B(n1930), .CI(
        C[2166]), .CO(C[2167]) );
  FA_6022 \FA_INST_0[4].FA_INST_1[119].FA_  ( .A(A[2167]), .B(n1929), .CI(
        C[2167]), .CO(C[2168]) );
  FA_6021 \FA_INST_0[4].FA_INST_1[120].FA_  ( .A(A[2168]), .B(n1928), .CI(
        C[2168]), .CO(C[2169]) );
  FA_6020 \FA_INST_0[4].FA_INST_1[121].FA_  ( .A(A[2169]), .B(n1927), .CI(
        C[2169]), .CO(C[2170]) );
  FA_6019 \FA_INST_0[4].FA_INST_1[122].FA_  ( .A(A[2170]), .B(n1926), .CI(
        C[2170]), .CO(C[2171]) );
  FA_6018 \FA_INST_0[4].FA_INST_1[123].FA_  ( .A(A[2171]), .B(n1925), .CI(
        C[2171]), .CO(C[2172]) );
  FA_6017 \FA_INST_0[4].FA_INST_1[124].FA_  ( .A(A[2172]), .B(n1924), .CI(
        C[2172]), .CO(C[2173]) );
  FA_6016 \FA_INST_0[4].FA_INST_1[125].FA_  ( .A(A[2173]), .B(n1923), .CI(
        C[2173]), .CO(C[2174]) );
  FA_6015 \FA_INST_0[4].FA_INST_1[126].FA_  ( .A(A[2174]), .B(n1922), .CI(
        C[2174]), .CO(C[2175]) );
  FA_6014 \FA_INST_0[4].FA_INST_1[127].FA_  ( .A(A[2175]), .B(n1921), .CI(
        C[2175]), .CO(C[2176]) );
  FA_6013 \FA_INST_0[4].FA_INST_1[128].FA_  ( .A(A[2176]), .B(n1920), .CI(
        C[2176]), .CO(C[2177]) );
  FA_6012 \FA_INST_0[4].FA_INST_1[129].FA_  ( .A(A[2177]), .B(n1919), .CI(
        C[2177]), .CO(C[2178]) );
  FA_6011 \FA_INST_0[4].FA_INST_1[130].FA_  ( .A(A[2178]), .B(n1918), .CI(
        C[2178]), .CO(C[2179]) );
  FA_6010 \FA_INST_0[4].FA_INST_1[131].FA_  ( .A(A[2179]), .B(n1917), .CI(
        C[2179]), .CO(C[2180]) );
  FA_6009 \FA_INST_0[4].FA_INST_1[132].FA_  ( .A(A[2180]), .B(n1916), .CI(
        C[2180]), .CO(C[2181]) );
  FA_6008 \FA_INST_0[4].FA_INST_1[133].FA_  ( .A(A[2181]), .B(n1915), .CI(
        C[2181]), .CO(C[2182]) );
  FA_6007 \FA_INST_0[4].FA_INST_1[134].FA_  ( .A(A[2182]), .B(n1914), .CI(
        C[2182]), .CO(C[2183]) );
  FA_6006 \FA_INST_0[4].FA_INST_1[135].FA_  ( .A(A[2183]), .B(n1913), .CI(
        C[2183]), .CO(C[2184]) );
  FA_6005 \FA_INST_0[4].FA_INST_1[136].FA_  ( .A(A[2184]), .B(n1912), .CI(
        C[2184]), .CO(C[2185]) );
  FA_6004 \FA_INST_0[4].FA_INST_1[137].FA_  ( .A(A[2185]), .B(n1911), .CI(
        C[2185]), .CO(C[2186]) );
  FA_6003 \FA_INST_0[4].FA_INST_1[138].FA_  ( .A(A[2186]), .B(n1910), .CI(
        C[2186]), .CO(C[2187]) );
  FA_6002 \FA_INST_0[4].FA_INST_1[139].FA_  ( .A(A[2187]), .B(n1909), .CI(
        C[2187]), .CO(C[2188]) );
  FA_6001 \FA_INST_0[4].FA_INST_1[140].FA_  ( .A(A[2188]), .B(n1908), .CI(
        C[2188]), .CO(C[2189]) );
  FA_6000 \FA_INST_0[4].FA_INST_1[141].FA_  ( .A(A[2189]), .B(n1907), .CI(
        C[2189]), .CO(C[2190]) );
  FA_5999 \FA_INST_0[4].FA_INST_1[142].FA_  ( .A(A[2190]), .B(n1906), .CI(
        C[2190]), .CO(C[2191]) );
  FA_5998 \FA_INST_0[4].FA_INST_1[143].FA_  ( .A(A[2191]), .B(n1905), .CI(
        C[2191]), .CO(C[2192]) );
  FA_5997 \FA_INST_0[4].FA_INST_1[144].FA_  ( .A(A[2192]), .B(n1904), .CI(
        C[2192]), .CO(C[2193]) );
  FA_5996 \FA_INST_0[4].FA_INST_1[145].FA_  ( .A(A[2193]), .B(n1903), .CI(
        C[2193]), .CO(C[2194]) );
  FA_5995 \FA_INST_0[4].FA_INST_1[146].FA_  ( .A(A[2194]), .B(n1902), .CI(
        C[2194]), .CO(C[2195]) );
  FA_5994 \FA_INST_0[4].FA_INST_1[147].FA_  ( .A(A[2195]), .B(n1901), .CI(
        C[2195]), .CO(C[2196]) );
  FA_5993 \FA_INST_0[4].FA_INST_1[148].FA_  ( .A(A[2196]), .B(n1900), .CI(
        C[2196]), .CO(C[2197]) );
  FA_5992 \FA_INST_0[4].FA_INST_1[149].FA_  ( .A(A[2197]), .B(n1899), .CI(
        C[2197]), .CO(C[2198]) );
  FA_5991 \FA_INST_0[4].FA_INST_1[150].FA_  ( .A(A[2198]), .B(n1898), .CI(
        C[2198]), .CO(C[2199]) );
  FA_5990 \FA_INST_0[4].FA_INST_1[151].FA_  ( .A(A[2199]), .B(n1897), .CI(
        C[2199]), .CO(C[2200]) );
  FA_5989 \FA_INST_0[4].FA_INST_1[152].FA_  ( .A(A[2200]), .B(n1896), .CI(
        C[2200]), .CO(C[2201]) );
  FA_5988 \FA_INST_0[4].FA_INST_1[153].FA_  ( .A(A[2201]), .B(n1895), .CI(
        C[2201]), .CO(C[2202]) );
  FA_5987 \FA_INST_0[4].FA_INST_1[154].FA_  ( .A(A[2202]), .B(n1894), .CI(
        C[2202]), .CO(C[2203]) );
  FA_5986 \FA_INST_0[4].FA_INST_1[155].FA_  ( .A(A[2203]), .B(n1893), .CI(
        C[2203]), .CO(C[2204]) );
  FA_5985 \FA_INST_0[4].FA_INST_1[156].FA_  ( .A(A[2204]), .B(n1892), .CI(
        C[2204]), .CO(C[2205]) );
  FA_5984 \FA_INST_0[4].FA_INST_1[157].FA_  ( .A(A[2205]), .B(n1891), .CI(
        C[2205]), .CO(C[2206]) );
  FA_5983 \FA_INST_0[4].FA_INST_1[158].FA_  ( .A(A[2206]), .B(n1890), .CI(
        C[2206]), .CO(C[2207]) );
  FA_5982 \FA_INST_0[4].FA_INST_1[159].FA_  ( .A(A[2207]), .B(n1889), .CI(
        C[2207]), .CO(C[2208]) );
  FA_5981 \FA_INST_0[4].FA_INST_1[160].FA_  ( .A(A[2208]), .B(n1888), .CI(
        C[2208]), .CO(C[2209]) );
  FA_5980 \FA_INST_0[4].FA_INST_1[161].FA_  ( .A(A[2209]), .B(n1887), .CI(
        C[2209]), .CO(C[2210]) );
  FA_5979 \FA_INST_0[4].FA_INST_1[162].FA_  ( .A(A[2210]), .B(n1886), .CI(
        C[2210]), .CO(C[2211]) );
  FA_5978 \FA_INST_0[4].FA_INST_1[163].FA_  ( .A(A[2211]), .B(n1885), .CI(
        C[2211]), .CO(C[2212]) );
  FA_5977 \FA_INST_0[4].FA_INST_1[164].FA_  ( .A(A[2212]), .B(n1884), .CI(
        C[2212]), .CO(C[2213]) );
  FA_5976 \FA_INST_0[4].FA_INST_1[165].FA_  ( .A(A[2213]), .B(n1883), .CI(
        C[2213]), .CO(C[2214]) );
  FA_5975 \FA_INST_0[4].FA_INST_1[166].FA_  ( .A(A[2214]), .B(n1882), .CI(
        C[2214]), .CO(C[2215]) );
  FA_5974 \FA_INST_0[4].FA_INST_1[167].FA_  ( .A(A[2215]), .B(n1881), .CI(
        C[2215]), .CO(C[2216]) );
  FA_5973 \FA_INST_0[4].FA_INST_1[168].FA_  ( .A(A[2216]), .B(n1880), .CI(
        C[2216]), .CO(C[2217]) );
  FA_5972 \FA_INST_0[4].FA_INST_1[169].FA_  ( .A(A[2217]), .B(n1879), .CI(
        C[2217]), .CO(C[2218]) );
  FA_5971 \FA_INST_0[4].FA_INST_1[170].FA_  ( .A(A[2218]), .B(n1878), .CI(
        C[2218]), .CO(C[2219]) );
  FA_5970 \FA_INST_0[4].FA_INST_1[171].FA_  ( .A(A[2219]), .B(n1877), .CI(
        C[2219]), .CO(C[2220]) );
  FA_5969 \FA_INST_0[4].FA_INST_1[172].FA_  ( .A(A[2220]), .B(n1876), .CI(
        C[2220]), .CO(C[2221]) );
  FA_5968 \FA_INST_0[4].FA_INST_1[173].FA_  ( .A(A[2221]), .B(n1875), .CI(
        C[2221]), .CO(C[2222]) );
  FA_5967 \FA_INST_0[4].FA_INST_1[174].FA_  ( .A(A[2222]), .B(n1874), .CI(
        C[2222]), .CO(C[2223]) );
  FA_5966 \FA_INST_0[4].FA_INST_1[175].FA_  ( .A(A[2223]), .B(n1873), .CI(
        C[2223]), .CO(C[2224]) );
  FA_5965 \FA_INST_0[4].FA_INST_1[176].FA_  ( .A(A[2224]), .B(n1872), .CI(
        C[2224]), .CO(C[2225]) );
  FA_5964 \FA_INST_0[4].FA_INST_1[177].FA_  ( .A(A[2225]), .B(n1871), .CI(
        C[2225]), .CO(C[2226]) );
  FA_5963 \FA_INST_0[4].FA_INST_1[178].FA_  ( .A(A[2226]), .B(n1870), .CI(
        C[2226]), .CO(C[2227]) );
  FA_5962 \FA_INST_0[4].FA_INST_1[179].FA_  ( .A(A[2227]), .B(n1869), .CI(
        C[2227]), .CO(C[2228]) );
  FA_5961 \FA_INST_0[4].FA_INST_1[180].FA_  ( .A(A[2228]), .B(n1868), .CI(
        C[2228]), .CO(C[2229]) );
  FA_5960 \FA_INST_0[4].FA_INST_1[181].FA_  ( .A(A[2229]), .B(n1867), .CI(
        C[2229]), .CO(C[2230]) );
  FA_5959 \FA_INST_0[4].FA_INST_1[182].FA_  ( .A(A[2230]), .B(n1866), .CI(
        C[2230]), .CO(C[2231]) );
  FA_5958 \FA_INST_0[4].FA_INST_1[183].FA_  ( .A(A[2231]), .B(n1865), .CI(
        C[2231]), .CO(C[2232]) );
  FA_5957 \FA_INST_0[4].FA_INST_1[184].FA_  ( .A(A[2232]), .B(n1864), .CI(
        C[2232]), .CO(C[2233]) );
  FA_5956 \FA_INST_0[4].FA_INST_1[185].FA_  ( .A(A[2233]), .B(n1863), .CI(
        C[2233]), .CO(C[2234]) );
  FA_5955 \FA_INST_0[4].FA_INST_1[186].FA_  ( .A(A[2234]), .B(n1862), .CI(
        C[2234]), .CO(C[2235]) );
  FA_5954 \FA_INST_0[4].FA_INST_1[187].FA_  ( .A(A[2235]), .B(n1861), .CI(
        C[2235]), .CO(C[2236]) );
  FA_5953 \FA_INST_0[4].FA_INST_1[188].FA_  ( .A(A[2236]), .B(n1860), .CI(
        C[2236]), .CO(C[2237]) );
  FA_5952 \FA_INST_0[4].FA_INST_1[189].FA_  ( .A(A[2237]), .B(n1859), .CI(
        C[2237]), .CO(C[2238]) );
  FA_5951 \FA_INST_0[4].FA_INST_1[190].FA_  ( .A(A[2238]), .B(n1858), .CI(
        C[2238]), .CO(C[2239]) );
  FA_5950 \FA_INST_0[4].FA_INST_1[191].FA_  ( .A(A[2239]), .B(n1857), .CI(
        C[2239]), .CO(C[2240]) );
  FA_5949 \FA_INST_0[4].FA_INST_1[192].FA_  ( .A(A[2240]), .B(n1856), .CI(
        C[2240]), .CO(C[2241]) );
  FA_5948 \FA_INST_0[4].FA_INST_1[193].FA_  ( .A(A[2241]), .B(n1855), .CI(
        C[2241]), .CO(C[2242]) );
  FA_5947 \FA_INST_0[4].FA_INST_1[194].FA_  ( .A(A[2242]), .B(n1854), .CI(
        C[2242]), .CO(C[2243]) );
  FA_5946 \FA_INST_0[4].FA_INST_1[195].FA_  ( .A(A[2243]), .B(n1853), .CI(
        C[2243]), .CO(C[2244]) );
  FA_5945 \FA_INST_0[4].FA_INST_1[196].FA_  ( .A(A[2244]), .B(n1852), .CI(
        C[2244]), .CO(C[2245]) );
  FA_5944 \FA_INST_0[4].FA_INST_1[197].FA_  ( .A(A[2245]), .B(n1851), .CI(
        C[2245]), .CO(C[2246]) );
  FA_5943 \FA_INST_0[4].FA_INST_1[198].FA_  ( .A(A[2246]), .B(n1850), .CI(
        C[2246]), .CO(C[2247]) );
  FA_5942 \FA_INST_0[4].FA_INST_1[199].FA_  ( .A(A[2247]), .B(n1849), .CI(
        C[2247]), .CO(C[2248]) );
  FA_5941 \FA_INST_0[4].FA_INST_1[200].FA_  ( .A(A[2248]), .B(n1848), .CI(
        C[2248]), .CO(C[2249]) );
  FA_5940 \FA_INST_0[4].FA_INST_1[201].FA_  ( .A(A[2249]), .B(n1847), .CI(
        C[2249]), .CO(C[2250]) );
  FA_5939 \FA_INST_0[4].FA_INST_1[202].FA_  ( .A(A[2250]), .B(n1846), .CI(
        C[2250]), .CO(C[2251]) );
  FA_5938 \FA_INST_0[4].FA_INST_1[203].FA_  ( .A(A[2251]), .B(n1845), .CI(
        C[2251]), .CO(C[2252]) );
  FA_5937 \FA_INST_0[4].FA_INST_1[204].FA_  ( .A(A[2252]), .B(n1844), .CI(
        C[2252]), .CO(C[2253]) );
  FA_5936 \FA_INST_0[4].FA_INST_1[205].FA_  ( .A(A[2253]), .B(n1843), .CI(
        C[2253]), .CO(C[2254]) );
  FA_5935 \FA_INST_0[4].FA_INST_1[206].FA_  ( .A(A[2254]), .B(n1842), .CI(
        C[2254]), .CO(C[2255]) );
  FA_5934 \FA_INST_0[4].FA_INST_1[207].FA_  ( .A(A[2255]), .B(n1841), .CI(
        C[2255]), .CO(C[2256]) );
  FA_5933 \FA_INST_0[4].FA_INST_1[208].FA_  ( .A(A[2256]), .B(n1840), .CI(
        C[2256]), .CO(C[2257]) );
  FA_5932 \FA_INST_0[4].FA_INST_1[209].FA_  ( .A(A[2257]), .B(n1839), .CI(
        C[2257]), .CO(C[2258]) );
  FA_5931 \FA_INST_0[4].FA_INST_1[210].FA_  ( .A(A[2258]), .B(n1838), .CI(
        C[2258]), .CO(C[2259]) );
  FA_5930 \FA_INST_0[4].FA_INST_1[211].FA_  ( .A(A[2259]), .B(n1837), .CI(
        C[2259]), .CO(C[2260]) );
  FA_5929 \FA_INST_0[4].FA_INST_1[212].FA_  ( .A(A[2260]), .B(n1836), .CI(
        C[2260]), .CO(C[2261]) );
  FA_5928 \FA_INST_0[4].FA_INST_1[213].FA_  ( .A(A[2261]), .B(n1835), .CI(
        C[2261]), .CO(C[2262]) );
  FA_5927 \FA_INST_0[4].FA_INST_1[214].FA_  ( .A(A[2262]), .B(n1834), .CI(
        C[2262]), .CO(C[2263]) );
  FA_5926 \FA_INST_0[4].FA_INST_1[215].FA_  ( .A(A[2263]), .B(n1833), .CI(
        C[2263]), .CO(C[2264]) );
  FA_5925 \FA_INST_0[4].FA_INST_1[216].FA_  ( .A(A[2264]), .B(n1832), .CI(
        C[2264]), .CO(C[2265]) );
  FA_5924 \FA_INST_0[4].FA_INST_1[217].FA_  ( .A(A[2265]), .B(n1831), .CI(
        C[2265]), .CO(C[2266]) );
  FA_5923 \FA_INST_0[4].FA_INST_1[218].FA_  ( .A(A[2266]), .B(n1830), .CI(
        C[2266]), .CO(C[2267]) );
  FA_5922 \FA_INST_0[4].FA_INST_1[219].FA_  ( .A(A[2267]), .B(n1829), .CI(
        C[2267]), .CO(C[2268]) );
  FA_5921 \FA_INST_0[4].FA_INST_1[220].FA_  ( .A(A[2268]), .B(n1828), .CI(
        C[2268]), .CO(C[2269]) );
  FA_5920 \FA_INST_0[4].FA_INST_1[221].FA_  ( .A(A[2269]), .B(n1827), .CI(
        C[2269]), .CO(C[2270]) );
  FA_5919 \FA_INST_0[4].FA_INST_1[222].FA_  ( .A(A[2270]), .B(n1826), .CI(
        C[2270]), .CO(C[2271]) );
  FA_5918 \FA_INST_0[4].FA_INST_1[223].FA_  ( .A(A[2271]), .B(n1825), .CI(
        C[2271]), .CO(C[2272]) );
  FA_5917 \FA_INST_0[4].FA_INST_1[224].FA_  ( .A(A[2272]), .B(n1824), .CI(
        C[2272]), .CO(C[2273]) );
  FA_5916 \FA_INST_0[4].FA_INST_1[225].FA_  ( .A(A[2273]), .B(n1823), .CI(
        C[2273]), .CO(C[2274]) );
  FA_5915 \FA_INST_0[4].FA_INST_1[226].FA_  ( .A(A[2274]), .B(n1822), .CI(
        C[2274]), .CO(C[2275]) );
  FA_5914 \FA_INST_0[4].FA_INST_1[227].FA_  ( .A(A[2275]), .B(n1821), .CI(
        C[2275]), .CO(C[2276]) );
  FA_5913 \FA_INST_0[4].FA_INST_1[228].FA_  ( .A(A[2276]), .B(n1820), .CI(
        C[2276]), .CO(C[2277]) );
  FA_5912 \FA_INST_0[4].FA_INST_1[229].FA_  ( .A(A[2277]), .B(n1819), .CI(
        C[2277]), .CO(C[2278]) );
  FA_5911 \FA_INST_0[4].FA_INST_1[230].FA_  ( .A(A[2278]), .B(n1818), .CI(
        C[2278]), .CO(C[2279]) );
  FA_5910 \FA_INST_0[4].FA_INST_1[231].FA_  ( .A(A[2279]), .B(n1817), .CI(
        C[2279]), .CO(C[2280]) );
  FA_5909 \FA_INST_0[4].FA_INST_1[232].FA_  ( .A(A[2280]), .B(n1816), .CI(
        C[2280]), .CO(C[2281]) );
  FA_5908 \FA_INST_0[4].FA_INST_1[233].FA_  ( .A(A[2281]), .B(n1815), .CI(
        C[2281]), .CO(C[2282]) );
  FA_5907 \FA_INST_0[4].FA_INST_1[234].FA_  ( .A(A[2282]), .B(n1814), .CI(
        C[2282]), .CO(C[2283]) );
  FA_5906 \FA_INST_0[4].FA_INST_1[235].FA_  ( .A(A[2283]), .B(n1813), .CI(
        C[2283]), .CO(C[2284]) );
  FA_5905 \FA_INST_0[4].FA_INST_1[236].FA_  ( .A(A[2284]), .B(n1812), .CI(
        C[2284]), .CO(C[2285]) );
  FA_5904 \FA_INST_0[4].FA_INST_1[237].FA_  ( .A(A[2285]), .B(n1811), .CI(
        C[2285]), .CO(C[2286]) );
  FA_5903 \FA_INST_0[4].FA_INST_1[238].FA_  ( .A(A[2286]), .B(n1810), .CI(
        C[2286]), .CO(C[2287]) );
  FA_5902 \FA_INST_0[4].FA_INST_1[239].FA_  ( .A(A[2287]), .B(n1809), .CI(
        C[2287]), .CO(C[2288]) );
  FA_5901 \FA_INST_0[4].FA_INST_1[240].FA_  ( .A(A[2288]), .B(n1808), .CI(
        C[2288]), .CO(C[2289]) );
  FA_5900 \FA_INST_0[4].FA_INST_1[241].FA_  ( .A(A[2289]), .B(n1807), .CI(
        C[2289]), .CO(C[2290]) );
  FA_5899 \FA_INST_0[4].FA_INST_1[242].FA_  ( .A(A[2290]), .B(n1806), .CI(
        C[2290]), .CO(C[2291]) );
  FA_5898 \FA_INST_0[4].FA_INST_1[243].FA_  ( .A(A[2291]), .B(n1805), .CI(
        C[2291]), .CO(C[2292]) );
  FA_5897 \FA_INST_0[4].FA_INST_1[244].FA_  ( .A(A[2292]), .B(n1804), .CI(
        C[2292]), .CO(C[2293]) );
  FA_5896 \FA_INST_0[4].FA_INST_1[245].FA_  ( .A(A[2293]), .B(n1803), .CI(
        C[2293]), .CO(C[2294]) );
  FA_5895 \FA_INST_0[4].FA_INST_1[246].FA_  ( .A(A[2294]), .B(n1802), .CI(
        C[2294]), .CO(C[2295]) );
  FA_5894 \FA_INST_0[4].FA_INST_1[247].FA_  ( .A(A[2295]), .B(n1801), .CI(
        C[2295]), .CO(C[2296]) );
  FA_5893 \FA_INST_0[4].FA_INST_1[248].FA_  ( .A(A[2296]), .B(n1800), .CI(
        C[2296]), .CO(C[2297]) );
  FA_5892 \FA_INST_0[4].FA_INST_1[249].FA_  ( .A(A[2297]), .B(n1799), .CI(
        C[2297]), .CO(C[2298]) );
  FA_5891 \FA_INST_0[4].FA_INST_1[250].FA_  ( .A(A[2298]), .B(n1798), .CI(
        C[2298]), .CO(C[2299]) );
  FA_5890 \FA_INST_0[4].FA_INST_1[251].FA_  ( .A(A[2299]), .B(n1797), .CI(
        C[2299]), .CO(C[2300]) );
  FA_5889 \FA_INST_0[4].FA_INST_1[252].FA_  ( .A(A[2300]), .B(n1796), .CI(
        C[2300]), .CO(C[2301]) );
  FA_5888 \FA_INST_0[4].FA_INST_1[253].FA_  ( .A(A[2301]), .B(n1795), .CI(
        C[2301]), .CO(C[2302]) );
  FA_5887 \FA_INST_0[4].FA_INST_1[254].FA_  ( .A(A[2302]), .B(n1794), .CI(
        C[2302]), .CO(C[2303]) );
  FA_5886 \FA_INST_0[4].FA_INST_1[255].FA_  ( .A(A[2303]), .B(n1793), .CI(
        C[2303]), .CO(C[2304]) );
  FA_5885 \FA_INST_0[4].FA_INST_1[256].FA_  ( .A(A[2304]), .B(n1792), .CI(
        C[2304]), .CO(C[2305]) );
  FA_5884 \FA_INST_0[4].FA_INST_1[257].FA_  ( .A(A[2305]), .B(n1791), .CI(
        C[2305]), .CO(C[2306]) );
  FA_5883 \FA_INST_0[4].FA_INST_1[258].FA_  ( .A(A[2306]), .B(n1790), .CI(
        C[2306]), .CO(C[2307]) );
  FA_5882 \FA_INST_0[4].FA_INST_1[259].FA_  ( .A(A[2307]), .B(n1789), .CI(
        C[2307]), .CO(C[2308]) );
  FA_5881 \FA_INST_0[4].FA_INST_1[260].FA_  ( .A(A[2308]), .B(n1788), .CI(
        C[2308]), .CO(C[2309]) );
  FA_5880 \FA_INST_0[4].FA_INST_1[261].FA_  ( .A(A[2309]), .B(n1787), .CI(
        C[2309]), .CO(C[2310]) );
  FA_5879 \FA_INST_0[4].FA_INST_1[262].FA_  ( .A(A[2310]), .B(n1786), .CI(
        C[2310]), .CO(C[2311]) );
  FA_5878 \FA_INST_0[4].FA_INST_1[263].FA_  ( .A(A[2311]), .B(n1785), .CI(
        C[2311]), .CO(C[2312]) );
  FA_5877 \FA_INST_0[4].FA_INST_1[264].FA_  ( .A(A[2312]), .B(n1784), .CI(
        C[2312]), .CO(C[2313]) );
  FA_5876 \FA_INST_0[4].FA_INST_1[265].FA_  ( .A(A[2313]), .B(n1783), .CI(
        C[2313]), .CO(C[2314]) );
  FA_5875 \FA_INST_0[4].FA_INST_1[266].FA_  ( .A(A[2314]), .B(n1782), .CI(
        C[2314]), .CO(C[2315]) );
  FA_5874 \FA_INST_0[4].FA_INST_1[267].FA_  ( .A(A[2315]), .B(n1781), .CI(
        C[2315]), .CO(C[2316]) );
  FA_5873 \FA_INST_0[4].FA_INST_1[268].FA_  ( .A(A[2316]), .B(n1780), .CI(
        C[2316]), .CO(C[2317]) );
  FA_5872 \FA_INST_0[4].FA_INST_1[269].FA_  ( .A(A[2317]), .B(n1779), .CI(
        C[2317]), .CO(C[2318]) );
  FA_5871 \FA_INST_0[4].FA_INST_1[270].FA_  ( .A(A[2318]), .B(n1778), .CI(
        C[2318]), .CO(C[2319]) );
  FA_5870 \FA_INST_0[4].FA_INST_1[271].FA_  ( .A(A[2319]), .B(n1777), .CI(
        C[2319]), .CO(C[2320]) );
  FA_5869 \FA_INST_0[4].FA_INST_1[272].FA_  ( .A(A[2320]), .B(n1776), .CI(
        C[2320]), .CO(C[2321]) );
  FA_5868 \FA_INST_0[4].FA_INST_1[273].FA_  ( .A(A[2321]), .B(n1775), .CI(
        C[2321]), .CO(C[2322]) );
  FA_5867 \FA_INST_0[4].FA_INST_1[274].FA_  ( .A(A[2322]), .B(n1774), .CI(
        C[2322]), .CO(C[2323]) );
  FA_5866 \FA_INST_0[4].FA_INST_1[275].FA_  ( .A(A[2323]), .B(n1773), .CI(
        C[2323]), .CO(C[2324]) );
  FA_5865 \FA_INST_0[4].FA_INST_1[276].FA_  ( .A(A[2324]), .B(n1772), .CI(
        C[2324]), .CO(C[2325]) );
  FA_5864 \FA_INST_0[4].FA_INST_1[277].FA_  ( .A(A[2325]), .B(n1771), .CI(
        C[2325]), .CO(C[2326]) );
  FA_5863 \FA_INST_0[4].FA_INST_1[278].FA_  ( .A(A[2326]), .B(n1770), .CI(
        C[2326]), .CO(C[2327]) );
  FA_5862 \FA_INST_0[4].FA_INST_1[279].FA_  ( .A(A[2327]), .B(n1769), .CI(
        C[2327]), .CO(C[2328]) );
  FA_5861 \FA_INST_0[4].FA_INST_1[280].FA_  ( .A(A[2328]), .B(n1768), .CI(
        C[2328]), .CO(C[2329]) );
  FA_5860 \FA_INST_0[4].FA_INST_1[281].FA_  ( .A(A[2329]), .B(n1767), .CI(
        C[2329]), .CO(C[2330]) );
  FA_5859 \FA_INST_0[4].FA_INST_1[282].FA_  ( .A(A[2330]), .B(n1766), .CI(
        C[2330]), .CO(C[2331]) );
  FA_5858 \FA_INST_0[4].FA_INST_1[283].FA_  ( .A(A[2331]), .B(n1765), .CI(
        C[2331]), .CO(C[2332]) );
  FA_5857 \FA_INST_0[4].FA_INST_1[284].FA_  ( .A(A[2332]), .B(n1764), .CI(
        C[2332]), .CO(C[2333]) );
  FA_5856 \FA_INST_0[4].FA_INST_1[285].FA_  ( .A(A[2333]), .B(n1763), .CI(
        C[2333]), .CO(C[2334]) );
  FA_5855 \FA_INST_0[4].FA_INST_1[286].FA_  ( .A(A[2334]), .B(n1762), .CI(
        C[2334]), .CO(C[2335]) );
  FA_5854 \FA_INST_0[4].FA_INST_1[287].FA_  ( .A(A[2335]), .B(n1761), .CI(
        C[2335]), .CO(C[2336]) );
  FA_5853 \FA_INST_0[4].FA_INST_1[288].FA_  ( .A(A[2336]), .B(n1760), .CI(
        C[2336]), .CO(C[2337]) );
  FA_5852 \FA_INST_0[4].FA_INST_1[289].FA_  ( .A(A[2337]), .B(n1759), .CI(
        C[2337]), .CO(C[2338]) );
  FA_5851 \FA_INST_0[4].FA_INST_1[290].FA_  ( .A(A[2338]), .B(n1758), .CI(
        C[2338]), .CO(C[2339]) );
  FA_5850 \FA_INST_0[4].FA_INST_1[291].FA_  ( .A(A[2339]), .B(n1757), .CI(
        C[2339]), .CO(C[2340]) );
  FA_5849 \FA_INST_0[4].FA_INST_1[292].FA_  ( .A(A[2340]), .B(n1756), .CI(
        C[2340]), .CO(C[2341]) );
  FA_5848 \FA_INST_0[4].FA_INST_1[293].FA_  ( .A(A[2341]), .B(n1755), .CI(
        C[2341]), .CO(C[2342]) );
  FA_5847 \FA_INST_0[4].FA_INST_1[294].FA_  ( .A(A[2342]), .B(n1754), .CI(
        C[2342]), .CO(C[2343]) );
  FA_5846 \FA_INST_0[4].FA_INST_1[295].FA_  ( .A(A[2343]), .B(n1753), .CI(
        C[2343]), .CO(C[2344]) );
  FA_5845 \FA_INST_0[4].FA_INST_1[296].FA_  ( .A(A[2344]), .B(n1752), .CI(
        C[2344]), .CO(C[2345]) );
  FA_5844 \FA_INST_0[4].FA_INST_1[297].FA_  ( .A(A[2345]), .B(n1751), .CI(
        C[2345]), .CO(C[2346]) );
  FA_5843 \FA_INST_0[4].FA_INST_1[298].FA_  ( .A(A[2346]), .B(n1750), .CI(
        C[2346]), .CO(C[2347]) );
  FA_5842 \FA_INST_0[4].FA_INST_1[299].FA_  ( .A(A[2347]), .B(n1749), .CI(
        C[2347]), .CO(C[2348]) );
  FA_5841 \FA_INST_0[4].FA_INST_1[300].FA_  ( .A(A[2348]), .B(n1748), .CI(
        C[2348]), .CO(C[2349]) );
  FA_5840 \FA_INST_0[4].FA_INST_1[301].FA_  ( .A(A[2349]), .B(n1747), .CI(
        C[2349]), .CO(C[2350]) );
  FA_5839 \FA_INST_0[4].FA_INST_1[302].FA_  ( .A(A[2350]), .B(n1746), .CI(
        C[2350]), .CO(C[2351]) );
  FA_5838 \FA_INST_0[4].FA_INST_1[303].FA_  ( .A(A[2351]), .B(n1745), .CI(
        C[2351]), .CO(C[2352]) );
  FA_5837 \FA_INST_0[4].FA_INST_1[304].FA_  ( .A(A[2352]), .B(n1744), .CI(
        C[2352]), .CO(C[2353]) );
  FA_5836 \FA_INST_0[4].FA_INST_1[305].FA_  ( .A(A[2353]), .B(n1743), .CI(
        C[2353]), .CO(C[2354]) );
  FA_5835 \FA_INST_0[4].FA_INST_1[306].FA_  ( .A(A[2354]), .B(n1742), .CI(
        C[2354]), .CO(C[2355]) );
  FA_5834 \FA_INST_0[4].FA_INST_1[307].FA_  ( .A(A[2355]), .B(n1741), .CI(
        C[2355]), .CO(C[2356]) );
  FA_5833 \FA_INST_0[4].FA_INST_1[308].FA_  ( .A(A[2356]), .B(n1740), .CI(
        C[2356]), .CO(C[2357]) );
  FA_5832 \FA_INST_0[4].FA_INST_1[309].FA_  ( .A(A[2357]), .B(n1739), .CI(
        C[2357]), .CO(C[2358]) );
  FA_5831 \FA_INST_0[4].FA_INST_1[310].FA_  ( .A(A[2358]), .B(n1738), .CI(
        C[2358]), .CO(C[2359]) );
  FA_5830 \FA_INST_0[4].FA_INST_1[311].FA_  ( .A(A[2359]), .B(n1737), .CI(
        C[2359]), .CO(C[2360]) );
  FA_5829 \FA_INST_0[4].FA_INST_1[312].FA_  ( .A(A[2360]), .B(n1736), .CI(
        C[2360]), .CO(C[2361]) );
  FA_5828 \FA_INST_0[4].FA_INST_1[313].FA_  ( .A(A[2361]), .B(n1735), .CI(
        C[2361]), .CO(C[2362]) );
  FA_5827 \FA_INST_0[4].FA_INST_1[314].FA_  ( .A(A[2362]), .B(n1734), .CI(
        C[2362]), .CO(C[2363]) );
  FA_5826 \FA_INST_0[4].FA_INST_1[315].FA_  ( .A(A[2363]), .B(n1733), .CI(
        C[2363]), .CO(C[2364]) );
  FA_5825 \FA_INST_0[4].FA_INST_1[316].FA_  ( .A(A[2364]), .B(n1732), .CI(
        C[2364]), .CO(C[2365]) );
  FA_5824 \FA_INST_0[4].FA_INST_1[317].FA_  ( .A(A[2365]), .B(n1731), .CI(
        C[2365]), .CO(C[2366]) );
  FA_5823 \FA_INST_0[4].FA_INST_1[318].FA_  ( .A(A[2366]), .B(n1730), .CI(
        C[2366]), .CO(C[2367]) );
  FA_5822 \FA_INST_0[4].FA_INST_1[319].FA_  ( .A(A[2367]), .B(n1729), .CI(
        C[2367]), .CO(C[2368]) );
  FA_5821 \FA_INST_0[4].FA_INST_1[320].FA_  ( .A(A[2368]), .B(n1728), .CI(
        C[2368]), .CO(C[2369]) );
  FA_5820 \FA_INST_0[4].FA_INST_1[321].FA_  ( .A(A[2369]), .B(n1727), .CI(
        C[2369]), .CO(C[2370]) );
  FA_5819 \FA_INST_0[4].FA_INST_1[322].FA_  ( .A(A[2370]), .B(n1726), .CI(
        C[2370]), .CO(C[2371]) );
  FA_5818 \FA_INST_0[4].FA_INST_1[323].FA_  ( .A(A[2371]), .B(n1725), .CI(
        C[2371]), .CO(C[2372]) );
  FA_5817 \FA_INST_0[4].FA_INST_1[324].FA_  ( .A(A[2372]), .B(n1724), .CI(
        C[2372]), .CO(C[2373]) );
  FA_5816 \FA_INST_0[4].FA_INST_1[325].FA_  ( .A(A[2373]), .B(n1723), .CI(
        C[2373]), .CO(C[2374]) );
  FA_5815 \FA_INST_0[4].FA_INST_1[326].FA_  ( .A(A[2374]), .B(n1722), .CI(
        C[2374]), .CO(C[2375]) );
  FA_5814 \FA_INST_0[4].FA_INST_1[327].FA_  ( .A(A[2375]), .B(n1721), .CI(
        C[2375]), .CO(C[2376]) );
  FA_5813 \FA_INST_0[4].FA_INST_1[328].FA_  ( .A(A[2376]), .B(n1720), .CI(
        C[2376]), .CO(C[2377]) );
  FA_5812 \FA_INST_0[4].FA_INST_1[329].FA_  ( .A(A[2377]), .B(n1719), .CI(
        C[2377]), .CO(C[2378]) );
  FA_5811 \FA_INST_0[4].FA_INST_1[330].FA_  ( .A(A[2378]), .B(n1718), .CI(
        C[2378]), .CO(C[2379]) );
  FA_5810 \FA_INST_0[4].FA_INST_1[331].FA_  ( .A(A[2379]), .B(n1717), .CI(
        C[2379]), .CO(C[2380]) );
  FA_5809 \FA_INST_0[4].FA_INST_1[332].FA_  ( .A(A[2380]), .B(n1716), .CI(
        C[2380]), .CO(C[2381]) );
  FA_5808 \FA_INST_0[4].FA_INST_1[333].FA_  ( .A(A[2381]), .B(n1715), .CI(
        C[2381]), .CO(C[2382]) );
  FA_5807 \FA_INST_0[4].FA_INST_1[334].FA_  ( .A(A[2382]), .B(n1714), .CI(
        C[2382]), .CO(C[2383]) );
  FA_5806 \FA_INST_0[4].FA_INST_1[335].FA_  ( .A(A[2383]), .B(n1713), .CI(
        C[2383]), .CO(C[2384]) );
  FA_5805 \FA_INST_0[4].FA_INST_1[336].FA_  ( .A(A[2384]), .B(n1712), .CI(
        C[2384]), .CO(C[2385]) );
  FA_5804 \FA_INST_0[4].FA_INST_1[337].FA_  ( .A(A[2385]), .B(n1711), .CI(
        C[2385]), .CO(C[2386]) );
  FA_5803 \FA_INST_0[4].FA_INST_1[338].FA_  ( .A(A[2386]), .B(n1710), .CI(
        C[2386]), .CO(C[2387]) );
  FA_5802 \FA_INST_0[4].FA_INST_1[339].FA_  ( .A(A[2387]), .B(n1709), .CI(
        C[2387]), .CO(C[2388]) );
  FA_5801 \FA_INST_0[4].FA_INST_1[340].FA_  ( .A(A[2388]), .B(n1708), .CI(
        C[2388]), .CO(C[2389]) );
  FA_5800 \FA_INST_0[4].FA_INST_1[341].FA_  ( .A(A[2389]), .B(n1707), .CI(
        C[2389]), .CO(C[2390]) );
  FA_5799 \FA_INST_0[4].FA_INST_1[342].FA_  ( .A(A[2390]), .B(n1706), .CI(
        C[2390]), .CO(C[2391]) );
  FA_5798 \FA_INST_0[4].FA_INST_1[343].FA_  ( .A(A[2391]), .B(n1705), .CI(
        C[2391]), .CO(C[2392]) );
  FA_5797 \FA_INST_0[4].FA_INST_1[344].FA_  ( .A(A[2392]), .B(n1704), .CI(
        C[2392]), .CO(C[2393]) );
  FA_5796 \FA_INST_0[4].FA_INST_1[345].FA_  ( .A(A[2393]), .B(n1703), .CI(
        C[2393]), .CO(C[2394]) );
  FA_5795 \FA_INST_0[4].FA_INST_1[346].FA_  ( .A(A[2394]), .B(n1702), .CI(
        C[2394]), .CO(C[2395]) );
  FA_5794 \FA_INST_0[4].FA_INST_1[347].FA_  ( .A(A[2395]), .B(n1701), .CI(
        C[2395]), .CO(C[2396]) );
  FA_5793 \FA_INST_0[4].FA_INST_1[348].FA_  ( .A(A[2396]), .B(n1700), .CI(
        C[2396]), .CO(C[2397]) );
  FA_5792 \FA_INST_0[4].FA_INST_1[349].FA_  ( .A(A[2397]), .B(n1699), .CI(
        C[2397]), .CO(C[2398]) );
  FA_5791 \FA_INST_0[4].FA_INST_1[350].FA_  ( .A(A[2398]), .B(n1698), .CI(
        C[2398]), .CO(C[2399]) );
  FA_5790 \FA_INST_0[4].FA_INST_1[351].FA_  ( .A(A[2399]), .B(n1697), .CI(
        C[2399]), .CO(C[2400]) );
  FA_5789 \FA_INST_0[4].FA_INST_1[352].FA_  ( .A(A[2400]), .B(n1696), .CI(
        C[2400]), .CO(C[2401]) );
  FA_5788 \FA_INST_0[4].FA_INST_1[353].FA_  ( .A(A[2401]), .B(n1695), .CI(
        C[2401]), .CO(C[2402]) );
  FA_5787 \FA_INST_0[4].FA_INST_1[354].FA_  ( .A(A[2402]), .B(n1694), .CI(
        C[2402]), .CO(C[2403]) );
  FA_5786 \FA_INST_0[4].FA_INST_1[355].FA_  ( .A(A[2403]), .B(n1693), .CI(
        C[2403]), .CO(C[2404]) );
  FA_5785 \FA_INST_0[4].FA_INST_1[356].FA_  ( .A(A[2404]), .B(n1692), .CI(
        C[2404]), .CO(C[2405]) );
  FA_5784 \FA_INST_0[4].FA_INST_1[357].FA_  ( .A(A[2405]), .B(n1691), .CI(
        C[2405]), .CO(C[2406]) );
  FA_5783 \FA_INST_0[4].FA_INST_1[358].FA_  ( .A(A[2406]), .B(n1690), .CI(
        C[2406]), .CO(C[2407]) );
  FA_5782 \FA_INST_0[4].FA_INST_1[359].FA_  ( .A(A[2407]), .B(n1689), .CI(
        C[2407]), .CO(C[2408]) );
  FA_5781 \FA_INST_0[4].FA_INST_1[360].FA_  ( .A(A[2408]), .B(n1688), .CI(
        C[2408]), .CO(C[2409]) );
  FA_5780 \FA_INST_0[4].FA_INST_1[361].FA_  ( .A(A[2409]), .B(n1687), .CI(
        C[2409]), .CO(C[2410]) );
  FA_5779 \FA_INST_0[4].FA_INST_1[362].FA_  ( .A(A[2410]), .B(n1686), .CI(
        C[2410]), .CO(C[2411]) );
  FA_5778 \FA_INST_0[4].FA_INST_1[363].FA_  ( .A(A[2411]), .B(n1685), .CI(
        C[2411]), .CO(C[2412]) );
  FA_5777 \FA_INST_0[4].FA_INST_1[364].FA_  ( .A(A[2412]), .B(n1684), .CI(
        C[2412]), .CO(C[2413]) );
  FA_5776 \FA_INST_0[4].FA_INST_1[365].FA_  ( .A(A[2413]), .B(n1683), .CI(
        C[2413]), .CO(C[2414]) );
  FA_5775 \FA_INST_0[4].FA_INST_1[366].FA_  ( .A(A[2414]), .B(n1682), .CI(
        C[2414]), .CO(C[2415]) );
  FA_5774 \FA_INST_0[4].FA_INST_1[367].FA_  ( .A(A[2415]), .B(n1681), .CI(
        C[2415]), .CO(C[2416]) );
  FA_5773 \FA_INST_0[4].FA_INST_1[368].FA_  ( .A(A[2416]), .B(n1680), .CI(
        C[2416]), .CO(C[2417]) );
  FA_5772 \FA_INST_0[4].FA_INST_1[369].FA_  ( .A(A[2417]), .B(n1679), .CI(
        C[2417]), .CO(C[2418]) );
  FA_5771 \FA_INST_0[4].FA_INST_1[370].FA_  ( .A(A[2418]), .B(n1678), .CI(
        C[2418]), .CO(C[2419]) );
  FA_5770 \FA_INST_0[4].FA_INST_1[371].FA_  ( .A(A[2419]), .B(n1677), .CI(
        C[2419]), .CO(C[2420]) );
  FA_5769 \FA_INST_0[4].FA_INST_1[372].FA_  ( .A(A[2420]), .B(n1676), .CI(
        C[2420]), .CO(C[2421]) );
  FA_5768 \FA_INST_0[4].FA_INST_1[373].FA_  ( .A(A[2421]), .B(n1675), .CI(
        C[2421]), .CO(C[2422]) );
  FA_5767 \FA_INST_0[4].FA_INST_1[374].FA_  ( .A(A[2422]), .B(n1674), .CI(
        C[2422]), .CO(C[2423]) );
  FA_5766 \FA_INST_0[4].FA_INST_1[375].FA_  ( .A(A[2423]), .B(n1673), .CI(
        C[2423]), .CO(C[2424]) );
  FA_5765 \FA_INST_0[4].FA_INST_1[376].FA_  ( .A(A[2424]), .B(n1672), .CI(
        C[2424]), .CO(C[2425]) );
  FA_5764 \FA_INST_0[4].FA_INST_1[377].FA_  ( .A(A[2425]), .B(n1671), .CI(
        C[2425]), .CO(C[2426]) );
  FA_5763 \FA_INST_0[4].FA_INST_1[378].FA_  ( .A(A[2426]), .B(n1670), .CI(
        C[2426]), .CO(C[2427]) );
  FA_5762 \FA_INST_0[4].FA_INST_1[379].FA_  ( .A(A[2427]), .B(n1669), .CI(
        C[2427]), .CO(C[2428]) );
  FA_5761 \FA_INST_0[4].FA_INST_1[380].FA_  ( .A(A[2428]), .B(n1668), .CI(
        C[2428]), .CO(C[2429]) );
  FA_5760 \FA_INST_0[4].FA_INST_1[381].FA_  ( .A(A[2429]), .B(n1667), .CI(
        C[2429]), .CO(C[2430]) );
  FA_5759 \FA_INST_0[4].FA_INST_1[382].FA_  ( .A(A[2430]), .B(n1666), .CI(
        C[2430]), .CO(C[2431]) );
  FA_5758 \FA_INST_0[4].FA_INST_1[383].FA_  ( .A(A[2431]), .B(n1665), .CI(
        C[2431]), .CO(C[2432]) );
  FA_5757 \FA_INST_0[4].FA_INST_1[384].FA_  ( .A(A[2432]), .B(n1664), .CI(
        C[2432]), .CO(C[2433]) );
  FA_5756 \FA_INST_0[4].FA_INST_1[385].FA_  ( .A(A[2433]), .B(n1663), .CI(
        C[2433]), .CO(C[2434]) );
  FA_5755 \FA_INST_0[4].FA_INST_1[386].FA_  ( .A(A[2434]), .B(n1662), .CI(
        C[2434]), .CO(C[2435]) );
  FA_5754 \FA_INST_0[4].FA_INST_1[387].FA_  ( .A(A[2435]), .B(n1661), .CI(
        C[2435]), .CO(C[2436]) );
  FA_5753 \FA_INST_0[4].FA_INST_1[388].FA_  ( .A(A[2436]), .B(n1660), .CI(
        C[2436]), .CO(C[2437]) );
  FA_5752 \FA_INST_0[4].FA_INST_1[389].FA_  ( .A(A[2437]), .B(n1659), .CI(
        C[2437]), .CO(C[2438]) );
  FA_5751 \FA_INST_0[4].FA_INST_1[390].FA_  ( .A(A[2438]), .B(n1658), .CI(
        C[2438]), .CO(C[2439]) );
  FA_5750 \FA_INST_0[4].FA_INST_1[391].FA_  ( .A(A[2439]), .B(n1657), .CI(
        C[2439]), .CO(C[2440]) );
  FA_5749 \FA_INST_0[4].FA_INST_1[392].FA_  ( .A(A[2440]), .B(n1656), .CI(
        C[2440]), .CO(C[2441]) );
  FA_5748 \FA_INST_0[4].FA_INST_1[393].FA_  ( .A(A[2441]), .B(n1655), .CI(
        C[2441]), .CO(C[2442]) );
  FA_5747 \FA_INST_0[4].FA_INST_1[394].FA_  ( .A(A[2442]), .B(n1654), .CI(
        C[2442]), .CO(C[2443]) );
  FA_5746 \FA_INST_0[4].FA_INST_1[395].FA_  ( .A(A[2443]), .B(n1653), .CI(
        C[2443]), .CO(C[2444]) );
  FA_5745 \FA_INST_0[4].FA_INST_1[396].FA_  ( .A(A[2444]), .B(n1652), .CI(
        C[2444]), .CO(C[2445]) );
  FA_5744 \FA_INST_0[4].FA_INST_1[397].FA_  ( .A(A[2445]), .B(n1651), .CI(
        C[2445]), .CO(C[2446]) );
  FA_5743 \FA_INST_0[4].FA_INST_1[398].FA_  ( .A(A[2446]), .B(n1650), .CI(
        C[2446]), .CO(C[2447]) );
  FA_5742 \FA_INST_0[4].FA_INST_1[399].FA_  ( .A(A[2447]), .B(n1649), .CI(
        C[2447]), .CO(C[2448]) );
  FA_5741 \FA_INST_0[4].FA_INST_1[400].FA_  ( .A(A[2448]), .B(n1648), .CI(
        C[2448]), .CO(C[2449]) );
  FA_5740 \FA_INST_0[4].FA_INST_1[401].FA_  ( .A(A[2449]), .B(n1647), .CI(
        C[2449]), .CO(C[2450]) );
  FA_5739 \FA_INST_0[4].FA_INST_1[402].FA_  ( .A(A[2450]), .B(n1646), .CI(
        C[2450]), .CO(C[2451]) );
  FA_5738 \FA_INST_0[4].FA_INST_1[403].FA_  ( .A(A[2451]), .B(n1645), .CI(
        C[2451]), .CO(C[2452]) );
  FA_5737 \FA_INST_0[4].FA_INST_1[404].FA_  ( .A(A[2452]), .B(n1644), .CI(
        C[2452]), .CO(C[2453]) );
  FA_5736 \FA_INST_0[4].FA_INST_1[405].FA_  ( .A(A[2453]), .B(n1643), .CI(
        C[2453]), .CO(C[2454]) );
  FA_5735 \FA_INST_0[4].FA_INST_1[406].FA_  ( .A(A[2454]), .B(n1642), .CI(
        C[2454]), .CO(C[2455]) );
  FA_5734 \FA_INST_0[4].FA_INST_1[407].FA_  ( .A(A[2455]), .B(n1641), .CI(
        C[2455]), .CO(C[2456]) );
  FA_5733 \FA_INST_0[4].FA_INST_1[408].FA_  ( .A(A[2456]), .B(n1640), .CI(
        C[2456]), .CO(C[2457]) );
  FA_5732 \FA_INST_0[4].FA_INST_1[409].FA_  ( .A(A[2457]), .B(n1639), .CI(
        C[2457]), .CO(C[2458]) );
  FA_5731 \FA_INST_0[4].FA_INST_1[410].FA_  ( .A(A[2458]), .B(n1638), .CI(
        C[2458]), .CO(C[2459]) );
  FA_5730 \FA_INST_0[4].FA_INST_1[411].FA_  ( .A(A[2459]), .B(n1637), .CI(
        C[2459]), .CO(C[2460]) );
  FA_5729 \FA_INST_0[4].FA_INST_1[412].FA_  ( .A(A[2460]), .B(n1636), .CI(
        C[2460]), .CO(C[2461]) );
  FA_5728 \FA_INST_0[4].FA_INST_1[413].FA_  ( .A(A[2461]), .B(n1635), .CI(
        C[2461]), .CO(C[2462]) );
  FA_5727 \FA_INST_0[4].FA_INST_1[414].FA_  ( .A(A[2462]), .B(n1634), .CI(
        C[2462]), .CO(C[2463]) );
  FA_5726 \FA_INST_0[4].FA_INST_1[415].FA_  ( .A(A[2463]), .B(n1633), .CI(
        C[2463]), .CO(C[2464]) );
  FA_5725 \FA_INST_0[4].FA_INST_1[416].FA_  ( .A(A[2464]), .B(n1632), .CI(
        C[2464]), .CO(C[2465]) );
  FA_5724 \FA_INST_0[4].FA_INST_1[417].FA_  ( .A(A[2465]), .B(n1631), .CI(
        C[2465]), .CO(C[2466]) );
  FA_5723 \FA_INST_0[4].FA_INST_1[418].FA_  ( .A(A[2466]), .B(n1630), .CI(
        C[2466]), .CO(C[2467]) );
  FA_5722 \FA_INST_0[4].FA_INST_1[419].FA_  ( .A(A[2467]), .B(n1629), .CI(
        C[2467]), .CO(C[2468]) );
  FA_5721 \FA_INST_0[4].FA_INST_1[420].FA_  ( .A(A[2468]), .B(n1628), .CI(
        C[2468]), .CO(C[2469]) );
  FA_5720 \FA_INST_0[4].FA_INST_1[421].FA_  ( .A(A[2469]), .B(n1627), .CI(
        C[2469]), .CO(C[2470]) );
  FA_5719 \FA_INST_0[4].FA_INST_1[422].FA_  ( .A(A[2470]), .B(n1626), .CI(
        C[2470]), .CO(C[2471]) );
  FA_5718 \FA_INST_0[4].FA_INST_1[423].FA_  ( .A(A[2471]), .B(n1625), .CI(
        C[2471]), .CO(C[2472]) );
  FA_5717 \FA_INST_0[4].FA_INST_1[424].FA_  ( .A(A[2472]), .B(n1624), .CI(
        C[2472]), .CO(C[2473]) );
  FA_5716 \FA_INST_0[4].FA_INST_1[425].FA_  ( .A(A[2473]), .B(n1623), .CI(
        C[2473]), .CO(C[2474]) );
  FA_5715 \FA_INST_0[4].FA_INST_1[426].FA_  ( .A(A[2474]), .B(n1622), .CI(
        C[2474]), .CO(C[2475]) );
  FA_5714 \FA_INST_0[4].FA_INST_1[427].FA_  ( .A(A[2475]), .B(n1621), .CI(
        C[2475]), .CO(C[2476]) );
  FA_5713 \FA_INST_0[4].FA_INST_1[428].FA_  ( .A(A[2476]), .B(n1620), .CI(
        C[2476]), .CO(C[2477]) );
  FA_5712 \FA_INST_0[4].FA_INST_1[429].FA_  ( .A(A[2477]), .B(n1619), .CI(
        C[2477]), .CO(C[2478]) );
  FA_5711 \FA_INST_0[4].FA_INST_1[430].FA_  ( .A(A[2478]), .B(n1618), .CI(
        C[2478]), .CO(C[2479]) );
  FA_5710 \FA_INST_0[4].FA_INST_1[431].FA_  ( .A(A[2479]), .B(n1617), .CI(
        C[2479]), .CO(C[2480]) );
  FA_5709 \FA_INST_0[4].FA_INST_1[432].FA_  ( .A(A[2480]), .B(n1616), .CI(
        C[2480]), .CO(C[2481]) );
  FA_5708 \FA_INST_0[4].FA_INST_1[433].FA_  ( .A(A[2481]), .B(n1615), .CI(
        C[2481]), .CO(C[2482]) );
  FA_5707 \FA_INST_0[4].FA_INST_1[434].FA_  ( .A(A[2482]), .B(n1614), .CI(
        C[2482]), .CO(C[2483]) );
  FA_5706 \FA_INST_0[4].FA_INST_1[435].FA_  ( .A(A[2483]), .B(n1613), .CI(
        C[2483]), .CO(C[2484]) );
  FA_5705 \FA_INST_0[4].FA_INST_1[436].FA_  ( .A(A[2484]), .B(n1612), .CI(
        C[2484]), .CO(C[2485]) );
  FA_5704 \FA_INST_0[4].FA_INST_1[437].FA_  ( .A(A[2485]), .B(n1611), .CI(
        C[2485]), .CO(C[2486]) );
  FA_5703 \FA_INST_0[4].FA_INST_1[438].FA_  ( .A(A[2486]), .B(n1610), .CI(
        C[2486]), .CO(C[2487]) );
  FA_5702 \FA_INST_0[4].FA_INST_1[439].FA_  ( .A(A[2487]), .B(n1609), .CI(
        C[2487]), .CO(C[2488]) );
  FA_5701 \FA_INST_0[4].FA_INST_1[440].FA_  ( .A(A[2488]), .B(n1608), .CI(
        C[2488]), .CO(C[2489]) );
  FA_5700 \FA_INST_0[4].FA_INST_1[441].FA_  ( .A(A[2489]), .B(n1607), .CI(
        C[2489]), .CO(C[2490]) );
  FA_5699 \FA_INST_0[4].FA_INST_1[442].FA_  ( .A(A[2490]), .B(n1606), .CI(
        C[2490]), .CO(C[2491]) );
  FA_5698 \FA_INST_0[4].FA_INST_1[443].FA_  ( .A(A[2491]), .B(n1605), .CI(
        C[2491]), .CO(C[2492]) );
  FA_5697 \FA_INST_0[4].FA_INST_1[444].FA_  ( .A(A[2492]), .B(n1604), .CI(
        C[2492]), .CO(C[2493]) );
  FA_5696 \FA_INST_0[4].FA_INST_1[445].FA_  ( .A(A[2493]), .B(n1603), .CI(
        C[2493]), .CO(C[2494]) );
  FA_5695 \FA_INST_0[4].FA_INST_1[446].FA_  ( .A(A[2494]), .B(n1602), .CI(
        C[2494]), .CO(C[2495]) );
  FA_5694 \FA_INST_0[4].FA_INST_1[447].FA_  ( .A(A[2495]), .B(n1601), .CI(
        C[2495]), .CO(C[2496]) );
  FA_5693 \FA_INST_0[4].FA_INST_1[448].FA_  ( .A(A[2496]), .B(n1600), .CI(
        C[2496]), .CO(C[2497]) );
  FA_5692 \FA_INST_0[4].FA_INST_1[449].FA_  ( .A(A[2497]), .B(n1599), .CI(
        C[2497]), .CO(C[2498]) );
  FA_5691 \FA_INST_0[4].FA_INST_1[450].FA_  ( .A(A[2498]), .B(n1598), .CI(
        C[2498]), .CO(C[2499]) );
  FA_5690 \FA_INST_0[4].FA_INST_1[451].FA_  ( .A(A[2499]), .B(n1597), .CI(
        C[2499]), .CO(C[2500]) );
  FA_5689 \FA_INST_0[4].FA_INST_1[452].FA_  ( .A(A[2500]), .B(n1596), .CI(
        C[2500]), .CO(C[2501]) );
  FA_5688 \FA_INST_0[4].FA_INST_1[453].FA_  ( .A(A[2501]), .B(n1595), .CI(
        C[2501]), .CO(C[2502]) );
  FA_5687 \FA_INST_0[4].FA_INST_1[454].FA_  ( .A(A[2502]), .B(n1594), .CI(
        C[2502]), .CO(C[2503]) );
  FA_5686 \FA_INST_0[4].FA_INST_1[455].FA_  ( .A(A[2503]), .B(n1593), .CI(
        C[2503]), .CO(C[2504]) );
  FA_5685 \FA_INST_0[4].FA_INST_1[456].FA_  ( .A(A[2504]), .B(n1592), .CI(
        C[2504]), .CO(C[2505]) );
  FA_5684 \FA_INST_0[4].FA_INST_1[457].FA_  ( .A(A[2505]), .B(n1591), .CI(
        C[2505]), .CO(C[2506]) );
  FA_5683 \FA_INST_0[4].FA_INST_1[458].FA_  ( .A(A[2506]), .B(n1590), .CI(
        C[2506]), .CO(C[2507]) );
  FA_5682 \FA_INST_0[4].FA_INST_1[459].FA_  ( .A(A[2507]), .B(n1589), .CI(
        C[2507]), .CO(C[2508]) );
  FA_5681 \FA_INST_0[4].FA_INST_1[460].FA_  ( .A(A[2508]), .B(n1588), .CI(
        C[2508]), .CO(C[2509]) );
  FA_5680 \FA_INST_0[4].FA_INST_1[461].FA_  ( .A(A[2509]), .B(n1587), .CI(
        C[2509]), .CO(C[2510]) );
  FA_5679 \FA_INST_0[4].FA_INST_1[462].FA_  ( .A(A[2510]), .B(n1586), .CI(
        C[2510]), .CO(C[2511]) );
  FA_5678 \FA_INST_0[4].FA_INST_1[463].FA_  ( .A(A[2511]), .B(n1585), .CI(
        C[2511]), .CO(C[2512]) );
  FA_5677 \FA_INST_0[4].FA_INST_1[464].FA_  ( .A(A[2512]), .B(n1584), .CI(
        C[2512]), .CO(C[2513]) );
  FA_5676 \FA_INST_0[4].FA_INST_1[465].FA_  ( .A(A[2513]), .B(n1583), .CI(
        C[2513]), .CO(C[2514]) );
  FA_5675 \FA_INST_0[4].FA_INST_1[466].FA_  ( .A(A[2514]), .B(n1582), .CI(
        C[2514]), .CO(C[2515]) );
  FA_5674 \FA_INST_0[4].FA_INST_1[467].FA_  ( .A(A[2515]), .B(n1581), .CI(
        C[2515]), .CO(C[2516]) );
  FA_5673 \FA_INST_0[4].FA_INST_1[468].FA_  ( .A(A[2516]), .B(n1580), .CI(
        C[2516]), .CO(C[2517]) );
  FA_5672 \FA_INST_0[4].FA_INST_1[469].FA_  ( .A(A[2517]), .B(n1579), .CI(
        C[2517]), .CO(C[2518]) );
  FA_5671 \FA_INST_0[4].FA_INST_1[470].FA_  ( .A(A[2518]), .B(n1578), .CI(
        C[2518]), .CO(C[2519]) );
  FA_5670 \FA_INST_0[4].FA_INST_1[471].FA_  ( .A(A[2519]), .B(n1577), .CI(
        C[2519]), .CO(C[2520]) );
  FA_5669 \FA_INST_0[4].FA_INST_1[472].FA_  ( .A(A[2520]), .B(n1576), .CI(
        C[2520]), .CO(C[2521]) );
  FA_5668 \FA_INST_0[4].FA_INST_1[473].FA_  ( .A(A[2521]), .B(n1575), .CI(
        C[2521]), .CO(C[2522]) );
  FA_5667 \FA_INST_0[4].FA_INST_1[474].FA_  ( .A(A[2522]), .B(n1574), .CI(
        C[2522]), .CO(C[2523]) );
  FA_5666 \FA_INST_0[4].FA_INST_1[475].FA_  ( .A(A[2523]), .B(n1573), .CI(
        C[2523]), .CO(C[2524]) );
  FA_5665 \FA_INST_0[4].FA_INST_1[476].FA_  ( .A(A[2524]), .B(n1572), .CI(
        C[2524]), .CO(C[2525]) );
  FA_5664 \FA_INST_0[4].FA_INST_1[477].FA_  ( .A(A[2525]), .B(n1571), .CI(
        C[2525]), .CO(C[2526]) );
  FA_5663 \FA_INST_0[4].FA_INST_1[478].FA_  ( .A(A[2526]), .B(n1570), .CI(
        C[2526]), .CO(C[2527]) );
  FA_5662 \FA_INST_0[4].FA_INST_1[479].FA_  ( .A(A[2527]), .B(n1569), .CI(
        C[2527]), .CO(C[2528]) );
  FA_5661 \FA_INST_0[4].FA_INST_1[480].FA_  ( .A(A[2528]), .B(n1568), .CI(
        C[2528]), .CO(C[2529]) );
  FA_5660 \FA_INST_0[4].FA_INST_1[481].FA_  ( .A(A[2529]), .B(n1567), .CI(
        C[2529]), .CO(C[2530]) );
  FA_5659 \FA_INST_0[4].FA_INST_1[482].FA_  ( .A(A[2530]), .B(n1566), .CI(
        C[2530]), .CO(C[2531]) );
  FA_5658 \FA_INST_0[4].FA_INST_1[483].FA_  ( .A(A[2531]), .B(n1565), .CI(
        C[2531]), .CO(C[2532]) );
  FA_5657 \FA_INST_0[4].FA_INST_1[484].FA_  ( .A(A[2532]), .B(n1564), .CI(
        C[2532]), .CO(C[2533]) );
  FA_5656 \FA_INST_0[4].FA_INST_1[485].FA_  ( .A(A[2533]), .B(n1563), .CI(
        C[2533]), .CO(C[2534]) );
  FA_5655 \FA_INST_0[4].FA_INST_1[486].FA_  ( .A(A[2534]), .B(n1562), .CI(
        C[2534]), .CO(C[2535]) );
  FA_5654 \FA_INST_0[4].FA_INST_1[487].FA_  ( .A(A[2535]), .B(n1561), .CI(
        C[2535]), .CO(C[2536]) );
  FA_5653 \FA_INST_0[4].FA_INST_1[488].FA_  ( .A(A[2536]), .B(n1560), .CI(
        C[2536]), .CO(C[2537]) );
  FA_5652 \FA_INST_0[4].FA_INST_1[489].FA_  ( .A(A[2537]), .B(n1559), .CI(
        C[2537]), .CO(C[2538]) );
  FA_5651 \FA_INST_0[4].FA_INST_1[490].FA_  ( .A(A[2538]), .B(n1558), .CI(
        C[2538]), .CO(C[2539]) );
  FA_5650 \FA_INST_0[4].FA_INST_1[491].FA_  ( .A(A[2539]), .B(n1557), .CI(
        C[2539]), .CO(C[2540]) );
  FA_5649 \FA_INST_0[4].FA_INST_1[492].FA_  ( .A(A[2540]), .B(n1556), .CI(
        C[2540]), .CO(C[2541]) );
  FA_5648 \FA_INST_0[4].FA_INST_1[493].FA_  ( .A(A[2541]), .B(n1555), .CI(
        C[2541]), .CO(C[2542]) );
  FA_5647 \FA_INST_0[4].FA_INST_1[494].FA_  ( .A(A[2542]), .B(n1554), .CI(
        C[2542]), .CO(C[2543]) );
  FA_5646 \FA_INST_0[4].FA_INST_1[495].FA_  ( .A(A[2543]), .B(n1553), .CI(
        C[2543]), .CO(C[2544]) );
  FA_5645 \FA_INST_0[4].FA_INST_1[496].FA_  ( .A(A[2544]), .B(n1552), .CI(
        C[2544]), .CO(C[2545]) );
  FA_5644 \FA_INST_0[4].FA_INST_1[497].FA_  ( .A(A[2545]), .B(n1551), .CI(
        C[2545]), .CO(C[2546]) );
  FA_5643 \FA_INST_0[4].FA_INST_1[498].FA_  ( .A(A[2546]), .B(n1550), .CI(
        C[2546]), .CO(C[2547]) );
  FA_5642 \FA_INST_0[4].FA_INST_1[499].FA_  ( .A(A[2547]), .B(n1549), .CI(
        C[2547]), .CO(C[2548]) );
  FA_5641 \FA_INST_0[4].FA_INST_1[500].FA_  ( .A(A[2548]), .B(n1548), .CI(
        C[2548]), .CO(C[2549]) );
  FA_5640 \FA_INST_0[4].FA_INST_1[501].FA_  ( .A(A[2549]), .B(n1547), .CI(
        C[2549]), .CO(C[2550]) );
  FA_5639 \FA_INST_0[4].FA_INST_1[502].FA_  ( .A(A[2550]), .B(n1546), .CI(
        C[2550]), .CO(C[2551]) );
  FA_5638 \FA_INST_0[4].FA_INST_1[503].FA_  ( .A(A[2551]), .B(n1545), .CI(
        C[2551]), .CO(C[2552]) );
  FA_5637 \FA_INST_0[4].FA_INST_1[504].FA_  ( .A(A[2552]), .B(n1544), .CI(
        C[2552]), .CO(C[2553]) );
  FA_5636 \FA_INST_0[4].FA_INST_1[505].FA_  ( .A(A[2553]), .B(n1543), .CI(
        C[2553]), .CO(C[2554]) );
  FA_5635 \FA_INST_0[4].FA_INST_1[506].FA_  ( .A(A[2554]), .B(n1542), .CI(
        C[2554]), .CO(C[2555]) );
  FA_5634 \FA_INST_0[4].FA_INST_1[507].FA_  ( .A(A[2555]), .B(n1541), .CI(
        C[2555]), .CO(C[2556]) );
  FA_5633 \FA_INST_0[4].FA_INST_1[508].FA_  ( .A(A[2556]), .B(n1540), .CI(
        C[2556]), .CO(C[2557]) );
  FA_5632 \FA_INST_0[4].FA_INST_1[509].FA_  ( .A(A[2557]), .B(n1539), .CI(
        C[2557]), .CO(C[2558]) );
  FA_5631 \FA_INST_0[4].FA_INST_1[510].FA_  ( .A(A[2558]), .B(n1538), .CI(
        C[2558]), .CO(C[2559]) );
  FA_5630 \FA_INST_0[4].FA_INST_1[511].FA_  ( .A(A[2559]), .B(n1537), .CI(
        C[2559]), .CO(C[2560]) );
  FA_5629 \FA_INST_0[5].FA_INST_1[0].FA_  ( .A(A[2560]), .B(n1536), .CI(
        C[2560]), .CO(C[2561]) );
  FA_5628 \FA_INST_0[5].FA_INST_1[1].FA_  ( .A(A[2561]), .B(n1535), .CI(
        C[2561]), .CO(C[2562]) );
  FA_5627 \FA_INST_0[5].FA_INST_1[2].FA_  ( .A(A[2562]), .B(n1534), .CI(
        C[2562]), .CO(C[2563]) );
  FA_5626 \FA_INST_0[5].FA_INST_1[3].FA_  ( .A(A[2563]), .B(n1533), .CI(
        C[2563]), .CO(C[2564]) );
  FA_5625 \FA_INST_0[5].FA_INST_1[4].FA_  ( .A(A[2564]), .B(n1532), .CI(
        C[2564]), .CO(C[2565]) );
  FA_5624 \FA_INST_0[5].FA_INST_1[5].FA_  ( .A(A[2565]), .B(n1531), .CI(
        C[2565]), .CO(C[2566]) );
  FA_5623 \FA_INST_0[5].FA_INST_1[6].FA_  ( .A(A[2566]), .B(n1530), .CI(
        C[2566]), .CO(C[2567]) );
  FA_5622 \FA_INST_0[5].FA_INST_1[7].FA_  ( .A(A[2567]), .B(n1529), .CI(
        C[2567]), .CO(C[2568]) );
  FA_5621 \FA_INST_0[5].FA_INST_1[8].FA_  ( .A(A[2568]), .B(n1528), .CI(
        C[2568]), .CO(C[2569]) );
  FA_5620 \FA_INST_0[5].FA_INST_1[9].FA_  ( .A(A[2569]), .B(n1527), .CI(
        C[2569]), .CO(C[2570]) );
  FA_5619 \FA_INST_0[5].FA_INST_1[10].FA_  ( .A(A[2570]), .B(n1526), .CI(
        C[2570]), .CO(C[2571]) );
  FA_5618 \FA_INST_0[5].FA_INST_1[11].FA_  ( .A(A[2571]), .B(n1525), .CI(
        C[2571]), .CO(C[2572]) );
  FA_5617 \FA_INST_0[5].FA_INST_1[12].FA_  ( .A(A[2572]), .B(n1524), .CI(
        C[2572]), .CO(C[2573]) );
  FA_5616 \FA_INST_0[5].FA_INST_1[13].FA_  ( .A(A[2573]), .B(n1523), .CI(
        C[2573]), .CO(C[2574]) );
  FA_5615 \FA_INST_0[5].FA_INST_1[14].FA_  ( .A(A[2574]), .B(n1522), .CI(
        C[2574]), .CO(C[2575]) );
  FA_5614 \FA_INST_0[5].FA_INST_1[15].FA_  ( .A(A[2575]), .B(n1521), .CI(
        C[2575]), .CO(C[2576]) );
  FA_5613 \FA_INST_0[5].FA_INST_1[16].FA_  ( .A(A[2576]), .B(n1520), .CI(
        C[2576]), .CO(C[2577]) );
  FA_5612 \FA_INST_0[5].FA_INST_1[17].FA_  ( .A(A[2577]), .B(n1519), .CI(
        C[2577]), .CO(C[2578]) );
  FA_5611 \FA_INST_0[5].FA_INST_1[18].FA_  ( .A(A[2578]), .B(n1518), .CI(
        C[2578]), .CO(C[2579]) );
  FA_5610 \FA_INST_0[5].FA_INST_1[19].FA_  ( .A(A[2579]), .B(n1517), .CI(
        C[2579]), .CO(C[2580]) );
  FA_5609 \FA_INST_0[5].FA_INST_1[20].FA_  ( .A(A[2580]), .B(n1516), .CI(
        C[2580]), .CO(C[2581]) );
  FA_5608 \FA_INST_0[5].FA_INST_1[21].FA_  ( .A(A[2581]), .B(n1515), .CI(
        C[2581]), .CO(C[2582]) );
  FA_5607 \FA_INST_0[5].FA_INST_1[22].FA_  ( .A(A[2582]), .B(n1514), .CI(
        C[2582]), .CO(C[2583]) );
  FA_5606 \FA_INST_0[5].FA_INST_1[23].FA_  ( .A(A[2583]), .B(n1513), .CI(
        C[2583]), .CO(C[2584]) );
  FA_5605 \FA_INST_0[5].FA_INST_1[24].FA_  ( .A(A[2584]), .B(n1512), .CI(
        C[2584]), .CO(C[2585]) );
  FA_5604 \FA_INST_0[5].FA_INST_1[25].FA_  ( .A(A[2585]), .B(n1511), .CI(
        C[2585]), .CO(C[2586]) );
  FA_5603 \FA_INST_0[5].FA_INST_1[26].FA_  ( .A(A[2586]), .B(n1510), .CI(
        C[2586]), .CO(C[2587]) );
  FA_5602 \FA_INST_0[5].FA_INST_1[27].FA_  ( .A(A[2587]), .B(n1509), .CI(
        C[2587]), .CO(C[2588]) );
  FA_5601 \FA_INST_0[5].FA_INST_1[28].FA_  ( .A(A[2588]), .B(n1508), .CI(
        C[2588]), .CO(C[2589]) );
  FA_5600 \FA_INST_0[5].FA_INST_1[29].FA_  ( .A(A[2589]), .B(n1507), .CI(
        C[2589]), .CO(C[2590]) );
  FA_5599 \FA_INST_0[5].FA_INST_1[30].FA_  ( .A(A[2590]), .B(n1506), .CI(
        C[2590]), .CO(C[2591]) );
  FA_5598 \FA_INST_0[5].FA_INST_1[31].FA_  ( .A(A[2591]), .B(n1505), .CI(
        C[2591]), .CO(C[2592]) );
  FA_5597 \FA_INST_0[5].FA_INST_1[32].FA_  ( .A(A[2592]), .B(n1504), .CI(
        C[2592]), .CO(C[2593]) );
  FA_5596 \FA_INST_0[5].FA_INST_1[33].FA_  ( .A(A[2593]), .B(n1503), .CI(
        C[2593]), .CO(C[2594]) );
  FA_5595 \FA_INST_0[5].FA_INST_1[34].FA_  ( .A(A[2594]), .B(n1502), .CI(
        C[2594]), .CO(C[2595]) );
  FA_5594 \FA_INST_0[5].FA_INST_1[35].FA_  ( .A(A[2595]), .B(n1501), .CI(
        C[2595]), .CO(C[2596]) );
  FA_5593 \FA_INST_0[5].FA_INST_1[36].FA_  ( .A(A[2596]), .B(n1500), .CI(
        C[2596]), .CO(C[2597]) );
  FA_5592 \FA_INST_0[5].FA_INST_1[37].FA_  ( .A(A[2597]), .B(n1499), .CI(
        C[2597]), .CO(C[2598]) );
  FA_5591 \FA_INST_0[5].FA_INST_1[38].FA_  ( .A(A[2598]), .B(n1498), .CI(
        C[2598]), .CO(C[2599]) );
  FA_5590 \FA_INST_0[5].FA_INST_1[39].FA_  ( .A(A[2599]), .B(n1497), .CI(
        C[2599]), .CO(C[2600]) );
  FA_5589 \FA_INST_0[5].FA_INST_1[40].FA_  ( .A(A[2600]), .B(n1496), .CI(
        C[2600]), .CO(C[2601]) );
  FA_5588 \FA_INST_0[5].FA_INST_1[41].FA_  ( .A(A[2601]), .B(n1495), .CI(
        C[2601]), .CO(C[2602]) );
  FA_5587 \FA_INST_0[5].FA_INST_1[42].FA_  ( .A(A[2602]), .B(n1494), .CI(
        C[2602]), .CO(C[2603]) );
  FA_5586 \FA_INST_0[5].FA_INST_1[43].FA_  ( .A(A[2603]), .B(n1493), .CI(
        C[2603]), .CO(C[2604]) );
  FA_5585 \FA_INST_0[5].FA_INST_1[44].FA_  ( .A(A[2604]), .B(n1492), .CI(
        C[2604]), .CO(C[2605]) );
  FA_5584 \FA_INST_0[5].FA_INST_1[45].FA_  ( .A(A[2605]), .B(n1491), .CI(
        C[2605]), .CO(C[2606]) );
  FA_5583 \FA_INST_0[5].FA_INST_1[46].FA_  ( .A(A[2606]), .B(n1490), .CI(
        C[2606]), .CO(C[2607]) );
  FA_5582 \FA_INST_0[5].FA_INST_1[47].FA_  ( .A(A[2607]), .B(n1489), .CI(
        C[2607]), .CO(C[2608]) );
  FA_5581 \FA_INST_0[5].FA_INST_1[48].FA_  ( .A(A[2608]), .B(n1488), .CI(
        C[2608]), .CO(C[2609]) );
  FA_5580 \FA_INST_0[5].FA_INST_1[49].FA_  ( .A(A[2609]), .B(n1487), .CI(
        C[2609]), .CO(C[2610]) );
  FA_5579 \FA_INST_0[5].FA_INST_1[50].FA_  ( .A(A[2610]), .B(n1486), .CI(
        C[2610]), .CO(C[2611]) );
  FA_5578 \FA_INST_0[5].FA_INST_1[51].FA_  ( .A(A[2611]), .B(n1485), .CI(
        C[2611]), .CO(C[2612]) );
  FA_5577 \FA_INST_0[5].FA_INST_1[52].FA_  ( .A(A[2612]), .B(n1484), .CI(
        C[2612]), .CO(C[2613]) );
  FA_5576 \FA_INST_0[5].FA_INST_1[53].FA_  ( .A(A[2613]), .B(n1483), .CI(
        C[2613]), .CO(C[2614]) );
  FA_5575 \FA_INST_0[5].FA_INST_1[54].FA_  ( .A(A[2614]), .B(n1482), .CI(
        C[2614]), .CO(C[2615]) );
  FA_5574 \FA_INST_0[5].FA_INST_1[55].FA_  ( .A(A[2615]), .B(n1481), .CI(
        C[2615]), .CO(C[2616]) );
  FA_5573 \FA_INST_0[5].FA_INST_1[56].FA_  ( .A(A[2616]), .B(n1480), .CI(
        C[2616]), .CO(C[2617]) );
  FA_5572 \FA_INST_0[5].FA_INST_1[57].FA_  ( .A(A[2617]), .B(n1479), .CI(
        C[2617]), .CO(C[2618]) );
  FA_5571 \FA_INST_0[5].FA_INST_1[58].FA_  ( .A(A[2618]), .B(n1478), .CI(
        C[2618]), .CO(C[2619]) );
  FA_5570 \FA_INST_0[5].FA_INST_1[59].FA_  ( .A(A[2619]), .B(n1477), .CI(
        C[2619]), .CO(C[2620]) );
  FA_5569 \FA_INST_0[5].FA_INST_1[60].FA_  ( .A(A[2620]), .B(n1476), .CI(
        C[2620]), .CO(C[2621]) );
  FA_5568 \FA_INST_0[5].FA_INST_1[61].FA_  ( .A(A[2621]), .B(n1475), .CI(
        C[2621]), .CO(C[2622]) );
  FA_5567 \FA_INST_0[5].FA_INST_1[62].FA_  ( .A(A[2622]), .B(n1474), .CI(
        C[2622]), .CO(C[2623]) );
  FA_5566 \FA_INST_0[5].FA_INST_1[63].FA_  ( .A(A[2623]), .B(n1473), .CI(
        C[2623]), .CO(C[2624]) );
  FA_5565 \FA_INST_0[5].FA_INST_1[64].FA_  ( .A(A[2624]), .B(n1472), .CI(
        C[2624]), .CO(C[2625]) );
  FA_5564 \FA_INST_0[5].FA_INST_1[65].FA_  ( .A(A[2625]), .B(n1471), .CI(
        C[2625]), .CO(C[2626]) );
  FA_5563 \FA_INST_0[5].FA_INST_1[66].FA_  ( .A(A[2626]), .B(n1470), .CI(
        C[2626]), .CO(C[2627]) );
  FA_5562 \FA_INST_0[5].FA_INST_1[67].FA_  ( .A(A[2627]), .B(n1469), .CI(
        C[2627]), .CO(C[2628]) );
  FA_5561 \FA_INST_0[5].FA_INST_1[68].FA_  ( .A(A[2628]), .B(n1468), .CI(
        C[2628]), .CO(C[2629]) );
  FA_5560 \FA_INST_0[5].FA_INST_1[69].FA_  ( .A(A[2629]), .B(n1467), .CI(
        C[2629]), .CO(C[2630]) );
  FA_5559 \FA_INST_0[5].FA_INST_1[70].FA_  ( .A(A[2630]), .B(n1466), .CI(
        C[2630]), .CO(C[2631]) );
  FA_5558 \FA_INST_0[5].FA_INST_1[71].FA_  ( .A(A[2631]), .B(n1465), .CI(
        C[2631]), .CO(C[2632]) );
  FA_5557 \FA_INST_0[5].FA_INST_1[72].FA_  ( .A(A[2632]), .B(n1464), .CI(
        C[2632]), .CO(C[2633]) );
  FA_5556 \FA_INST_0[5].FA_INST_1[73].FA_  ( .A(A[2633]), .B(n1463), .CI(
        C[2633]), .CO(C[2634]) );
  FA_5555 \FA_INST_0[5].FA_INST_1[74].FA_  ( .A(A[2634]), .B(n1462), .CI(
        C[2634]), .CO(C[2635]) );
  FA_5554 \FA_INST_0[5].FA_INST_1[75].FA_  ( .A(A[2635]), .B(n1461), .CI(
        C[2635]), .CO(C[2636]) );
  FA_5553 \FA_INST_0[5].FA_INST_1[76].FA_  ( .A(A[2636]), .B(n1460), .CI(
        C[2636]), .CO(C[2637]) );
  FA_5552 \FA_INST_0[5].FA_INST_1[77].FA_  ( .A(A[2637]), .B(n1459), .CI(
        C[2637]), .CO(C[2638]) );
  FA_5551 \FA_INST_0[5].FA_INST_1[78].FA_  ( .A(A[2638]), .B(n1458), .CI(
        C[2638]), .CO(C[2639]) );
  FA_5550 \FA_INST_0[5].FA_INST_1[79].FA_  ( .A(A[2639]), .B(n1457), .CI(
        C[2639]), .CO(C[2640]) );
  FA_5549 \FA_INST_0[5].FA_INST_1[80].FA_  ( .A(A[2640]), .B(n1456), .CI(
        C[2640]), .CO(C[2641]) );
  FA_5548 \FA_INST_0[5].FA_INST_1[81].FA_  ( .A(A[2641]), .B(n1455), .CI(
        C[2641]), .CO(C[2642]) );
  FA_5547 \FA_INST_0[5].FA_INST_1[82].FA_  ( .A(A[2642]), .B(n1454), .CI(
        C[2642]), .CO(C[2643]) );
  FA_5546 \FA_INST_0[5].FA_INST_1[83].FA_  ( .A(A[2643]), .B(n1453), .CI(
        C[2643]), .CO(C[2644]) );
  FA_5545 \FA_INST_0[5].FA_INST_1[84].FA_  ( .A(A[2644]), .B(n1452), .CI(
        C[2644]), .CO(C[2645]) );
  FA_5544 \FA_INST_0[5].FA_INST_1[85].FA_  ( .A(A[2645]), .B(n1451), .CI(
        C[2645]), .CO(C[2646]) );
  FA_5543 \FA_INST_0[5].FA_INST_1[86].FA_  ( .A(A[2646]), .B(n1450), .CI(
        C[2646]), .CO(C[2647]) );
  FA_5542 \FA_INST_0[5].FA_INST_1[87].FA_  ( .A(A[2647]), .B(n1449), .CI(
        C[2647]), .CO(C[2648]) );
  FA_5541 \FA_INST_0[5].FA_INST_1[88].FA_  ( .A(A[2648]), .B(n1448), .CI(
        C[2648]), .CO(C[2649]) );
  FA_5540 \FA_INST_0[5].FA_INST_1[89].FA_  ( .A(A[2649]), .B(n1447), .CI(
        C[2649]), .CO(C[2650]) );
  FA_5539 \FA_INST_0[5].FA_INST_1[90].FA_  ( .A(A[2650]), .B(n1446), .CI(
        C[2650]), .CO(C[2651]) );
  FA_5538 \FA_INST_0[5].FA_INST_1[91].FA_  ( .A(A[2651]), .B(n1445), .CI(
        C[2651]), .CO(C[2652]) );
  FA_5537 \FA_INST_0[5].FA_INST_1[92].FA_  ( .A(A[2652]), .B(n1444), .CI(
        C[2652]), .CO(C[2653]) );
  FA_5536 \FA_INST_0[5].FA_INST_1[93].FA_  ( .A(A[2653]), .B(n1443), .CI(
        C[2653]), .CO(C[2654]) );
  FA_5535 \FA_INST_0[5].FA_INST_1[94].FA_  ( .A(A[2654]), .B(n1442), .CI(
        C[2654]), .CO(C[2655]) );
  FA_5534 \FA_INST_0[5].FA_INST_1[95].FA_  ( .A(A[2655]), .B(n1441), .CI(
        C[2655]), .CO(C[2656]) );
  FA_5533 \FA_INST_0[5].FA_INST_1[96].FA_  ( .A(A[2656]), .B(n1440), .CI(
        C[2656]), .CO(C[2657]) );
  FA_5532 \FA_INST_0[5].FA_INST_1[97].FA_  ( .A(A[2657]), .B(n1439), .CI(
        C[2657]), .CO(C[2658]) );
  FA_5531 \FA_INST_0[5].FA_INST_1[98].FA_  ( .A(A[2658]), .B(n1438), .CI(
        C[2658]), .CO(C[2659]) );
  FA_5530 \FA_INST_0[5].FA_INST_1[99].FA_  ( .A(A[2659]), .B(n1437), .CI(
        C[2659]), .CO(C[2660]) );
  FA_5529 \FA_INST_0[5].FA_INST_1[100].FA_  ( .A(A[2660]), .B(n1436), .CI(
        C[2660]), .CO(C[2661]) );
  FA_5528 \FA_INST_0[5].FA_INST_1[101].FA_  ( .A(A[2661]), .B(n1435), .CI(
        C[2661]), .CO(C[2662]) );
  FA_5527 \FA_INST_0[5].FA_INST_1[102].FA_  ( .A(A[2662]), .B(n1434), .CI(
        C[2662]), .CO(C[2663]) );
  FA_5526 \FA_INST_0[5].FA_INST_1[103].FA_  ( .A(A[2663]), .B(n1433), .CI(
        C[2663]), .CO(C[2664]) );
  FA_5525 \FA_INST_0[5].FA_INST_1[104].FA_  ( .A(A[2664]), .B(n1432), .CI(
        C[2664]), .CO(C[2665]) );
  FA_5524 \FA_INST_0[5].FA_INST_1[105].FA_  ( .A(A[2665]), .B(n1431), .CI(
        C[2665]), .CO(C[2666]) );
  FA_5523 \FA_INST_0[5].FA_INST_1[106].FA_  ( .A(A[2666]), .B(n1430), .CI(
        C[2666]), .CO(C[2667]) );
  FA_5522 \FA_INST_0[5].FA_INST_1[107].FA_  ( .A(A[2667]), .B(n1429), .CI(
        C[2667]), .CO(C[2668]) );
  FA_5521 \FA_INST_0[5].FA_INST_1[108].FA_  ( .A(A[2668]), .B(n1428), .CI(
        C[2668]), .CO(C[2669]) );
  FA_5520 \FA_INST_0[5].FA_INST_1[109].FA_  ( .A(A[2669]), .B(n1427), .CI(
        C[2669]), .CO(C[2670]) );
  FA_5519 \FA_INST_0[5].FA_INST_1[110].FA_  ( .A(A[2670]), .B(n1426), .CI(
        C[2670]), .CO(C[2671]) );
  FA_5518 \FA_INST_0[5].FA_INST_1[111].FA_  ( .A(A[2671]), .B(n1425), .CI(
        C[2671]), .CO(C[2672]) );
  FA_5517 \FA_INST_0[5].FA_INST_1[112].FA_  ( .A(A[2672]), .B(n1424), .CI(
        C[2672]), .CO(C[2673]) );
  FA_5516 \FA_INST_0[5].FA_INST_1[113].FA_  ( .A(A[2673]), .B(n1423), .CI(
        C[2673]), .CO(C[2674]) );
  FA_5515 \FA_INST_0[5].FA_INST_1[114].FA_  ( .A(A[2674]), .B(n1422), .CI(
        C[2674]), .CO(C[2675]) );
  FA_5514 \FA_INST_0[5].FA_INST_1[115].FA_  ( .A(A[2675]), .B(n1421), .CI(
        C[2675]), .CO(C[2676]) );
  FA_5513 \FA_INST_0[5].FA_INST_1[116].FA_  ( .A(A[2676]), .B(n1420), .CI(
        C[2676]), .CO(C[2677]) );
  FA_5512 \FA_INST_0[5].FA_INST_1[117].FA_  ( .A(A[2677]), .B(n1419), .CI(
        C[2677]), .CO(C[2678]) );
  FA_5511 \FA_INST_0[5].FA_INST_1[118].FA_  ( .A(A[2678]), .B(n1418), .CI(
        C[2678]), .CO(C[2679]) );
  FA_5510 \FA_INST_0[5].FA_INST_1[119].FA_  ( .A(A[2679]), .B(n1417), .CI(
        C[2679]), .CO(C[2680]) );
  FA_5509 \FA_INST_0[5].FA_INST_1[120].FA_  ( .A(A[2680]), .B(n1416), .CI(
        C[2680]), .CO(C[2681]) );
  FA_5508 \FA_INST_0[5].FA_INST_1[121].FA_  ( .A(A[2681]), .B(n1415), .CI(
        C[2681]), .CO(C[2682]) );
  FA_5507 \FA_INST_0[5].FA_INST_1[122].FA_  ( .A(A[2682]), .B(n1414), .CI(
        C[2682]), .CO(C[2683]) );
  FA_5506 \FA_INST_0[5].FA_INST_1[123].FA_  ( .A(A[2683]), .B(n1413), .CI(
        C[2683]), .CO(C[2684]) );
  FA_5505 \FA_INST_0[5].FA_INST_1[124].FA_  ( .A(A[2684]), .B(n1412), .CI(
        C[2684]), .CO(C[2685]) );
  FA_5504 \FA_INST_0[5].FA_INST_1[125].FA_  ( .A(A[2685]), .B(n1411), .CI(
        C[2685]), .CO(C[2686]) );
  FA_5503 \FA_INST_0[5].FA_INST_1[126].FA_  ( .A(A[2686]), .B(n1410), .CI(
        C[2686]), .CO(C[2687]) );
  FA_5502 \FA_INST_0[5].FA_INST_1[127].FA_  ( .A(A[2687]), .B(n1409), .CI(
        C[2687]), .CO(C[2688]) );
  FA_5501 \FA_INST_0[5].FA_INST_1[128].FA_  ( .A(A[2688]), .B(n1408), .CI(
        C[2688]), .CO(C[2689]) );
  FA_5500 \FA_INST_0[5].FA_INST_1[129].FA_  ( .A(A[2689]), .B(n1407), .CI(
        C[2689]), .CO(C[2690]) );
  FA_5499 \FA_INST_0[5].FA_INST_1[130].FA_  ( .A(A[2690]), .B(n1406), .CI(
        C[2690]), .CO(C[2691]) );
  FA_5498 \FA_INST_0[5].FA_INST_1[131].FA_  ( .A(A[2691]), .B(n1405), .CI(
        C[2691]), .CO(C[2692]) );
  FA_5497 \FA_INST_0[5].FA_INST_1[132].FA_  ( .A(A[2692]), .B(n1404), .CI(
        C[2692]), .CO(C[2693]) );
  FA_5496 \FA_INST_0[5].FA_INST_1[133].FA_  ( .A(A[2693]), .B(n1403), .CI(
        C[2693]), .CO(C[2694]) );
  FA_5495 \FA_INST_0[5].FA_INST_1[134].FA_  ( .A(A[2694]), .B(n1402), .CI(
        C[2694]), .CO(C[2695]) );
  FA_5494 \FA_INST_0[5].FA_INST_1[135].FA_  ( .A(A[2695]), .B(n1401), .CI(
        C[2695]), .CO(C[2696]) );
  FA_5493 \FA_INST_0[5].FA_INST_1[136].FA_  ( .A(A[2696]), .B(n1400), .CI(
        C[2696]), .CO(C[2697]) );
  FA_5492 \FA_INST_0[5].FA_INST_1[137].FA_  ( .A(A[2697]), .B(n1399), .CI(
        C[2697]), .CO(C[2698]) );
  FA_5491 \FA_INST_0[5].FA_INST_1[138].FA_  ( .A(A[2698]), .B(n1398), .CI(
        C[2698]), .CO(C[2699]) );
  FA_5490 \FA_INST_0[5].FA_INST_1[139].FA_  ( .A(A[2699]), .B(n1397), .CI(
        C[2699]), .CO(C[2700]) );
  FA_5489 \FA_INST_0[5].FA_INST_1[140].FA_  ( .A(A[2700]), .B(n1396), .CI(
        C[2700]), .CO(C[2701]) );
  FA_5488 \FA_INST_0[5].FA_INST_1[141].FA_  ( .A(A[2701]), .B(n1395), .CI(
        C[2701]), .CO(C[2702]) );
  FA_5487 \FA_INST_0[5].FA_INST_1[142].FA_  ( .A(A[2702]), .B(n1394), .CI(
        C[2702]), .CO(C[2703]) );
  FA_5486 \FA_INST_0[5].FA_INST_1[143].FA_  ( .A(A[2703]), .B(n1393), .CI(
        C[2703]), .CO(C[2704]) );
  FA_5485 \FA_INST_0[5].FA_INST_1[144].FA_  ( .A(A[2704]), .B(n1392), .CI(
        C[2704]), .CO(C[2705]) );
  FA_5484 \FA_INST_0[5].FA_INST_1[145].FA_  ( .A(A[2705]), .B(n1391), .CI(
        C[2705]), .CO(C[2706]) );
  FA_5483 \FA_INST_0[5].FA_INST_1[146].FA_  ( .A(A[2706]), .B(n1390), .CI(
        C[2706]), .CO(C[2707]) );
  FA_5482 \FA_INST_0[5].FA_INST_1[147].FA_  ( .A(A[2707]), .B(n1389), .CI(
        C[2707]), .CO(C[2708]) );
  FA_5481 \FA_INST_0[5].FA_INST_1[148].FA_  ( .A(A[2708]), .B(n1388), .CI(
        C[2708]), .CO(C[2709]) );
  FA_5480 \FA_INST_0[5].FA_INST_1[149].FA_  ( .A(A[2709]), .B(n1387), .CI(
        C[2709]), .CO(C[2710]) );
  FA_5479 \FA_INST_0[5].FA_INST_1[150].FA_  ( .A(A[2710]), .B(n1386), .CI(
        C[2710]), .CO(C[2711]) );
  FA_5478 \FA_INST_0[5].FA_INST_1[151].FA_  ( .A(A[2711]), .B(n1385), .CI(
        C[2711]), .CO(C[2712]) );
  FA_5477 \FA_INST_0[5].FA_INST_1[152].FA_  ( .A(A[2712]), .B(n1384), .CI(
        C[2712]), .CO(C[2713]) );
  FA_5476 \FA_INST_0[5].FA_INST_1[153].FA_  ( .A(A[2713]), .B(n1383), .CI(
        C[2713]), .CO(C[2714]) );
  FA_5475 \FA_INST_0[5].FA_INST_1[154].FA_  ( .A(A[2714]), .B(n1382), .CI(
        C[2714]), .CO(C[2715]) );
  FA_5474 \FA_INST_0[5].FA_INST_1[155].FA_  ( .A(A[2715]), .B(n1381), .CI(
        C[2715]), .CO(C[2716]) );
  FA_5473 \FA_INST_0[5].FA_INST_1[156].FA_  ( .A(A[2716]), .B(n1380), .CI(
        C[2716]), .CO(C[2717]) );
  FA_5472 \FA_INST_0[5].FA_INST_1[157].FA_  ( .A(A[2717]), .B(n1379), .CI(
        C[2717]), .CO(C[2718]) );
  FA_5471 \FA_INST_0[5].FA_INST_1[158].FA_  ( .A(A[2718]), .B(n1378), .CI(
        C[2718]), .CO(C[2719]) );
  FA_5470 \FA_INST_0[5].FA_INST_1[159].FA_  ( .A(A[2719]), .B(n1377), .CI(
        C[2719]), .CO(C[2720]) );
  FA_5469 \FA_INST_0[5].FA_INST_1[160].FA_  ( .A(A[2720]), .B(n1376), .CI(
        C[2720]), .CO(C[2721]) );
  FA_5468 \FA_INST_0[5].FA_INST_1[161].FA_  ( .A(A[2721]), .B(n1375), .CI(
        C[2721]), .CO(C[2722]) );
  FA_5467 \FA_INST_0[5].FA_INST_1[162].FA_  ( .A(A[2722]), .B(n1374), .CI(
        C[2722]), .CO(C[2723]) );
  FA_5466 \FA_INST_0[5].FA_INST_1[163].FA_  ( .A(A[2723]), .B(n1373), .CI(
        C[2723]), .CO(C[2724]) );
  FA_5465 \FA_INST_0[5].FA_INST_1[164].FA_  ( .A(A[2724]), .B(n1372), .CI(
        C[2724]), .CO(C[2725]) );
  FA_5464 \FA_INST_0[5].FA_INST_1[165].FA_  ( .A(A[2725]), .B(n1371), .CI(
        C[2725]), .CO(C[2726]) );
  FA_5463 \FA_INST_0[5].FA_INST_1[166].FA_  ( .A(A[2726]), .B(n1370), .CI(
        C[2726]), .CO(C[2727]) );
  FA_5462 \FA_INST_0[5].FA_INST_1[167].FA_  ( .A(A[2727]), .B(n1369), .CI(
        C[2727]), .CO(C[2728]) );
  FA_5461 \FA_INST_0[5].FA_INST_1[168].FA_  ( .A(A[2728]), .B(n1368), .CI(
        C[2728]), .CO(C[2729]) );
  FA_5460 \FA_INST_0[5].FA_INST_1[169].FA_  ( .A(A[2729]), .B(n1367), .CI(
        C[2729]), .CO(C[2730]) );
  FA_5459 \FA_INST_0[5].FA_INST_1[170].FA_  ( .A(A[2730]), .B(n1366), .CI(
        C[2730]), .CO(C[2731]) );
  FA_5458 \FA_INST_0[5].FA_INST_1[171].FA_  ( .A(A[2731]), .B(n1365), .CI(
        C[2731]), .CO(C[2732]) );
  FA_5457 \FA_INST_0[5].FA_INST_1[172].FA_  ( .A(A[2732]), .B(n1364), .CI(
        C[2732]), .CO(C[2733]) );
  FA_5456 \FA_INST_0[5].FA_INST_1[173].FA_  ( .A(A[2733]), .B(n1363), .CI(
        C[2733]), .CO(C[2734]) );
  FA_5455 \FA_INST_0[5].FA_INST_1[174].FA_  ( .A(A[2734]), .B(n1362), .CI(
        C[2734]), .CO(C[2735]) );
  FA_5454 \FA_INST_0[5].FA_INST_1[175].FA_  ( .A(A[2735]), .B(n1361), .CI(
        C[2735]), .CO(C[2736]) );
  FA_5453 \FA_INST_0[5].FA_INST_1[176].FA_  ( .A(A[2736]), .B(n1360), .CI(
        C[2736]), .CO(C[2737]) );
  FA_5452 \FA_INST_0[5].FA_INST_1[177].FA_  ( .A(A[2737]), .B(n1359), .CI(
        C[2737]), .CO(C[2738]) );
  FA_5451 \FA_INST_0[5].FA_INST_1[178].FA_  ( .A(A[2738]), .B(n1358), .CI(
        C[2738]), .CO(C[2739]) );
  FA_5450 \FA_INST_0[5].FA_INST_1[179].FA_  ( .A(A[2739]), .B(n1357), .CI(
        C[2739]), .CO(C[2740]) );
  FA_5449 \FA_INST_0[5].FA_INST_1[180].FA_  ( .A(A[2740]), .B(n1356), .CI(
        C[2740]), .CO(C[2741]) );
  FA_5448 \FA_INST_0[5].FA_INST_1[181].FA_  ( .A(A[2741]), .B(n1355), .CI(
        C[2741]), .CO(C[2742]) );
  FA_5447 \FA_INST_0[5].FA_INST_1[182].FA_  ( .A(A[2742]), .B(n1354), .CI(
        C[2742]), .CO(C[2743]) );
  FA_5446 \FA_INST_0[5].FA_INST_1[183].FA_  ( .A(A[2743]), .B(n1353), .CI(
        C[2743]), .CO(C[2744]) );
  FA_5445 \FA_INST_0[5].FA_INST_1[184].FA_  ( .A(A[2744]), .B(n1352), .CI(
        C[2744]), .CO(C[2745]) );
  FA_5444 \FA_INST_0[5].FA_INST_1[185].FA_  ( .A(A[2745]), .B(n1351), .CI(
        C[2745]), .CO(C[2746]) );
  FA_5443 \FA_INST_0[5].FA_INST_1[186].FA_  ( .A(A[2746]), .B(n1350), .CI(
        C[2746]), .CO(C[2747]) );
  FA_5442 \FA_INST_0[5].FA_INST_1[187].FA_  ( .A(A[2747]), .B(n1349), .CI(
        C[2747]), .CO(C[2748]) );
  FA_5441 \FA_INST_0[5].FA_INST_1[188].FA_  ( .A(A[2748]), .B(n1348), .CI(
        C[2748]), .CO(C[2749]) );
  FA_5440 \FA_INST_0[5].FA_INST_1[189].FA_  ( .A(A[2749]), .B(n1347), .CI(
        C[2749]), .CO(C[2750]) );
  FA_5439 \FA_INST_0[5].FA_INST_1[190].FA_  ( .A(A[2750]), .B(n1346), .CI(
        C[2750]), .CO(C[2751]) );
  FA_5438 \FA_INST_0[5].FA_INST_1[191].FA_  ( .A(A[2751]), .B(n1345), .CI(
        C[2751]), .CO(C[2752]) );
  FA_5437 \FA_INST_0[5].FA_INST_1[192].FA_  ( .A(A[2752]), .B(n1344), .CI(
        C[2752]), .CO(C[2753]) );
  FA_5436 \FA_INST_0[5].FA_INST_1[193].FA_  ( .A(A[2753]), .B(n1343), .CI(
        C[2753]), .CO(C[2754]) );
  FA_5435 \FA_INST_0[5].FA_INST_1[194].FA_  ( .A(A[2754]), .B(n1342), .CI(
        C[2754]), .CO(C[2755]) );
  FA_5434 \FA_INST_0[5].FA_INST_1[195].FA_  ( .A(A[2755]), .B(n1341), .CI(
        C[2755]), .CO(C[2756]) );
  FA_5433 \FA_INST_0[5].FA_INST_1[196].FA_  ( .A(A[2756]), .B(n1340), .CI(
        C[2756]), .CO(C[2757]) );
  FA_5432 \FA_INST_0[5].FA_INST_1[197].FA_  ( .A(A[2757]), .B(n1339), .CI(
        C[2757]), .CO(C[2758]) );
  FA_5431 \FA_INST_0[5].FA_INST_1[198].FA_  ( .A(A[2758]), .B(n1338), .CI(
        C[2758]), .CO(C[2759]) );
  FA_5430 \FA_INST_0[5].FA_INST_1[199].FA_  ( .A(A[2759]), .B(n1337), .CI(
        C[2759]), .CO(C[2760]) );
  FA_5429 \FA_INST_0[5].FA_INST_1[200].FA_  ( .A(A[2760]), .B(n1336), .CI(
        C[2760]), .CO(C[2761]) );
  FA_5428 \FA_INST_0[5].FA_INST_1[201].FA_  ( .A(A[2761]), .B(n1335), .CI(
        C[2761]), .CO(C[2762]) );
  FA_5427 \FA_INST_0[5].FA_INST_1[202].FA_  ( .A(A[2762]), .B(n1334), .CI(
        C[2762]), .CO(C[2763]) );
  FA_5426 \FA_INST_0[5].FA_INST_1[203].FA_  ( .A(A[2763]), .B(n1333), .CI(
        C[2763]), .CO(C[2764]) );
  FA_5425 \FA_INST_0[5].FA_INST_1[204].FA_  ( .A(A[2764]), .B(n1332), .CI(
        C[2764]), .CO(C[2765]) );
  FA_5424 \FA_INST_0[5].FA_INST_1[205].FA_  ( .A(A[2765]), .B(n1331), .CI(
        C[2765]), .CO(C[2766]) );
  FA_5423 \FA_INST_0[5].FA_INST_1[206].FA_  ( .A(A[2766]), .B(n1330), .CI(
        C[2766]), .CO(C[2767]) );
  FA_5422 \FA_INST_0[5].FA_INST_1[207].FA_  ( .A(A[2767]), .B(n1329), .CI(
        C[2767]), .CO(C[2768]) );
  FA_5421 \FA_INST_0[5].FA_INST_1[208].FA_  ( .A(A[2768]), .B(n1328), .CI(
        C[2768]), .CO(C[2769]) );
  FA_5420 \FA_INST_0[5].FA_INST_1[209].FA_  ( .A(A[2769]), .B(n1327), .CI(
        C[2769]), .CO(C[2770]) );
  FA_5419 \FA_INST_0[5].FA_INST_1[210].FA_  ( .A(A[2770]), .B(n1326), .CI(
        C[2770]), .CO(C[2771]) );
  FA_5418 \FA_INST_0[5].FA_INST_1[211].FA_  ( .A(A[2771]), .B(n1325), .CI(
        C[2771]), .CO(C[2772]) );
  FA_5417 \FA_INST_0[5].FA_INST_1[212].FA_  ( .A(A[2772]), .B(n1324), .CI(
        C[2772]), .CO(C[2773]) );
  FA_5416 \FA_INST_0[5].FA_INST_1[213].FA_  ( .A(A[2773]), .B(n1323), .CI(
        C[2773]), .CO(C[2774]) );
  FA_5415 \FA_INST_0[5].FA_INST_1[214].FA_  ( .A(A[2774]), .B(n1322), .CI(
        C[2774]), .CO(C[2775]) );
  FA_5414 \FA_INST_0[5].FA_INST_1[215].FA_  ( .A(A[2775]), .B(n1321), .CI(
        C[2775]), .CO(C[2776]) );
  FA_5413 \FA_INST_0[5].FA_INST_1[216].FA_  ( .A(A[2776]), .B(n1320), .CI(
        C[2776]), .CO(C[2777]) );
  FA_5412 \FA_INST_0[5].FA_INST_1[217].FA_  ( .A(A[2777]), .B(n1319), .CI(
        C[2777]), .CO(C[2778]) );
  FA_5411 \FA_INST_0[5].FA_INST_1[218].FA_  ( .A(A[2778]), .B(n1318), .CI(
        C[2778]), .CO(C[2779]) );
  FA_5410 \FA_INST_0[5].FA_INST_1[219].FA_  ( .A(A[2779]), .B(n1317), .CI(
        C[2779]), .CO(C[2780]) );
  FA_5409 \FA_INST_0[5].FA_INST_1[220].FA_  ( .A(A[2780]), .B(n1316), .CI(
        C[2780]), .CO(C[2781]) );
  FA_5408 \FA_INST_0[5].FA_INST_1[221].FA_  ( .A(A[2781]), .B(n1315), .CI(
        C[2781]), .CO(C[2782]) );
  FA_5407 \FA_INST_0[5].FA_INST_1[222].FA_  ( .A(A[2782]), .B(n1314), .CI(
        C[2782]), .CO(C[2783]) );
  FA_5406 \FA_INST_0[5].FA_INST_1[223].FA_  ( .A(A[2783]), .B(n1313), .CI(
        C[2783]), .CO(C[2784]) );
  FA_5405 \FA_INST_0[5].FA_INST_1[224].FA_  ( .A(A[2784]), .B(n1312), .CI(
        C[2784]), .CO(C[2785]) );
  FA_5404 \FA_INST_0[5].FA_INST_1[225].FA_  ( .A(A[2785]), .B(n1311), .CI(
        C[2785]), .CO(C[2786]) );
  FA_5403 \FA_INST_0[5].FA_INST_1[226].FA_  ( .A(A[2786]), .B(n1310), .CI(
        C[2786]), .CO(C[2787]) );
  FA_5402 \FA_INST_0[5].FA_INST_1[227].FA_  ( .A(A[2787]), .B(n1309), .CI(
        C[2787]), .CO(C[2788]) );
  FA_5401 \FA_INST_0[5].FA_INST_1[228].FA_  ( .A(A[2788]), .B(n1308), .CI(
        C[2788]), .CO(C[2789]) );
  FA_5400 \FA_INST_0[5].FA_INST_1[229].FA_  ( .A(A[2789]), .B(n1307), .CI(
        C[2789]), .CO(C[2790]) );
  FA_5399 \FA_INST_0[5].FA_INST_1[230].FA_  ( .A(A[2790]), .B(n1306), .CI(
        C[2790]), .CO(C[2791]) );
  FA_5398 \FA_INST_0[5].FA_INST_1[231].FA_  ( .A(A[2791]), .B(n1305), .CI(
        C[2791]), .CO(C[2792]) );
  FA_5397 \FA_INST_0[5].FA_INST_1[232].FA_  ( .A(A[2792]), .B(n1304), .CI(
        C[2792]), .CO(C[2793]) );
  FA_5396 \FA_INST_0[5].FA_INST_1[233].FA_  ( .A(A[2793]), .B(n1303), .CI(
        C[2793]), .CO(C[2794]) );
  FA_5395 \FA_INST_0[5].FA_INST_1[234].FA_  ( .A(A[2794]), .B(n1302), .CI(
        C[2794]), .CO(C[2795]) );
  FA_5394 \FA_INST_0[5].FA_INST_1[235].FA_  ( .A(A[2795]), .B(n1301), .CI(
        C[2795]), .CO(C[2796]) );
  FA_5393 \FA_INST_0[5].FA_INST_1[236].FA_  ( .A(A[2796]), .B(n1300), .CI(
        C[2796]), .CO(C[2797]) );
  FA_5392 \FA_INST_0[5].FA_INST_1[237].FA_  ( .A(A[2797]), .B(n1299), .CI(
        C[2797]), .CO(C[2798]) );
  FA_5391 \FA_INST_0[5].FA_INST_1[238].FA_  ( .A(A[2798]), .B(n1298), .CI(
        C[2798]), .CO(C[2799]) );
  FA_5390 \FA_INST_0[5].FA_INST_1[239].FA_  ( .A(A[2799]), .B(n1297), .CI(
        C[2799]), .CO(C[2800]) );
  FA_5389 \FA_INST_0[5].FA_INST_1[240].FA_  ( .A(A[2800]), .B(n1296), .CI(
        C[2800]), .CO(C[2801]) );
  FA_5388 \FA_INST_0[5].FA_INST_1[241].FA_  ( .A(A[2801]), .B(n1295), .CI(
        C[2801]), .CO(C[2802]) );
  FA_5387 \FA_INST_0[5].FA_INST_1[242].FA_  ( .A(A[2802]), .B(n1294), .CI(
        C[2802]), .CO(C[2803]) );
  FA_5386 \FA_INST_0[5].FA_INST_1[243].FA_  ( .A(A[2803]), .B(n1293), .CI(
        C[2803]), .CO(C[2804]) );
  FA_5385 \FA_INST_0[5].FA_INST_1[244].FA_  ( .A(A[2804]), .B(n1292), .CI(
        C[2804]), .CO(C[2805]) );
  FA_5384 \FA_INST_0[5].FA_INST_1[245].FA_  ( .A(A[2805]), .B(n1291), .CI(
        C[2805]), .CO(C[2806]) );
  FA_5383 \FA_INST_0[5].FA_INST_1[246].FA_  ( .A(A[2806]), .B(n1290), .CI(
        C[2806]), .CO(C[2807]) );
  FA_5382 \FA_INST_0[5].FA_INST_1[247].FA_  ( .A(A[2807]), .B(n1289), .CI(
        C[2807]), .CO(C[2808]) );
  FA_5381 \FA_INST_0[5].FA_INST_1[248].FA_  ( .A(A[2808]), .B(n1288), .CI(
        C[2808]), .CO(C[2809]) );
  FA_5380 \FA_INST_0[5].FA_INST_1[249].FA_  ( .A(A[2809]), .B(n1287), .CI(
        C[2809]), .CO(C[2810]) );
  FA_5379 \FA_INST_0[5].FA_INST_1[250].FA_  ( .A(A[2810]), .B(n1286), .CI(
        C[2810]), .CO(C[2811]) );
  FA_5378 \FA_INST_0[5].FA_INST_1[251].FA_  ( .A(A[2811]), .B(n1285), .CI(
        C[2811]), .CO(C[2812]) );
  FA_5377 \FA_INST_0[5].FA_INST_1[252].FA_  ( .A(A[2812]), .B(n1284), .CI(
        C[2812]), .CO(C[2813]) );
  FA_5376 \FA_INST_0[5].FA_INST_1[253].FA_  ( .A(A[2813]), .B(n1283), .CI(
        C[2813]), .CO(C[2814]) );
  FA_5375 \FA_INST_0[5].FA_INST_1[254].FA_  ( .A(A[2814]), .B(n1282), .CI(
        C[2814]), .CO(C[2815]) );
  FA_5374 \FA_INST_0[5].FA_INST_1[255].FA_  ( .A(A[2815]), .B(n1281), .CI(
        C[2815]), .CO(C[2816]) );
  FA_5373 \FA_INST_0[5].FA_INST_1[256].FA_  ( .A(A[2816]), .B(n1280), .CI(
        C[2816]), .CO(C[2817]) );
  FA_5372 \FA_INST_0[5].FA_INST_1[257].FA_  ( .A(A[2817]), .B(n1279), .CI(
        C[2817]), .CO(C[2818]) );
  FA_5371 \FA_INST_0[5].FA_INST_1[258].FA_  ( .A(A[2818]), .B(n1278), .CI(
        C[2818]), .CO(C[2819]) );
  FA_5370 \FA_INST_0[5].FA_INST_1[259].FA_  ( .A(A[2819]), .B(n1277), .CI(
        C[2819]), .CO(C[2820]) );
  FA_5369 \FA_INST_0[5].FA_INST_1[260].FA_  ( .A(A[2820]), .B(n1276), .CI(
        C[2820]), .CO(C[2821]) );
  FA_5368 \FA_INST_0[5].FA_INST_1[261].FA_  ( .A(A[2821]), .B(n1275), .CI(
        C[2821]), .CO(C[2822]) );
  FA_5367 \FA_INST_0[5].FA_INST_1[262].FA_  ( .A(A[2822]), .B(n1274), .CI(
        C[2822]), .CO(C[2823]) );
  FA_5366 \FA_INST_0[5].FA_INST_1[263].FA_  ( .A(A[2823]), .B(n1273), .CI(
        C[2823]), .CO(C[2824]) );
  FA_5365 \FA_INST_0[5].FA_INST_1[264].FA_  ( .A(A[2824]), .B(n1272), .CI(
        C[2824]), .CO(C[2825]) );
  FA_5364 \FA_INST_0[5].FA_INST_1[265].FA_  ( .A(A[2825]), .B(n1271), .CI(
        C[2825]), .CO(C[2826]) );
  FA_5363 \FA_INST_0[5].FA_INST_1[266].FA_  ( .A(A[2826]), .B(n1270), .CI(
        C[2826]), .CO(C[2827]) );
  FA_5362 \FA_INST_0[5].FA_INST_1[267].FA_  ( .A(A[2827]), .B(n1269), .CI(
        C[2827]), .CO(C[2828]) );
  FA_5361 \FA_INST_0[5].FA_INST_1[268].FA_  ( .A(A[2828]), .B(n1268), .CI(
        C[2828]), .CO(C[2829]) );
  FA_5360 \FA_INST_0[5].FA_INST_1[269].FA_  ( .A(A[2829]), .B(n1267), .CI(
        C[2829]), .CO(C[2830]) );
  FA_5359 \FA_INST_0[5].FA_INST_1[270].FA_  ( .A(A[2830]), .B(n1266), .CI(
        C[2830]), .CO(C[2831]) );
  FA_5358 \FA_INST_0[5].FA_INST_1[271].FA_  ( .A(A[2831]), .B(n1265), .CI(
        C[2831]), .CO(C[2832]) );
  FA_5357 \FA_INST_0[5].FA_INST_1[272].FA_  ( .A(A[2832]), .B(n1264), .CI(
        C[2832]), .CO(C[2833]) );
  FA_5356 \FA_INST_0[5].FA_INST_1[273].FA_  ( .A(A[2833]), .B(n1263), .CI(
        C[2833]), .CO(C[2834]) );
  FA_5355 \FA_INST_0[5].FA_INST_1[274].FA_  ( .A(A[2834]), .B(n1262), .CI(
        C[2834]), .CO(C[2835]) );
  FA_5354 \FA_INST_0[5].FA_INST_1[275].FA_  ( .A(A[2835]), .B(n1261), .CI(
        C[2835]), .CO(C[2836]) );
  FA_5353 \FA_INST_0[5].FA_INST_1[276].FA_  ( .A(A[2836]), .B(n1260), .CI(
        C[2836]), .CO(C[2837]) );
  FA_5352 \FA_INST_0[5].FA_INST_1[277].FA_  ( .A(A[2837]), .B(n1259), .CI(
        C[2837]), .CO(C[2838]) );
  FA_5351 \FA_INST_0[5].FA_INST_1[278].FA_  ( .A(A[2838]), .B(n1258), .CI(
        C[2838]), .CO(C[2839]) );
  FA_5350 \FA_INST_0[5].FA_INST_1[279].FA_  ( .A(A[2839]), .B(n1257), .CI(
        C[2839]), .CO(C[2840]) );
  FA_5349 \FA_INST_0[5].FA_INST_1[280].FA_  ( .A(A[2840]), .B(n1256), .CI(
        C[2840]), .CO(C[2841]) );
  FA_5348 \FA_INST_0[5].FA_INST_1[281].FA_  ( .A(A[2841]), .B(n1255), .CI(
        C[2841]), .CO(C[2842]) );
  FA_5347 \FA_INST_0[5].FA_INST_1[282].FA_  ( .A(A[2842]), .B(n1254), .CI(
        C[2842]), .CO(C[2843]) );
  FA_5346 \FA_INST_0[5].FA_INST_1[283].FA_  ( .A(A[2843]), .B(n1253), .CI(
        C[2843]), .CO(C[2844]) );
  FA_5345 \FA_INST_0[5].FA_INST_1[284].FA_  ( .A(A[2844]), .B(n1252), .CI(
        C[2844]), .CO(C[2845]) );
  FA_5344 \FA_INST_0[5].FA_INST_1[285].FA_  ( .A(A[2845]), .B(n1251), .CI(
        C[2845]), .CO(C[2846]) );
  FA_5343 \FA_INST_0[5].FA_INST_1[286].FA_  ( .A(A[2846]), .B(n1250), .CI(
        C[2846]), .CO(C[2847]) );
  FA_5342 \FA_INST_0[5].FA_INST_1[287].FA_  ( .A(A[2847]), .B(n1249), .CI(
        C[2847]), .CO(C[2848]) );
  FA_5341 \FA_INST_0[5].FA_INST_1[288].FA_  ( .A(A[2848]), .B(n1248), .CI(
        C[2848]), .CO(C[2849]) );
  FA_5340 \FA_INST_0[5].FA_INST_1[289].FA_  ( .A(A[2849]), .B(n1247), .CI(
        C[2849]), .CO(C[2850]) );
  FA_5339 \FA_INST_0[5].FA_INST_1[290].FA_  ( .A(A[2850]), .B(n1246), .CI(
        C[2850]), .CO(C[2851]) );
  FA_5338 \FA_INST_0[5].FA_INST_1[291].FA_  ( .A(A[2851]), .B(n1245), .CI(
        C[2851]), .CO(C[2852]) );
  FA_5337 \FA_INST_0[5].FA_INST_1[292].FA_  ( .A(A[2852]), .B(n1244), .CI(
        C[2852]), .CO(C[2853]) );
  FA_5336 \FA_INST_0[5].FA_INST_1[293].FA_  ( .A(A[2853]), .B(n1243), .CI(
        C[2853]), .CO(C[2854]) );
  FA_5335 \FA_INST_0[5].FA_INST_1[294].FA_  ( .A(A[2854]), .B(n1242), .CI(
        C[2854]), .CO(C[2855]) );
  FA_5334 \FA_INST_0[5].FA_INST_1[295].FA_  ( .A(A[2855]), .B(n1241), .CI(
        C[2855]), .CO(C[2856]) );
  FA_5333 \FA_INST_0[5].FA_INST_1[296].FA_  ( .A(A[2856]), .B(n1240), .CI(
        C[2856]), .CO(C[2857]) );
  FA_5332 \FA_INST_0[5].FA_INST_1[297].FA_  ( .A(A[2857]), .B(n1239), .CI(
        C[2857]), .CO(C[2858]) );
  FA_5331 \FA_INST_0[5].FA_INST_1[298].FA_  ( .A(A[2858]), .B(n1238), .CI(
        C[2858]), .CO(C[2859]) );
  FA_5330 \FA_INST_0[5].FA_INST_1[299].FA_  ( .A(A[2859]), .B(n1237), .CI(
        C[2859]), .CO(C[2860]) );
  FA_5329 \FA_INST_0[5].FA_INST_1[300].FA_  ( .A(A[2860]), .B(n1236), .CI(
        C[2860]), .CO(C[2861]) );
  FA_5328 \FA_INST_0[5].FA_INST_1[301].FA_  ( .A(A[2861]), .B(n1235), .CI(
        C[2861]), .CO(C[2862]) );
  FA_5327 \FA_INST_0[5].FA_INST_1[302].FA_  ( .A(A[2862]), .B(n1234), .CI(
        C[2862]), .CO(C[2863]) );
  FA_5326 \FA_INST_0[5].FA_INST_1[303].FA_  ( .A(A[2863]), .B(n1233), .CI(
        C[2863]), .CO(C[2864]) );
  FA_5325 \FA_INST_0[5].FA_INST_1[304].FA_  ( .A(A[2864]), .B(n1232), .CI(
        C[2864]), .CO(C[2865]) );
  FA_5324 \FA_INST_0[5].FA_INST_1[305].FA_  ( .A(A[2865]), .B(n1231), .CI(
        C[2865]), .CO(C[2866]) );
  FA_5323 \FA_INST_0[5].FA_INST_1[306].FA_  ( .A(A[2866]), .B(n1230), .CI(
        C[2866]), .CO(C[2867]) );
  FA_5322 \FA_INST_0[5].FA_INST_1[307].FA_  ( .A(A[2867]), .B(n1229), .CI(
        C[2867]), .CO(C[2868]) );
  FA_5321 \FA_INST_0[5].FA_INST_1[308].FA_  ( .A(A[2868]), .B(n1228), .CI(
        C[2868]), .CO(C[2869]) );
  FA_5320 \FA_INST_0[5].FA_INST_1[309].FA_  ( .A(A[2869]), .B(n1227), .CI(
        C[2869]), .CO(C[2870]) );
  FA_5319 \FA_INST_0[5].FA_INST_1[310].FA_  ( .A(A[2870]), .B(n1226), .CI(
        C[2870]), .CO(C[2871]) );
  FA_5318 \FA_INST_0[5].FA_INST_1[311].FA_  ( .A(A[2871]), .B(n1225), .CI(
        C[2871]), .CO(C[2872]) );
  FA_5317 \FA_INST_0[5].FA_INST_1[312].FA_  ( .A(A[2872]), .B(n1224), .CI(
        C[2872]), .CO(C[2873]) );
  FA_5316 \FA_INST_0[5].FA_INST_1[313].FA_  ( .A(A[2873]), .B(n1223), .CI(
        C[2873]), .CO(C[2874]) );
  FA_5315 \FA_INST_0[5].FA_INST_1[314].FA_  ( .A(A[2874]), .B(n1222), .CI(
        C[2874]), .CO(C[2875]) );
  FA_5314 \FA_INST_0[5].FA_INST_1[315].FA_  ( .A(A[2875]), .B(n1221), .CI(
        C[2875]), .CO(C[2876]) );
  FA_5313 \FA_INST_0[5].FA_INST_1[316].FA_  ( .A(A[2876]), .B(n1220), .CI(
        C[2876]), .CO(C[2877]) );
  FA_5312 \FA_INST_0[5].FA_INST_1[317].FA_  ( .A(A[2877]), .B(n1219), .CI(
        C[2877]), .CO(C[2878]) );
  FA_5311 \FA_INST_0[5].FA_INST_1[318].FA_  ( .A(A[2878]), .B(n1218), .CI(
        C[2878]), .CO(C[2879]) );
  FA_5310 \FA_INST_0[5].FA_INST_1[319].FA_  ( .A(A[2879]), .B(n1217), .CI(
        C[2879]), .CO(C[2880]) );
  FA_5309 \FA_INST_0[5].FA_INST_1[320].FA_  ( .A(A[2880]), .B(n1216), .CI(
        C[2880]), .CO(C[2881]) );
  FA_5308 \FA_INST_0[5].FA_INST_1[321].FA_  ( .A(A[2881]), .B(n1215), .CI(
        C[2881]), .CO(C[2882]) );
  FA_5307 \FA_INST_0[5].FA_INST_1[322].FA_  ( .A(A[2882]), .B(n1214), .CI(
        C[2882]), .CO(C[2883]) );
  FA_5306 \FA_INST_0[5].FA_INST_1[323].FA_  ( .A(A[2883]), .B(n1213), .CI(
        C[2883]), .CO(C[2884]) );
  FA_5305 \FA_INST_0[5].FA_INST_1[324].FA_  ( .A(A[2884]), .B(n1212), .CI(
        C[2884]), .CO(C[2885]) );
  FA_5304 \FA_INST_0[5].FA_INST_1[325].FA_  ( .A(A[2885]), .B(n1211), .CI(
        C[2885]), .CO(C[2886]) );
  FA_5303 \FA_INST_0[5].FA_INST_1[326].FA_  ( .A(A[2886]), .B(n1210), .CI(
        C[2886]), .CO(C[2887]) );
  FA_5302 \FA_INST_0[5].FA_INST_1[327].FA_  ( .A(A[2887]), .B(n1209), .CI(
        C[2887]), .CO(C[2888]) );
  FA_5301 \FA_INST_0[5].FA_INST_1[328].FA_  ( .A(A[2888]), .B(n1208), .CI(
        C[2888]), .CO(C[2889]) );
  FA_5300 \FA_INST_0[5].FA_INST_1[329].FA_  ( .A(A[2889]), .B(n1207), .CI(
        C[2889]), .CO(C[2890]) );
  FA_5299 \FA_INST_0[5].FA_INST_1[330].FA_  ( .A(A[2890]), .B(n1206), .CI(
        C[2890]), .CO(C[2891]) );
  FA_5298 \FA_INST_0[5].FA_INST_1[331].FA_  ( .A(A[2891]), .B(n1205), .CI(
        C[2891]), .CO(C[2892]) );
  FA_5297 \FA_INST_0[5].FA_INST_1[332].FA_  ( .A(A[2892]), .B(n1204), .CI(
        C[2892]), .CO(C[2893]) );
  FA_5296 \FA_INST_0[5].FA_INST_1[333].FA_  ( .A(A[2893]), .B(n1203), .CI(
        C[2893]), .CO(C[2894]) );
  FA_5295 \FA_INST_0[5].FA_INST_1[334].FA_  ( .A(A[2894]), .B(n1202), .CI(
        C[2894]), .CO(C[2895]) );
  FA_5294 \FA_INST_0[5].FA_INST_1[335].FA_  ( .A(A[2895]), .B(n1201), .CI(
        C[2895]), .CO(C[2896]) );
  FA_5293 \FA_INST_0[5].FA_INST_1[336].FA_  ( .A(A[2896]), .B(n1200), .CI(
        C[2896]), .CO(C[2897]) );
  FA_5292 \FA_INST_0[5].FA_INST_1[337].FA_  ( .A(A[2897]), .B(n1199), .CI(
        C[2897]), .CO(C[2898]) );
  FA_5291 \FA_INST_0[5].FA_INST_1[338].FA_  ( .A(A[2898]), .B(n1198), .CI(
        C[2898]), .CO(C[2899]) );
  FA_5290 \FA_INST_0[5].FA_INST_1[339].FA_  ( .A(A[2899]), .B(n1197), .CI(
        C[2899]), .CO(C[2900]) );
  FA_5289 \FA_INST_0[5].FA_INST_1[340].FA_  ( .A(A[2900]), .B(n1196), .CI(
        C[2900]), .CO(C[2901]) );
  FA_5288 \FA_INST_0[5].FA_INST_1[341].FA_  ( .A(A[2901]), .B(n1195), .CI(
        C[2901]), .CO(C[2902]) );
  FA_5287 \FA_INST_0[5].FA_INST_1[342].FA_  ( .A(A[2902]), .B(n1194), .CI(
        C[2902]), .CO(C[2903]) );
  FA_5286 \FA_INST_0[5].FA_INST_1[343].FA_  ( .A(A[2903]), .B(n1193), .CI(
        C[2903]), .CO(C[2904]) );
  FA_5285 \FA_INST_0[5].FA_INST_1[344].FA_  ( .A(A[2904]), .B(n1192), .CI(
        C[2904]), .CO(C[2905]) );
  FA_5284 \FA_INST_0[5].FA_INST_1[345].FA_  ( .A(A[2905]), .B(n1191), .CI(
        C[2905]), .CO(C[2906]) );
  FA_5283 \FA_INST_0[5].FA_INST_1[346].FA_  ( .A(A[2906]), .B(n1190), .CI(
        C[2906]), .CO(C[2907]) );
  FA_5282 \FA_INST_0[5].FA_INST_1[347].FA_  ( .A(A[2907]), .B(n1189), .CI(
        C[2907]), .CO(C[2908]) );
  FA_5281 \FA_INST_0[5].FA_INST_1[348].FA_  ( .A(A[2908]), .B(n1188), .CI(
        C[2908]), .CO(C[2909]) );
  FA_5280 \FA_INST_0[5].FA_INST_1[349].FA_  ( .A(A[2909]), .B(n1187), .CI(
        C[2909]), .CO(C[2910]) );
  FA_5279 \FA_INST_0[5].FA_INST_1[350].FA_  ( .A(A[2910]), .B(n1186), .CI(
        C[2910]), .CO(C[2911]) );
  FA_5278 \FA_INST_0[5].FA_INST_1[351].FA_  ( .A(A[2911]), .B(n1185), .CI(
        C[2911]), .CO(C[2912]) );
  FA_5277 \FA_INST_0[5].FA_INST_1[352].FA_  ( .A(A[2912]), .B(n1184), .CI(
        C[2912]), .CO(C[2913]) );
  FA_5276 \FA_INST_0[5].FA_INST_1[353].FA_  ( .A(A[2913]), .B(n1183), .CI(
        C[2913]), .CO(C[2914]) );
  FA_5275 \FA_INST_0[5].FA_INST_1[354].FA_  ( .A(A[2914]), .B(n1182), .CI(
        C[2914]), .CO(C[2915]) );
  FA_5274 \FA_INST_0[5].FA_INST_1[355].FA_  ( .A(A[2915]), .B(n1181), .CI(
        C[2915]), .CO(C[2916]) );
  FA_5273 \FA_INST_0[5].FA_INST_1[356].FA_  ( .A(A[2916]), .B(n1180), .CI(
        C[2916]), .CO(C[2917]) );
  FA_5272 \FA_INST_0[5].FA_INST_1[357].FA_  ( .A(A[2917]), .B(n1179), .CI(
        C[2917]), .CO(C[2918]) );
  FA_5271 \FA_INST_0[5].FA_INST_1[358].FA_  ( .A(A[2918]), .B(n1178), .CI(
        C[2918]), .CO(C[2919]) );
  FA_5270 \FA_INST_0[5].FA_INST_1[359].FA_  ( .A(A[2919]), .B(n1177), .CI(
        C[2919]), .CO(C[2920]) );
  FA_5269 \FA_INST_0[5].FA_INST_1[360].FA_  ( .A(A[2920]), .B(n1176), .CI(
        C[2920]), .CO(C[2921]) );
  FA_5268 \FA_INST_0[5].FA_INST_1[361].FA_  ( .A(A[2921]), .B(n1175), .CI(
        C[2921]), .CO(C[2922]) );
  FA_5267 \FA_INST_0[5].FA_INST_1[362].FA_  ( .A(A[2922]), .B(n1174), .CI(
        C[2922]), .CO(C[2923]) );
  FA_5266 \FA_INST_0[5].FA_INST_1[363].FA_  ( .A(A[2923]), .B(n1173), .CI(
        C[2923]), .CO(C[2924]) );
  FA_5265 \FA_INST_0[5].FA_INST_1[364].FA_  ( .A(A[2924]), .B(n1172), .CI(
        C[2924]), .CO(C[2925]) );
  FA_5264 \FA_INST_0[5].FA_INST_1[365].FA_  ( .A(A[2925]), .B(n1171), .CI(
        C[2925]), .CO(C[2926]) );
  FA_5263 \FA_INST_0[5].FA_INST_1[366].FA_  ( .A(A[2926]), .B(n1170), .CI(
        C[2926]), .CO(C[2927]) );
  FA_5262 \FA_INST_0[5].FA_INST_1[367].FA_  ( .A(A[2927]), .B(n1169), .CI(
        C[2927]), .CO(C[2928]) );
  FA_5261 \FA_INST_0[5].FA_INST_1[368].FA_  ( .A(A[2928]), .B(n1168), .CI(
        C[2928]), .CO(C[2929]) );
  FA_5260 \FA_INST_0[5].FA_INST_1[369].FA_  ( .A(A[2929]), .B(n1167), .CI(
        C[2929]), .CO(C[2930]) );
  FA_5259 \FA_INST_0[5].FA_INST_1[370].FA_  ( .A(A[2930]), .B(n1166), .CI(
        C[2930]), .CO(C[2931]) );
  FA_5258 \FA_INST_0[5].FA_INST_1[371].FA_  ( .A(A[2931]), .B(n1165), .CI(
        C[2931]), .CO(C[2932]) );
  FA_5257 \FA_INST_0[5].FA_INST_1[372].FA_  ( .A(A[2932]), .B(n1164), .CI(
        C[2932]), .CO(C[2933]) );
  FA_5256 \FA_INST_0[5].FA_INST_1[373].FA_  ( .A(A[2933]), .B(n1163), .CI(
        C[2933]), .CO(C[2934]) );
  FA_5255 \FA_INST_0[5].FA_INST_1[374].FA_  ( .A(A[2934]), .B(n1162), .CI(
        C[2934]), .CO(C[2935]) );
  FA_5254 \FA_INST_0[5].FA_INST_1[375].FA_  ( .A(A[2935]), .B(n1161), .CI(
        C[2935]), .CO(C[2936]) );
  FA_5253 \FA_INST_0[5].FA_INST_1[376].FA_  ( .A(A[2936]), .B(n1160), .CI(
        C[2936]), .CO(C[2937]) );
  FA_5252 \FA_INST_0[5].FA_INST_1[377].FA_  ( .A(A[2937]), .B(n1159), .CI(
        C[2937]), .CO(C[2938]) );
  FA_5251 \FA_INST_0[5].FA_INST_1[378].FA_  ( .A(A[2938]), .B(n1158), .CI(
        C[2938]), .CO(C[2939]) );
  FA_5250 \FA_INST_0[5].FA_INST_1[379].FA_  ( .A(A[2939]), .B(n1157), .CI(
        C[2939]), .CO(C[2940]) );
  FA_5249 \FA_INST_0[5].FA_INST_1[380].FA_  ( .A(A[2940]), .B(n1156), .CI(
        C[2940]), .CO(C[2941]) );
  FA_5248 \FA_INST_0[5].FA_INST_1[381].FA_  ( .A(A[2941]), .B(n1155), .CI(
        C[2941]), .CO(C[2942]) );
  FA_5247 \FA_INST_0[5].FA_INST_1[382].FA_  ( .A(A[2942]), .B(n1154), .CI(
        C[2942]), .CO(C[2943]) );
  FA_5246 \FA_INST_0[5].FA_INST_1[383].FA_  ( .A(A[2943]), .B(n1153), .CI(
        C[2943]), .CO(C[2944]) );
  FA_5245 \FA_INST_0[5].FA_INST_1[384].FA_  ( .A(A[2944]), .B(n1152), .CI(
        C[2944]), .CO(C[2945]) );
  FA_5244 \FA_INST_0[5].FA_INST_1[385].FA_  ( .A(A[2945]), .B(n1151), .CI(
        C[2945]), .CO(C[2946]) );
  FA_5243 \FA_INST_0[5].FA_INST_1[386].FA_  ( .A(A[2946]), .B(n1150), .CI(
        C[2946]), .CO(C[2947]) );
  FA_5242 \FA_INST_0[5].FA_INST_1[387].FA_  ( .A(A[2947]), .B(n1149), .CI(
        C[2947]), .CO(C[2948]) );
  FA_5241 \FA_INST_0[5].FA_INST_1[388].FA_  ( .A(A[2948]), .B(n1148), .CI(
        C[2948]), .CO(C[2949]) );
  FA_5240 \FA_INST_0[5].FA_INST_1[389].FA_  ( .A(A[2949]), .B(n1147), .CI(
        C[2949]), .CO(C[2950]) );
  FA_5239 \FA_INST_0[5].FA_INST_1[390].FA_  ( .A(A[2950]), .B(n1146), .CI(
        C[2950]), .CO(C[2951]) );
  FA_5238 \FA_INST_0[5].FA_INST_1[391].FA_  ( .A(A[2951]), .B(n1145), .CI(
        C[2951]), .CO(C[2952]) );
  FA_5237 \FA_INST_0[5].FA_INST_1[392].FA_  ( .A(A[2952]), .B(n1144), .CI(
        C[2952]), .CO(C[2953]) );
  FA_5236 \FA_INST_0[5].FA_INST_1[393].FA_  ( .A(A[2953]), .B(n1143), .CI(
        C[2953]), .CO(C[2954]) );
  FA_5235 \FA_INST_0[5].FA_INST_1[394].FA_  ( .A(A[2954]), .B(n1142), .CI(
        C[2954]), .CO(C[2955]) );
  FA_5234 \FA_INST_0[5].FA_INST_1[395].FA_  ( .A(A[2955]), .B(n1141), .CI(
        C[2955]), .CO(C[2956]) );
  FA_5233 \FA_INST_0[5].FA_INST_1[396].FA_  ( .A(A[2956]), .B(n1140), .CI(
        C[2956]), .CO(C[2957]) );
  FA_5232 \FA_INST_0[5].FA_INST_1[397].FA_  ( .A(A[2957]), .B(n1139), .CI(
        C[2957]), .CO(C[2958]) );
  FA_5231 \FA_INST_0[5].FA_INST_1[398].FA_  ( .A(A[2958]), .B(n1138), .CI(
        C[2958]), .CO(C[2959]) );
  FA_5230 \FA_INST_0[5].FA_INST_1[399].FA_  ( .A(A[2959]), .B(n1137), .CI(
        C[2959]), .CO(C[2960]) );
  FA_5229 \FA_INST_0[5].FA_INST_1[400].FA_  ( .A(A[2960]), .B(n1136), .CI(
        C[2960]), .CO(C[2961]) );
  FA_5228 \FA_INST_0[5].FA_INST_1[401].FA_  ( .A(A[2961]), .B(n1135), .CI(
        C[2961]), .CO(C[2962]) );
  FA_5227 \FA_INST_0[5].FA_INST_1[402].FA_  ( .A(A[2962]), .B(n1134), .CI(
        C[2962]), .CO(C[2963]) );
  FA_5226 \FA_INST_0[5].FA_INST_1[403].FA_  ( .A(A[2963]), .B(n1133), .CI(
        C[2963]), .CO(C[2964]) );
  FA_5225 \FA_INST_0[5].FA_INST_1[404].FA_  ( .A(A[2964]), .B(n1132), .CI(
        C[2964]), .CO(C[2965]) );
  FA_5224 \FA_INST_0[5].FA_INST_1[405].FA_  ( .A(A[2965]), .B(n1131), .CI(
        C[2965]), .CO(C[2966]) );
  FA_5223 \FA_INST_0[5].FA_INST_1[406].FA_  ( .A(A[2966]), .B(n1130), .CI(
        C[2966]), .CO(C[2967]) );
  FA_5222 \FA_INST_0[5].FA_INST_1[407].FA_  ( .A(A[2967]), .B(n1129), .CI(
        C[2967]), .CO(C[2968]) );
  FA_5221 \FA_INST_0[5].FA_INST_1[408].FA_  ( .A(A[2968]), .B(n1128), .CI(
        C[2968]), .CO(C[2969]) );
  FA_5220 \FA_INST_0[5].FA_INST_1[409].FA_  ( .A(A[2969]), .B(n1127), .CI(
        C[2969]), .CO(C[2970]) );
  FA_5219 \FA_INST_0[5].FA_INST_1[410].FA_  ( .A(A[2970]), .B(n1126), .CI(
        C[2970]), .CO(C[2971]) );
  FA_5218 \FA_INST_0[5].FA_INST_1[411].FA_  ( .A(A[2971]), .B(n1125), .CI(
        C[2971]), .CO(C[2972]) );
  FA_5217 \FA_INST_0[5].FA_INST_1[412].FA_  ( .A(A[2972]), .B(n1124), .CI(
        C[2972]), .CO(C[2973]) );
  FA_5216 \FA_INST_0[5].FA_INST_1[413].FA_  ( .A(A[2973]), .B(n1123), .CI(
        C[2973]), .CO(C[2974]) );
  FA_5215 \FA_INST_0[5].FA_INST_1[414].FA_  ( .A(A[2974]), .B(n1122), .CI(
        C[2974]), .CO(C[2975]) );
  FA_5214 \FA_INST_0[5].FA_INST_1[415].FA_  ( .A(A[2975]), .B(n1121), .CI(
        C[2975]), .CO(C[2976]) );
  FA_5213 \FA_INST_0[5].FA_INST_1[416].FA_  ( .A(A[2976]), .B(n1120), .CI(
        C[2976]), .CO(C[2977]) );
  FA_5212 \FA_INST_0[5].FA_INST_1[417].FA_  ( .A(A[2977]), .B(n1119), .CI(
        C[2977]), .CO(C[2978]) );
  FA_5211 \FA_INST_0[5].FA_INST_1[418].FA_  ( .A(A[2978]), .B(n1118), .CI(
        C[2978]), .CO(C[2979]) );
  FA_5210 \FA_INST_0[5].FA_INST_1[419].FA_  ( .A(A[2979]), .B(n1117), .CI(
        C[2979]), .CO(C[2980]) );
  FA_5209 \FA_INST_0[5].FA_INST_1[420].FA_  ( .A(A[2980]), .B(n1116), .CI(
        C[2980]), .CO(C[2981]) );
  FA_5208 \FA_INST_0[5].FA_INST_1[421].FA_  ( .A(A[2981]), .B(n1115), .CI(
        C[2981]), .CO(C[2982]) );
  FA_5207 \FA_INST_0[5].FA_INST_1[422].FA_  ( .A(A[2982]), .B(n1114), .CI(
        C[2982]), .CO(C[2983]) );
  FA_5206 \FA_INST_0[5].FA_INST_1[423].FA_  ( .A(A[2983]), .B(n1113), .CI(
        C[2983]), .CO(C[2984]) );
  FA_5205 \FA_INST_0[5].FA_INST_1[424].FA_  ( .A(A[2984]), .B(n1112), .CI(
        C[2984]), .CO(C[2985]) );
  FA_5204 \FA_INST_0[5].FA_INST_1[425].FA_  ( .A(A[2985]), .B(n1111), .CI(
        C[2985]), .CO(C[2986]) );
  FA_5203 \FA_INST_0[5].FA_INST_1[426].FA_  ( .A(A[2986]), .B(n1110), .CI(
        C[2986]), .CO(C[2987]) );
  FA_5202 \FA_INST_0[5].FA_INST_1[427].FA_  ( .A(A[2987]), .B(n1109), .CI(
        C[2987]), .CO(C[2988]) );
  FA_5201 \FA_INST_0[5].FA_INST_1[428].FA_  ( .A(A[2988]), .B(n1108), .CI(
        C[2988]), .CO(C[2989]) );
  FA_5200 \FA_INST_0[5].FA_INST_1[429].FA_  ( .A(A[2989]), .B(n1107), .CI(
        C[2989]), .CO(C[2990]) );
  FA_5199 \FA_INST_0[5].FA_INST_1[430].FA_  ( .A(A[2990]), .B(n1106), .CI(
        C[2990]), .CO(C[2991]) );
  FA_5198 \FA_INST_0[5].FA_INST_1[431].FA_  ( .A(A[2991]), .B(n1105), .CI(
        C[2991]), .CO(C[2992]) );
  FA_5197 \FA_INST_0[5].FA_INST_1[432].FA_  ( .A(A[2992]), .B(n1104), .CI(
        C[2992]), .CO(C[2993]) );
  FA_5196 \FA_INST_0[5].FA_INST_1[433].FA_  ( .A(A[2993]), .B(n1103), .CI(
        C[2993]), .CO(C[2994]) );
  FA_5195 \FA_INST_0[5].FA_INST_1[434].FA_  ( .A(A[2994]), .B(n1102), .CI(
        C[2994]), .CO(C[2995]) );
  FA_5194 \FA_INST_0[5].FA_INST_1[435].FA_  ( .A(A[2995]), .B(n1101), .CI(
        C[2995]), .CO(C[2996]) );
  FA_5193 \FA_INST_0[5].FA_INST_1[436].FA_  ( .A(A[2996]), .B(n1100), .CI(
        C[2996]), .CO(C[2997]) );
  FA_5192 \FA_INST_0[5].FA_INST_1[437].FA_  ( .A(A[2997]), .B(n1099), .CI(
        C[2997]), .CO(C[2998]) );
  FA_5191 \FA_INST_0[5].FA_INST_1[438].FA_  ( .A(A[2998]), .B(n1098), .CI(
        C[2998]), .CO(C[2999]) );
  FA_5190 \FA_INST_0[5].FA_INST_1[439].FA_  ( .A(A[2999]), .B(n1097), .CI(
        C[2999]), .CO(C[3000]) );
  FA_5189 \FA_INST_0[5].FA_INST_1[440].FA_  ( .A(A[3000]), .B(n1096), .CI(
        C[3000]), .CO(C[3001]) );
  FA_5188 \FA_INST_0[5].FA_INST_1[441].FA_  ( .A(A[3001]), .B(n1095), .CI(
        C[3001]), .CO(C[3002]) );
  FA_5187 \FA_INST_0[5].FA_INST_1[442].FA_  ( .A(A[3002]), .B(n1094), .CI(
        C[3002]), .CO(C[3003]) );
  FA_5186 \FA_INST_0[5].FA_INST_1[443].FA_  ( .A(A[3003]), .B(n1093), .CI(
        C[3003]), .CO(C[3004]) );
  FA_5185 \FA_INST_0[5].FA_INST_1[444].FA_  ( .A(A[3004]), .B(n1092), .CI(
        C[3004]), .CO(C[3005]) );
  FA_5184 \FA_INST_0[5].FA_INST_1[445].FA_  ( .A(A[3005]), .B(n1091), .CI(
        C[3005]), .CO(C[3006]) );
  FA_5183 \FA_INST_0[5].FA_INST_1[446].FA_  ( .A(A[3006]), .B(n1090), .CI(
        C[3006]), .CO(C[3007]) );
  FA_5182 \FA_INST_0[5].FA_INST_1[447].FA_  ( .A(A[3007]), .B(n1089), .CI(
        C[3007]), .CO(C[3008]) );
  FA_5181 \FA_INST_0[5].FA_INST_1[448].FA_  ( .A(A[3008]), .B(n1088), .CI(
        C[3008]), .CO(C[3009]) );
  FA_5180 \FA_INST_0[5].FA_INST_1[449].FA_  ( .A(A[3009]), .B(n1087), .CI(
        C[3009]), .CO(C[3010]) );
  FA_5179 \FA_INST_0[5].FA_INST_1[450].FA_  ( .A(A[3010]), .B(n1086), .CI(
        C[3010]), .CO(C[3011]) );
  FA_5178 \FA_INST_0[5].FA_INST_1[451].FA_  ( .A(A[3011]), .B(n1085), .CI(
        C[3011]), .CO(C[3012]) );
  FA_5177 \FA_INST_0[5].FA_INST_1[452].FA_  ( .A(A[3012]), .B(n1084), .CI(
        C[3012]), .CO(C[3013]) );
  FA_5176 \FA_INST_0[5].FA_INST_1[453].FA_  ( .A(A[3013]), .B(n1083), .CI(
        C[3013]), .CO(C[3014]) );
  FA_5175 \FA_INST_0[5].FA_INST_1[454].FA_  ( .A(A[3014]), .B(n1082), .CI(
        C[3014]), .CO(C[3015]) );
  FA_5174 \FA_INST_0[5].FA_INST_1[455].FA_  ( .A(A[3015]), .B(n1081), .CI(
        C[3015]), .CO(C[3016]) );
  FA_5173 \FA_INST_0[5].FA_INST_1[456].FA_  ( .A(A[3016]), .B(n1080), .CI(
        C[3016]), .CO(C[3017]) );
  FA_5172 \FA_INST_0[5].FA_INST_1[457].FA_  ( .A(A[3017]), .B(n1079), .CI(
        C[3017]), .CO(C[3018]) );
  FA_5171 \FA_INST_0[5].FA_INST_1[458].FA_  ( .A(A[3018]), .B(n1078), .CI(
        C[3018]), .CO(C[3019]) );
  FA_5170 \FA_INST_0[5].FA_INST_1[459].FA_  ( .A(A[3019]), .B(n1077), .CI(
        C[3019]), .CO(C[3020]) );
  FA_5169 \FA_INST_0[5].FA_INST_1[460].FA_  ( .A(A[3020]), .B(n1076), .CI(
        C[3020]), .CO(C[3021]) );
  FA_5168 \FA_INST_0[5].FA_INST_1[461].FA_  ( .A(A[3021]), .B(n1075), .CI(
        C[3021]), .CO(C[3022]) );
  FA_5167 \FA_INST_0[5].FA_INST_1[462].FA_  ( .A(A[3022]), .B(n1074), .CI(
        C[3022]), .CO(C[3023]) );
  FA_5166 \FA_INST_0[5].FA_INST_1[463].FA_  ( .A(A[3023]), .B(n1073), .CI(
        C[3023]), .CO(C[3024]) );
  FA_5165 \FA_INST_0[5].FA_INST_1[464].FA_  ( .A(A[3024]), .B(n1072), .CI(
        C[3024]), .CO(C[3025]) );
  FA_5164 \FA_INST_0[5].FA_INST_1[465].FA_  ( .A(A[3025]), .B(n1071), .CI(
        C[3025]), .CO(C[3026]) );
  FA_5163 \FA_INST_0[5].FA_INST_1[466].FA_  ( .A(A[3026]), .B(n1070), .CI(
        C[3026]), .CO(C[3027]) );
  FA_5162 \FA_INST_0[5].FA_INST_1[467].FA_  ( .A(A[3027]), .B(n1069), .CI(
        C[3027]), .CO(C[3028]) );
  FA_5161 \FA_INST_0[5].FA_INST_1[468].FA_  ( .A(A[3028]), .B(n1068), .CI(
        C[3028]), .CO(C[3029]) );
  FA_5160 \FA_INST_0[5].FA_INST_1[469].FA_  ( .A(A[3029]), .B(n1067), .CI(
        C[3029]), .CO(C[3030]) );
  FA_5159 \FA_INST_0[5].FA_INST_1[470].FA_  ( .A(A[3030]), .B(n1066), .CI(
        C[3030]), .CO(C[3031]) );
  FA_5158 \FA_INST_0[5].FA_INST_1[471].FA_  ( .A(A[3031]), .B(n1065), .CI(
        C[3031]), .CO(C[3032]) );
  FA_5157 \FA_INST_0[5].FA_INST_1[472].FA_  ( .A(A[3032]), .B(n1064), .CI(
        C[3032]), .CO(C[3033]) );
  FA_5156 \FA_INST_0[5].FA_INST_1[473].FA_  ( .A(A[3033]), .B(n1063), .CI(
        C[3033]), .CO(C[3034]) );
  FA_5155 \FA_INST_0[5].FA_INST_1[474].FA_  ( .A(A[3034]), .B(n1062), .CI(
        C[3034]), .CO(C[3035]) );
  FA_5154 \FA_INST_0[5].FA_INST_1[475].FA_  ( .A(A[3035]), .B(n1061), .CI(
        C[3035]), .CO(C[3036]) );
  FA_5153 \FA_INST_0[5].FA_INST_1[476].FA_  ( .A(A[3036]), .B(n1060), .CI(
        C[3036]), .CO(C[3037]) );
  FA_5152 \FA_INST_0[5].FA_INST_1[477].FA_  ( .A(A[3037]), .B(n1059), .CI(
        C[3037]), .CO(C[3038]) );
  FA_5151 \FA_INST_0[5].FA_INST_1[478].FA_  ( .A(A[3038]), .B(n1058), .CI(
        C[3038]), .CO(C[3039]) );
  FA_5150 \FA_INST_0[5].FA_INST_1[479].FA_  ( .A(A[3039]), .B(n1057), .CI(
        C[3039]), .CO(C[3040]) );
  FA_5149 \FA_INST_0[5].FA_INST_1[480].FA_  ( .A(A[3040]), .B(n1056), .CI(
        C[3040]), .CO(C[3041]) );
  FA_5148 \FA_INST_0[5].FA_INST_1[481].FA_  ( .A(A[3041]), .B(n1055), .CI(
        C[3041]), .CO(C[3042]) );
  FA_5147 \FA_INST_0[5].FA_INST_1[482].FA_  ( .A(A[3042]), .B(n1054), .CI(
        C[3042]), .CO(C[3043]) );
  FA_5146 \FA_INST_0[5].FA_INST_1[483].FA_  ( .A(A[3043]), .B(n1053), .CI(
        C[3043]), .CO(C[3044]) );
  FA_5145 \FA_INST_0[5].FA_INST_1[484].FA_  ( .A(A[3044]), .B(n1052), .CI(
        C[3044]), .CO(C[3045]) );
  FA_5144 \FA_INST_0[5].FA_INST_1[485].FA_  ( .A(A[3045]), .B(n1051), .CI(
        C[3045]), .CO(C[3046]) );
  FA_5143 \FA_INST_0[5].FA_INST_1[486].FA_  ( .A(A[3046]), .B(n1050), .CI(
        C[3046]), .CO(C[3047]) );
  FA_5142 \FA_INST_0[5].FA_INST_1[487].FA_  ( .A(A[3047]), .B(n1049), .CI(
        C[3047]), .CO(C[3048]) );
  FA_5141 \FA_INST_0[5].FA_INST_1[488].FA_  ( .A(A[3048]), .B(n1048), .CI(
        C[3048]), .CO(C[3049]) );
  FA_5140 \FA_INST_0[5].FA_INST_1[489].FA_  ( .A(A[3049]), .B(n1047), .CI(
        C[3049]), .CO(C[3050]) );
  FA_5139 \FA_INST_0[5].FA_INST_1[490].FA_  ( .A(A[3050]), .B(n1046), .CI(
        C[3050]), .CO(C[3051]) );
  FA_5138 \FA_INST_0[5].FA_INST_1[491].FA_  ( .A(A[3051]), .B(n1045), .CI(
        C[3051]), .CO(C[3052]) );
  FA_5137 \FA_INST_0[5].FA_INST_1[492].FA_  ( .A(A[3052]), .B(n1044), .CI(
        C[3052]), .CO(C[3053]) );
  FA_5136 \FA_INST_0[5].FA_INST_1[493].FA_  ( .A(A[3053]), .B(n1043), .CI(
        C[3053]), .CO(C[3054]) );
  FA_5135 \FA_INST_0[5].FA_INST_1[494].FA_  ( .A(A[3054]), .B(n1042), .CI(
        C[3054]), .CO(C[3055]) );
  FA_5134 \FA_INST_0[5].FA_INST_1[495].FA_  ( .A(A[3055]), .B(n1041), .CI(
        C[3055]), .CO(C[3056]) );
  FA_5133 \FA_INST_0[5].FA_INST_1[496].FA_  ( .A(A[3056]), .B(n1040), .CI(
        C[3056]), .CO(C[3057]) );
  FA_5132 \FA_INST_0[5].FA_INST_1[497].FA_  ( .A(A[3057]), .B(n1039), .CI(
        C[3057]), .CO(C[3058]) );
  FA_5131 \FA_INST_0[5].FA_INST_1[498].FA_  ( .A(A[3058]), .B(n1038), .CI(
        C[3058]), .CO(C[3059]) );
  FA_5130 \FA_INST_0[5].FA_INST_1[499].FA_  ( .A(A[3059]), .B(n1037), .CI(
        C[3059]), .CO(C[3060]) );
  FA_5129 \FA_INST_0[5].FA_INST_1[500].FA_  ( .A(A[3060]), .B(n1036), .CI(
        C[3060]), .CO(C[3061]) );
  FA_5128 \FA_INST_0[5].FA_INST_1[501].FA_  ( .A(A[3061]), .B(n1035), .CI(
        C[3061]), .CO(C[3062]) );
  FA_5127 \FA_INST_0[5].FA_INST_1[502].FA_  ( .A(A[3062]), .B(n1034), .CI(
        C[3062]), .CO(C[3063]) );
  FA_5126 \FA_INST_0[5].FA_INST_1[503].FA_  ( .A(A[3063]), .B(n1033), .CI(
        C[3063]), .CO(C[3064]) );
  FA_5125 \FA_INST_0[5].FA_INST_1[504].FA_  ( .A(A[3064]), .B(n1032), .CI(
        C[3064]), .CO(C[3065]) );
  FA_5124 \FA_INST_0[5].FA_INST_1[505].FA_  ( .A(A[3065]), .B(n1031), .CI(
        C[3065]), .CO(C[3066]) );
  FA_5123 \FA_INST_0[5].FA_INST_1[506].FA_  ( .A(A[3066]), .B(n1030), .CI(
        C[3066]), .CO(C[3067]) );
  FA_5122 \FA_INST_0[5].FA_INST_1[507].FA_  ( .A(A[3067]), .B(n1029), .CI(
        C[3067]), .CO(C[3068]) );
  FA_5121 \FA_INST_0[5].FA_INST_1[508].FA_  ( .A(A[3068]), .B(n1028), .CI(
        C[3068]), .CO(C[3069]) );
  FA_5120 \FA_INST_0[5].FA_INST_1[509].FA_  ( .A(A[3069]), .B(n1027), .CI(
        C[3069]), .CO(C[3070]) );
  FA_5119 \FA_INST_0[5].FA_INST_1[510].FA_  ( .A(A[3070]), .B(n1026), .CI(
        C[3070]), .CO(C[3071]) );
  FA_5118 \FA_INST_0[5].FA_INST_1[511].FA_  ( .A(A[3071]), .B(n1025), .CI(
        C[3071]), .CO(C[3072]) );
  FA_5117 \FA_INST_0[6].FA_INST_1[0].FA_  ( .A(A[3072]), .B(n1024), .CI(
        C[3072]), .CO(C[3073]) );
  FA_5116 \FA_INST_0[6].FA_INST_1[1].FA_  ( .A(A[3073]), .B(n1023), .CI(
        C[3073]), .CO(C[3074]) );
  FA_5115 \FA_INST_0[6].FA_INST_1[2].FA_  ( .A(A[3074]), .B(n1022), .CI(
        C[3074]), .CO(C[3075]) );
  FA_5114 \FA_INST_0[6].FA_INST_1[3].FA_  ( .A(A[3075]), .B(n1021), .CI(
        C[3075]), .CO(C[3076]) );
  FA_5113 \FA_INST_0[6].FA_INST_1[4].FA_  ( .A(A[3076]), .B(n1020), .CI(
        C[3076]), .CO(C[3077]) );
  FA_5112 \FA_INST_0[6].FA_INST_1[5].FA_  ( .A(A[3077]), .B(n1019), .CI(
        C[3077]), .CO(C[3078]) );
  FA_5111 \FA_INST_0[6].FA_INST_1[6].FA_  ( .A(A[3078]), .B(n1018), .CI(
        C[3078]), .CO(C[3079]) );
  FA_5110 \FA_INST_0[6].FA_INST_1[7].FA_  ( .A(A[3079]), .B(n1017), .CI(
        C[3079]), .CO(C[3080]) );
  FA_5109 \FA_INST_0[6].FA_INST_1[8].FA_  ( .A(A[3080]), .B(n1016), .CI(
        C[3080]), .CO(C[3081]) );
  FA_5108 \FA_INST_0[6].FA_INST_1[9].FA_  ( .A(A[3081]), .B(n1015), .CI(
        C[3081]), .CO(C[3082]) );
  FA_5107 \FA_INST_0[6].FA_INST_1[10].FA_  ( .A(A[3082]), .B(n1014), .CI(
        C[3082]), .CO(C[3083]) );
  FA_5106 \FA_INST_0[6].FA_INST_1[11].FA_  ( .A(A[3083]), .B(n1013), .CI(
        C[3083]), .CO(C[3084]) );
  FA_5105 \FA_INST_0[6].FA_INST_1[12].FA_  ( .A(A[3084]), .B(n1012), .CI(
        C[3084]), .CO(C[3085]) );
  FA_5104 \FA_INST_0[6].FA_INST_1[13].FA_  ( .A(A[3085]), .B(n1011), .CI(
        C[3085]), .CO(C[3086]) );
  FA_5103 \FA_INST_0[6].FA_INST_1[14].FA_  ( .A(A[3086]), .B(n1010), .CI(
        C[3086]), .CO(C[3087]) );
  FA_5102 \FA_INST_0[6].FA_INST_1[15].FA_  ( .A(A[3087]), .B(n1009), .CI(
        C[3087]), .CO(C[3088]) );
  FA_5101 \FA_INST_0[6].FA_INST_1[16].FA_  ( .A(A[3088]), .B(n1008), .CI(
        C[3088]), .CO(C[3089]) );
  FA_5100 \FA_INST_0[6].FA_INST_1[17].FA_  ( .A(A[3089]), .B(n1007), .CI(
        C[3089]), .CO(C[3090]) );
  FA_5099 \FA_INST_0[6].FA_INST_1[18].FA_  ( .A(A[3090]), .B(n1006), .CI(
        C[3090]), .CO(C[3091]) );
  FA_5098 \FA_INST_0[6].FA_INST_1[19].FA_  ( .A(A[3091]), .B(n1005), .CI(
        C[3091]), .CO(C[3092]) );
  FA_5097 \FA_INST_0[6].FA_INST_1[20].FA_  ( .A(A[3092]), .B(n1004), .CI(
        C[3092]), .CO(C[3093]) );
  FA_5096 \FA_INST_0[6].FA_INST_1[21].FA_  ( .A(A[3093]), .B(n1003), .CI(
        C[3093]), .CO(C[3094]) );
  FA_5095 \FA_INST_0[6].FA_INST_1[22].FA_  ( .A(A[3094]), .B(n1002), .CI(
        C[3094]), .CO(C[3095]) );
  FA_5094 \FA_INST_0[6].FA_INST_1[23].FA_  ( .A(A[3095]), .B(n1001), .CI(
        C[3095]), .CO(C[3096]) );
  FA_5093 \FA_INST_0[6].FA_INST_1[24].FA_  ( .A(A[3096]), .B(n1000), .CI(
        C[3096]), .CO(C[3097]) );
  FA_5092 \FA_INST_0[6].FA_INST_1[25].FA_  ( .A(A[3097]), .B(n999), .CI(
        C[3097]), .CO(C[3098]) );
  FA_5091 \FA_INST_0[6].FA_INST_1[26].FA_  ( .A(A[3098]), .B(n998), .CI(
        C[3098]), .CO(C[3099]) );
  FA_5090 \FA_INST_0[6].FA_INST_1[27].FA_  ( .A(A[3099]), .B(n997), .CI(
        C[3099]), .CO(C[3100]) );
  FA_5089 \FA_INST_0[6].FA_INST_1[28].FA_  ( .A(A[3100]), .B(n996), .CI(
        C[3100]), .CO(C[3101]) );
  FA_5088 \FA_INST_0[6].FA_INST_1[29].FA_  ( .A(A[3101]), .B(n995), .CI(
        C[3101]), .CO(C[3102]) );
  FA_5087 \FA_INST_0[6].FA_INST_1[30].FA_  ( .A(A[3102]), .B(n994), .CI(
        C[3102]), .CO(C[3103]) );
  FA_5086 \FA_INST_0[6].FA_INST_1[31].FA_  ( .A(A[3103]), .B(n993), .CI(
        C[3103]), .CO(C[3104]) );
  FA_5085 \FA_INST_0[6].FA_INST_1[32].FA_  ( .A(A[3104]), .B(n992), .CI(
        C[3104]), .CO(C[3105]) );
  FA_5084 \FA_INST_0[6].FA_INST_1[33].FA_  ( .A(A[3105]), .B(n991), .CI(
        C[3105]), .CO(C[3106]) );
  FA_5083 \FA_INST_0[6].FA_INST_1[34].FA_  ( .A(A[3106]), .B(n990), .CI(
        C[3106]), .CO(C[3107]) );
  FA_5082 \FA_INST_0[6].FA_INST_1[35].FA_  ( .A(A[3107]), .B(n989), .CI(
        C[3107]), .CO(C[3108]) );
  FA_5081 \FA_INST_0[6].FA_INST_1[36].FA_  ( .A(A[3108]), .B(n988), .CI(
        C[3108]), .CO(C[3109]) );
  FA_5080 \FA_INST_0[6].FA_INST_1[37].FA_  ( .A(A[3109]), .B(n987), .CI(
        C[3109]), .CO(C[3110]) );
  FA_5079 \FA_INST_0[6].FA_INST_1[38].FA_  ( .A(A[3110]), .B(n986), .CI(
        C[3110]), .CO(C[3111]) );
  FA_5078 \FA_INST_0[6].FA_INST_1[39].FA_  ( .A(A[3111]), .B(n985), .CI(
        C[3111]), .CO(C[3112]) );
  FA_5077 \FA_INST_0[6].FA_INST_1[40].FA_  ( .A(A[3112]), .B(n984), .CI(
        C[3112]), .CO(C[3113]) );
  FA_5076 \FA_INST_0[6].FA_INST_1[41].FA_  ( .A(A[3113]), .B(n983), .CI(
        C[3113]), .CO(C[3114]) );
  FA_5075 \FA_INST_0[6].FA_INST_1[42].FA_  ( .A(A[3114]), .B(n982), .CI(
        C[3114]), .CO(C[3115]) );
  FA_5074 \FA_INST_0[6].FA_INST_1[43].FA_  ( .A(A[3115]), .B(n981), .CI(
        C[3115]), .CO(C[3116]) );
  FA_5073 \FA_INST_0[6].FA_INST_1[44].FA_  ( .A(A[3116]), .B(n980), .CI(
        C[3116]), .CO(C[3117]) );
  FA_5072 \FA_INST_0[6].FA_INST_1[45].FA_  ( .A(A[3117]), .B(n979), .CI(
        C[3117]), .CO(C[3118]) );
  FA_5071 \FA_INST_0[6].FA_INST_1[46].FA_  ( .A(A[3118]), .B(n978), .CI(
        C[3118]), .CO(C[3119]) );
  FA_5070 \FA_INST_0[6].FA_INST_1[47].FA_  ( .A(A[3119]), .B(n977), .CI(
        C[3119]), .CO(C[3120]) );
  FA_5069 \FA_INST_0[6].FA_INST_1[48].FA_  ( .A(A[3120]), .B(n976), .CI(
        C[3120]), .CO(C[3121]) );
  FA_5068 \FA_INST_0[6].FA_INST_1[49].FA_  ( .A(A[3121]), .B(n975), .CI(
        C[3121]), .CO(C[3122]) );
  FA_5067 \FA_INST_0[6].FA_INST_1[50].FA_  ( .A(A[3122]), .B(n974), .CI(
        C[3122]), .CO(C[3123]) );
  FA_5066 \FA_INST_0[6].FA_INST_1[51].FA_  ( .A(A[3123]), .B(n973), .CI(
        C[3123]), .CO(C[3124]) );
  FA_5065 \FA_INST_0[6].FA_INST_1[52].FA_  ( .A(A[3124]), .B(n972), .CI(
        C[3124]), .CO(C[3125]) );
  FA_5064 \FA_INST_0[6].FA_INST_1[53].FA_  ( .A(A[3125]), .B(n971), .CI(
        C[3125]), .CO(C[3126]) );
  FA_5063 \FA_INST_0[6].FA_INST_1[54].FA_  ( .A(A[3126]), .B(n970), .CI(
        C[3126]), .CO(C[3127]) );
  FA_5062 \FA_INST_0[6].FA_INST_1[55].FA_  ( .A(A[3127]), .B(n969), .CI(
        C[3127]), .CO(C[3128]) );
  FA_5061 \FA_INST_0[6].FA_INST_1[56].FA_  ( .A(A[3128]), .B(n968), .CI(
        C[3128]), .CO(C[3129]) );
  FA_5060 \FA_INST_0[6].FA_INST_1[57].FA_  ( .A(A[3129]), .B(n967), .CI(
        C[3129]), .CO(C[3130]) );
  FA_5059 \FA_INST_0[6].FA_INST_1[58].FA_  ( .A(A[3130]), .B(n966), .CI(
        C[3130]), .CO(C[3131]) );
  FA_5058 \FA_INST_0[6].FA_INST_1[59].FA_  ( .A(A[3131]), .B(n965), .CI(
        C[3131]), .CO(C[3132]) );
  FA_5057 \FA_INST_0[6].FA_INST_1[60].FA_  ( .A(A[3132]), .B(n964), .CI(
        C[3132]), .CO(C[3133]) );
  FA_5056 \FA_INST_0[6].FA_INST_1[61].FA_  ( .A(A[3133]), .B(n963), .CI(
        C[3133]), .CO(C[3134]) );
  FA_5055 \FA_INST_0[6].FA_INST_1[62].FA_  ( .A(A[3134]), .B(n962), .CI(
        C[3134]), .CO(C[3135]) );
  FA_5054 \FA_INST_0[6].FA_INST_1[63].FA_  ( .A(A[3135]), .B(n961), .CI(
        C[3135]), .CO(C[3136]) );
  FA_5053 \FA_INST_0[6].FA_INST_1[64].FA_  ( .A(A[3136]), .B(n960), .CI(
        C[3136]), .CO(C[3137]) );
  FA_5052 \FA_INST_0[6].FA_INST_1[65].FA_  ( .A(A[3137]), .B(n959), .CI(
        C[3137]), .CO(C[3138]) );
  FA_5051 \FA_INST_0[6].FA_INST_1[66].FA_  ( .A(A[3138]), .B(n958), .CI(
        C[3138]), .CO(C[3139]) );
  FA_5050 \FA_INST_0[6].FA_INST_1[67].FA_  ( .A(A[3139]), .B(n957), .CI(
        C[3139]), .CO(C[3140]) );
  FA_5049 \FA_INST_0[6].FA_INST_1[68].FA_  ( .A(A[3140]), .B(n956), .CI(
        C[3140]), .CO(C[3141]) );
  FA_5048 \FA_INST_0[6].FA_INST_1[69].FA_  ( .A(A[3141]), .B(n955), .CI(
        C[3141]), .CO(C[3142]) );
  FA_5047 \FA_INST_0[6].FA_INST_1[70].FA_  ( .A(A[3142]), .B(n954), .CI(
        C[3142]), .CO(C[3143]) );
  FA_5046 \FA_INST_0[6].FA_INST_1[71].FA_  ( .A(A[3143]), .B(n953), .CI(
        C[3143]), .CO(C[3144]) );
  FA_5045 \FA_INST_0[6].FA_INST_1[72].FA_  ( .A(A[3144]), .B(n952), .CI(
        C[3144]), .CO(C[3145]) );
  FA_5044 \FA_INST_0[6].FA_INST_1[73].FA_  ( .A(A[3145]), .B(n951), .CI(
        C[3145]), .CO(C[3146]) );
  FA_5043 \FA_INST_0[6].FA_INST_1[74].FA_  ( .A(A[3146]), .B(n950), .CI(
        C[3146]), .CO(C[3147]) );
  FA_5042 \FA_INST_0[6].FA_INST_1[75].FA_  ( .A(A[3147]), .B(n949), .CI(
        C[3147]), .CO(C[3148]) );
  FA_5041 \FA_INST_0[6].FA_INST_1[76].FA_  ( .A(A[3148]), .B(n948), .CI(
        C[3148]), .CO(C[3149]) );
  FA_5040 \FA_INST_0[6].FA_INST_1[77].FA_  ( .A(A[3149]), .B(n947), .CI(
        C[3149]), .CO(C[3150]) );
  FA_5039 \FA_INST_0[6].FA_INST_1[78].FA_  ( .A(A[3150]), .B(n946), .CI(
        C[3150]), .CO(C[3151]) );
  FA_5038 \FA_INST_0[6].FA_INST_1[79].FA_  ( .A(A[3151]), .B(n945), .CI(
        C[3151]), .CO(C[3152]) );
  FA_5037 \FA_INST_0[6].FA_INST_1[80].FA_  ( .A(A[3152]), .B(n944), .CI(
        C[3152]), .CO(C[3153]) );
  FA_5036 \FA_INST_0[6].FA_INST_1[81].FA_  ( .A(A[3153]), .B(n943), .CI(
        C[3153]), .CO(C[3154]) );
  FA_5035 \FA_INST_0[6].FA_INST_1[82].FA_  ( .A(A[3154]), .B(n942), .CI(
        C[3154]), .CO(C[3155]) );
  FA_5034 \FA_INST_0[6].FA_INST_1[83].FA_  ( .A(A[3155]), .B(n941), .CI(
        C[3155]), .CO(C[3156]) );
  FA_5033 \FA_INST_0[6].FA_INST_1[84].FA_  ( .A(A[3156]), .B(n940), .CI(
        C[3156]), .CO(C[3157]) );
  FA_5032 \FA_INST_0[6].FA_INST_1[85].FA_  ( .A(A[3157]), .B(n939), .CI(
        C[3157]), .CO(C[3158]) );
  FA_5031 \FA_INST_0[6].FA_INST_1[86].FA_  ( .A(A[3158]), .B(n938), .CI(
        C[3158]), .CO(C[3159]) );
  FA_5030 \FA_INST_0[6].FA_INST_1[87].FA_  ( .A(A[3159]), .B(n937), .CI(
        C[3159]), .CO(C[3160]) );
  FA_5029 \FA_INST_0[6].FA_INST_1[88].FA_  ( .A(A[3160]), .B(n936), .CI(
        C[3160]), .CO(C[3161]) );
  FA_5028 \FA_INST_0[6].FA_INST_1[89].FA_  ( .A(A[3161]), .B(n935), .CI(
        C[3161]), .CO(C[3162]) );
  FA_5027 \FA_INST_0[6].FA_INST_1[90].FA_  ( .A(A[3162]), .B(n934), .CI(
        C[3162]), .CO(C[3163]) );
  FA_5026 \FA_INST_0[6].FA_INST_1[91].FA_  ( .A(A[3163]), .B(n933), .CI(
        C[3163]), .CO(C[3164]) );
  FA_5025 \FA_INST_0[6].FA_INST_1[92].FA_  ( .A(A[3164]), .B(n932), .CI(
        C[3164]), .CO(C[3165]) );
  FA_5024 \FA_INST_0[6].FA_INST_1[93].FA_  ( .A(A[3165]), .B(n931), .CI(
        C[3165]), .CO(C[3166]) );
  FA_5023 \FA_INST_0[6].FA_INST_1[94].FA_  ( .A(A[3166]), .B(n930), .CI(
        C[3166]), .CO(C[3167]) );
  FA_5022 \FA_INST_0[6].FA_INST_1[95].FA_  ( .A(A[3167]), .B(n929), .CI(
        C[3167]), .CO(C[3168]) );
  FA_5021 \FA_INST_0[6].FA_INST_1[96].FA_  ( .A(A[3168]), .B(n928), .CI(
        C[3168]), .CO(C[3169]) );
  FA_5020 \FA_INST_0[6].FA_INST_1[97].FA_  ( .A(A[3169]), .B(n927), .CI(
        C[3169]), .CO(C[3170]) );
  FA_5019 \FA_INST_0[6].FA_INST_1[98].FA_  ( .A(A[3170]), .B(n926), .CI(
        C[3170]), .CO(C[3171]) );
  FA_5018 \FA_INST_0[6].FA_INST_1[99].FA_  ( .A(A[3171]), .B(n925), .CI(
        C[3171]), .CO(C[3172]) );
  FA_5017 \FA_INST_0[6].FA_INST_1[100].FA_  ( .A(A[3172]), .B(n924), .CI(
        C[3172]), .CO(C[3173]) );
  FA_5016 \FA_INST_0[6].FA_INST_1[101].FA_  ( .A(A[3173]), .B(n923), .CI(
        C[3173]), .CO(C[3174]) );
  FA_5015 \FA_INST_0[6].FA_INST_1[102].FA_  ( .A(A[3174]), .B(n922), .CI(
        C[3174]), .CO(C[3175]) );
  FA_5014 \FA_INST_0[6].FA_INST_1[103].FA_  ( .A(A[3175]), .B(n921), .CI(
        C[3175]), .CO(C[3176]) );
  FA_5013 \FA_INST_0[6].FA_INST_1[104].FA_  ( .A(A[3176]), .B(n920), .CI(
        C[3176]), .CO(C[3177]) );
  FA_5012 \FA_INST_0[6].FA_INST_1[105].FA_  ( .A(A[3177]), .B(n919), .CI(
        C[3177]), .CO(C[3178]) );
  FA_5011 \FA_INST_0[6].FA_INST_1[106].FA_  ( .A(A[3178]), .B(n918), .CI(
        C[3178]), .CO(C[3179]) );
  FA_5010 \FA_INST_0[6].FA_INST_1[107].FA_  ( .A(A[3179]), .B(n917), .CI(
        C[3179]), .CO(C[3180]) );
  FA_5009 \FA_INST_0[6].FA_INST_1[108].FA_  ( .A(A[3180]), .B(n916), .CI(
        C[3180]), .CO(C[3181]) );
  FA_5008 \FA_INST_0[6].FA_INST_1[109].FA_  ( .A(A[3181]), .B(n915), .CI(
        C[3181]), .CO(C[3182]) );
  FA_5007 \FA_INST_0[6].FA_INST_1[110].FA_  ( .A(A[3182]), .B(n914), .CI(
        C[3182]), .CO(C[3183]) );
  FA_5006 \FA_INST_0[6].FA_INST_1[111].FA_  ( .A(A[3183]), .B(n913), .CI(
        C[3183]), .CO(C[3184]) );
  FA_5005 \FA_INST_0[6].FA_INST_1[112].FA_  ( .A(A[3184]), .B(n912), .CI(
        C[3184]), .CO(C[3185]) );
  FA_5004 \FA_INST_0[6].FA_INST_1[113].FA_  ( .A(A[3185]), .B(n911), .CI(
        C[3185]), .CO(C[3186]) );
  FA_5003 \FA_INST_0[6].FA_INST_1[114].FA_  ( .A(A[3186]), .B(n910), .CI(
        C[3186]), .CO(C[3187]) );
  FA_5002 \FA_INST_0[6].FA_INST_1[115].FA_  ( .A(A[3187]), .B(n909), .CI(
        C[3187]), .CO(C[3188]) );
  FA_5001 \FA_INST_0[6].FA_INST_1[116].FA_  ( .A(A[3188]), .B(n908), .CI(
        C[3188]), .CO(C[3189]) );
  FA_5000 \FA_INST_0[6].FA_INST_1[117].FA_  ( .A(A[3189]), .B(n907), .CI(
        C[3189]), .CO(C[3190]) );
  FA_4999 \FA_INST_0[6].FA_INST_1[118].FA_  ( .A(A[3190]), .B(n906), .CI(
        C[3190]), .CO(C[3191]) );
  FA_4998 \FA_INST_0[6].FA_INST_1[119].FA_  ( .A(A[3191]), .B(n905), .CI(
        C[3191]), .CO(C[3192]) );
  FA_4997 \FA_INST_0[6].FA_INST_1[120].FA_  ( .A(A[3192]), .B(n904), .CI(
        C[3192]), .CO(C[3193]) );
  FA_4996 \FA_INST_0[6].FA_INST_1[121].FA_  ( .A(A[3193]), .B(n903), .CI(
        C[3193]), .CO(C[3194]) );
  FA_4995 \FA_INST_0[6].FA_INST_1[122].FA_  ( .A(A[3194]), .B(n902), .CI(
        C[3194]), .CO(C[3195]) );
  FA_4994 \FA_INST_0[6].FA_INST_1[123].FA_  ( .A(A[3195]), .B(n901), .CI(
        C[3195]), .CO(C[3196]) );
  FA_4993 \FA_INST_0[6].FA_INST_1[124].FA_  ( .A(A[3196]), .B(n900), .CI(
        C[3196]), .CO(C[3197]) );
  FA_4992 \FA_INST_0[6].FA_INST_1[125].FA_  ( .A(A[3197]), .B(n899), .CI(
        C[3197]), .CO(C[3198]) );
  FA_4991 \FA_INST_0[6].FA_INST_1[126].FA_  ( .A(A[3198]), .B(n898), .CI(
        C[3198]), .CO(C[3199]) );
  FA_4990 \FA_INST_0[6].FA_INST_1[127].FA_  ( .A(A[3199]), .B(n897), .CI(
        C[3199]), .CO(C[3200]) );
  FA_4989 \FA_INST_0[6].FA_INST_1[128].FA_  ( .A(A[3200]), .B(n896), .CI(
        C[3200]), .CO(C[3201]) );
  FA_4988 \FA_INST_0[6].FA_INST_1[129].FA_  ( .A(A[3201]), .B(n895), .CI(
        C[3201]), .CO(C[3202]) );
  FA_4987 \FA_INST_0[6].FA_INST_1[130].FA_  ( .A(A[3202]), .B(n894), .CI(
        C[3202]), .CO(C[3203]) );
  FA_4986 \FA_INST_0[6].FA_INST_1[131].FA_  ( .A(A[3203]), .B(n893), .CI(
        C[3203]), .CO(C[3204]) );
  FA_4985 \FA_INST_0[6].FA_INST_1[132].FA_  ( .A(A[3204]), .B(n892), .CI(
        C[3204]), .CO(C[3205]) );
  FA_4984 \FA_INST_0[6].FA_INST_1[133].FA_  ( .A(A[3205]), .B(n891), .CI(
        C[3205]), .CO(C[3206]) );
  FA_4983 \FA_INST_0[6].FA_INST_1[134].FA_  ( .A(A[3206]), .B(n890), .CI(
        C[3206]), .CO(C[3207]) );
  FA_4982 \FA_INST_0[6].FA_INST_1[135].FA_  ( .A(A[3207]), .B(n889), .CI(
        C[3207]), .CO(C[3208]) );
  FA_4981 \FA_INST_0[6].FA_INST_1[136].FA_  ( .A(A[3208]), .B(n888), .CI(
        C[3208]), .CO(C[3209]) );
  FA_4980 \FA_INST_0[6].FA_INST_1[137].FA_  ( .A(A[3209]), .B(n887), .CI(
        C[3209]), .CO(C[3210]) );
  FA_4979 \FA_INST_0[6].FA_INST_1[138].FA_  ( .A(A[3210]), .B(n886), .CI(
        C[3210]), .CO(C[3211]) );
  FA_4978 \FA_INST_0[6].FA_INST_1[139].FA_  ( .A(A[3211]), .B(n885), .CI(
        C[3211]), .CO(C[3212]) );
  FA_4977 \FA_INST_0[6].FA_INST_1[140].FA_  ( .A(A[3212]), .B(n884), .CI(
        C[3212]), .CO(C[3213]) );
  FA_4976 \FA_INST_0[6].FA_INST_1[141].FA_  ( .A(A[3213]), .B(n883), .CI(
        C[3213]), .CO(C[3214]) );
  FA_4975 \FA_INST_0[6].FA_INST_1[142].FA_  ( .A(A[3214]), .B(n882), .CI(
        C[3214]), .CO(C[3215]) );
  FA_4974 \FA_INST_0[6].FA_INST_1[143].FA_  ( .A(A[3215]), .B(n881), .CI(
        C[3215]), .CO(C[3216]) );
  FA_4973 \FA_INST_0[6].FA_INST_1[144].FA_  ( .A(A[3216]), .B(n880), .CI(
        C[3216]), .CO(C[3217]) );
  FA_4972 \FA_INST_0[6].FA_INST_1[145].FA_  ( .A(A[3217]), .B(n879), .CI(
        C[3217]), .CO(C[3218]) );
  FA_4971 \FA_INST_0[6].FA_INST_1[146].FA_  ( .A(A[3218]), .B(n878), .CI(
        C[3218]), .CO(C[3219]) );
  FA_4970 \FA_INST_0[6].FA_INST_1[147].FA_  ( .A(A[3219]), .B(n877), .CI(
        C[3219]), .CO(C[3220]) );
  FA_4969 \FA_INST_0[6].FA_INST_1[148].FA_  ( .A(A[3220]), .B(n876), .CI(
        C[3220]), .CO(C[3221]) );
  FA_4968 \FA_INST_0[6].FA_INST_1[149].FA_  ( .A(A[3221]), .B(n875), .CI(
        C[3221]), .CO(C[3222]) );
  FA_4967 \FA_INST_0[6].FA_INST_1[150].FA_  ( .A(A[3222]), .B(n874), .CI(
        C[3222]), .CO(C[3223]) );
  FA_4966 \FA_INST_0[6].FA_INST_1[151].FA_  ( .A(A[3223]), .B(n873), .CI(
        C[3223]), .CO(C[3224]) );
  FA_4965 \FA_INST_0[6].FA_INST_1[152].FA_  ( .A(A[3224]), .B(n872), .CI(
        C[3224]), .CO(C[3225]) );
  FA_4964 \FA_INST_0[6].FA_INST_1[153].FA_  ( .A(A[3225]), .B(n871), .CI(
        C[3225]), .CO(C[3226]) );
  FA_4963 \FA_INST_0[6].FA_INST_1[154].FA_  ( .A(A[3226]), .B(n870), .CI(
        C[3226]), .CO(C[3227]) );
  FA_4962 \FA_INST_0[6].FA_INST_1[155].FA_  ( .A(A[3227]), .B(n869), .CI(
        C[3227]), .CO(C[3228]) );
  FA_4961 \FA_INST_0[6].FA_INST_1[156].FA_  ( .A(A[3228]), .B(n868), .CI(
        C[3228]), .CO(C[3229]) );
  FA_4960 \FA_INST_0[6].FA_INST_1[157].FA_  ( .A(A[3229]), .B(n867), .CI(
        C[3229]), .CO(C[3230]) );
  FA_4959 \FA_INST_0[6].FA_INST_1[158].FA_  ( .A(A[3230]), .B(n866), .CI(
        C[3230]), .CO(C[3231]) );
  FA_4958 \FA_INST_0[6].FA_INST_1[159].FA_  ( .A(A[3231]), .B(n865), .CI(
        C[3231]), .CO(C[3232]) );
  FA_4957 \FA_INST_0[6].FA_INST_1[160].FA_  ( .A(A[3232]), .B(n864), .CI(
        C[3232]), .CO(C[3233]) );
  FA_4956 \FA_INST_0[6].FA_INST_1[161].FA_  ( .A(A[3233]), .B(n863), .CI(
        C[3233]), .CO(C[3234]) );
  FA_4955 \FA_INST_0[6].FA_INST_1[162].FA_  ( .A(A[3234]), .B(n862), .CI(
        C[3234]), .CO(C[3235]) );
  FA_4954 \FA_INST_0[6].FA_INST_1[163].FA_  ( .A(A[3235]), .B(n861), .CI(
        C[3235]), .CO(C[3236]) );
  FA_4953 \FA_INST_0[6].FA_INST_1[164].FA_  ( .A(A[3236]), .B(n860), .CI(
        C[3236]), .CO(C[3237]) );
  FA_4952 \FA_INST_0[6].FA_INST_1[165].FA_  ( .A(A[3237]), .B(n859), .CI(
        C[3237]), .CO(C[3238]) );
  FA_4951 \FA_INST_0[6].FA_INST_1[166].FA_  ( .A(A[3238]), .B(n858), .CI(
        C[3238]), .CO(C[3239]) );
  FA_4950 \FA_INST_0[6].FA_INST_1[167].FA_  ( .A(A[3239]), .B(n857), .CI(
        C[3239]), .CO(C[3240]) );
  FA_4949 \FA_INST_0[6].FA_INST_1[168].FA_  ( .A(A[3240]), .B(n856), .CI(
        C[3240]), .CO(C[3241]) );
  FA_4948 \FA_INST_0[6].FA_INST_1[169].FA_  ( .A(A[3241]), .B(n855), .CI(
        C[3241]), .CO(C[3242]) );
  FA_4947 \FA_INST_0[6].FA_INST_1[170].FA_  ( .A(A[3242]), .B(n854), .CI(
        C[3242]), .CO(C[3243]) );
  FA_4946 \FA_INST_0[6].FA_INST_1[171].FA_  ( .A(A[3243]), .B(n853), .CI(
        C[3243]), .CO(C[3244]) );
  FA_4945 \FA_INST_0[6].FA_INST_1[172].FA_  ( .A(A[3244]), .B(n852), .CI(
        C[3244]), .CO(C[3245]) );
  FA_4944 \FA_INST_0[6].FA_INST_1[173].FA_  ( .A(A[3245]), .B(n851), .CI(
        C[3245]), .CO(C[3246]) );
  FA_4943 \FA_INST_0[6].FA_INST_1[174].FA_  ( .A(A[3246]), .B(n850), .CI(
        C[3246]), .CO(C[3247]) );
  FA_4942 \FA_INST_0[6].FA_INST_1[175].FA_  ( .A(A[3247]), .B(n849), .CI(
        C[3247]), .CO(C[3248]) );
  FA_4941 \FA_INST_0[6].FA_INST_1[176].FA_  ( .A(A[3248]), .B(n848), .CI(
        C[3248]), .CO(C[3249]) );
  FA_4940 \FA_INST_0[6].FA_INST_1[177].FA_  ( .A(A[3249]), .B(n847), .CI(
        C[3249]), .CO(C[3250]) );
  FA_4939 \FA_INST_0[6].FA_INST_1[178].FA_  ( .A(A[3250]), .B(n846), .CI(
        C[3250]), .CO(C[3251]) );
  FA_4938 \FA_INST_0[6].FA_INST_1[179].FA_  ( .A(A[3251]), .B(n845), .CI(
        C[3251]), .CO(C[3252]) );
  FA_4937 \FA_INST_0[6].FA_INST_1[180].FA_  ( .A(A[3252]), .B(n844), .CI(
        C[3252]), .CO(C[3253]) );
  FA_4936 \FA_INST_0[6].FA_INST_1[181].FA_  ( .A(A[3253]), .B(n843), .CI(
        C[3253]), .CO(C[3254]) );
  FA_4935 \FA_INST_0[6].FA_INST_1[182].FA_  ( .A(A[3254]), .B(n842), .CI(
        C[3254]), .CO(C[3255]) );
  FA_4934 \FA_INST_0[6].FA_INST_1[183].FA_  ( .A(A[3255]), .B(n841), .CI(
        C[3255]), .CO(C[3256]) );
  FA_4933 \FA_INST_0[6].FA_INST_1[184].FA_  ( .A(A[3256]), .B(n840), .CI(
        C[3256]), .CO(C[3257]) );
  FA_4932 \FA_INST_0[6].FA_INST_1[185].FA_  ( .A(A[3257]), .B(n839), .CI(
        C[3257]), .CO(C[3258]) );
  FA_4931 \FA_INST_0[6].FA_INST_1[186].FA_  ( .A(A[3258]), .B(n838), .CI(
        C[3258]), .CO(C[3259]) );
  FA_4930 \FA_INST_0[6].FA_INST_1[187].FA_  ( .A(A[3259]), .B(n837), .CI(
        C[3259]), .CO(C[3260]) );
  FA_4929 \FA_INST_0[6].FA_INST_1[188].FA_  ( .A(A[3260]), .B(n836), .CI(
        C[3260]), .CO(C[3261]) );
  FA_4928 \FA_INST_0[6].FA_INST_1[189].FA_  ( .A(A[3261]), .B(n835), .CI(
        C[3261]), .CO(C[3262]) );
  FA_4927 \FA_INST_0[6].FA_INST_1[190].FA_  ( .A(A[3262]), .B(n834), .CI(
        C[3262]), .CO(C[3263]) );
  FA_4926 \FA_INST_0[6].FA_INST_1[191].FA_  ( .A(A[3263]), .B(n833), .CI(
        C[3263]), .CO(C[3264]) );
  FA_4925 \FA_INST_0[6].FA_INST_1[192].FA_  ( .A(A[3264]), .B(n832), .CI(
        C[3264]), .CO(C[3265]) );
  FA_4924 \FA_INST_0[6].FA_INST_1[193].FA_  ( .A(A[3265]), .B(n831), .CI(
        C[3265]), .CO(C[3266]) );
  FA_4923 \FA_INST_0[6].FA_INST_1[194].FA_  ( .A(A[3266]), .B(n830), .CI(
        C[3266]), .CO(C[3267]) );
  FA_4922 \FA_INST_0[6].FA_INST_1[195].FA_  ( .A(A[3267]), .B(n829), .CI(
        C[3267]), .CO(C[3268]) );
  FA_4921 \FA_INST_0[6].FA_INST_1[196].FA_  ( .A(A[3268]), .B(n828), .CI(
        C[3268]), .CO(C[3269]) );
  FA_4920 \FA_INST_0[6].FA_INST_1[197].FA_  ( .A(A[3269]), .B(n827), .CI(
        C[3269]), .CO(C[3270]) );
  FA_4919 \FA_INST_0[6].FA_INST_1[198].FA_  ( .A(A[3270]), .B(n826), .CI(
        C[3270]), .CO(C[3271]) );
  FA_4918 \FA_INST_0[6].FA_INST_1[199].FA_  ( .A(A[3271]), .B(n825), .CI(
        C[3271]), .CO(C[3272]) );
  FA_4917 \FA_INST_0[6].FA_INST_1[200].FA_  ( .A(A[3272]), .B(n824), .CI(
        C[3272]), .CO(C[3273]) );
  FA_4916 \FA_INST_0[6].FA_INST_1[201].FA_  ( .A(A[3273]), .B(n823), .CI(
        C[3273]), .CO(C[3274]) );
  FA_4915 \FA_INST_0[6].FA_INST_1[202].FA_  ( .A(A[3274]), .B(n822), .CI(
        C[3274]), .CO(C[3275]) );
  FA_4914 \FA_INST_0[6].FA_INST_1[203].FA_  ( .A(A[3275]), .B(n821), .CI(
        C[3275]), .CO(C[3276]) );
  FA_4913 \FA_INST_0[6].FA_INST_1[204].FA_  ( .A(A[3276]), .B(n820), .CI(
        C[3276]), .CO(C[3277]) );
  FA_4912 \FA_INST_0[6].FA_INST_1[205].FA_  ( .A(A[3277]), .B(n819), .CI(
        C[3277]), .CO(C[3278]) );
  FA_4911 \FA_INST_0[6].FA_INST_1[206].FA_  ( .A(A[3278]), .B(n818), .CI(
        C[3278]), .CO(C[3279]) );
  FA_4910 \FA_INST_0[6].FA_INST_1[207].FA_  ( .A(A[3279]), .B(n817), .CI(
        C[3279]), .CO(C[3280]) );
  FA_4909 \FA_INST_0[6].FA_INST_1[208].FA_  ( .A(A[3280]), .B(n816), .CI(
        C[3280]), .CO(C[3281]) );
  FA_4908 \FA_INST_0[6].FA_INST_1[209].FA_  ( .A(A[3281]), .B(n815), .CI(
        C[3281]), .CO(C[3282]) );
  FA_4907 \FA_INST_0[6].FA_INST_1[210].FA_  ( .A(A[3282]), .B(n814), .CI(
        C[3282]), .CO(C[3283]) );
  FA_4906 \FA_INST_0[6].FA_INST_1[211].FA_  ( .A(A[3283]), .B(n813), .CI(
        C[3283]), .CO(C[3284]) );
  FA_4905 \FA_INST_0[6].FA_INST_1[212].FA_  ( .A(A[3284]), .B(n812), .CI(
        C[3284]), .CO(C[3285]) );
  FA_4904 \FA_INST_0[6].FA_INST_1[213].FA_  ( .A(A[3285]), .B(n811), .CI(
        C[3285]), .CO(C[3286]) );
  FA_4903 \FA_INST_0[6].FA_INST_1[214].FA_  ( .A(A[3286]), .B(n810), .CI(
        C[3286]), .CO(C[3287]) );
  FA_4902 \FA_INST_0[6].FA_INST_1[215].FA_  ( .A(A[3287]), .B(n809), .CI(
        C[3287]), .CO(C[3288]) );
  FA_4901 \FA_INST_0[6].FA_INST_1[216].FA_  ( .A(A[3288]), .B(n808), .CI(
        C[3288]), .CO(C[3289]) );
  FA_4900 \FA_INST_0[6].FA_INST_1[217].FA_  ( .A(A[3289]), .B(n807), .CI(
        C[3289]), .CO(C[3290]) );
  FA_4899 \FA_INST_0[6].FA_INST_1[218].FA_  ( .A(A[3290]), .B(n806), .CI(
        C[3290]), .CO(C[3291]) );
  FA_4898 \FA_INST_0[6].FA_INST_1[219].FA_  ( .A(A[3291]), .B(n805), .CI(
        C[3291]), .CO(C[3292]) );
  FA_4897 \FA_INST_0[6].FA_INST_1[220].FA_  ( .A(A[3292]), .B(n804), .CI(
        C[3292]), .CO(C[3293]) );
  FA_4896 \FA_INST_0[6].FA_INST_1[221].FA_  ( .A(A[3293]), .B(n803), .CI(
        C[3293]), .CO(C[3294]) );
  FA_4895 \FA_INST_0[6].FA_INST_1[222].FA_  ( .A(A[3294]), .B(n802), .CI(
        C[3294]), .CO(C[3295]) );
  FA_4894 \FA_INST_0[6].FA_INST_1[223].FA_  ( .A(A[3295]), .B(n801), .CI(
        C[3295]), .CO(C[3296]) );
  FA_4893 \FA_INST_0[6].FA_INST_1[224].FA_  ( .A(A[3296]), .B(n800), .CI(
        C[3296]), .CO(C[3297]) );
  FA_4892 \FA_INST_0[6].FA_INST_1[225].FA_  ( .A(A[3297]), .B(n799), .CI(
        C[3297]), .CO(C[3298]) );
  FA_4891 \FA_INST_0[6].FA_INST_1[226].FA_  ( .A(A[3298]), .B(n798), .CI(
        C[3298]), .CO(C[3299]) );
  FA_4890 \FA_INST_0[6].FA_INST_1[227].FA_  ( .A(A[3299]), .B(n797), .CI(
        C[3299]), .CO(C[3300]) );
  FA_4889 \FA_INST_0[6].FA_INST_1[228].FA_  ( .A(A[3300]), .B(n796), .CI(
        C[3300]), .CO(C[3301]) );
  FA_4888 \FA_INST_0[6].FA_INST_1[229].FA_  ( .A(A[3301]), .B(n795), .CI(
        C[3301]), .CO(C[3302]) );
  FA_4887 \FA_INST_0[6].FA_INST_1[230].FA_  ( .A(A[3302]), .B(n794), .CI(
        C[3302]), .CO(C[3303]) );
  FA_4886 \FA_INST_0[6].FA_INST_1[231].FA_  ( .A(A[3303]), .B(n793), .CI(
        C[3303]), .CO(C[3304]) );
  FA_4885 \FA_INST_0[6].FA_INST_1[232].FA_  ( .A(A[3304]), .B(n792), .CI(
        C[3304]), .CO(C[3305]) );
  FA_4884 \FA_INST_0[6].FA_INST_1[233].FA_  ( .A(A[3305]), .B(n791), .CI(
        C[3305]), .CO(C[3306]) );
  FA_4883 \FA_INST_0[6].FA_INST_1[234].FA_  ( .A(A[3306]), .B(n790), .CI(
        C[3306]), .CO(C[3307]) );
  FA_4882 \FA_INST_0[6].FA_INST_1[235].FA_  ( .A(A[3307]), .B(n789), .CI(
        C[3307]), .CO(C[3308]) );
  FA_4881 \FA_INST_0[6].FA_INST_1[236].FA_  ( .A(A[3308]), .B(n788), .CI(
        C[3308]), .CO(C[3309]) );
  FA_4880 \FA_INST_0[6].FA_INST_1[237].FA_  ( .A(A[3309]), .B(n787), .CI(
        C[3309]), .CO(C[3310]) );
  FA_4879 \FA_INST_0[6].FA_INST_1[238].FA_  ( .A(A[3310]), .B(n786), .CI(
        C[3310]), .CO(C[3311]) );
  FA_4878 \FA_INST_0[6].FA_INST_1[239].FA_  ( .A(A[3311]), .B(n785), .CI(
        C[3311]), .CO(C[3312]) );
  FA_4877 \FA_INST_0[6].FA_INST_1[240].FA_  ( .A(A[3312]), .B(n784), .CI(
        C[3312]), .CO(C[3313]) );
  FA_4876 \FA_INST_0[6].FA_INST_1[241].FA_  ( .A(A[3313]), .B(n783), .CI(
        C[3313]), .CO(C[3314]) );
  FA_4875 \FA_INST_0[6].FA_INST_1[242].FA_  ( .A(A[3314]), .B(n782), .CI(
        C[3314]), .CO(C[3315]) );
  FA_4874 \FA_INST_0[6].FA_INST_1[243].FA_  ( .A(A[3315]), .B(n781), .CI(
        C[3315]), .CO(C[3316]) );
  FA_4873 \FA_INST_0[6].FA_INST_1[244].FA_  ( .A(A[3316]), .B(n780), .CI(
        C[3316]), .CO(C[3317]) );
  FA_4872 \FA_INST_0[6].FA_INST_1[245].FA_  ( .A(A[3317]), .B(n779), .CI(
        C[3317]), .CO(C[3318]) );
  FA_4871 \FA_INST_0[6].FA_INST_1[246].FA_  ( .A(A[3318]), .B(n778), .CI(
        C[3318]), .CO(C[3319]) );
  FA_4870 \FA_INST_0[6].FA_INST_1[247].FA_  ( .A(A[3319]), .B(n777), .CI(
        C[3319]), .CO(C[3320]) );
  FA_4869 \FA_INST_0[6].FA_INST_1[248].FA_  ( .A(A[3320]), .B(n776), .CI(
        C[3320]), .CO(C[3321]) );
  FA_4868 \FA_INST_0[6].FA_INST_1[249].FA_  ( .A(A[3321]), .B(n775), .CI(
        C[3321]), .CO(C[3322]) );
  FA_4867 \FA_INST_0[6].FA_INST_1[250].FA_  ( .A(A[3322]), .B(n774), .CI(
        C[3322]), .CO(C[3323]) );
  FA_4866 \FA_INST_0[6].FA_INST_1[251].FA_  ( .A(A[3323]), .B(n773), .CI(
        C[3323]), .CO(C[3324]) );
  FA_4865 \FA_INST_0[6].FA_INST_1[252].FA_  ( .A(A[3324]), .B(n772), .CI(
        C[3324]), .CO(C[3325]) );
  FA_4864 \FA_INST_0[6].FA_INST_1[253].FA_  ( .A(A[3325]), .B(n771), .CI(
        C[3325]), .CO(C[3326]) );
  FA_4863 \FA_INST_0[6].FA_INST_1[254].FA_  ( .A(A[3326]), .B(n770), .CI(
        C[3326]), .CO(C[3327]) );
  FA_4862 \FA_INST_0[6].FA_INST_1[255].FA_  ( .A(A[3327]), .B(n769), .CI(
        C[3327]), .CO(C[3328]) );
  FA_4861 \FA_INST_0[6].FA_INST_1[256].FA_  ( .A(A[3328]), .B(n768), .CI(
        C[3328]), .CO(C[3329]) );
  FA_4860 \FA_INST_0[6].FA_INST_1[257].FA_  ( .A(A[3329]), .B(n767), .CI(
        C[3329]), .CO(C[3330]) );
  FA_4859 \FA_INST_0[6].FA_INST_1[258].FA_  ( .A(A[3330]), .B(n766), .CI(
        C[3330]), .CO(C[3331]) );
  FA_4858 \FA_INST_0[6].FA_INST_1[259].FA_  ( .A(A[3331]), .B(n765), .CI(
        C[3331]), .CO(C[3332]) );
  FA_4857 \FA_INST_0[6].FA_INST_1[260].FA_  ( .A(A[3332]), .B(n764), .CI(
        C[3332]), .CO(C[3333]) );
  FA_4856 \FA_INST_0[6].FA_INST_1[261].FA_  ( .A(A[3333]), .B(n763), .CI(
        C[3333]), .CO(C[3334]) );
  FA_4855 \FA_INST_0[6].FA_INST_1[262].FA_  ( .A(A[3334]), .B(n762), .CI(
        C[3334]), .CO(C[3335]) );
  FA_4854 \FA_INST_0[6].FA_INST_1[263].FA_  ( .A(A[3335]), .B(n761), .CI(
        C[3335]), .CO(C[3336]) );
  FA_4853 \FA_INST_0[6].FA_INST_1[264].FA_  ( .A(A[3336]), .B(n760), .CI(
        C[3336]), .CO(C[3337]) );
  FA_4852 \FA_INST_0[6].FA_INST_1[265].FA_  ( .A(A[3337]), .B(n759), .CI(
        C[3337]), .CO(C[3338]) );
  FA_4851 \FA_INST_0[6].FA_INST_1[266].FA_  ( .A(A[3338]), .B(n758), .CI(
        C[3338]), .CO(C[3339]) );
  FA_4850 \FA_INST_0[6].FA_INST_1[267].FA_  ( .A(A[3339]), .B(n757), .CI(
        C[3339]), .CO(C[3340]) );
  FA_4849 \FA_INST_0[6].FA_INST_1[268].FA_  ( .A(A[3340]), .B(n756), .CI(
        C[3340]), .CO(C[3341]) );
  FA_4848 \FA_INST_0[6].FA_INST_1[269].FA_  ( .A(A[3341]), .B(n755), .CI(
        C[3341]), .CO(C[3342]) );
  FA_4847 \FA_INST_0[6].FA_INST_1[270].FA_  ( .A(A[3342]), .B(n754), .CI(
        C[3342]), .CO(C[3343]) );
  FA_4846 \FA_INST_0[6].FA_INST_1[271].FA_  ( .A(A[3343]), .B(n753), .CI(
        C[3343]), .CO(C[3344]) );
  FA_4845 \FA_INST_0[6].FA_INST_1[272].FA_  ( .A(A[3344]), .B(n752), .CI(
        C[3344]), .CO(C[3345]) );
  FA_4844 \FA_INST_0[6].FA_INST_1[273].FA_  ( .A(A[3345]), .B(n751), .CI(
        C[3345]), .CO(C[3346]) );
  FA_4843 \FA_INST_0[6].FA_INST_1[274].FA_  ( .A(A[3346]), .B(n750), .CI(
        C[3346]), .CO(C[3347]) );
  FA_4842 \FA_INST_0[6].FA_INST_1[275].FA_  ( .A(A[3347]), .B(n749), .CI(
        C[3347]), .CO(C[3348]) );
  FA_4841 \FA_INST_0[6].FA_INST_1[276].FA_  ( .A(A[3348]), .B(n748), .CI(
        C[3348]), .CO(C[3349]) );
  FA_4840 \FA_INST_0[6].FA_INST_1[277].FA_  ( .A(A[3349]), .B(n747), .CI(
        C[3349]), .CO(C[3350]) );
  FA_4839 \FA_INST_0[6].FA_INST_1[278].FA_  ( .A(A[3350]), .B(n746), .CI(
        C[3350]), .CO(C[3351]) );
  FA_4838 \FA_INST_0[6].FA_INST_1[279].FA_  ( .A(A[3351]), .B(n745), .CI(
        C[3351]), .CO(C[3352]) );
  FA_4837 \FA_INST_0[6].FA_INST_1[280].FA_  ( .A(A[3352]), .B(n744), .CI(
        C[3352]), .CO(C[3353]) );
  FA_4836 \FA_INST_0[6].FA_INST_1[281].FA_  ( .A(A[3353]), .B(n743), .CI(
        C[3353]), .CO(C[3354]) );
  FA_4835 \FA_INST_0[6].FA_INST_1[282].FA_  ( .A(A[3354]), .B(n742), .CI(
        C[3354]), .CO(C[3355]) );
  FA_4834 \FA_INST_0[6].FA_INST_1[283].FA_  ( .A(A[3355]), .B(n741), .CI(
        C[3355]), .CO(C[3356]) );
  FA_4833 \FA_INST_0[6].FA_INST_1[284].FA_  ( .A(A[3356]), .B(n740), .CI(
        C[3356]), .CO(C[3357]) );
  FA_4832 \FA_INST_0[6].FA_INST_1[285].FA_  ( .A(A[3357]), .B(n739), .CI(
        C[3357]), .CO(C[3358]) );
  FA_4831 \FA_INST_0[6].FA_INST_1[286].FA_  ( .A(A[3358]), .B(n738), .CI(
        C[3358]), .CO(C[3359]) );
  FA_4830 \FA_INST_0[6].FA_INST_1[287].FA_  ( .A(A[3359]), .B(n737), .CI(
        C[3359]), .CO(C[3360]) );
  FA_4829 \FA_INST_0[6].FA_INST_1[288].FA_  ( .A(A[3360]), .B(n736), .CI(
        C[3360]), .CO(C[3361]) );
  FA_4828 \FA_INST_0[6].FA_INST_1[289].FA_  ( .A(A[3361]), .B(n735), .CI(
        C[3361]), .CO(C[3362]) );
  FA_4827 \FA_INST_0[6].FA_INST_1[290].FA_  ( .A(A[3362]), .B(n734), .CI(
        C[3362]), .CO(C[3363]) );
  FA_4826 \FA_INST_0[6].FA_INST_1[291].FA_  ( .A(A[3363]), .B(n733), .CI(
        C[3363]), .CO(C[3364]) );
  FA_4825 \FA_INST_0[6].FA_INST_1[292].FA_  ( .A(A[3364]), .B(n732), .CI(
        C[3364]), .CO(C[3365]) );
  FA_4824 \FA_INST_0[6].FA_INST_1[293].FA_  ( .A(A[3365]), .B(n731), .CI(
        C[3365]), .CO(C[3366]) );
  FA_4823 \FA_INST_0[6].FA_INST_1[294].FA_  ( .A(A[3366]), .B(n730), .CI(
        C[3366]), .CO(C[3367]) );
  FA_4822 \FA_INST_0[6].FA_INST_1[295].FA_  ( .A(A[3367]), .B(n729), .CI(
        C[3367]), .CO(C[3368]) );
  FA_4821 \FA_INST_0[6].FA_INST_1[296].FA_  ( .A(A[3368]), .B(n728), .CI(
        C[3368]), .CO(C[3369]) );
  FA_4820 \FA_INST_0[6].FA_INST_1[297].FA_  ( .A(A[3369]), .B(n727), .CI(
        C[3369]), .CO(C[3370]) );
  FA_4819 \FA_INST_0[6].FA_INST_1[298].FA_  ( .A(A[3370]), .B(n726), .CI(
        C[3370]), .CO(C[3371]) );
  FA_4818 \FA_INST_0[6].FA_INST_1[299].FA_  ( .A(A[3371]), .B(n725), .CI(
        C[3371]), .CO(C[3372]) );
  FA_4817 \FA_INST_0[6].FA_INST_1[300].FA_  ( .A(A[3372]), .B(n724), .CI(
        C[3372]), .CO(C[3373]) );
  FA_4816 \FA_INST_0[6].FA_INST_1[301].FA_  ( .A(A[3373]), .B(n723), .CI(
        C[3373]), .CO(C[3374]) );
  FA_4815 \FA_INST_0[6].FA_INST_1[302].FA_  ( .A(A[3374]), .B(n722), .CI(
        C[3374]), .CO(C[3375]) );
  FA_4814 \FA_INST_0[6].FA_INST_1[303].FA_  ( .A(A[3375]), .B(n721), .CI(
        C[3375]), .CO(C[3376]) );
  FA_4813 \FA_INST_0[6].FA_INST_1[304].FA_  ( .A(A[3376]), .B(n720), .CI(
        C[3376]), .CO(C[3377]) );
  FA_4812 \FA_INST_0[6].FA_INST_1[305].FA_  ( .A(A[3377]), .B(n719), .CI(
        C[3377]), .CO(C[3378]) );
  FA_4811 \FA_INST_0[6].FA_INST_1[306].FA_  ( .A(A[3378]), .B(n718), .CI(
        C[3378]), .CO(C[3379]) );
  FA_4810 \FA_INST_0[6].FA_INST_1[307].FA_  ( .A(A[3379]), .B(n717), .CI(
        C[3379]), .CO(C[3380]) );
  FA_4809 \FA_INST_0[6].FA_INST_1[308].FA_  ( .A(A[3380]), .B(n716), .CI(
        C[3380]), .CO(C[3381]) );
  FA_4808 \FA_INST_0[6].FA_INST_1[309].FA_  ( .A(A[3381]), .B(n715), .CI(
        C[3381]), .CO(C[3382]) );
  FA_4807 \FA_INST_0[6].FA_INST_1[310].FA_  ( .A(A[3382]), .B(n714), .CI(
        C[3382]), .CO(C[3383]) );
  FA_4806 \FA_INST_0[6].FA_INST_1[311].FA_  ( .A(A[3383]), .B(n713), .CI(
        C[3383]), .CO(C[3384]) );
  FA_4805 \FA_INST_0[6].FA_INST_1[312].FA_  ( .A(A[3384]), .B(n712), .CI(
        C[3384]), .CO(C[3385]) );
  FA_4804 \FA_INST_0[6].FA_INST_1[313].FA_  ( .A(A[3385]), .B(n711), .CI(
        C[3385]), .CO(C[3386]) );
  FA_4803 \FA_INST_0[6].FA_INST_1[314].FA_  ( .A(A[3386]), .B(n710), .CI(
        C[3386]), .CO(C[3387]) );
  FA_4802 \FA_INST_0[6].FA_INST_1[315].FA_  ( .A(A[3387]), .B(n709), .CI(
        C[3387]), .CO(C[3388]) );
  FA_4801 \FA_INST_0[6].FA_INST_1[316].FA_  ( .A(A[3388]), .B(n708), .CI(
        C[3388]), .CO(C[3389]) );
  FA_4800 \FA_INST_0[6].FA_INST_1[317].FA_  ( .A(A[3389]), .B(n707), .CI(
        C[3389]), .CO(C[3390]) );
  FA_4799 \FA_INST_0[6].FA_INST_1[318].FA_  ( .A(A[3390]), .B(n706), .CI(
        C[3390]), .CO(C[3391]) );
  FA_4798 \FA_INST_0[6].FA_INST_1[319].FA_  ( .A(A[3391]), .B(n705), .CI(
        C[3391]), .CO(C[3392]) );
  FA_4797 \FA_INST_0[6].FA_INST_1[320].FA_  ( .A(A[3392]), .B(n704), .CI(
        C[3392]), .CO(C[3393]) );
  FA_4796 \FA_INST_0[6].FA_INST_1[321].FA_  ( .A(A[3393]), .B(n703), .CI(
        C[3393]), .CO(C[3394]) );
  FA_4795 \FA_INST_0[6].FA_INST_1[322].FA_  ( .A(A[3394]), .B(n702), .CI(
        C[3394]), .CO(C[3395]) );
  FA_4794 \FA_INST_0[6].FA_INST_1[323].FA_  ( .A(A[3395]), .B(n701), .CI(
        C[3395]), .CO(C[3396]) );
  FA_4793 \FA_INST_0[6].FA_INST_1[324].FA_  ( .A(A[3396]), .B(n700), .CI(
        C[3396]), .CO(C[3397]) );
  FA_4792 \FA_INST_0[6].FA_INST_1[325].FA_  ( .A(A[3397]), .B(n699), .CI(
        C[3397]), .CO(C[3398]) );
  FA_4791 \FA_INST_0[6].FA_INST_1[326].FA_  ( .A(A[3398]), .B(n698), .CI(
        C[3398]), .CO(C[3399]) );
  FA_4790 \FA_INST_0[6].FA_INST_1[327].FA_  ( .A(A[3399]), .B(n697), .CI(
        C[3399]), .CO(C[3400]) );
  FA_4789 \FA_INST_0[6].FA_INST_1[328].FA_  ( .A(A[3400]), .B(n696), .CI(
        C[3400]), .CO(C[3401]) );
  FA_4788 \FA_INST_0[6].FA_INST_1[329].FA_  ( .A(A[3401]), .B(n695), .CI(
        C[3401]), .CO(C[3402]) );
  FA_4787 \FA_INST_0[6].FA_INST_1[330].FA_  ( .A(A[3402]), .B(n694), .CI(
        C[3402]), .CO(C[3403]) );
  FA_4786 \FA_INST_0[6].FA_INST_1[331].FA_  ( .A(A[3403]), .B(n693), .CI(
        C[3403]), .CO(C[3404]) );
  FA_4785 \FA_INST_0[6].FA_INST_1[332].FA_  ( .A(A[3404]), .B(n692), .CI(
        C[3404]), .CO(C[3405]) );
  FA_4784 \FA_INST_0[6].FA_INST_1[333].FA_  ( .A(A[3405]), .B(n691), .CI(
        C[3405]), .CO(C[3406]) );
  FA_4783 \FA_INST_0[6].FA_INST_1[334].FA_  ( .A(A[3406]), .B(n690), .CI(
        C[3406]), .CO(C[3407]) );
  FA_4782 \FA_INST_0[6].FA_INST_1[335].FA_  ( .A(A[3407]), .B(n689), .CI(
        C[3407]), .CO(C[3408]) );
  FA_4781 \FA_INST_0[6].FA_INST_1[336].FA_  ( .A(A[3408]), .B(n688), .CI(
        C[3408]), .CO(C[3409]) );
  FA_4780 \FA_INST_0[6].FA_INST_1[337].FA_  ( .A(A[3409]), .B(n687), .CI(
        C[3409]), .CO(C[3410]) );
  FA_4779 \FA_INST_0[6].FA_INST_1[338].FA_  ( .A(A[3410]), .B(n686), .CI(
        C[3410]), .CO(C[3411]) );
  FA_4778 \FA_INST_0[6].FA_INST_1[339].FA_  ( .A(A[3411]), .B(n685), .CI(
        C[3411]), .CO(C[3412]) );
  FA_4777 \FA_INST_0[6].FA_INST_1[340].FA_  ( .A(A[3412]), .B(n684), .CI(
        C[3412]), .CO(C[3413]) );
  FA_4776 \FA_INST_0[6].FA_INST_1[341].FA_  ( .A(A[3413]), .B(n683), .CI(
        C[3413]), .CO(C[3414]) );
  FA_4775 \FA_INST_0[6].FA_INST_1[342].FA_  ( .A(A[3414]), .B(n682), .CI(
        C[3414]), .CO(C[3415]) );
  FA_4774 \FA_INST_0[6].FA_INST_1[343].FA_  ( .A(A[3415]), .B(n681), .CI(
        C[3415]), .CO(C[3416]) );
  FA_4773 \FA_INST_0[6].FA_INST_1[344].FA_  ( .A(A[3416]), .B(n680), .CI(
        C[3416]), .CO(C[3417]) );
  FA_4772 \FA_INST_0[6].FA_INST_1[345].FA_  ( .A(A[3417]), .B(n679), .CI(
        C[3417]), .CO(C[3418]) );
  FA_4771 \FA_INST_0[6].FA_INST_1[346].FA_  ( .A(A[3418]), .B(n678), .CI(
        C[3418]), .CO(C[3419]) );
  FA_4770 \FA_INST_0[6].FA_INST_1[347].FA_  ( .A(A[3419]), .B(n677), .CI(
        C[3419]), .CO(C[3420]) );
  FA_4769 \FA_INST_0[6].FA_INST_1[348].FA_  ( .A(A[3420]), .B(n676), .CI(
        C[3420]), .CO(C[3421]) );
  FA_4768 \FA_INST_0[6].FA_INST_1[349].FA_  ( .A(A[3421]), .B(n675), .CI(
        C[3421]), .CO(C[3422]) );
  FA_4767 \FA_INST_0[6].FA_INST_1[350].FA_  ( .A(A[3422]), .B(n674), .CI(
        C[3422]), .CO(C[3423]) );
  FA_4766 \FA_INST_0[6].FA_INST_1[351].FA_  ( .A(A[3423]), .B(n673), .CI(
        C[3423]), .CO(C[3424]) );
  FA_4765 \FA_INST_0[6].FA_INST_1[352].FA_  ( .A(A[3424]), .B(n672), .CI(
        C[3424]), .CO(C[3425]) );
  FA_4764 \FA_INST_0[6].FA_INST_1[353].FA_  ( .A(A[3425]), .B(n671), .CI(
        C[3425]), .CO(C[3426]) );
  FA_4763 \FA_INST_0[6].FA_INST_1[354].FA_  ( .A(A[3426]), .B(n670), .CI(
        C[3426]), .CO(C[3427]) );
  FA_4762 \FA_INST_0[6].FA_INST_1[355].FA_  ( .A(A[3427]), .B(n669), .CI(
        C[3427]), .CO(C[3428]) );
  FA_4761 \FA_INST_0[6].FA_INST_1[356].FA_  ( .A(A[3428]), .B(n668), .CI(
        C[3428]), .CO(C[3429]) );
  FA_4760 \FA_INST_0[6].FA_INST_1[357].FA_  ( .A(A[3429]), .B(n667), .CI(
        C[3429]), .CO(C[3430]) );
  FA_4759 \FA_INST_0[6].FA_INST_1[358].FA_  ( .A(A[3430]), .B(n666), .CI(
        C[3430]), .CO(C[3431]) );
  FA_4758 \FA_INST_0[6].FA_INST_1[359].FA_  ( .A(A[3431]), .B(n665), .CI(
        C[3431]), .CO(C[3432]) );
  FA_4757 \FA_INST_0[6].FA_INST_1[360].FA_  ( .A(A[3432]), .B(n664), .CI(
        C[3432]), .CO(C[3433]) );
  FA_4756 \FA_INST_0[6].FA_INST_1[361].FA_  ( .A(A[3433]), .B(n663), .CI(
        C[3433]), .CO(C[3434]) );
  FA_4755 \FA_INST_0[6].FA_INST_1[362].FA_  ( .A(A[3434]), .B(n662), .CI(
        C[3434]), .CO(C[3435]) );
  FA_4754 \FA_INST_0[6].FA_INST_1[363].FA_  ( .A(A[3435]), .B(n661), .CI(
        C[3435]), .CO(C[3436]) );
  FA_4753 \FA_INST_0[6].FA_INST_1[364].FA_  ( .A(A[3436]), .B(n660), .CI(
        C[3436]), .CO(C[3437]) );
  FA_4752 \FA_INST_0[6].FA_INST_1[365].FA_  ( .A(A[3437]), .B(n659), .CI(
        C[3437]), .CO(C[3438]) );
  FA_4751 \FA_INST_0[6].FA_INST_1[366].FA_  ( .A(A[3438]), .B(n658), .CI(
        C[3438]), .CO(C[3439]) );
  FA_4750 \FA_INST_0[6].FA_INST_1[367].FA_  ( .A(A[3439]), .B(n657), .CI(
        C[3439]), .CO(C[3440]) );
  FA_4749 \FA_INST_0[6].FA_INST_1[368].FA_  ( .A(A[3440]), .B(n656), .CI(
        C[3440]), .CO(C[3441]) );
  FA_4748 \FA_INST_0[6].FA_INST_1[369].FA_  ( .A(A[3441]), .B(n655), .CI(
        C[3441]), .CO(C[3442]) );
  FA_4747 \FA_INST_0[6].FA_INST_1[370].FA_  ( .A(A[3442]), .B(n654), .CI(
        C[3442]), .CO(C[3443]) );
  FA_4746 \FA_INST_0[6].FA_INST_1[371].FA_  ( .A(A[3443]), .B(n653), .CI(
        C[3443]), .CO(C[3444]) );
  FA_4745 \FA_INST_0[6].FA_INST_1[372].FA_  ( .A(A[3444]), .B(n652), .CI(
        C[3444]), .CO(C[3445]) );
  FA_4744 \FA_INST_0[6].FA_INST_1[373].FA_  ( .A(A[3445]), .B(n651), .CI(
        C[3445]), .CO(C[3446]) );
  FA_4743 \FA_INST_0[6].FA_INST_1[374].FA_  ( .A(A[3446]), .B(n650), .CI(
        C[3446]), .CO(C[3447]) );
  FA_4742 \FA_INST_0[6].FA_INST_1[375].FA_  ( .A(A[3447]), .B(n649), .CI(
        C[3447]), .CO(C[3448]) );
  FA_4741 \FA_INST_0[6].FA_INST_1[376].FA_  ( .A(A[3448]), .B(n648), .CI(
        C[3448]), .CO(C[3449]) );
  FA_4740 \FA_INST_0[6].FA_INST_1[377].FA_  ( .A(A[3449]), .B(n647), .CI(
        C[3449]), .CO(C[3450]) );
  FA_4739 \FA_INST_0[6].FA_INST_1[378].FA_  ( .A(A[3450]), .B(n646), .CI(
        C[3450]), .CO(C[3451]) );
  FA_4738 \FA_INST_0[6].FA_INST_1[379].FA_  ( .A(A[3451]), .B(n645), .CI(
        C[3451]), .CO(C[3452]) );
  FA_4737 \FA_INST_0[6].FA_INST_1[380].FA_  ( .A(A[3452]), .B(n644), .CI(
        C[3452]), .CO(C[3453]) );
  FA_4736 \FA_INST_0[6].FA_INST_1[381].FA_  ( .A(A[3453]), .B(n643), .CI(
        C[3453]), .CO(C[3454]) );
  FA_4735 \FA_INST_0[6].FA_INST_1[382].FA_  ( .A(A[3454]), .B(n642), .CI(
        C[3454]), .CO(C[3455]) );
  FA_4734 \FA_INST_0[6].FA_INST_1[383].FA_  ( .A(A[3455]), .B(n641), .CI(
        C[3455]), .CO(C[3456]) );
  FA_4733 \FA_INST_0[6].FA_INST_1[384].FA_  ( .A(A[3456]), .B(n640), .CI(
        C[3456]), .CO(C[3457]) );
  FA_4732 \FA_INST_0[6].FA_INST_1[385].FA_  ( .A(A[3457]), .B(n639), .CI(
        C[3457]), .CO(C[3458]) );
  FA_4731 \FA_INST_0[6].FA_INST_1[386].FA_  ( .A(A[3458]), .B(n638), .CI(
        C[3458]), .CO(C[3459]) );
  FA_4730 \FA_INST_0[6].FA_INST_1[387].FA_  ( .A(A[3459]), .B(n637), .CI(
        C[3459]), .CO(C[3460]) );
  FA_4729 \FA_INST_0[6].FA_INST_1[388].FA_  ( .A(A[3460]), .B(n636), .CI(
        C[3460]), .CO(C[3461]) );
  FA_4728 \FA_INST_0[6].FA_INST_1[389].FA_  ( .A(A[3461]), .B(n635), .CI(
        C[3461]), .CO(C[3462]) );
  FA_4727 \FA_INST_0[6].FA_INST_1[390].FA_  ( .A(A[3462]), .B(n634), .CI(
        C[3462]), .CO(C[3463]) );
  FA_4726 \FA_INST_0[6].FA_INST_1[391].FA_  ( .A(A[3463]), .B(n633), .CI(
        C[3463]), .CO(C[3464]) );
  FA_4725 \FA_INST_0[6].FA_INST_1[392].FA_  ( .A(A[3464]), .B(n632), .CI(
        C[3464]), .CO(C[3465]) );
  FA_4724 \FA_INST_0[6].FA_INST_1[393].FA_  ( .A(A[3465]), .B(n631), .CI(
        C[3465]), .CO(C[3466]) );
  FA_4723 \FA_INST_0[6].FA_INST_1[394].FA_  ( .A(A[3466]), .B(n630), .CI(
        C[3466]), .CO(C[3467]) );
  FA_4722 \FA_INST_0[6].FA_INST_1[395].FA_  ( .A(A[3467]), .B(n629), .CI(
        C[3467]), .CO(C[3468]) );
  FA_4721 \FA_INST_0[6].FA_INST_1[396].FA_  ( .A(A[3468]), .B(n628), .CI(
        C[3468]), .CO(C[3469]) );
  FA_4720 \FA_INST_0[6].FA_INST_1[397].FA_  ( .A(A[3469]), .B(n627), .CI(
        C[3469]), .CO(C[3470]) );
  FA_4719 \FA_INST_0[6].FA_INST_1[398].FA_  ( .A(A[3470]), .B(n626), .CI(
        C[3470]), .CO(C[3471]) );
  FA_4718 \FA_INST_0[6].FA_INST_1[399].FA_  ( .A(A[3471]), .B(n625), .CI(
        C[3471]), .CO(C[3472]) );
  FA_4717 \FA_INST_0[6].FA_INST_1[400].FA_  ( .A(A[3472]), .B(n624), .CI(
        C[3472]), .CO(C[3473]) );
  FA_4716 \FA_INST_0[6].FA_INST_1[401].FA_  ( .A(A[3473]), .B(n623), .CI(
        C[3473]), .CO(C[3474]) );
  FA_4715 \FA_INST_0[6].FA_INST_1[402].FA_  ( .A(A[3474]), .B(n622), .CI(
        C[3474]), .CO(C[3475]) );
  FA_4714 \FA_INST_0[6].FA_INST_1[403].FA_  ( .A(A[3475]), .B(n621), .CI(
        C[3475]), .CO(C[3476]) );
  FA_4713 \FA_INST_0[6].FA_INST_1[404].FA_  ( .A(A[3476]), .B(n620), .CI(
        C[3476]), .CO(C[3477]) );
  FA_4712 \FA_INST_0[6].FA_INST_1[405].FA_  ( .A(A[3477]), .B(n619), .CI(
        C[3477]), .CO(C[3478]) );
  FA_4711 \FA_INST_0[6].FA_INST_1[406].FA_  ( .A(A[3478]), .B(n618), .CI(
        C[3478]), .CO(C[3479]) );
  FA_4710 \FA_INST_0[6].FA_INST_1[407].FA_  ( .A(A[3479]), .B(n617), .CI(
        C[3479]), .CO(C[3480]) );
  FA_4709 \FA_INST_0[6].FA_INST_1[408].FA_  ( .A(A[3480]), .B(n616), .CI(
        C[3480]), .CO(C[3481]) );
  FA_4708 \FA_INST_0[6].FA_INST_1[409].FA_  ( .A(A[3481]), .B(n615), .CI(
        C[3481]), .CO(C[3482]) );
  FA_4707 \FA_INST_0[6].FA_INST_1[410].FA_  ( .A(A[3482]), .B(n614), .CI(
        C[3482]), .CO(C[3483]) );
  FA_4706 \FA_INST_0[6].FA_INST_1[411].FA_  ( .A(A[3483]), .B(n613), .CI(
        C[3483]), .CO(C[3484]) );
  FA_4705 \FA_INST_0[6].FA_INST_1[412].FA_  ( .A(A[3484]), .B(n612), .CI(
        C[3484]), .CO(C[3485]) );
  FA_4704 \FA_INST_0[6].FA_INST_1[413].FA_  ( .A(A[3485]), .B(n611), .CI(
        C[3485]), .CO(C[3486]) );
  FA_4703 \FA_INST_0[6].FA_INST_1[414].FA_  ( .A(A[3486]), .B(n610), .CI(
        C[3486]), .CO(C[3487]) );
  FA_4702 \FA_INST_0[6].FA_INST_1[415].FA_  ( .A(A[3487]), .B(n609), .CI(
        C[3487]), .CO(C[3488]) );
  FA_4701 \FA_INST_0[6].FA_INST_1[416].FA_  ( .A(A[3488]), .B(n608), .CI(
        C[3488]), .CO(C[3489]) );
  FA_4700 \FA_INST_0[6].FA_INST_1[417].FA_  ( .A(A[3489]), .B(n607), .CI(
        C[3489]), .CO(C[3490]) );
  FA_4699 \FA_INST_0[6].FA_INST_1[418].FA_  ( .A(A[3490]), .B(n606), .CI(
        C[3490]), .CO(C[3491]) );
  FA_4698 \FA_INST_0[6].FA_INST_1[419].FA_  ( .A(A[3491]), .B(n605), .CI(
        C[3491]), .CO(C[3492]) );
  FA_4697 \FA_INST_0[6].FA_INST_1[420].FA_  ( .A(A[3492]), .B(n604), .CI(
        C[3492]), .CO(C[3493]) );
  FA_4696 \FA_INST_0[6].FA_INST_1[421].FA_  ( .A(A[3493]), .B(n603), .CI(
        C[3493]), .CO(C[3494]) );
  FA_4695 \FA_INST_0[6].FA_INST_1[422].FA_  ( .A(A[3494]), .B(n602), .CI(
        C[3494]), .CO(C[3495]) );
  FA_4694 \FA_INST_0[6].FA_INST_1[423].FA_  ( .A(A[3495]), .B(n601), .CI(
        C[3495]), .CO(C[3496]) );
  FA_4693 \FA_INST_0[6].FA_INST_1[424].FA_  ( .A(A[3496]), .B(n600), .CI(
        C[3496]), .CO(C[3497]) );
  FA_4692 \FA_INST_0[6].FA_INST_1[425].FA_  ( .A(A[3497]), .B(n599), .CI(
        C[3497]), .CO(C[3498]) );
  FA_4691 \FA_INST_0[6].FA_INST_1[426].FA_  ( .A(A[3498]), .B(n598), .CI(
        C[3498]), .CO(C[3499]) );
  FA_4690 \FA_INST_0[6].FA_INST_1[427].FA_  ( .A(A[3499]), .B(n597), .CI(
        C[3499]), .CO(C[3500]) );
  FA_4689 \FA_INST_0[6].FA_INST_1[428].FA_  ( .A(A[3500]), .B(n596), .CI(
        C[3500]), .CO(C[3501]) );
  FA_4688 \FA_INST_0[6].FA_INST_1[429].FA_  ( .A(A[3501]), .B(n595), .CI(
        C[3501]), .CO(C[3502]) );
  FA_4687 \FA_INST_0[6].FA_INST_1[430].FA_  ( .A(A[3502]), .B(n594), .CI(
        C[3502]), .CO(C[3503]) );
  FA_4686 \FA_INST_0[6].FA_INST_1[431].FA_  ( .A(A[3503]), .B(n593), .CI(
        C[3503]), .CO(C[3504]) );
  FA_4685 \FA_INST_0[6].FA_INST_1[432].FA_  ( .A(A[3504]), .B(n592), .CI(
        C[3504]), .CO(C[3505]) );
  FA_4684 \FA_INST_0[6].FA_INST_1[433].FA_  ( .A(A[3505]), .B(n591), .CI(
        C[3505]), .CO(C[3506]) );
  FA_4683 \FA_INST_0[6].FA_INST_1[434].FA_  ( .A(A[3506]), .B(n590), .CI(
        C[3506]), .CO(C[3507]) );
  FA_4682 \FA_INST_0[6].FA_INST_1[435].FA_  ( .A(A[3507]), .B(n589), .CI(
        C[3507]), .CO(C[3508]) );
  FA_4681 \FA_INST_0[6].FA_INST_1[436].FA_  ( .A(A[3508]), .B(n588), .CI(
        C[3508]), .CO(C[3509]) );
  FA_4680 \FA_INST_0[6].FA_INST_1[437].FA_  ( .A(A[3509]), .B(n587), .CI(
        C[3509]), .CO(C[3510]) );
  FA_4679 \FA_INST_0[6].FA_INST_1[438].FA_  ( .A(A[3510]), .B(n586), .CI(
        C[3510]), .CO(C[3511]) );
  FA_4678 \FA_INST_0[6].FA_INST_1[439].FA_  ( .A(A[3511]), .B(n585), .CI(
        C[3511]), .CO(C[3512]) );
  FA_4677 \FA_INST_0[6].FA_INST_1[440].FA_  ( .A(A[3512]), .B(n584), .CI(
        C[3512]), .CO(C[3513]) );
  FA_4676 \FA_INST_0[6].FA_INST_1[441].FA_  ( .A(A[3513]), .B(n583), .CI(
        C[3513]), .CO(C[3514]) );
  FA_4675 \FA_INST_0[6].FA_INST_1[442].FA_  ( .A(A[3514]), .B(n582), .CI(
        C[3514]), .CO(C[3515]) );
  FA_4674 \FA_INST_0[6].FA_INST_1[443].FA_  ( .A(A[3515]), .B(n581), .CI(
        C[3515]), .CO(C[3516]) );
  FA_4673 \FA_INST_0[6].FA_INST_1[444].FA_  ( .A(A[3516]), .B(n580), .CI(
        C[3516]), .CO(C[3517]) );
  FA_4672 \FA_INST_0[6].FA_INST_1[445].FA_  ( .A(A[3517]), .B(n579), .CI(
        C[3517]), .CO(C[3518]) );
  FA_4671 \FA_INST_0[6].FA_INST_1[446].FA_  ( .A(A[3518]), .B(n578), .CI(
        C[3518]), .CO(C[3519]) );
  FA_4670 \FA_INST_0[6].FA_INST_1[447].FA_  ( .A(A[3519]), .B(n577), .CI(
        C[3519]), .CO(C[3520]) );
  FA_4669 \FA_INST_0[6].FA_INST_1[448].FA_  ( .A(A[3520]), .B(n576), .CI(
        C[3520]), .CO(C[3521]) );
  FA_4668 \FA_INST_0[6].FA_INST_1[449].FA_  ( .A(A[3521]), .B(n575), .CI(
        C[3521]), .CO(C[3522]) );
  FA_4667 \FA_INST_0[6].FA_INST_1[450].FA_  ( .A(A[3522]), .B(n574), .CI(
        C[3522]), .CO(C[3523]) );
  FA_4666 \FA_INST_0[6].FA_INST_1[451].FA_  ( .A(A[3523]), .B(n573), .CI(
        C[3523]), .CO(C[3524]) );
  FA_4665 \FA_INST_0[6].FA_INST_1[452].FA_  ( .A(A[3524]), .B(n572), .CI(
        C[3524]), .CO(C[3525]) );
  FA_4664 \FA_INST_0[6].FA_INST_1[453].FA_  ( .A(A[3525]), .B(n571), .CI(
        C[3525]), .CO(C[3526]) );
  FA_4663 \FA_INST_0[6].FA_INST_1[454].FA_  ( .A(A[3526]), .B(n570), .CI(
        C[3526]), .CO(C[3527]) );
  FA_4662 \FA_INST_0[6].FA_INST_1[455].FA_  ( .A(A[3527]), .B(n569), .CI(
        C[3527]), .CO(C[3528]) );
  FA_4661 \FA_INST_0[6].FA_INST_1[456].FA_  ( .A(A[3528]), .B(n568), .CI(
        C[3528]), .CO(C[3529]) );
  FA_4660 \FA_INST_0[6].FA_INST_1[457].FA_  ( .A(A[3529]), .B(n567), .CI(
        C[3529]), .CO(C[3530]) );
  FA_4659 \FA_INST_0[6].FA_INST_1[458].FA_  ( .A(A[3530]), .B(n566), .CI(
        C[3530]), .CO(C[3531]) );
  FA_4658 \FA_INST_0[6].FA_INST_1[459].FA_  ( .A(A[3531]), .B(n565), .CI(
        C[3531]), .CO(C[3532]) );
  FA_4657 \FA_INST_0[6].FA_INST_1[460].FA_  ( .A(A[3532]), .B(n564), .CI(
        C[3532]), .CO(C[3533]) );
  FA_4656 \FA_INST_0[6].FA_INST_1[461].FA_  ( .A(A[3533]), .B(n563), .CI(
        C[3533]), .CO(C[3534]) );
  FA_4655 \FA_INST_0[6].FA_INST_1[462].FA_  ( .A(A[3534]), .B(n562), .CI(
        C[3534]), .CO(C[3535]) );
  FA_4654 \FA_INST_0[6].FA_INST_1[463].FA_  ( .A(A[3535]), .B(n561), .CI(
        C[3535]), .CO(C[3536]) );
  FA_4653 \FA_INST_0[6].FA_INST_1[464].FA_  ( .A(A[3536]), .B(n560), .CI(
        C[3536]), .CO(C[3537]) );
  FA_4652 \FA_INST_0[6].FA_INST_1[465].FA_  ( .A(A[3537]), .B(n559), .CI(
        C[3537]), .CO(C[3538]) );
  FA_4651 \FA_INST_0[6].FA_INST_1[466].FA_  ( .A(A[3538]), .B(n558), .CI(
        C[3538]), .CO(C[3539]) );
  FA_4650 \FA_INST_0[6].FA_INST_1[467].FA_  ( .A(A[3539]), .B(n557), .CI(
        C[3539]), .CO(C[3540]) );
  FA_4649 \FA_INST_0[6].FA_INST_1[468].FA_  ( .A(A[3540]), .B(n556), .CI(
        C[3540]), .CO(C[3541]) );
  FA_4648 \FA_INST_0[6].FA_INST_1[469].FA_  ( .A(A[3541]), .B(n555), .CI(
        C[3541]), .CO(C[3542]) );
  FA_4647 \FA_INST_0[6].FA_INST_1[470].FA_  ( .A(A[3542]), .B(n554), .CI(
        C[3542]), .CO(C[3543]) );
  FA_4646 \FA_INST_0[6].FA_INST_1[471].FA_  ( .A(A[3543]), .B(n553), .CI(
        C[3543]), .CO(C[3544]) );
  FA_4645 \FA_INST_0[6].FA_INST_1[472].FA_  ( .A(A[3544]), .B(n552), .CI(
        C[3544]), .CO(C[3545]) );
  FA_4644 \FA_INST_0[6].FA_INST_1[473].FA_  ( .A(A[3545]), .B(n551), .CI(
        C[3545]), .CO(C[3546]) );
  FA_4643 \FA_INST_0[6].FA_INST_1[474].FA_  ( .A(A[3546]), .B(n550), .CI(
        C[3546]), .CO(C[3547]) );
  FA_4642 \FA_INST_0[6].FA_INST_1[475].FA_  ( .A(A[3547]), .B(n549), .CI(
        C[3547]), .CO(C[3548]) );
  FA_4641 \FA_INST_0[6].FA_INST_1[476].FA_  ( .A(A[3548]), .B(n548), .CI(
        C[3548]), .CO(C[3549]) );
  FA_4640 \FA_INST_0[6].FA_INST_1[477].FA_  ( .A(A[3549]), .B(n547), .CI(
        C[3549]), .CO(C[3550]) );
  FA_4639 \FA_INST_0[6].FA_INST_1[478].FA_  ( .A(A[3550]), .B(n546), .CI(
        C[3550]), .CO(C[3551]) );
  FA_4638 \FA_INST_0[6].FA_INST_1[479].FA_  ( .A(A[3551]), .B(n545), .CI(
        C[3551]), .CO(C[3552]) );
  FA_4637 \FA_INST_0[6].FA_INST_1[480].FA_  ( .A(A[3552]), .B(n544), .CI(
        C[3552]), .CO(C[3553]) );
  FA_4636 \FA_INST_0[6].FA_INST_1[481].FA_  ( .A(A[3553]), .B(n543), .CI(
        C[3553]), .CO(C[3554]) );
  FA_4635 \FA_INST_0[6].FA_INST_1[482].FA_  ( .A(A[3554]), .B(n542), .CI(
        C[3554]), .CO(C[3555]) );
  FA_4634 \FA_INST_0[6].FA_INST_1[483].FA_  ( .A(A[3555]), .B(n541), .CI(
        C[3555]), .CO(C[3556]) );
  FA_4633 \FA_INST_0[6].FA_INST_1[484].FA_  ( .A(A[3556]), .B(n540), .CI(
        C[3556]), .CO(C[3557]) );
  FA_4632 \FA_INST_0[6].FA_INST_1[485].FA_  ( .A(A[3557]), .B(n539), .CI(
        C[3557]), .CO(C[3558]) );
  FA_4631 \FA_INST_0[6].FA_INST_1[486].FA_  ( .A(A[3558]), .B(n538), .CI(
        C[3558]), .CO(C[3559]) );
  FA_4630 \FA_INST_0[6].FA_INST_1[487].FA_  ( .A(A[3559]), .B(n537), .CI(
        C[3559]), .CO(C[3560]) );
  FA_4629 \FA_INST_0[6].FA_INST_1[488].FA_  ( .A(A[3560]), .B(n536), .CI(
        C[3560]), .CO(C[3561]) );
  FA_4628 \FA_INST_0[6].FA_INST_1[489].FA_  ( .A(A[3561]), .B(n535), .CI(
        C[3561]), .CO(C[3562]) );
  FA_4627 \FA_INST_0[6].FA_INST_1[490].FA_  ( .A(A[3562]), .B(n534), .CI(
        C[3562]), .CO(C[3563]) );
  FA_4626 \FA_INST_0[6].FA_INST_1[491].FA_  ( .A(A[3563]), .B(n533), .CI(
        C[3563]), .CO(C[3564]) );
  FA_4625 \FA_INST_0[6].FA_INST_1[492].FA_  ( .A(A[3564]), .B(n532), .CI(
        C[3564]), .CO(C[3565]) );
  FA_4624 \FA_INST_0[6].FA_INST_1[493].FA_  ( .A(A[3565]), .B(n531), .CI(
        C[3565]), .CO(C[3566]) );
  FA_4623 \FA_INST_0[6].FA_INST_1[494].FA_  ( .A(A[3566]), .B(n530), .CI(
        C[3566]), .CO(C[3567]) );
  FA_4622 \FA_INST_0[6].FA_INST_1[495].FA_  ( .A(A[3567]), .B(n529), .CI(
        C[3567]), .CO(C[3568]) );
  FA_4621 \FA_INST_0[6].FA_INST_1[496].FA_  ( .A(A[3568]), .B(n528), .CI(
        C[3568]), .CO(C[3569]) );
  FA_4620 \FA_INST_0[6].FA_INST_1[497].FA_  ( .A(A[3569]), .B(n527), .CI(
        C[3569]), .CO(C[3570]) );
  FA_4619 \FA_INST_0[6].FA_INST_1[498].FA_  ( .A(A[3570]), .B(n526), .CI(
        C[3570]), .CO(C[3571]) );
  FA_4618 \FA_INST_0[6].FA_INST_1[499].FA_  ( .A(A[3571]), .B(n525), .CI(
        C[3571]), .CO(C[3572]) );
  FA_4617 \FA_INST_0[6].FA_INST_1[500].FA_  ( .A(A[3572]), .B(n524), .CI(
        C[3572]), .CO(C[3573]) );
  FA_4616 \FA_INST_0[6].FA_INST_1[501].FA_  ( .A(A[3573]), .B(n523), .CI(
        C[3573]), .CO(C[3574]) );
  FA_4615 \FA_INST_0[6].FA_INST_1[502].FA_  ( .A(A[3574]), .B(n522), .CI(
        C[3574]), .CO(C[3575]) );
  FA_4614 \FA_INST_0[6].FA_INST_1[503].FA_  ( .A(A[3575]), .B(n521), .CI(
        C[3575]), .CO(C[3576]) );
  FA_4613 \FA_INST_0[6].FA_INST_1[504].FA_  ( .A(A[3576]), .B(n520), .CI(
        C[3576]), .CO(C[3577]) );
  FA_4612 \FA_INST_0[6].FA_INST_1[505].FA_  ( .A(A[3577]), .B(n519), .CI(
        C[3577]), .CO(C[3578]) );
  FA_4611 \FA_INST_0[6].FA_INST_1[506].FA_  ( .A(A[3578]), .B(n518), .CI(
        C[3578]), .CO(C[3579]) );
  FA_4610 \FA_INST_0[6].FA_INST_1[507].FA_  ( .A(A[3579]), .B(n517), .CI(
        C[3579]), .CO(C[3580]) );
  FA_4609 \FA_INST_0[6].FA_INST_1[508].FA_  ( .A(A[3580]), .B(n516), .CI(
        C[3580]), .CO(C[3581]) );
  FA_4608 \FA_INST_0[6].FA_INST_1[509].FA_  ( .A(A[3581]), .B(n515), .CI(
        C[3581]), .CO(C[3582]) );
  FA_4607 \FA_INST_0[6].FA_INST_1[510].FA_  ( .A(A[3582]), .B(n514), .CI(
        C[3582]), .CO(C[3583]) );
  FA_4606 \FA_INST_0[6].FA_INST_1[511].FA_  ( .A(A[3583]), .B(n513), .CI(
        C[3583]), .CO(C[3584]) );
  FA_4605 \FA_INST_0[7].FA_INST_1[0].FA_  ( .A(A[3584]), .B(n512), .CI(C[3584]), .CO(C[3585]) );
  FA_4604 \FA_INST_0[7].FA_INST_1[1].FA_  ( .A(A[3585]), .B(n511), .CI(C[3585]), .CO(C[3586]) );
  FA_4603 \FA_INST_0[7].FA_INST_1[2].FA_  ( .A(A[3586]), .B(n510), .CI(C[3586]), .CO(C[3587]) );
  FA_4602 \FA_INST_0[7].FA_INST_1[3].FA_  ( .A(A[3587]), .B(n509), .CI(C[3587]), .CO(C[3588]) );
  FA_4601 \FA_INST_0[7].FA_INST_1[4].FA_  ( .A(A[3588]), .B(n508), .CI(C[3588]), .CO(C[3589]) );
  FA_4600 \FA_INST_0[7].FA_INST_1[5].FA_  ( .A(A[3589]), .B(n507), .CI(C[3589]), .CO(C[3590]) );
  FA_4599 \FA_INST_0[7].FA_INST_1[6].FA_  ( .A(A[3590]), .B(n506), .CI(C[3590]), .CO(C[3591]) );
  FA_4598 \FA_INST_0[7].FA_INST_1[7].FA_  ( .A(A[3591]), .B(n505), .CI(C[3591]), .CO(C[3592]) );
  FA_4597 \FA_INST_0[7].FA_INST_1[8].FA_  ( .A(A[3592]), .B(n504), .CI(C[3592]), .CO(C[3593]) );
  FA_4596 \FA_INST_0[7].FA_INST_1[9].FA_  ( .A(A[3593]), .B(n503), .CI(C[3593]), .CO(C[3594]) );
  FA_4595 \FA_INST_0[7].FA_INST_1[10].FA_  ( .A(A[3594]), .B(n502), .CI(
        C[3594]), .CO(C[3595]) );
  FA_4594 \FA_INST_0[7].FA_INST_1[11].FA_  ( .A(A[3595]), .B(n501), .CI(
        C[3595]), .CO(C[3596]) );
  FA_4593 \FA_INST_0[7].FA_INST_1[12].FA_  ( .A(A[3596]), .B(n500), .CI(
        C[3596]), .CO(C[3597]) );
  FA_4592 \FA_INST_0[7].FA_INST_1[13].FA_  ( .A(A[3597]), .B(n499), .CI(
        C[3597]), .CO(C[3598]) );
  FA_4591 \FA_INST_0[7].FA_INST_1[14].FA_  ( .A(A[3598]), .B(n498), .CI(
        C[3598]), .CO(C[3599]) );
  FA_4590 \FA_INST_0[7].FA_INST_1[15].FA_  ( .A(A[3599]), .B(n497), .CI(
        C[3599]), .CO(C[3600]) );
  FA_4589 \FA_INST_0[7].FA_INST_1[16].FA_  ( .A(A[3600]), .B(n496), .CI(
        C[3600]), .CO(C[3601]) );
  FA_4588 \FA_INST_0[7].FA_INST_1[17].FA_  ( .A(A[3601]), .B(n495), .CI(
        C[3601]), .CO(C[3602]) );
  FA_4587 \FA_INST_0[7].FA_INST_1[18].FA_  ( .A(A[3602]), .B(n494), .CI(
        C[3602]), .CO(C[3603]) );
  FA_4586 \FA_INST_0[7].FA_INST_1[19].FA_  ( .A(A[3603]), .B(n493), .CI(
        C[3603]), .CO(C[3604]) );
  FA_4585 \FA_INST_0[7].FA_INST_1[20].FA_  ( .A(A[3604]), .B(n492), .CI(
        C[3604]), .CO(C[3605]) );
  FA_4584 \FA_INST_0[7].FA_INST_1[21].FA_  ( .A(A[3605]), .B(n491), .CI(
        C[3605]), .CO(C[3606]) );
  FA_4583 \FA_INST_0[7].FA_INST_1[22].FA_  ( .A(A[3606]), .B(n490), .CI(
        C[3606]), .CO(C[3607]) );
  FA_4582 \FA_INST_0[7].FA_INST_1[23].FA_  ( .A(A[3607]), .B(n489), .CI(
        C[3607]), .CO(C[3608]) );
  FA_4581 \FA_INST_0[7].FA_INST_1[24].FA_  ( .A(A[3608]), .B(n488), .CI(
        C[3608]), .CO(C[3609]) );
  FA_4580 \FA_INST_0[7].FA_INST_1[25].FA_  ( .A(A[3609]), .B(n487), .CI(
        C[3609]), .CO(C[3610]) );
  FA_4579 \FA_INST_0[7].FA_INST_1[26].FA_  ( .A(A[3610]), .B(n486), .CI(
        C[3610]), .CO(C[3611]) );
  FA_4578 \FA_INST_0[7].FA_INST_1[27].FA_  ( .A(A[3611]), .B(n485), .CI(
        C[3611]), .CO(C[3612]) );
  FA_4577 \FA_INST_0[7].FA_INST_1[28].FA_  ( .A(A[3612]), .B(n484), .CI(
        C[3612]), .CO(C[3613]) );
  FA_4576 \FA_INST_0[7].FA_INST_1[29].FA_  ( .A(A[3613]), .B(n483), .CI(
        C[3613]), .CO(C[3614]) );
  FA_4575 \FA_INST_0[7].FA_INST_1[30].FA_  ( .A(A[3614]), .B(n482), .CI(
        C[3614]), .CO(C[3615]) );
  FA_4574 \FA_INST_0[7].FA_INST_1[31].FA_  ( .A(A[3615]), .B(n481), .CI(
        C[3615]), .CO(C[3616]) );
  FA_4573 \FA_INST_0[7].FA_INST_1[32].FA_  ( .A(A[3616]), .B(n480), .CI(
        C[3616]), .CO(C[3617]) );
  FA_4572 \FA_INST_0[7].FA_INST_1[33].FA_  ( .A(A[3617]), .B(n479), .CI(
        C[3617]), .CO(C[3618]) );
  FA_4571 \FA_INST_0[7].FA_INST_1[34].FA_  ( .A(A[3618]), .B(n478), .CI(
        C[3618]), .CO(C[3619]) );
  FA_4570 \FA_INST_0[7].FA_INST_1[35].FA_  ( .A(A[3619]), .B(n477), .CI(
        C[3619]), .CO(C[3620]) );
  FA_4569 \FA_INST_0[7].FA_INST_1[36].FA_  ( .A(A[3620]), .B(n476), .CI(
        C[3620]), .CO(C[3621]) );
  FA_4568 \FA_INST_0[7].FA_INST_1[37].FA_  ( .A(A[3621]), .B(n475), .CI(
        C[3621]), .CO(C[3622]) );
  FA_4567 \FA_INST_0[7].FA_INST_1[38].FA_  ( .A(A[3622]), .B(n474), .CI(
        C[3622]), .CO(C[3623]) );
  FA_4566 \FA_INST_0[7].FA_INST_1[39].FA_  ( .A(A[3623]), .B(n473), .CI(
        C[3623]), .CO(C[3624]) );
  FA_4565 \FA_INST_0[7].FA_INST_1[40].FA_  ( .A(A[3624]), .B(n472), .CI(
        C[3624]), .CO(C[3625]) );
  FA_4564 \FA_INST_0[7].FA_INST_1[41].FA_  ( .A(A[3625]), .B(n471), .CI(
        C[3625]), .CO(C[3626]) );
  FA_4563 \FA_INST_0[7].FA_INST_1[42].FA_  ( .A(A[3626]), .B(n470), .CI(
        C[3626]), .CO(C[3627]) );
  FA_4562 \FA_INST_0[7].FA_INST_1[43].FA_  ( .A(A[3627]), .B(n469), .CI(
        C[3627]), .CO(C[3628]) );
  FA_4561 \FA_INST_0[7].FA_INST_1[44].FA_  ( .A(A[3628]), .B(n468), .CI(
        C[3628]), .CO(C[3629]) );
  FA_4560 \FA_INST_0[7].FA_INST_1[45].FA_  ( .A(A[3629]), .B(n467), .CI(
        C[3629]), .CO(C[3630]) );
  FA_4559 \FA_INST_0[7].FA_INST_1[46].FA_  ( .A(A[3630]), .B(n466), .CI(
        C[3630]), .CO(C[3631]) );
  FA_4558 \FA_INST_0[7].FA_INST_1[47].FA_  ( .A(A[3631]), .B(n465), .CI(
        C[3631]), .CO(C[3632]) );
  FA_4557 \FA_INST_0[7].FA_INST_1[48].FA_  ( .A(A[3632]), .B(n464), .CI(
        C[3632]), .CO(C[3633]) );
  FA_4556 \FA_INST_0[7].FA_INST_1[49].FA_  ( .A(A[3633]), .B(n463), .CI(
        C[3633]), .CO(C[3634]) );
  FA_4555 \FA_INST_0[7].FA_INST_1[50].FA_  ( .A(A[3634]), .B(n462), .CI(
        C[3634]), .CO(C[3635]) );
  FA_4554 \FA_INST_0[7].FA_INST_1[51].FA_  ( .A(A[3635]), .B(n461), .CI(
        C[3635]), .CO(C[3636]) );
  FA_4553 \FA_INST_0[7].FA_INST_1[52].FA_  ( .A(A[3636]), .B(n460), .CI(
        C[3636]), .CO(C[3637]) );
  FA_4552 \FA_INST_0[7].FA_INST_1[53].FA_  ( .A(A[3637]), .B(n459), .CI(
        C[3637]), .CO(C[3638]) );
  FA_4551 \FA_INST_0[7].FA_INST_1[54].FA_  ( .A(A[3638]), .B(n458), .CI(
        C[3638]), .CO(C[3639]) );
  FA_4550 \FA_INST_0[7].FA_INST_1[55].FA_  ( .A(A[3639]), .B(n457), .CI(
        C[3639]), .CO(C[3640]) );
  FA_4549 \FA_INST_0[7].FA_INST_1[56].FA_  ( .A(A[3640]), .B(n456), .CI(
        C[3640]), .CO(C[3641]) );
  FA_4548 \FA_INST_0[7].FA_INST_1[57].FA_  ( .A(A[3641]), .B(n455), .CI(
        C[3641]), .CO(C[3642]) );
  FA_4547 \FA_INST_0[7].FA_INST_1[58].FA_  ( .A(A[3642]), .B(n454), .CI(
        C[3642]), .CO(C[3643]) );
  FA_4546 \FA_INST_0[7].FA_INST_1[59].FA_  ( .A(A[3643]), .B(n453), .CI(
        C[3643]), .CO(C[3644]) );
  FA_4545 \FA_INST_0[7].FA_INST_1[60].FA_  ( .A(A[3644]), .B(n452), .CI(
        C[3644]), .CO(C[3645]) );
  FA_4544 \FA_INST_0[7].FA_INST_1[61].FA_  ( .A(A[3645]), .B(n451), .CI(
        C[3645]), .CO(C[3646]) );
  FA_4543 \FA_INST_0[7].FA_INST_1[62].FA_  ( .A(A[3646]), .B(n450), .CI(
        C[3646]), .CO(C[3647]) );
  FA_4542 \FA_INST_0[7].FA_INST_1[63].FA_  ( .A(A[3647]), .B(n449), .CI(
        C[3647]), .CO(C[3648]) );
  FA_4541 \FA_INST_0[7].FA_INST_1[64].FA_  ( .A(A[3648]), .B(n448), .CI(
        C[3648]), .CO(C[3649]) );
  FA_4540 \FA_INST_0[7].FA_INST_1[65].FA_  ( .A(A[3649]), .B(n447), .CI(
        C[3649]), .CO(C[3650]) );
  FA_4539 \FA_INST_0[7].FA_INST_1[66].FA_  ( .A(A[3650]), .B(n446), .CI(
        C[3650]), .CO(C[3651]) );
  FA_4538 \FA_INST_0[7].FA_INST_1[67].FA_  ( .A(A[3651]), .B(n445), .CI(
        C[3651]), .CO(C[3652]) );
  FA_4537 \FA_INST_0[7].FA_INST_1[68].FA_  ( .A(A[3652]), .B(n444), .CI(
        C[3652]), .CO(C[3653]) );
  FA_4536 \FA_INST_0[7].FA_INST_1[69].FA_  ( .A(A[3653]), .B(n443), .CI(
        C[3653]), .CO(C[3654]) );
  FA_4535 \FA_INST_0[7].FA_INST_1[70].FA_  ( .A(A[3654]), .B(n442), .CI(
        C[3654]), .CO(C[3655]) );
  FA_4534 \FA_INST_0[7].FA_INST_1[71].FA_  ( .A(A[3655]), .B(n441), .CI(
        C[3655]), .CO(C[3656]) );
  FA_4533 \FA_INST_0[7].FA_INST_1[72].FA_  ( .A(A[3656]), .B(n440), .CI(
        C[3656]), .CO(C[3657]) );
  FA_4532 \FA_INST_0[7].FA_INST_1[73].FA_  ( .A(A[3657]), .B(n439), .CI(
        C[3657]), .CO(C[3658]) );
  FA_4531 \FA_INST_0[7].FA_INST_1[74].FA_  ( .A(A[3658]), .B(n438), .CI(
        C[3658]), .CO(C[3659]) );
  FA_4530 \FA_INST_0[7].FA_INST_1[75].FA_  ( .A(A[3659]), .B(n437), .CI(
        C[3659]), .CO(C[3660]) );
  FA_4529 \FA_INST_0[7].FA_INST_1[76].FA_  ( .A(A[3660]), .B(n436), .CI(
        C[3660]), .CO(C[3661]) );
  FA_4528 \FA_INST_0[7].FA_INST_1[77].FA_  ( .A(A[3661]), .B(n435), .CI(
        C[3661]), .CO(C[3662]) );
  FA_4527 \FA_INST_0[7].FA_INST_1[78].FA_  ( .A(A[3662]), .B(n434), .CI(
        C[3662]), .CO(C[3663]) );
  FA_4526 \FA_INST_0[7].FA_INST_1[79].FA_  ( .A(A[3663]), .B(n433), .CI(
        C[3663]), .CO(C[3664]) );
  FA_4525 \FA_INST_0[7].FA_INST_1[80].FA_  ( .A(A[3664]), .B(n432), .CI(
        C[3664]), .CO(C[3665]) );
  FA_4524 \FA_INST_0[7].FA_INST_1[81].FA_  ( .A(A[3665]), .B(n431), .CI(
        C[3665]), .CO(C[3666]) );
  FA_4523 \FA_INST_0[7].FA_INST_1[82].FA_  ( .A(A[3666]), .B(n430), .CI(
        C[3666]), .CO(C[3667]) );
  FA_4522 \FA_INST_0[7].FA_INST_1[83].FA_  ( .A(A[3667]), .B(n429), .CI(
        C[3667]), .CO(C[3668]) );
  FA_4521 \FA_INST_0[7].FA_INST_1[84].FA_  ( .A(A[3668]), .B(n428), .CI(
        C[3668]), .CO(C[3669]) );
  FA_4520 \FA_INST_0[7].FA_INST_1[85].FA_  ( .A(A[3669]), .B(n427), .CI(
        C[3669]), .CO(C[3670]) );
  FA_4519 \FA_INST_0[7].FA_INST_1[86].FA_  ( .A(A[3670]), .B(n426), .CI(
        C[3670]), .CO(C[3671]) );
  FA_4518 \FA_INST_0[7].FA_INST_1[87].FA_  ( .A(A[3671]), .B(n425), .CI(
        C[3671]), .CO(C[3672]) );
  FA_4517 \FA_INST_0[7].FA_INST_1[88].FA_  ( .A(A[3672]), .B(n424), .CI(
        C[3672]), .CO(C[3673]) );
  FA_4516 \FA_INST_0[7].FA_INST_1[89].FA_  ( .A(A[3673]), .B(n423), .CI(
        C[3673]), .CO(C[3674]) );
  FA_4515 \FA_INST_0[7].FA_INST_1[90].FA_  ( .A(A[3674]), .B(n422), .CI(
        C[3674]), .CO(C[3675]) );
  FA_4514 \FA_INST_0[7].FA_INST_1[91].FA_  ( .A(A[3675]), .B(n421), .CI(
        C[3675]), .CO(C[3676]) );
  FA_4513 \FA_INST_0[7].FA_INST_1[92].FA_  ( .A(A[3676]), .B(n420), .CI(
        C[3676]), .CO(C[3677]) );
  FA_4512 \FA_INST_0[7].FA_INST_1[93].FA_  ( .A(A[3677]), .B(n419), .CI(
        C[3677]), .CO(C[3678]) );
  FA_4511 \FA_INST_0[7].FA_INST_1[94].FA_  ( .A(A[3678]), .B(n418), .CI(
        C[3678]), .CO(C[3679]) );
  FA_4510 \FA_INST_0[7].FA_INST_1[95].FA_  ( .A(A[3679]), .B(n417), .CI(
        C[3679]), .CO(C[3680]) );
  FA_4509 \FA_INST_0[7].FA_INST_1[96].FA_  ( .A(A[3680]), .B(n416), .CI(
        C[3680]), .CO(C[3681]) );
  FA_4508 \FA_INST_0[7].FA_INST_1[97].FA_  ( .A(A[3681]), .B(n415), .CI(
        C[3681]), .CO(C[3682]) );
  FA_4507 \FA_INST_0[7].FA_INST_1[98].FA_  ( .A(A[3682]), .B(n414), .CI(
        C[3682]), .CO(C[3683]) );
  FA_4506 \FA_INST_0[7].FA_INST_1[99].FA_  ( .A(A[3683]), .B(n413), .CI(
        C[3683]), .CO(C[3684]) );
  FA_4505 \FA_INST_0[7].FA_INST_1[100].FA_  ( .A(A[3684]), .B(n412), .CI(
        C[3684]), .CO(C[3685]) );
  FA_4504 \FA_INST_0[7].FA_INST_1[101].FA_  ( .A(A[3685]), .B(n411), .CI(
        C[3685]), .CO(C[3686]) );
  FA_4503 \FA_INST_0[7].FA_INST_1[102].FA_  ( .A(A[3686]), .B(n410), .CI(
        C[3686]), .CO(C[3687]) );
  FA_4502 \FA_INST_0[7].FA_INST_1[103].FA_  ( .A(A[3687]), .B(n409), .CI(
        C[3687]), .CO(C[3688]) );
  FA_4501 \FA_INST_0[7].FA_INST_1[104].FA_  ( .A(A[3688]), .B(n408), .CI(
        C[3688]), .CO(C[3689]) );
  FA_4500 \FA_INST_0[7].FA_INST_1[105].FA_  ( .A(A[3689]), .B(n407), .CI(
        C[3689]), .CO(C[3690]) );
  FA_4499 \FA_INST_0[7].FA_INST_1[106].FA_  ( .A(A[3690]), .B(n406), .CI(
        C[3690]), .CO(C[3691]) );
  FA_4498 \FA_INST_0[7].FA_INST_1[107].FA_  ( .A(A[3691]), .B(n405), .CI(
        C[3691]), .CO(C[3692]) );
  FA_4497 \FA_INST_0[7].FA_INST_1[108].FA_  ( .A(A[3692]), .B(n404), .CI(
        C[3692]), .CO(C[3693]) );
  FA_4496 \FA_INST_0[7].FA_INST_1[109].FA_  ( .A(A[3693]), .B(n403), .CI(
        C[3693]), .CO(C[3694]) );
  FA_4495 \FA_INST_0[7].FA_INST_1[110].FA_  ( .A(A[3694]), .B(n402), .CI(
        C[3694]), .CO(C[3695]) );
  FA_4494 \FA_INST_0[7].FA_INST_1[111].FA_  ( .A(A[3695]), .B(n401), .CI(
        C[3695]), .CO(C[3696]) );
  FA_4493 \FA_INST_0[7].FA_INST_1[112].FA_  ( .A(A[3696]), .B(n400), .CI(
        C[3696]), .CO(C[3697]) );
  FA_4492 \FA_INST_0[7].FA_INST_1[113].FA_  ( .A(A[3697]), .B(n399), .CI(
        C[3697]), .CO(C[3698]) );
  FA_4491 \FA_INST_0[7].FA_INST_1[114].FA_  ( .A(A[3698]), .B(n398), .CI(
        C[3698]), .CO(C[3699]) );
  FA_4490 \FA_INST_0[7].FA_INST_1[115].FA_  ( .A(A[3699]), .B(n397), .CI(
        C[3699]), .CO(C[3700]) );
  FA_4489 \FA_INST_0[7].FA_INST_1[116].FA_  ( .A(A[3700]), .B(n396), .CI(
        C[3700]), .CO(C[3701]) );
  FA_4488 \FA_INST_0[7].FA_INST_1[117].FA_  ( .A(A[3701]), .B(n395), .CI(
        C[3701]), .CO(C[3702]) );
  FA_4487 \FA_INST_0[7].FA_INST_1[118].FA_  ( .A(A[3702]), .B(n394), .CI(
        C[3702]), .CO(C[3703]) );
  FA_4486 \FA_INST_0[7].FA_INST_1[119].FA_  ( .A(A[3703]), .B(n393), .CI(
        C[3703]), .CO(C[3704]) );
  FA_4485 \FA_INST_0[7].FA_INST_1[120].FA_  ( .A(A[3704]), .B(n392), .CI(
        C[3704]), .CO(C[3705]) );
  FA_4484 \FA_INST_0[7].FA_INST_1[121].FA_  ( .A(A[3705]), .B(n391), .CI(
        C[3705]), .CO(C[3706]) );
  FA_4483 \FA_INST_0[7].FA_INST_1[122].FA_  ( .A(A[3706]), .B(n390), .CI(
        C[3706]), .CO(C[3707]) );
  FA_4482 \FA_INST_0[7].FA_INST_1[123].FA_  ( .A(A[3707]), .B(n389), .CI(
        C[3707]), .CO(C[3708]) );
  FA_4481 \FA_INST_0[7].FA_INST_1[124].FA_  ( .A(A[3708]), .B(n388), .CI(
        C[3708]), .CO(C[3709]) );
  FA_4480 \FA_INST_0[7].FA_INST_1[125].FA_  ( .A(A[3709]), .B(n387), .CI(
        C[3709]), .CO(C[3710]) );
  FA_4479 \FA_INST_0[7].FA_INST_1[126].FA_  ( .A(A[3710]), .B(n386), .CI(
        C[3710]), .CO(C[3711]) );
  FA_4478 \FA_INST_0[7].FA_INST_1[127].FA_  ( .A(A[3711]), .B(n385), .CI(
        C[3711]), .CO(C[3712]) );
  FA_4477 \FA_INST_0[7].FA_INST_1[128].FA_  ( .A(A[3712]), .B(n384), .CI(
        C[3712]), .CO(C[3713]) );
  FA_4476 \FA_INST_0[7].FA_INST_1[129].FA_  ( .A(A[3713]), .B(n383), .CI(
        C[3713]), .CO(C[3714]) );
  FA_4475 \FA_INST_0[7].FA_INST_1[130].FA_  ( .A(A[3714]), .B(n382), .CI(
        C[3714]), .CO(C[3715]) );
  FA_4474 \FA_INST_0[7].FA_INST_1[131].FA_  ( .A(A[3715]), .B(n381), .CI(
        C[3715]), .CO(C[3716]) );
  FA_4473 \FA_INST_0[7].FA_INST_1[132].FA_  ( .A(A[3716]), .B(n380), .CI(
        C[3716]), .CO(C[3717]) );
  FA_4472 \FA_INST_0[7].FA_INST_1[133].FA_  ( .A(A[3717]), .B(n379), .CI(
        C[3717]), .CO(C[3718]) );
  FA_4471 \FA_INST_0[7].FA_INST_1[134].FA_  ( .A(A[3718]), .B(n378), .CI(
        C[3718]), .CO(C[3719]) );
  FA_4470 \FA_INST_0[7].FA_INST_1[135].FA_  ( .A(A[3719]), .B(n377), .CI(
        C[3719]), .CO(C[3720]) );
  FA_4469 \FA_INST_0[7].FA_INST_1[136].FA_  ( .A(A[3720]), .B(n376), .CI(
        C[3720]), .CO(C[3721]) );
  FA_4468 \FA_INST_0[7].FA_INST_1[137].FA_  ( .A(A[3721]), .B(n375), .CI(
        C[3721]), .CO(C[3722]) );
  FA_4467 \FA_INST_0[7].FA_INST_1[138].FA_  ( .A(A[3722]), .B(n374), .CI(
        C[3722]), .CO(C[3723]) );
  FA_4466 \FA_INST_0[7].FA_INST_1[139].FA_  ( .A(A[3723]), .B(n373), .CI(
        C[3723]), .CO(C[3724]) );
  FA_4465 \FA_INST_0[7].FA_INST_1[140].FA_  ( .A(A[3724]), .B(n372), .CI(
        C[3724]), .CO(C[3725]) );
  FA_4464 \FA_INST_0[7].FA_INST_1[141].FA_  ( .A(A[3725]), .B(n371), .CI(
        C[3725]), .CO(C[3726]) );
  FA_4463 \FA_INST_0[7].FA_INST_1[142].FA_  ( .A(A[3726]), .B(n370), .CI(
        C[3726]), .CO(C[3727]) );
  FA_4462 \FA_INST_0[7].FA_INST_1[143].FA_  ( .A(A[3727]), .B(n369), .CI(
        C[3727]), .CO(C[3728]) );
  FA_4461 \FA_INST_0[7].FA_INST_1[144].FA_  ( .A(A[3728]), .B(n368), .CI(
        C[3728]), .CO(C[3729]) );
  FA_4460 \FA_INST_0[7].FA_INST_1[145].FA_  ( .A(A[3729]), .B(n367), .CI(
        C[3729]), .CO(C[3730]) );
  FA_4459 \FA_INST_0[7].FA_INST_1[146].FA_  ( .A(A[3730]), .B(n366), .CI(
        C[3730]), .CO(C[3731]) );
  FA_4458 \FA_INST_0[7].FA_INST_1[147].FA_  ( .A(A[3731]), .B(n365), .CI(
        C[3731]), .CO(C[3732]) );
  FA_4457 \FA_INST_0[7].FA_INST_1[148].FA_  ( .A(A[3732]), .B(n364), .CI(
        C[3732]), .CO(C[3733]) );
  FA_4456 \FA_INST_0[7].FA_INST_1[149].FA_  ( .A(A[3733]), .B(n363), .CI(
        C[3733]), .CO(C[3734]) );
  FA_4455 \FA_INST_0[7].FA_INST_1[150].FA_  ( .A(A[3734]), .B(n362), .CI(
        C[3734]), .CO(C[3735]) );
  FA_4454 \FA_INST_0[7].FA_INST_1[151].FA_  ( .A(A[3735]), .B(n361), .CI(
        C[3735]), .CO(C[3736]) );
  FA_4453 \FA_INST_0[7].FA_INST_1[152].FA_  ( .A(A[3736]), .B(n360), .CI(
        C[3736]), .CO(C[3737]) );
  FA_4452 \FA_INST_0[7].FA_INST_1[153].FA_  ( .A(A[3737]), .B(n359), .CI(
        C[3737]), .CO(C[3738]) );
  FA_4451 \FA_INST_0[7].FA_INST_1[154].FA_  ( .A(A[3738]), .B(n358), .CI(
        C[3738]), .CO(C[3739]) );
  FA_4450 \FA_INST_0[7].FA_INST_1[155].FA_  ( .A(A[3739]), .B(n357), .CI(
        C[3739]), .CO(C[3740]) );
  FA_4449 \FA_INST_0[7].FA_INST_1[156].FA_  ( .A(A[3740]), .B(n356), .CI(
        C[3740]), .CO(C[3741]) );
  FA_4448 \FA_INST_0[7].FA_INST_1[157].FA_  ( .A(A[3741]), .B(n355), .CI(
        C[3741]), .CO(C[3742]) );
  FA_4447 \FA_INST_0[7].FA_INST_1[158].FA_  ( .A(A[3742]), .B(n354), .CI(
        C[3742]), .CO(C[3743]) );
  FA_4446 \FA_INST_0[7].FA_INST_1[159].FA_  ( .A(A[3743]), .B(n353), .CI(
        C[3743]), .CO(C[3744]) );
  FA_4445 \FA_INST_0[7].FA_INST_1[160].FA_  ( .A(A[3744]), .B(n352), .CI(
        C[3744]), .CO(C[3745]) );
  FA_4444 \FA_INST_0[7].FA_INST_1[161].FA_  ( .A(A[3745]), .B(n351), .CI(
        C[3745]), .CO(C[3746]) );
  FA_4443 \FA_INST_0[7].FA_INST_1[162].FA_  ( .A(A[3746]), .B(n350), .CI(
        C[3746]), .CO(C[3747]) );
  FA_4442 \FA_INST_0[7].FA_INST_1[163].FA_  ( .A(A[3747]), .B(n349), .CI(
        C[3747]), .CO(C[3748]) );
  FA_4441 \FA_INST_0[7].FA_INST_1[164].FA_  ( .A(A[3748]), .B(n348), .CI(
        C[3748]), .CO(C[3749]) );
  FA_4440 \FA_INST_0[7].FA_INST_1[165].FA_  ( .A(A[3749]), .B(n347), .CI(
        C[3749]), .CO(C[3750]) );
  FA_4439 \FA_INST_0[7].FA_INST_1[166].FA_  ( .A(A[3750]), .B(n346), .CI(
        C[3750]), .CO(C[3751]) );
  FA_4438 \FA_INST_0[7].FA_INST_1[167].FA_  ( .A(A[3751]), .B(n345), .CI(
        C[3751]), .CO(C[3752]) );
  FA_4437 \FA_INST_0[7].FA_INST_1[168].FA_  ( .A(A[3752]), .B(n344), .CI(
        C[3752]), .CO(C[3753]) );
  FA_4436 \FA_INST_0[7].FA_INST_1[169].FA_  ( .A(A[3753]), .B(n343), .CI(
        C[3753]), .CO(C[3754]) );
  FA_4435 \FA_INST_0[7].FA_INST_1[170].FA_  ( .A(A[3754]), .B(n342), .CI(
        C[3754]), .CO(C[3755]) );
  FA_4434 \FA_INST_0[7].FA_INST_1[171].FA_  ( .A(A[3755]), .B(n341), .CI(
        C[3755]), .CO(C[3756]) );
  FA_4433 \FA_INST_0[7].FA_INST_1[172].FA_  ( .A(A[3756]), .B(n340), .CI(
        C[3756]), .CO(C[3757]) );
  FA_4432 \FA_INST_0[7].FA_INST_1[173].FA_  ( .A(A[3757]), .B(n339), .CI(
        C[3757]), .CO(C[3758]) );
  FA_4431 \FA_INST_0[7].FA_INST_1[174].FA_  ( .A(A[3758]), .B(n338), .CI(
        C[3758]), .CO(C[3759]) );
  FA_4430 \FA_INST_0[7].FA_INST_1[175].FA_  ( .A(A[3759]), .B(n337), .CI(
        C[3759]), .CO(C[3760]) );
  FA_4429 \FA_INST_0[7].FA_INST_1[176].FA_  ( .A(A[3760]), .B(n336), .CI(
        C[3760]), .CO(C[3761]) );
  FA_4428 \FA_INST_0[7].FA_INST_1[177].FA_  ( .A(A[3761]), .B(n335), .CI(
        C[3761]), .CO(C[3762]) );
  FA_4427 \FA_INST_0[7].FA_INST_1[178].FA_  ( .A(A[3762]), .B(n334), .CI(
        C[3762]), .CO(C[3763]) );
  FA_4426 \FA_INST_0[7].FA_INST_1[179].FA_  ( .A(A[3763]), .B(n333), .CI(
        C[3763]), .CO(C[3764]) );
  FA_4425 \FA_INST_0[7].FA_INST_1[180].FA_  ( .A(A[3764]), .B(n332), .CI(
        C[3764]), .CO(C[3765]) );
  FA_4424 \FA_INST_0[7].FA_INST_1[181].FA_  ( .A(A[3765]), .B(n331), .CI(
        C[3765]), .CO(C[3766]) );
  FA_4423 \FA_INST_0[7].FA_INST_1[182].FA_  ( .A(A[3766]), .B(n330), .CI(
        C[3766]), .CO(C[3767]) );
  FA_4422 \FA_INST_0[7].FA_INST_1[183].FA_  ( .A(A[3767]), .B(n329), .CI(
        C[3767]), .CO(C[3768]) );
  FA_4421 \FA_INST_0[7].FA_INST_1[184].FA_  ( .A(A[3768]), .B(n328), .CI(
        C[3768]), .CO(C[3769]) );
  FA_4420 \FA_INST_0[7].FA_INST_1[185].FA_  ( .A(A[3769]), .B(n327), .CI(
        C[3769]), .CO(C[3770]) );
  FA_4419 \FA_INST_0[7].FA_INST_1[186].FA_  ( .A(A[3770]), .B(n326), .CI(
        C[3770]), .CO(C[3771]) );
  FA_4418 \FA_INST_0[7].FA_INST_1[187].FA_  ( .A(A[3771]), .B(n325), .CI(
        C[3771]), .CO(C[3772]) );
  FA_4417 \FA_INST_0[7].FA_INST_1[188].FA_  ( .A(A[3772]), .B(n324), .CI(
        C[3772]), .CO(C[3773]) );
  FA_4416 \FA_INST_0[7].FA_INST_1[189].FA_  ( .A(A[3773]), .B(n323), .CI(
        C[3773]), .CO(C[3774]) );
  FA_4415 \FA_INST_0[7].FA_INST_1[190].FA_  ( .A(A[3774]), .B(n322), .CI(
        C[3774]), .CO(C[3775]) );
  FA_4414 \FA_INST_0[7].FA_INST_1[191].FA_  ( .A(A[3775]), .B(n321), .CI(
        C[3775]), .CO(C[3776]) );
  FA_4413 \FA_INST_0[7].FA_INST_1[192].FA_  ( .A(A[3776]), .B(n320), .CI(
        C[3776]), .CO(C[3777]) );
  FA_4412 \FA_INST_0[7].FA_INST_1[193].FA_  ( .A(A[3777]), .B(n319), .CI(
        C[3777]), .CO(C[3778]) );
  FA_4411 \FA_INST_0[7].FA_INST_1[194].FA_  ( .A(A[3778]), .B(n318), .CI(
        C[3778]), .CO(C[3779]) );
  FA_4410 \FA_INST_0[7].FA_INST_1[195].FA_  ( .A(A[3779]), .B(n317), .CI(
        C[3779]), .CO(C[3780]) );
  FA_4409 \FA_INST_0[7].FA_INST_1[196].FA_  ( .A(A[3780]), .B(n316), .CI(
        C[3780]), .CO(C[3781]) );
  FA_4408 \FA_INST_0[7].FA_INST_1[197].FA_  ( .A(A[3781]), .B(n315), .CI(
        C[3781]), .CO(C[3782]) );
  FA_4407 \FA_INST_0[7].FA_INST_1[198].FA_  ( .A(A[3782]), .B(n314), .CI(
        C[3782]), .CO(C[3783]) );
  FA_4406 \FA_INST_0[7].FA_INST_1[199].FA_  ( .A(A[3783]), .B(n313), .CI(
        C[3783]), .CO(C[3784]) );
  FA_4405 \FA_INST_0[7].FA_INST_1[200].FA_  ( .A(A[3784]), .B(n312), .CI(
        C[3784]), .CO(C[3785]) );
  FA_4404 \FA_INST_0[7].FA_INST_1[201].FA_  ( .A(A[3785]), .B(n311), .CI(
        C[3785]), .CO(C[3786]) );
  FA_4403 \FA_INST_0[7].FA_INST_1[202].FA_  ( .A(A[3786]), .B(n310), .CI(
        C[3786]), .CO(C[3787]) );
  FA_4402 \FA_INST_0[7].FA_INST_1[203].FA_  ( .A(A[3787]), .B(n309), .CI(
        C[3787]), .CO(C[3788]) );
  FA_4401 \FA_INST_0[7].FA_INST_1[204].FA_  ( .A(A[3788]), .B(n308), .CI(
        C[3788]), .CO(C[3789]) );
  FA_4400 \FA_INST_0[7].FA_INST_1[205].FA_  ( .A(A[3789]), .B(n307), .CI(
        C[3789]), .CO(C[3790]) );
  FA_4399 \FA_INST_0[7].FA_INST_1[206].FA_  ( .A(A[3790]), .B(n306), .CI(
        C[3790]), .CO(C[3791]) );
  FA_4398 \FA_INST_0[7].FA_INST_1[207].FA_  ( .A(A[3791]), .B(n305), .CI(
        C[3791]), .CO(C[3792]) );
  FA_4397 \FA_INST_0[7].FA_INST_1[208].FA_  ( .A(A[3792]), .B(n304), .CI(
        C[3792]), .CO(C[3793]) );
  FA_4396 \FA_INST_0[7].FA_INST_1[209].FA_  ( .A(A[3793]), .B(n303), .CI(
        C[3793]), .CO(C[3794]) );
  FA_4395 \FA_INST_0[7].FA_INST_1[210].FA_  ( .A(A[3794]), .B(n302), .CI(
        C[3794]), .CO(C[3795]) );
  FA_4394 \FA_INST_0[7].FA_INST_1[211].FA_  ( .A(A[3795]), .B(n301), .CI(
        C[3795]), .CO(C[3796]) );
  FA_4393 \FA_INST_0[7].FA_INST_1[212].FA_  ( .A(A[3796]), .B(n300), .CI(
        C[3796]), .CO(C[3797]) );
  FA_4392 \FA_INST_0[7].FA_INST_1[213].FA_  ( .A(A[3797]), .B(n299), .CI(
        C[3797]), .CO(C[3798]) );
  FA_4391 \FA_INST_0[7].FA_INST_1[214].FA_  ( .A(A[3798]), .B(n298), .CI(
        C[3798]), .CO(C[3799]) );
  FA_4390 \FA_INST_0[7].FA_INST_1[215].FA_  ( .A(A[3799]), .B(n297), .CI(
        C[3799]), .CO(C[3800]) );
  FA_4389 \FA_INST_0[7].FA_INST_1[216].FA_  ( .A(A[3800]), .B(n296), .CI(
        C[3800]), .CO(C[3801]) );
  FA_4388 \FA_INST_0[7].FA_INST_1[217].FA_  ( .A(A[3801]), .B(n295), .CI(
        C[3801]), .CO(C[3802]) );
  FA_4387 \FA_INST_0[7].FA_INST_1[218].FA_  ( .A(A[3802]), .B(n294), .CI(
        C[3802]), .CO(C[3803]) );
  FA_4386 \FA_INST_0[7].FA_INST_1[219].FA_  ( .A(A[3803]), .B(n293), .CI(
        C[3803]), .CO(C[3804]) );
  FA_4385 \FA_INST_0[7].FA_INST_1[220].FA_  ( .A(A[3804]), .B(n292), .CI(
        C[3804]), .CO(C[3805]) );
  FA_4384 \FA_INST_0[7].FA_INST_1[221].FA_  ( .A(A[3805]), .B(n291), .CI(
        C[3805]), .CO(C[3806]) );
  FA_4383 \FA_INST_0[7].FA_INST_1[222].FA_  ( .A(A[3806]), .B(n290), .CI(
        C[3806]), .CO(C[3807]) );
  FA_4382 \FA_INST_0[7].FA_INST_1[223].FA_  ( .A(A[3807]), .B(n289), .CI(
        C[3807]), .CO(C[3808]) );
  FA_4381 \FA_INST_0[7].FA_INST_1[224].FA_  ( .A(A[3808]), .B(n288), .CI(
        C[3808]), .CO(C[3809]) );
  FA_4380 \FA_INST_0[7].FA_INST_1[225].FA_  ( .A(A[3809]), .B(n287), .CI(
        C[3809]), .CO(C[3810]) );
  FA_4379 \FA_INST_0[7].FA_INST_1[226].FA_  ( .A(A[3810]), .B(n286), .CI(
        C[3810]), .CO(C[3811]) );
  FA_4378 \FA_INST_0[7].FA_INST_1[227].FA_  ( .A(A[3811]), .B(n285), .CI(
        C[3811]), .CO(C[3812]) );
  FA_4377 \FA_INST_0[7].FA_INST_1[228].FA_  ( .A(A[3812]), .B(n284), .CI(
        C[3812]), .CO(C[3813]) );
  FA_4376 \FA_INST_0[7].FA_INST_1[229].FA_  ( .A(A[3813]), .B(n283), .CI(
        C[3813]), .CO(C[3814]) );
  FA_4375 \FA_INST_0[7].FA_INST_1[230].FA_  ( .A(A[3814]), .B(n282), .CI(
        C[3814]), .CO(C[3815]) );
  FA_4374 \FA_INST_0[7].FA_INST_1[231].FA_  ( .A(A[3815]), .B(n281), .CI(
        C[3815]), .CO(C[3816]) );
  FA_4373 \FA_INST_0[7].FA_INST_1[232].FA_  ( .A(A[3816]), .B(n280), .CI(
        C[3816]), .CO(C[3817]) );
  FA_4372 \FA_INST_0[7].FA_INST_1[233].FA_  ( .A(A[3817]), .B(n279), .CI(
        C[3817]), .CO(C[3818]) );
  FA_4371 \FA_INST_0[7].FA_INST_1[234].FA_  ( .A(A[3818]), .B(n278), .CI(
        C[3818]), .CO(C[3819]) );
  FA_4370 \FA_INST_0[7].FA_INST_1[235].FA_  ( .A(A[3819]), .B(n277), .CI(
        C[3819]), .CO(C[3820]) );
  FA_4369 \FA_INST_0[7].FA_INST_1[236].FA_  ( .A(A[3820]), .B(n276), .CI(
        C[3820]), .CO(C[3821]) );
  FA_4368 \FA_INST_0[7].FA_INST_1[237].FA_  ( .A(A[3821]), .B(n275), .CI(
        C[3821]), .CO(C[3822]) );
  FA_4367 \FA_INST_0[7].FA_INST_1[238].FA_  ( .A(A[3822]), .B(n274), .CI(
        C[3822]), .CO(C[3823]) );
  FA_4366 \FA_INST_0[7].FA_INST_1[239].FA_  ( .A(A[3823]), .B(n273), .CI(
        C[3823]), .CO(C[3824]) );
  FA_4365 \FA_INST_0[7].FA_INST_1[240].FA_  ( .A(A[3824]), .B(n272), .CI(
        C[3824]), .CO(C[3825]) );
  FA_4364 \FA_INST_0[7].FA_INST_1[241].FA_  ( .A(A[3825]), .B(n271), .CI(
        C[3825]), .CO(C[3826]) );
  FA_4363 \FA_INST_0[7].FA_INST_1[242].FA_  ( .A(A[3826]), .B(n270), .CI(
        C[3826]), .CO(C[3827]) );
  FA_4362 \FA_INST_0[7].FA_INST_1[243].FA_  ( .A(A[3827]), .B(n269), .CI(
        C[3827]), .CO(C[3828]) );
  FA_4361 \FA_INST_0[7].FA_INST_1[244].FA_  ( .A(A[3828]), .B(n268), .CI(
        C[3828]), .CO(C[3829]) );
  FA_4360 \FA_INST_0[7].FA_INST_1[245].FA_  ( .A(A[3829]), .B(n267), .CI(
        C[3829]), .CO(C[3830]) );
  FA_4359 \FA_INST_0[7].FA_INST_1[246].FA_  ( .A(A[3830]), .B(n266), .CI(
        C[3830]), .CO(C[3831]) );
  FA_4358 \FA_INST_0[7].FA_INST_1[247].FA_  ( .A(A[3831]), .B(n265), .CI(
        C[3831]), .CO(C[3832]) );
  FA_4357 \FA_INST_0[7].FA_INST_1[248].FA_  ( .A(A[3832]), .B(n264), .CI(
        C[3832]), .CO(C[3833]) );
  FA_4356 \FA_INST_0[7].FA_INST_1[249].FA_  ( .A(A[3833]), .B(n263), .CI(
        C[3833]), .CO(C[3834]) );
  FA_4355 \FA_INST_0[7].FA_INST_1[250].FA_  ( .A(A[3834]), .B(n262), .CI(
        C[3834]), .CO(C[3835]) );
  FA_4354 \FA_INST_0[7].FA_INST_1[251].FA_  ( .A(A[3835]), .B(n261), .CI(
        C[3835]), .CO(C[3836]) );
  FA_4353 \FA_INST_0[7].FA_INST_1[252].FA_  ( .A(A[3836]), .B(n260), .CI(
        C[3836]), .CO(C[3837]) );
  FA_4352 \FA_INST_0[7].FA_INST_1[253].FA_  ( .A(A[3837]), .B(n259), .CI(
        C[3837]), .CO(C[3838]) );
  FA_4351 \FA_INST_0[7].FA_INST_1[254].FA_  ( .A(A[3838]), .B(n258), .CI(
        C[3838]), .CO(C[3839]) );
  FA_4350 \FA_INST_0[7].FA_INST_1[255].FA_  ( .A(A[3839]), .B(n257), .CI(
        C[3839]), .CO(C[3840]) );
  FA_4349 \FA_INST_0[7].FA_INST_1[256].FA_  ( .A(A[3840]), .B(n256), .CI(
        C[3840]), .CO(C[3841]) );
  FA_4348 \FA_INST_0[7].FA_INST_1[257].FA_  ( .A(A[3841]), .B(n255), .CI(
        C[3841]), .CO(C[3842]) );
  FA_4347 \FA_INST_0[7].FA_INST_1[258].FA_  ( .A(A[3842]), .B(n254), .CI(
        C[3842]), .CO(C[3843]) );
  FA_4346 \FA_INST_0[7].FA_INST_1[259].FA_  ( .A(A[3843]), .B(n253), .CI(
        C[3843]), .CO(C[3844]) );
  FA_4345 \FA_INST_0[7].FA_INST_1[260].FA_  ( .A(A[3844]), .B(n252), .CI(
        C[3844]), .CO(C[3845]) );
  FA_4344 \FA_INST_0[7].FA_INST_1[261].FA_  ( .A(A[3845]), .B(n251), .CI(
        C[3845]), .CO(C[3846]) );
  FA_4343 \FA_INST_0[7].FA_INST_1[262].FA_  ( .A(A[3846]), .B(n250), .CI(
        C[3846]), .CO(C[3847]) );
  FA_4342 \FA_INST_0[7].FA_INST_1[263].FA_  ( .A(A[3847]), .B(n249), .CI(
        C[3847]), .CO(C[3848]) );
  FA_4341 \FA_INST_0[7].FA_INST_1[264].FA_  ( .A(A[3848]), .B(n248), .CI(
        C[3848]), .CO(C[3849]) );
  FA_4340 \FA_INST_0[7].FA_INST_1[265].FA_  ( .A(A[3849]), .B(n247), .CI(
        C[3849]), .CO(C[3850]) );
  FA_4339 \FA_INST_0[7].FA_INST_1[266].FA_  ( .A(A[3850]), .B(n246), .CI(
        C[3850]), .CO(C[3851]) );
  FA_4338 \FA_INST_0[7].FA_INST_1[267].FA_  ( .A(A[3851]), .B(n245), .CI(
        C[3851]), .CO(C[3852]) );
  FA_4337 \FA_INST_0[7].FA_INST_1[268].FA_  ( .A(A[3852]), .B(n244), .CI(
        C[3852]), .CO(C[3853]) );
  FA_4336 \FA_INST_0[7].FA_INST_1[269].FA_  ( .A(A[3853]), .B(n243), .CI(
        C[3853]), .CO(C[3854]) );
  FA_4335 \FA_INST_0[7].FA_INST_1[270].FA_  ( .A(A[3854]), .B(n242), .CI(
        C[3854]), .CO(C[3855]) );
  FA_4334 \FA_INST_0[7].FA_INST_1[271].FA_  ( .A(A[3855]), .B(n241), .CI(
        C[3855]), .CO(C[3856]) );
  FA_4333 \FA_INST_0[7].FA_INST_1[272].FA_  ( .A(A[3856]), .B(n240), .CI(
        C[3856]), .CO(C[3857]) );
  FA_4332 \FA_INST_0[7].FA_INST_1[273].FA_  ( .A(A[3857]), .B(n239), .CI(
        C[3857]), .CO(C[3858]) );
  FA_4331 \FA_INST_0[7].FA_INST_1[274].FA_  ( .A(A[3858]), .B(n238), .CI(
        C[3858]), .CO(C[3859]) );
  FA_4330 \FA_INST_0[7].FA_INST_1[275].FA_  ( .A(A[3859]), .B(n237), .CI(
        C[3859]), .CO(C[3860]) );
  FA_4329 \FA_INST_0[7].FA_INST_1[276].FA_  ( .A(A[3860]), .B(n236), .CI(
        C[3860]), .CO(C[3861]) );
  FA_4328 \FA_INST_0[7].FA_INST_1[277].FA_  ( .A(A[3861]), .B(n235), .CI(
        C[3861]), .CO(C[3862]) );
  FA_4327 \FA_INST_0[7].FA_INST_1[278].FA_  ( .A(A[3862]), .B(n234), .CI(
        C[3862]), .CO(C[3863]) );
  FA_4326 \FA_INST_0[7].FA_INST_1[279].FA_  ( .A(A[3863]), .B(n233), .CI(
        C[3863]), .CO(C[3864]) );
  FA_4325 \FA_INST_0[7].FA_INST_1[280].FA_  ( .A(A[3864]), .B(n232), .CI(
        C[3864]), .CO(C[3865]) );
  FA_4324 \FA_INST_0[7].FA_INST_1[281].FA_  ( .A(A[3865]), .B(n231), .CI(
        C[3865]), .CO(C[3866]) );
  FA_4323 \FA_INST_0[7].FA_INST_1[282].FA_  ( .A(A[3866]), .B(n230), .CI(
        C[3866]), .CO(C[3867]) );
  FA_4322 \FA_INST_0[7].FA_INST_1[283].FA_  ( .A(A[3867]), .B(n229), .CI(
        C[3867]), .CO(C[3868]) );
  FA_4321 \FA_INST_0[7].FA_INST_1[284].FA_  ( .A(A[3868]), .B(n228), .CI(
        C[3868]), .CO(C[3869]) );
  FA_4320 \FA_INST_0[7].FA_INST_1[285].FA_  ( .A(A[3869]), .B(n227), .CI(
        C[3869]), .CO(C[3870]) );
  FA_4319 \FA_INST_0[7].FA_INST_1[286].FA_  ( .A(A[3870]), .B(n226), .CI(
        C[3870]), .CO(C[3871]) );
  FA_4318 \FA_INST_0[7].FA_INST_1[287].FA_  ( .A(A[3871]), .B(n225), .CI(
        C[3871]), .CO(C[3872]) );
  FA_4317 \FA_INST_0[7].FA_INST_1[288].FA_  ( .A(A[3872]), .B(n224), .CI(
        C[3872]), .CO(C[3873]) );
  FA_4316 \FA_INST_0[7].FA_INST_1[289].FA_  ( .A(A[3873]), .B(n223), .CI(
        C[3873]), .CO(C[3874]) );
  FA_4315 \FA_INST_0[7].FA_INST_1[290].FA_  ( .A(A[3874]), .B(n222), .CI(
        C[3874]), .CO(C[3875]) );
  FA_4314 \FA_INST_0[7].FA_INST_1[291].FA_  ( .A(A[3875]), .B(n221), .CI(
        C[3875]), .CO(C[3876]) );
  FA_4313 \FA_INST_0[7].FA_INST_1[292].FA_  ( .A(A[3876]), .B(n220), .CI(
        C[3876]), .CO(C[3877]) );
  FA_4312 \FA_INST_0[7].FA_INST_1[293].FA_  ( .A(A[3877]), .B(n219), .CI(
        C[3877]), .CO(C[3878]) );
  FA_4311 \FA_INST_0[7].FA_INST_1[294].FA_  ( .A(A[3878]), .B(n218), .CI(
        C[3878]), .CO(C[3879]) );
  FA_4310 \FA_INST_0[7].FA_INST_1[295].FA_  ( .A(A[3879]), .B(n217), .CI(
        C[3879]), .CO(C[3880]) );
  FA_4309 \FA_INST_0[7].FA_INST_1[296].FA_  ( .A(A[3880]), .B(n216), .CI(
        C[3880]), .CO(C[3881]) );
  FA_4308 \FA_INST_0[7].FA_INST_1[297].FA_  ( .A(A[3881]), .B(n215), .CI(
        C[3881]), .CO(C[3882]) );
  FA_4307 \FA_INST_0[7].FA_INST_1[298].FA_  ( .A(A[3882]), .B(n214), .CI(
        C[3882]), .CO(C[3883]) );
  FA_4306 \FA_INST_0[7].FA_INST_1[299].FA_  ( .A(A[3883]), .B(n213), .CI(
        C[3883]), .CO(C[3884]) );
  FA_4305 \FA_INST_0[7].FA_INST_1[300].FA_  ( .A(A[3884]), .B(n212), .CI(
        C[3884]), .CO(C[3885]) );
  FA_4304 \FA_INST_0[7].FA_INST_1[301].FA_  ( .A(A[3885]), .B(n211), .CI(
        C[3885]), .CO(C[3886]) );
  FA_4303 \FA_INST_0[7].FA_INST_1[302].FA_  ( .A(A[3886]), .B(n210), .CI(
        C[3886]), .CO(C[3887]) );
  FA_4302 \FA_INST_0[7].FA_INST_1[303].FA_  ( .A(A[3887]), .B(n209), .CI(
        C[3887]), .CO(C[3888]) );
  FA_4301 \FA_INST_0[7].FA_INST_1[304].FA_  ( .A(A[3888]), .B(n208), .CI(
        C[3888]), .CO(C[3889]) );
  FA_4300 \FA_INST_0[7].FA_INST_1[305].FA_  ( .A(A[3889]), .B(n207), .CI(
        C[3889]), .CO(C[3890]) );
  FA_4299 \FA_INST_0[7].FA_INST_1[306].FA_  ( .A(A[3890]), .B(n206), .CI(
        C[3890]), .CO(C[3891]) );
  FA_4298 \FA_INST_0[7].FA_INST_1[307].FA_  ( .A(A[3891]), .B(n205), .CI(
        C[3891]), .CO(C[3892]) );
  FA_4297 \FA_INST_0[7].FA_INST_1[308].FA_  ( .A(A[3892]), .B(n204), .CI(
        C[3892]), .CO(C[3893]) );
  FA_4296 \FA_INST_0[7].FA_INST_1[309].FA_  ( .A(A[3893]), .B(n203), .CI(
        C[3893]), .CO(C[3894]) );
  FA_4295 \FA_INST_0[7].FA_INST_1[310].FA_  ( .A(A[3894]), .B(n202), .CI(
        C[3894]), .CO(C[3895]) );
  FA_4294 \FA_INST_0[7].FA_INST_1[311].FA_  ( .A(A[3895]), .B(n201), .CI(
        C[3895]), .CO(C[3896]) );
  FA_4293 \FA_INST_0[7].FA_INST_1[312].FA_  ( .A(A[3896]), .B(n200), .CI(
        C[3896]), .CO(C[3897]) );
  FA_4292 \FA_INST_0[7].FA_INST_1[313].FA_  ( .A(A[3897]), .B(n199), .CI(
        C[3897]), .CO(C[3898]) );
  FA_4291 \FA_INST_0[7].FA_INST_1[314].FA_  ( .A(A[3898]), .B(n198), .CI(
        C[3898]), .CO(C[3899]) );
  FA_4290 \FA_INST_0[7].FA_INST_1[315].FA_  ( .A(A[3899]), .B(n197), .CI(
        C[3899]), .CO(C[3900]) );
  FA_4289 \FA_INST_0[7].FA_INST_1[316].FA_  ( .A(A[3900]), .B(n196), .CI(
        C[3900]), .CO(C[3901]) );
  FA_4288 \FA_INST_0[7].FA_INST_1[317].FA_  ( .A(A[3901]), .B(n195), .CI(
        C[3901]), .CO(C[3902]) );
  FA_4287 \FA_INST_0[7].FA_INST_1[318].FA_  ( .A(A[3902]), .B(n194), .CI(
        C[3902]), .CO(C[3903]) );
  FA_4286 \FA_INST_0[7].FA_INST_1[319].FA_  ( .A(A[3903]), .B(n193), .CI(
        C[3903]), .CO(C[3904]) );
  FA_4285 \FA_INST_0[7].FA_INST_1[320].FA_  ( .A(A[3904]), .B(n192), .CI(
        C[3904]), .CO(C[3905]) );
  FA_4284 \FA_INST_0[7].FA_INST_1[321].FA_  ( .A(A[3905]), .B(n191), .CI(
        C[3905]), .CO(C[3906]) );
  FA_4283 \FA_INST_0[7].FA_INST_1[322].FA_  ( .A(A[3906]), .B(n190), .CI(
        C[3906]), .CO(C[3907]) );
  FA_4282 \FA_INST_0[7].FA_INST_1[323].FA_  ( .A(A[3907]), .B(n189), .CI(
        C[3907]), .CO(C[3908]) );
  FA_4281 \FA_INST_0[7].FA_INST_1[324].FA_  ( .A(A[3908]), .B(n188), .CI(
        C[3908]), .CO(C[3909]) );
  FA_4280 \FA_INST_0[7].FA_INST_1[325].FA_  ( .A(A[3909]), .B(n187), .CI(
        C[3909]), .CO(C[3910]) );
  FA_4279 \FA_INST_0[7].FA_INST_1[326].FA_  ( .A(A[3910]), .B(n186), .CI(
        C[3910]), .CO(C[3911]) );
  FA_4278 \FA_INST_0[7].FA_INST_1[327].FA_  ( .A(A[3911]), .B(n185), .CI(
        C[3911]), .CO(C[3912]) );
  FA_4277 \FA_INST_0[7].FA_INST_1[328].FA_  ( .A(A[3912]), .B(n184), .CI(
        C[3912]), .CO(C[3913]) );
  FA_4276 \FA_INST_0[7].FA_INST_1[329].FA_  ( .A(A[3913]), .B(n183), .CI(
        C[3913]), .CO(C[3914]) );
  FA_4275 \FA_INST_0[7].FA_INST_1[330].FA_  ( .A(A[3914]), .B(n182), .CI(
        C[3914]), .CO(C[3915]) );
  FA_4274 \FA_INST_0[7].FA_INST_1[331].FA_  ( .A(A[3915]), .B(n181), .CI(
        C[3915]), .CO(C[3916]) );
  FA_4273 \FA_INST_0[7].FA_INST_1[332].FA_  ( .A(A[3916]), .B(n180), .CI(
        C[3916]), .CO(C[3917]) );
  FA_4272 \FA_INST_0[7].FA_INST_1[333].FA_  ( .A(A[3917]), .B(n179), .CI(
        C[3917]), .CO(C[3918]) );
  FA_4271 \FA_INST_0[7].FA_INST_1[334].FA_  ( .A(A[3918]), .B(n178), .CI(
        C[3918]), .CO(C[3919]) );
  FA_4270 \FA_INST_0[7].FA_INST_1[335].FA_  ( .A(A[3919]), .B(n177), .CI(
        C[3919]), .CO(C[3920]) );
  FA_4269 \FA_INST_0[7].FA_INST_1[336].FA_  ( .A(A[3920]), .B(n176), .CI(
        C[3920]), .CO(C[3921]) );
  FA_4268 \FA_INST_0[7].FA_INST_1[337].FA_  ( .A(A[3921]), .B(n175), .CI(
        C[3921]), .CO(C[3922]) );
  FA_4267 \FA_INST_0[7].FA_INST_1[338].FA_  ( .A(A[3922]), .B(n174), .CI(
        C[3922]), .CO(C[3923]) );
  FA_4266 \FA_INST_0[7].FA_INST_1[339].FA_  ( .A(A[3923]), .B(n173), .CI(
        C[3923]), .CO(C[3924]) );
  FA_4265 \FA_INST_0[7].FA_INST_1[340].FA_  ( .A(A[3924]), .B(n172), .CI(
        C[3924]), .CO(C[3925]) );
  FA_4264 \FA_INST_0[7].FA_INST_1[341].FA_  ( .A(A[3925]), .B(n171), .CI(
        C[3925]), .CO(C[3926]) );
  FA_4263 \FA_INST_0[7].FA_INST_1[342].FA_  ( .A(A[3926]), .B(n170), .CI(
        C[3926]), .CO(C[3927]) );
  FA_4262 \FA_INST_0[7].FA_INST_1[343].FA_  ( .A(A[3927]), .B(n169), .CI(
        C[3927]), .CO(C[3928]) );
  FA_4261 \FA_INST_0[7].FA_INST_1[344].FA_  ( .A(A[3928]), .B(n168), .CI(
        C[3928]), .CO(C[3929]) );
  FA_4260 \FA_INST_0[7].FA_INST_1[345].FA_  ( .A(A[3929]), .B(n167), .CI(
        C[3929]), .CO(C[3930]) );
  FA_4259 \FA_INST_0[7].FA_INST_1[346].FA_  ( .A(A[3930]), .B(n166), .CI(
        C[3930]), .CO(C[3931]) );
  FA_4258 \FA_INST_0[7].FA_INST_1[347].FA_  ( .A(A[3931]), .B(n165), .CI(
        C[3931]), .CO(C[3932]) );
  FA_4257 \FA_INST_0[7].FA_INST_1[348].FA_  ( .A(A[3932]), .B(n164), .CI(
        C[3932]), .CO(C[3933]) );
  FA_4256 \FA_INST_0[7].FA_INST_1[349].FA_  ( .A(A[3933]), .B(n163), .CI(
        C[3933]), .CO(C[3934]) );
  FA_4255 \FA_INST_0[7].FA_INST_1[350].FA_  ( .A(A[3934]), .B(n162), .CI(
        C[3934]), .CO(C[3935]) );
  FA_4254 \FA_INST_0[7].FA_INST_1[351].FA_  ( .A(A[3935]), .B(n161), .CI(
        C[3935]), .CO(C[3936]) );
  FA_4253 \FA_INST_0[7].FA_INST_1[352].FA_  ( .A(A[3936]), .B(n160), .CI(
        C[3936]), .CO(C[3937]) );
  FA_4252 \FA_INST_0[7].FA_INST_1[353].FA_  ( .A(A[3937]), .B(n159), .CI(
        C[3937]), .CO(C[3938]) );
  FA_4251 \FA_INST_0[7].FA_INST_1[354].FA_  ( .A(A[3938]), .B(n158), .CI(
        C[3938]), .CO(C[3939]) );
  FA_4250 \FA_INST_0[7].FA_INST_1[355].FA_  ( .A(A[3939]), .B(n157), .CI(
        C[3939]), .CO(C[3940]) );
  FA_4249 \FA_INST_0[7].FA_INST_1[356].FA_  ( .A(A[3940]), .B(n156), .CI(
        C[3940]), .CO(C[3941]) );
  FA_4248 \FA_INST_0[7].FA_INST_1[357].FA_  ( .A(A[3941]), .B(n155), .CI(
        C[3941]), .CO(C[3942]) );
  FA_4247 \FA_INST_0[7].FA_INST_1[358].FA_  ( .A(A[3942]), .B(n154), .CI(
        C[3942]), .CO(C[3943]) );
  FA_4246 \FA_INST_0[7].FA_INST_1[359].FA_  ( .A(A[3943]), .B(n153), .CI(
        C[3943]), .CO(C[3944]) );
  FA_4245 \FA_INST_0[7].FA_INST_1[360].FA_  ( .A(A[3944]), .B(n152), .CI(
        C[3944]), .CO(C[3945]) );
  FA_4244 \FA_INST_0[7].FA_INST_1[361].FA_  ( .A(A[3945]), .B(n151), .CI(
        C[3945]), .CO(C[3946]) );
  FA_4243 \FA_INST_0[7].FA_INST_1[362].FA_  ( .A(A[3946]), .B(n150), .CI(
        C[3946]), .CO(C[3947]) );
  FA_4242 \FA_INST_0[7].FA_INST_1[363].FA_  ( .A(A[3947]), .B(n149), .CI(
        C[3947]), .CO(C[3948]) );
  FA_4241 \FA_INST_0[7].FA_INST_1[364].FA_  ( .A(A[3948]), .B(n148), .CI(
        C[3948]), .CO(C[3949]) );
  FA_4240 \FA_INST_0[7].FA_INST_1[365].FA_  ( .A(A[3949]), .B(n147), .CI(
        C[3949]), .CO(C[3950]) );
  FA_4239 \FA_INST_0[7].FA_INST_1[366].FA_  ( .A(A[3950]), .B(n146), .CI(
        C[3950]), .CO(C[3951]) );
  FA_4238 \FA_INST_0[7].FA_INST_1[367].FA_  ( .A(A[3951]), .B(n145), .CI(
        C[3951]), .CO(C[3952]) );
  FA_4237 \FA_INST_0[7].FA_INST_1[368].FA_  ( .A(A[3952]), .B(n144), .CI(
        C[3952]), .CO(C[3953]) );
  FA_4236 \FA_INST_0[7].FA_INST_1[369].FA_  ( .A(A[3953]), .B(n143), .CI(
        C[3953]), .CO(C[3954]) );
  FA_4235 \FA_INST_0[7].FA_INST_1[370].FA_  ( .A(A[3954]), .B(n142), .CI(
        C[3954]), .CO(C[3955]) );
  FA_4234 \FA_INST_0[7].FA_INST_1[371].FA_  ( .A(A[3955]), .B(n141), .CI(
        C[3955]), .CO(C[3956]) );
  FA_4233 \FA_INST_0[7].FA_INST_1[372].FA_  ( .A(A[3956]), .B(n140), .CI(
        C[3956]), .CO(C[3957]) );
  FA_4232 \FA_INST_0[7].FA_INST_1[373].FA_  ( .A(A[3957]), .B(n139), .CI(
        C[3957]), .CO(C[3958]) );
  FA_4231 \FA_INST_0[7].FA_INST_1[374].FA_  ( .A(A[3958]), .B(n138), .CI(
        C[3958]), .CO(C[3959]) );
  FA_4230 \FA_INST_0[7].FA_INST_1[375].FA_  ( .A(A[3959]), .B(n137), .CI(
        C[3959]), .CO(C[3960]) );
  FA_4229 \FA_INST_0[7].FA_INST_1[376].FA_  ( .A(A[3960]), .B(n136), .CI(
        C[3960]), .CO(C[3961]) );
  FA_4228 \FA_INST_0[7].FA_INST_1[377].FA_  ( .A(A[3961]), .B(n135), .CI(
        C[3961]), .CO(C[3962]) );
  FA_4227 \FA_INST_0[7].FA_INST_1[378].FA_  ( .A(A[3962]), .B(n134), .CI(
        C[3962]), .CO(C[3963]) );
  FA_4226 \FA_INST_0[7].FA_INST_1[379].FA_  ( .A(A[3963]), .B(n133), .CI(
        C[3963]), .CO(C[3964]) );
  FA_4225 \FA_INST_0[7].FA_INST_1[380].FA_  ( .A(A[3964]), .B(n132), .CI(
        C[3964]), .CO(C[3965]) );
  FA_4224 \FA_INST_0[7].FA_INST_1[381].FA_  ( .A(A[3965]), .B(n131), .CI(
        C[3965]), .CO(C[3966]) );
  FA_4223 \FA_INST_0[7].FA_INST_1[382].FA_  ( .A(A[3966]), .B(n130), .CI(
        C[3966]), .CO(C[3967]) );
  FA_4222 \FA_INST_0[7].FA_INST_1[383].FA_  ( .A(A[3967]), .B(n129), .CI(
        C[3967]), .CO(C[3968]) );
  FA_4221 \FA_INST_0[7].FA_INST_1[384].FA_  ( .A(A[3968]), .B(n128), .CI(
        C[3968]), .CO(C[3969]) );
  FA_4220 \FA_INST_0[7].FA_INST_1[385].FA_  ( .A(A[3969]), .B(n127), .CI(
        C[3969]), .CO(C[3970]) );
  FA_4219 \FA_INST_0[7].FA_INST_1[386].FA_  ( .A(A[3970]), .B(n126), .CI(
        C[3970]), .CO(C[3971]) );
  FA_4218 \FA_INST_0[7].FA_INST_1[387].FA_  ( .A(A[3971]), .B(n125), .CI(
        C[3971]), .CO(C[3972]) );
  FA_4217 \FA_INST_0[7].FA_INST_1[388].FA_  ( .A(A[3972]), .B(n124), .CI(
        C[3972]), .CO(C[3973]) );
  FA_4216 \FA_INST_0[7].FA_INST_1[389].FA_  ( .A(A[3973]), .B(n123), .CI(
        C[3973]), .CO(C[3974]) );
  FA_4215 \FA_INST_0[7].FA_INST_1[390].FA_  ( .A(A[3974]), .B(n122), .CI(
        C[3974]), .CO(C[3975]) );
  FA_4214 \FA_INST_0[7].FA_INST_1[391].FA_  ( .A(A[3975]), .B(n121), .CI(
        C[3975]), .CO(C[3976]) );
  FA_4213 \FA_INST_0[7].FA_INST_1[392].FA_  ( .A(A[3976]), .B(n120), .CI(
        C[3976]), .CO(C[3977]) );
  FA_4212 \FA_INST_0[7].FA_INST_1[393].FA_  ( .A(A[3977]), .B(n119), .CI(
        C[3977]), .CO(C[3978]) );
  FA_4211 \FA_INST_0[7].FA_INST_1[394].FA_  ( .A(A[3978]), .B(n118), .CI(
        C[3978]), .CO(C[3979]) );
  FA_4210 \FA_INST_0[7].FA_INST_1[395].FA_  ( .A(A[3979]), .B(n117), .CI(
        C[3979]), .CO(C[3980]) );
  FA_4209 \FA_INST_0[7].FA_INST_1[396].FA_  ( .A(A[3980]), .B(n116), .CI(
        C[3980]), .CO(C[3981]) );
  FA_4208 \FA_INST_0[7].FA_INST_1[397].FA_  ( .A(A[3981]), .B(n115), .CI(
        C[3981]), .CO(C[3982]) );
  FA_4207 \FA_INST_0[7].FA_INST_1[398].FA_  ( .A(A[3982]), .B(n114), .CI(
        C[3982]), .CO(C[3983]) );
  FA_4206 \FA_INST_0[7].FA_INST_1[399].FA_  ( .A(A[3983]), .B(n113), .CI(
        C[3983]), .CO(C[3984]) );
  FA_4205 \FA_INST_0[7].FA_INST_1[400].FA_  ( .A(A[3984]), .B(n112), .CI(
        C[3984]), .CO(C[3985]) );
  FA_4204 \FA_INST_0[7].FA_INST_1[401].FA_  ( .A(A[3985]), .B(n111), .CI(
        C[3985]), .CO(C[3986]) );
  FA_4203 \FA_INST_0[7].FA_INST_1[402].FA_  ( .A(A[3986]), .B(n110), .CI(
        C[3986]), .CO(C[3987]) );
  FA_4202 \FA_INST_0[7].FA_INST_1[403].FA_  ( .A(A[3987]), .B(n109), .CI(
        C[3987]), .CO(C[3988]) );
  FA_4201 \FA_INST_0[7].FA_INST_1[404].FA_  ( .A(A[3988]), .B(n108), .CI(
        C[3988]), .CO(C[3989]) );
  FA_4200 \FA_INST_0[7].FA_INST_1[405].FA_  ( .A(A[3989]), .B(n107), .CI(
        C[3989]), .CO(C[3990]) );
  FA_4199 \FA_INST_0[7].FA_INST_1[406].FA_  ( .A(A[3990]), .B(n106), .CI(
        C[3990]), .CO(C[3991]) );
  FA_4198 \FA_INST_0[7].FA_INST_1[407].FA_  ( .A(A[3991]), .B(n105), .CI(
        C[3991]), .CO(C[3992]) );
  FA_4197 \FA_INST_0[7].FA_INST_1[408].FA_  ( .A(A[3992]), .B(n104), .CI(
        C[3992]), .CO(C[3993]) );
  FA_4196 \FA_INST_0[7].FA_INST_1[409].FA_  ( .A(A[3993]), .B(n103), .CI(
        C[3993]), .CO(C[3994]) );
  FA_4195 \FA_INST_0[7].FA_INST_1[410].FA_  ( .A(A[3994]), .B(n102), .CI(
        C[3994]), .CO(C[3995]) );
  FA_4194 \FA_INST_0[7].FA_INST_1[411].FA_  ( .A(A[3995]), .B(n101), .CI(
        C[3995]), .CO(C[3996]) );
  FA_4193 \FA_INST_0[7].FA_INST_1[412].FA_  ( .A(A[3996]), .B(n100), .CI(
        C[3996]), .CO(C[3997]) );
  FA_4192 \FA_INST_0[7].FA_INST_1[413].FA_  ( .A(A[3997]), .B(n99), .CI(
        C[3997]), .CO(C[3998]) );
  FA_4191 \FA_INST_0[7].FA_INST_1[414].FA_  ( .A(A[3998]), .B(n98), .CI(
        C[3998]), .CO(C[3999]) );
  FA_4190 \FA_INST_0[7].FA_INST_1[415].FA_  ( .A(A[3999]), .B(n97), .CI(
        C[3999]), .CO(C[4000]) );
  FA_4189 \FA_INST_0[7].FA_INST_1[416].FA_  ( .A(A[4000]), .B(n96), .CI(
        C[4000]), .CO(C[4001]) );
  FA_4188 \FA_INST_0[7].FA_INST_1[417].FA_  ( .A(A[4001]), .B(n95), .CI(
        C[4001]), .CO(C[4002]) );
  FA_4187 \FA_INST_0[7].FA_INST_1[418].FA_  ( .A(A[4002]), .B(n94), .CI(
        C[4002]), .CO(C[4003]) );
  FA_4186 \FA_INST_0[7].FA_INST_1[419].FA_  ( .A(A[4003]), .B(n93), .CI(
        C[4003]), .CO(C[4004]) );
  FA_4185 \FA_INST_0[7].FA_INST_1[420].FA_  ( .A(A[4004]), .B(n92), .CI(
        C[4004]), .CO(C[4005]) );
  FA_4184 \FA_INST_0[7].FA_INST_1[421].FA_  ( .A(A[4005]), .B(n91), .CI(
        C[4005]), .CO(C[4006]) );
  FA_4183 \FA_INST_0[7].FA_INST_1[422].FA_  ( .A(A[4006]), .B(n90), .CI(
        C[4006]), .CO(C[4007]) );
  FA_4182 \FA_INST_0[7].FA_INST_1[423].FA_  ( .A(A[4007]), .B(n89), .CI(
        C[4007]), .CO(C[4008]) );
  FA_4181 \FA_INST_0[7].FA_INST_1[424].FA_  ( .A(A[4008]), .B(n88), .CI(
        C[4008]), .CO(C[4009]) );
  FA_4180 \FA_INST_0[7].FA_INST_1[425].FA_  ( .A(A[4009]), .B(n87), .CI(
        C[4009]), .CO(C[4010]) );
  FA_4179 \FA_INST_0[7].FA_INST_1[426].FA_  ( .A(A[4010]), .B(n86), .CI(
        C[4010]), .CO(C[4011]) );
  FA_4178 \FA_INST_0[7].FA_INST_1[427].FA_  ( .A(A[4011]), .B(n85), .CI(
        C[4011]), .CO(C[4012]) );
  FA_4177 \FA_INST_0[7].FA_INST_1[428].FA_  ( .A(A[4012]), .B(n84), .CI(
        C[4012]), .CO(C[4013]) );
  FA_4176 \FA_INST_0[7].FA_INST_1[429].FA_  ( .A(A[4013]), .B(n83), .CI(
        C[4013]), .CO(C[4014]) );
  FA_4175 \FA_INST_0[7].FA_INST_1[430].FA_  ( .A(A[4014]), .B(n82), .CI(
        C[4014]), .CO(C[4015]) );
  FA_4174 \FA_INST_0[7].FA_INST_1[431].FA_  ( .A(A[4015]), .B(n81), .CI(
        C[4015]), .CO(C[4016]) );
  FA_4173 \FA_INST_0[7].FA_INST_1[432].FA_  ( .A(A[4016]), .B(n80), .CI(
        C[4016]), .CO(C[4017]) );
  FA_4172 \FA_INST_0[7].FA_INST_1[433].FA_  ( .A(A[4017]), .B(n79), .CI(
        C[4017]), .CO(C[4018]) );
  FA_4171 \FA_INST_0[7].FA_INST_1[434].FA_  ( .A(A[4018]), .B(n78), .CI(
        C[4018]), .CO(C[4019]) );
  FA_4170 \FA_INST_0[7].FA_INST_1[435].FA_  ( .A(A[4019]), .B(n77), .CI(
        C[4019]), .CO(C[4020]) );
  FA_4169 \FA_INST_0[7].FA_INST_1[436].FA_  ( .A(A[4020]), .B(n76), .CI(
        C[4020]), .CO(C[4021]) );
  FA_4168 \FA_INST_0[7].FA_INST_1[437].FA_  ( .A(A[4021]), .B(n75), .CI(
        C[4021]), .CO(C[4022]) );
  FA_4167 \FA_INST_0[7].FA_INST_1[438].FA_  ( .A(A[4022]), .B(n74), .CI(
        C[4022]), .CO(C[4023]) );
  FA_4166 \FA_INST_0[7].FA_INST_1[439].FA_  ( .A(A[4023]), .B(n73), .CI(
        C[4023]), .CO(C[4024]) );
  FA_4165 \FA_INST_0[7].FA_INST_1[440].FA_  ( .A(A[4024]), .B(n72), .CI(
        C[4024]), .CO(C[4025]) );
  FA_4164 \FA_INST_0[7].FA_INST_1[441].FA_  ( .A(A[4025]), .B(n71), .CI(
        C[4025]), .CO(C[4026]) );
  FA_4163 \FA_INST_0[7].FA_INST_1[442].FA_  ( .A(A[4026]), .B(n70), .CI(
        C[4026]), .CO(C[4027]) );
  FA_4162 \FA_INST_0[7].FA_INST_1[443].FA_  ( .A(A[4027]), .B(n69), .CI(
        C[4027]), .CO(C[4028]) );
  FA_4161 \FA_INST_0[7].FA_INST_1[444].FA_  ( .A(A[4028]), .B(n68), .CI(
        C[4028]), .CO(C[4029]) );
  FA_4160 \FA_INST_0[7].FA_INST_1[445].FA_  ( .A(A[4029]), .B(n67), .CI(
        C[4029]), .CO(C[4030]) );
  FA_4159 \FA_INST_0[7].FA_INST_1[446].FA_  ( .A(A[4030]), .B(n66), .CI(
        C[4030]), .CO(C[4031]) );
  FA_4158 \FA_INST_0[7].FA_INST_1[447].FA_  ( .A(A[4031]), .B(n65), .CI(
        C[4031]), .CO(C[4032]) );
  FA_4157 \FA_INST_0[7].FA_INST_1[448].FA_  ( .A(A[4032]), .B(n64), .CI(
        C[4032]), .CO(C[4033]) );
  FA_4156 \FA_INST_0[7].FA_INST_1[449].FA_  ( .A(A[4033]), .B(n63), .CI(
        C[4033]), .CO(C[4034]) );
  FA_4155 \FA_INST_0[7].FA_INST_1[450].FA_  ( .A(A[4034]), .B(n62), .CI(
        C[4034]), .CO(C[4035]) );
  FA_4154 \FA_INST_0[7].FA_INST_1[451].FA_  ( .A(A[4035]), .B(n61), .CI(
        C[4035]), .CO(C[4036]) );
  FA_4153 \FA_INST_0[7].FA_INST_1[452].FA_  ( .A(A[4036]), .B(n60), .CI(
        C[4036]), .CO(C[4037]) );
  FA_4152 \FA_INST_0[7].FA_INST_1[453].FA_  ( .A(A[4037]), .B(n59), .CI(
        C[4037]), .CO(C[4038]) );
  FA_4151 \FA_INST_0[7].FA_INST_1[454].FA_  ( .A(A[4038]), .B(n58), .CI(
        C[4038]), .CO(C[4039]) );
  FA_4150 \FA_INST_0[7].FA_INST_1[455].FA_  ( .A(A[4039]), .B(n57), .CI(
        C[4039]), .CO(C[4040]) );
  FA_4149 \FA_INST_0[7].FA_INST_1[456].FA_  ( .A(A[4040]), .B(n56), .CI(
        C[4040]), .CO(C[4041]) );
  FA_4148 \FA_INST_0[7].FA_INST_1[457].FA_  ( .A(A[4041]), .B(n55), .CI(
        C[4041]), .CO(C[4042]) );
  FA_4147 \FA_INST_0[7].FA_INST_1[458].FA_  ( .A(A[4042]), .B(n54), .CI(
        C[4042]), .CO(C[4043]) );
  FA_4146 \FA_INST_0[7].FA_INST_1[459].FA_  ( .A(A[4043]), .B(n53), .CI(
        C[4043]), .CO(C[4044]) );
  FA_4145 \FA_INST_0[7].FA_INST_1[460].FA_  ( .A(A[4044]), .B(n52), .CI(
        C[4044]), .CO(C[4045]) );
  FA_4144 \FA_INST_0[7].FA_INST_1[461].FA_  ( .A(A[4045]), .B(n51), .CI(
        C[4045]), .CO(C[4046]) );
  FA_4143 \FA_INST_0[7].FA_INST_1[462].FA_  ( .A(A[4046]), .B(n50), .CI(
        C[4046]), .CO(C[4047]) );
  FA_4142 \FA_INST_0[7].FA_INST_1[463].FA_  ( .A(A[4047]), .B(n49), .CI(
        C[4047]), .CO(C[4048]) );
  FA_4141 \FA_INST_0[7].FA_INST_1[464].FA_  ( .A(A[4048]), .B(n48), .CI(
        C[4048]), .CO(C[4049]) );
  FA_4140 \FA_INST_0[7].FA_INST_1[465].FA_  ( .A(A[4049]), .B(n47), .CI(
        C[4049]), .CO(C[4050]) );
  FA_4139 \FA_INST_0[7].FA_INST_1[466].FA_  ( .A(A[4050]), .B(n46), .CI(
        C[4050]), .CO(C[4051]) );
  FA_4138 \FA_INST_0[7].FA_INST_1[467].FA_  ( .A(A[4051]), .B(n45), .CI(
        C[4051]), .CO(C[4052]) );
  FA_4137 \FA_INST_0[7].FA_INST_1[468].FA_  ( .A(A[4052]), .B(n44), .CI(
        C[4052]), .CO(C[4053]) );
  FA_4136 \FA_INST_0[7].FA_INST_1[469].FA_  ( .A(A[4053]), .B(n43), .CI(
        C[4053]), .CO(C[4054]) );
  FA_4135 \FA_INST_0[7].FA_INST_1[470].FA_  ( .A(A[4054]), .B(n42), .CI(
        C[4054]), .CO(C[4055]) );
  FA_4134 \FA_INST_0[7].FA_INST_1[471].FA_  ( .A(A[4055]), .B(n41), .CI(
        C[4055]), .CO(C[4056]) );
  FA_4133 \FA_INST_0[7].FA_INST_1[472].FA_  ( .A(A[4056]), .B(n40), .CI(
        C[4056]), .CO(C[4057]) );
  FA_4132 \FA_INST_0[7].FA_INST_1[473].FA_  ( .A(A[4057]), .B(n39), .CI(
        C[4057]), .CO(C[4058]) );
  FA_4131 \FA_INST_0[7].FA_INST_1[474].FA_  ( .A(A[4058]), .B(n38), .CI(
        C[4058]), .CO(C[4059]) );
  FA_4130 \FA_INST_0[7].FA_INST_1[475].FA_  ( .A(A[4059]), .B(n37), .CI(
        C[4059]), .CO(C[4060]) );
  FA_4129 \FA_INST_0[7].FA_INST_1[476].FA_  ( .A(A[4060]), .B(n36), .CI(
        C[4060]), .CO(C[4061]) );
  FA_4128 \FA_INST_0[7].FA_INST_1[477].FA_  ( .A(A[4061]), .B(n35), .CI(
        C[4061]), .CO(C[4062]) );
  FA_4127 \FA_INST_0[7].FA_INST_1[478].FA_  ( .A(A[4062]), .B(n34), .CI(
        C[4062]), .CO(C[4063]) );
  FA_4126 \FA_INST_0[7].FA_INST_1[479].FA_  ( .A(A[4063]), .B(n33), .CI(
        C[4063]), .CO(C[4064]) );
  FA_4125 \FA_INST_0[7].FA_INST_1[480].FA_  ( .A(A[4064]), .B(n32), .CI(
        C[4064]), .CO(C[4065]) );
  FA_4124 \FA_INST_0[7].FA_INST_1[481].FA_  ( .A(A[4065]), .B(n31), .CI(
        C[4065]), .CO(C[4066]) );
  FA_4123 \FA_INST_0[7].FA_INST_1[482].FA_  ( .A(A[4066]), .B(n30), .CI(
        C[4066]), .CO(C[4067]) );
  FA_4122 \FA_INST_0[7].FA_INST_1[483].FA_  ( .A(A[4067]), .B(n29), .CI(
        C[4067]), .CO(C[4068]) );
  FA_4121 \FA_INST_0[7].FA_INST_1[484].FA_  ( .A(A[4068]), .B(n28), .CI(
        C[4068]), .CO(C[4069]) );
  FA_4120 \FA_INST_0[7].FA_INST_1[485].FA_  ( .A(A[4069]), .B(n27), .CI(
        C[4069]), .CO(C[4070]) );
  FA_4119 \FA_INST_0[7].FA_INST_1[486].FA_  ( .A(A[4070]), .B(n26), .CI(
        C[4070]), .CO(C[4071]) );
  FA_4118 \FA_INST_0[7].FA_INST_1[487].FA_  ( .A(A[4071]), .B(n25), .CI(
        C[4071]), .CO(C[4072]) );
  FA_4117 \FA_INST_0[7].FA_INST_1[488].FA_  ( .A(A[4072]), .B(n24), .CI(
        C[4072]), .CO(C[4073]) );
  FA_4116 \FA_INST_0[7].FA_INST_1[489].FA_  ( .A(A[4073]), .B(n23), .CI(
        C[4073]), .CO(C[4074]) );
  FA_4115 \FA_INST_0[7].FA_INST_1[490].FA_  ( .A(A[4074]), .B(n22), .CI(
        C[4074]), .CO(C[4075]) );
  FA_4114 \FA_INST_0[7].FA_INST_1[491].FA_  ( .A(A[4075]), .B(n21), .CI(
        C[4075]), .CO(C[4076]) );
  FA_4113 \FA_INST_0[7].FA_INST_1[492].FA_  ( .A(A[4076]), .B(n20), .CI(
        C[4076]), .CO(C[4077]) );
  FA_4112 \FA_INST_0[7].FA_INST_1[493].FA_  ( .A(A[4077]), .B(n19), .CI(
        C[4077]), .CO(C[4078]) );
  FA_4111 \FA_INST_0[7].FA_INST_1[494].FA_  ( .A(A[4078]), .B(n18), .CI(
        C[4078]), .CO(C[4079]) );
  FA_4110 \FA_INST_0[7].FA_INST_1[495].FA_  ( .A(A[4079]), .B(n17), .CI(
        C[4079]), .CO(C[4080]) );
  FA_4109 \FA_INST_0[7].FA_INST_1[496].FA_  ( .A(A[4080]), .B(n16), .CI(
        C[4080]), .CO(C[4081]) );
  FA_4108 \FA_INST_0[7].FA_INST_1[497].FA_  ( .A(A[4081]), .B(n15), .CI(
        C[4081]), .CO(C[4082]) );
  FA_4107 \FA_INST_0[7].FA_INST_1[498].FA_  ( .A(A[4082]), .B(n14), .CI(
        C[4082]), .CO(C[4083]) );
  FA_4106 \FA_INST_0[7].FA_INST_1[499].FA_  ( .A(A[4083]), .B(n13), .CI(
        C[4083]), .CO(C[4084]) );
  FA_4105 \FA_INST_0[7].FA_INST_1[500].FA_  ( .A(A[4084]), .B(n12), .CI(
        C[4084]), .CO(C[4085]) );
  FA_4104 \FA_INST_0[7].FA_INST_1[501].FA_  ( .A(A[4085]), .B(n11), .CI(
        C[4085]), .CO(C[4086]) );
  FA_4103 \FA_INST_0[7].FA_INST_1[502].FA_  ( .A(A[4086]), .B(n10), .CI(
        C[4086]), .CO(C[4087]) );
  FA_4102 \FA_INST_0[7].FA_INST_1[503].FA_  ( .A(A[4087]), .B(n9), .CI(C[4087]), .CO(C[4088]) );
  FA_4101 \FA_INST_0[7].FA_INST_1[504].FA_  ( .A(A[4088]), .B(n8), .CI(C[4088]), .CO(C[4089]) );
  FA_4100 \FA_INST_0[7].FA_INST_1[505].FA_  ( .A(A[4089]), .B(n7), .CI(C[4089]), .CO(C[4090]) );
  FA_4099 \FA_INST_0[7].FA_INST_1[506].FA_  ( .A(A[4090]), .B(n6), .CI(C[4090]), .CO(C[4091]) );
  FA_4098 \FA_INST_0[7].FA_INST_1[507].FA_  ( .A(A[4091]), .B(n5), .CI(C[4091]), .CO(C[4092]) );
  FA_4097 \FA_INST_0[7].FA_INST_1[508].FA_  ( .A(A[4092]), .B(n4), .CI(C[4092]), .CO(C[4093]) );
  FA_4096 \FA_INST_0[7].FA_INST_1[509].FA_  ( .A(A[4093]), .B(n3), .CI(C[4093]), .CO(C[4094]) );
  FA_4095 \FA_INST_0[7].FA_INST_1[510].FA_  ( .A(A[4094]), .B(n2), .CI(C[4094]), .CO(C[4095]) );
  FA_4094 \FA_INST_0[7].FA_INST_1[511].FA_  ( .A(A[4095]), .B(n1), .CI(C[4095]), .CO(O) );
  IV U2 ( .A(B[3097]), .Z(n999) );
  IV U3 ( .A(B[3098]), .Z(n998) );
  IV U4 ( .A(B[3099]), .Z(n997) );
  IV U5 ( .A(B[3100]), .Z(n996) );
  IV U6 ( .A(B[3101]), .Z(n995) );
  IV U7 ( .A(B[3102]), .Z(n994) );
  IV U8 ( .A(B[3103]), .Z(n993) );
  IV U9 ( .A(B[3104]), .Z(n992) );
  IV U10 ( .A(B[3105]), .Z(n991) );
  IV U11 ( .A(B[3106]), .Z(n990) );
  IV U12 ( .A(B[3997]), .Z(n99) );
  IV U13 ( .A(B[3107]), .Z(n989) );
  IV U14 ( .A(B[3108]), .Z(n988) );
  IV U15 ( .A(B[3109]), .Z(n987) );
  IV U16 ( .A(B[3110]), .Z(n986) );
  IV U17 ( .A(B[3111]), .Z(n985) );
  IV U18 ( .A(B[3112]), .Z(n984) );
  IV U19 ( .A(B[3113]), .Z(n983) );
  IV U20 ( .A(B[3114]), .Z(n982) );
  IV U21 ( .A(B[3115]), .Z(n981) );
  IV U22 ( .A(B[3116]), .Z(n980) );
  IV U23 ( .A(B[3998]), .Z(n98) );
  IV U24 ( .A(B[3117]), .Z(n979) );
  IV U25 ( .A(B[3118]), .Z(n978) );
  IV U26 ( .A(B[3119]), .Z(n977) );
  IV U27 ( .A(B[3120]), .Z(n976) );
  IV U28 ( .A(B[3121]), .Z(n975) );
  IV U29 ( .A(B[3122]), .Z(n974) );
  IV U30 ( .A(B[3123]), .Z(n973) );
  IV U31 ( .A(B[3124]), .Z(n972) );
  IV U32 ( .A(B[3125]), .Z(n971) );
  IV U33 ( .A(B[3126]), .Z(n970) );
  IV U34 ( .A(B[3999]), .Z(n97) );
  IV U35 ( .A(B[3127]), .Z(n969) );
  IV U36 ( .A(B[3128]), .Z(n968) );
  IV U37 ( .A(B[3129]), .Z(n967) );
  IV U38 ( .A(B[3130]), .Z(n966) );
  IV U39 ( .A(B[3131]), .Z(n965) );
  IV U40 ( .A(B[3132]), .Z(n964) );
  IV U41 ( .A(B[3133]), .Z(n963) );
  IV U42 ( .A(B[3134]), .Z(n962) );
  IV U43 ( .A(B[3135]), .Z(n961) );
  IV U44 ( .A(B[3136]), .Z(n960) );
  IV U45 ( .A(B[4000]), .Z(n96) );
  IV U46 ( .A(B[3137]), .Z(n959) );
  IV U47 ( .A(B[3138]), .Z(n958) );
  IV U48 ( .A(B[3139]), .Z(n957) );
  IV U49 ( .A(B[3140]), .Z(n956) );
  IV U50 ( .A(B[3141]), .Z(n955) );
  IV U51 ( .A(B[3142]), .Z(n954) );
  IV U52 ( .A(B[3143]), .Z(n953) );
  IV U53 ( .A(B[3144]), .Z(n952) );
  IV U54 ( .A(B[3145]), .Z(n951) );
  IV U55 ( .A(B[3146]), .Z(n950) );
  IV U56 ( .A(B[4001]), .Z(n95) );
  IV U57 ( .A(B[3147]), .Z(n949) );
  IV U58 ( .A(B[3148]), .Z(n948) );
  IV U59 ( .A(B[3149]), .Z(n947) );
  IV U60 ( .A(B[3150]), .Z(n946) );
  IV U61 ( .A(B[3151]), .Z(n945) );
  IV U62 ( .A(B[3152]), .Z(n944) );
  IV U63 ( .A(B[3153]), .Z(n943) );
  IV U64 ( .A(B[3154]), .Z(n942) );
  IV U65 ( .A(B[3155]), .Z(n941) );
  IV U66 ( .A(B[3156]), .Z(n940) );
  IV U67 ( .A(B[4002]), .Z(n94) );
  IV U68 ( .A(B[3157]), .Z(n939) );
  IV U69 ( .A(B[3158]), .Z(n938) );
  IV U70 ( .A(B[3159]), .Z(n937) );
  IV U71 ( .A(B[3160]), .Z(n936) );
  IV U72 ( .A(B[3161]), .Z(n935) );
  IV U73 ( .A(B[3162]), .Z(n934) );
  IV U74 ( .A(B[3163]), .Z(n933) );
  IV U75 ( .A(B[3164]), .Z(n932) );
  IV U76 ( .A(B[3165]), .Z(n931) );
  IV U77 ( .A(B[3166]), .Z(n930) );
  IV U78 ( .A(B[4003]), .Z(n93) );
  IV U79 ( .A(B[3167]), .Z(n929) );
  IV U80 ( .A(B[3168]), .Z(n928) );
  IV U81 ( .A(B[3169]), .Z(n927) );
  IV U82 ( .A(B[3170]), .Z(n926) );
  IV U83 ( .A(B[3171]), .Z(n925) );
  IV U84 ( .A(B[3172]), .Z(n924) );
  IV U85 ( .A(B[3173]), .Z(n923) );
  IV U86 ( .A(B[3174]), .Z(n922) );
  IV U87 ( .A(B[3175]), .Z(n921) );
  IV U88 ( .A(B[3176]), .Z(n920) );
  IV U89 ( .A(B[4004]), .Z(n92) );
  IV U90 ( .A(B[3177]), .Z(n919) );
  IV U91 ( .A(B[3178]), .Z(n918) );
  IV U92 ( .A(B[3179]), .Z(n917) );
  IV U93 ( .A(B[3180]), .Z(n916) );
  IV U94 ( .A(B[3181]), .Z(n915) );
  IV U95 ( .A(B[3182]), .Z(n914) );
  IV U96 ( .A(B[3183]), .Z(n913) );
  IV U97 ( .A(B[3184]), .Z(n912) );
  IV U98 ( .A(B[3185]), .Z(n911) );
  IV U99 ( .A(B[3186]), .Z(n910) );
  IV U100 ( .A(B[4005]), .Z(n91) );
  IV U101 ( .A(B[3187]), .Z(n909) );
  IV U102 ( .A(B[3188]), .Z(n908) );
  IV U103 ( .A(B[3189]), .Z(n907) );
  IV U104 ( .A(B[3190]), .Z(n906) );
  IV U105 ( .A(B[3191]), .Z(n905) );
  IV U106 ( .A(B[3192]), .Z(n904) );
  IV U107 ( .A(B[3193]), .Z(n903) );
  IV U108 ( .A(B[3194]), .Z(n902) );
  IV U109 ( .A(B[3195]), .Z(n901) );
  IV U110 ( .A(B[3196]), .Z(n900) );
  IV U111 ( .A(B[4006]), .Z(n90) );
  IV U112 ( .A(B[4087]), .Z(n9) );
  IV U113 ( .A(B[3197]), .Z(n899) );
  IV U114 ( .A(B[3198]), .Z(n898) );
  IV U115 ( .A(B[3199]), .Z(n897) );
  IV U116 ( .A(B[3200]), .Z(n896) );
  IV U117 ( .A(B[3201]), .Z(n895) );
  IV U118 ( .A(B[3202]), .Z(n894) );
  IV U119 ( .A(B[3203]), .Z(n893) );
  IV U120 ( .A(B[3204]), .Z(n892) );
  IV U121 ( .A(B[3205]), .Z(n891) );
  IV U122 ( .A(B[3206]), .Z(n890) );
  IV U123 ( .A(B[4007]), .Z(n89) );
  IV U124 ( .A(B[3207]), .Z(n889) );
  IV U125 ( .A(B[3208]), .Z(n888) );
  IV U126 ( .A(B[3209]), .Z(n887) );
  IV U127 ( .A(B[3210]), .Z(n886) );
  IV U128 ( .A(B[3211]), .Z(n885) );
  IV U129 ( .A(B[3212]), .Z(n884) );
  IV U130 ( .A(B[3213]), .Z(n883) );
  IV U131 ( .A(B[3214]), .Z(n882) );
  IV U132 ( .A(B[3215]), .Z(n881) );
  IV U133 ( .A(B[3216]), .Z(n880) );
  IV U134 ( .A(B[4008]), .Z(n88) );
  IV U135 ( .A(B[3217]), .Z(n879) );
  IV U136 ( .A(B[3218]), .Z(n878) );
  IV U137 ( .A(B[3219]), .Z(n877) );
  IV U138 ( .A(B[3220]), .Z(n876) );
  IV U139 ( .A(B[3221]), .Z(n875) );
  IV U140 ( .A(B[3222]), .Z(n874) );
  IV U141 ( .A(B[3223]), .Z(n873) );
  IV U142 ( .A(B[3224]), .Z(n872) );
  IV U143 ( .A(B[3225]), .Z(n871) );
  IV U144 ( .A(B[3226]), .Z(n870) );
  IV U145 ( .A(B[4009]), .Z(n87) );
  IV U146 ( .A(B[3227]), .Z(n869) );
  IV U147 ( .A(B[3228]), .Z(n868) );
  IV U148 ( .A(B[3229]), .Z(n867) );
  IV U149 ( .A(B[3230]), .Z(n866) );
  IV U150 ( .A(B[3231]), .Z(n865) );
  IV U151 ( .A(B[3232]), .Z(n864) );
  IV U152 ( .A(B[3233]), .Z(n863) );
  IV U153 ( .A(B[3234]), .Z(n862) );
  IV U154 ( .A(B[3235]), .Z(n861) );
  IV U155 ( .A(B[3236]), .Z(n860) );
  IV U156 ( .A(B[4010]), .Z(n86) );
  IV U157 ( .A(B[3237]), .Z(n859) );
  IV U158 ( .A(B[3238]), .Z(n858) );
  IV U159 ( .A(B[3239]), .Z(n857) );
  IV U160 ( .A(B[3240]), .Z(n856) );
  IV U161 ( .A(B[3241]), .Z(n855) );
  IV U162 ( .A(B[3242]), .Z(n854) );
  IV U163 ( .A(B[3243]), .Z(n853) );
  IV U164 ( .A(B[3244]), .Z(n852) );
  IV U165 ( .A(B[3245]), .Z(n851) );
  IV U166 ( .A(B[3246]), .Z(n850) );
  IV U167 ( .A(B[4011]), .Z(n85) );
  IV U168 ( .A(B[3247]), .Z(n849) );
  IV U169 ( .A(B[3248]), .Z(n848) );
  IV U170 ( .A(B[3249]), .Z(n847) );
  IV U171 ( .A(B[3250]), .Z(n846) );
  IV U172 ( .A(B[3251]), .Z(n845) );
  IV U173 ( .A(B[3252]), .Z(n844) );
  IV U174 ( .A(B[3253]), .Z(n843) );
  IV U175 ( .A(B[3254]), .Z(n842) );
  IV U176 ( .A(B[3255]), .Z(n841) );
  IV U177 ( .A(B[3256]), .Z(n840) );
  IV U178 ( .A(B[4012]), .Z(n84) );
  IV U179 ( .A(B[3257]), .Z(n839) );
  IV U180 ( .A(B[3258]), .Z(n838) );
  IV U181 ( .A(B[3259]), .Z(n837) );
  IV U182 ( .A(B[3260]), .Z(n836) );
  IV U183 ( .A(B[3261]), .Z(n835) );
  IV U184 ( .A(B[3262]), .Z(n834) );
  IV U185 ( .A(B[3263]), .Z(n833) );
  IV U186 ( .A(B[3264]), .Z(n832) );
  IV U187 ( .A(B[3265]), .Z(n831) );
  IV U188 ( .A(B[3266]), .Z(n830) );
  IV U189 ( .A(B[4013]), .Z(n83) );
  IV U190 ( .A(B[3267]), .Z(n829) );
  IV U191 ( .A(B[3268]), .Z(n828) );
  IV U192 ( .A(B[3269]), .Z(n827) );
  IV U193 ( .A(B[3270]), .Z(n826) );
  IV U194 ( .A(B[3271]), .Z(n825) );
  IV U195 ( .A(B[3272]), .Z(n824) );
  IV U196 ( .A(B[3273]), .Z(n823) );
  IV U197 ( .A(B[3274]), .Z(n822) );
  IV U198 ( .A(B[3275]), .Z(n821) );
  IV U199 ( .A(B[3276]), .Z(n820) );
  IV U200 ( .A(B[4014]), .Z(n82) );
  IV U201 ( .A(B[3277]), .Z(n819) );
  IV U202 ( .A(B[3278]), .Z(n818) );
  IV U203 ( .A(B[3279]), .Z(n817) );
  IV U204 ( .A(B[3280]), .Z(n816) );
  IV U205 ( .A(B[3281]), .Z(n815) );
  IV U206 ( .A(B[3282]), .Z(n814) );
  IV U207 ( .A(B[3283]), .Z(n813) );
  IV U208 ( .A(B[3284]), .Z(n812) );
  IV U209 ( .A(B[3285]), .Z(n811) );
  IV U210 ( .A(B[3286]), .Z(n810) );
  IV U211 ( .A(B[4015]), .Z(n81) );
  IV U212 ( .A(B[3287]), .Z(n809) );
  IV U213 ( .A(B[3288]), .Z(n808) );
  IV U214 ( .A(B[3289]), .Z(n807) );
  IV U215 ( .A(B[3290]), .Z(n806) );
  IV U216 ( .A(B[3291]), .Z(n805) );
  IV U217 ( .A(B[3292]), .Z(n804) );
  IV U218 ( .A(B[3293]), .Z(n803) );
  IV U219 ( .A(B[3294]), .Z(n802) );
  IV U220 ( .A(B[3295]), .Z(n801) );
  IV U221 ( .A(B[3296]), .Z(n800) );
  IV U222 ( .A(B[4016]), .Z(n80) );
  IV U223 ( .A(B[4088]), .Z(n8) );
  IV U224 ( .A(B[3297]), .Z(n799) );
  IV U225 ( .A(B[3298]), .Z(n798) );
  IV U226 ( .A(B[3299]), .Z(n797) );
  IV U227 ( .A(B[3300]), .Z(n796) );
  IV U228 ( .A(B[3301]), .Z(n795) );
  IV U229 ( .A(B[3302]), .Z(n794) );
  IV U230 ( .A(B[3303]), .Z(n793) );
  IV U231 ( .A(B[3304]), .Z(n792) );
  IV U232 ( .A(B[3305]), .Z(n791) );
  IV U233 ( .A(B[3306]), .Z(n790) );
  IV U234 ( .A(B[4017]), .Z(n79) );
  IV U235 ( .A(B[3307]), .Z(n789) );
  IV U236 ( .A(B[3308]), .Z(n788) );
  IV U237 ( .A(B[3309]), .Z(n787) );
  IV U238 ( .A(B[3310]), .Z(n786) );
  IV U239 ( .A(B[3311]), .Z(n785) );
  IV U240 ( .A(B[3312]), .Z(n784) );
  IV U241 ( .A(B[3313]), .Z(n783) );
  IV U242 ( .A(B[3314]), .Z(n782) );
  IV U243 ( .A(B[3315]), .Z(n781) );
  IV U244 ( .A(B[3316]), .Z(n780) );
  IV U245 ( .A(B[4018]), .Z(n78) );
  IV U246 ( .A(B[3317]), .Z(n779) );
  IV U247 ( .A(B[3318]), .Z(n778) );
  IV U248 ( .A(B[3319]), .Z(n777) );
  IV U249 ( .A(B[3320]), .Z(n776) );
  IV U250 ( .A(B[3321]), .Z(n775) );
  IV U251 ( .A(B[3322]), .Z(n774) );
  IV U252 ( .A(B[3323]), .Z(n773) );
  IV U253 ( .A(B[3324]), .Z(n772) );
  IV U254 ( .A(B[3325]), .Z(n771) );
  IV U255 ( .A(B[3326]), .Z(n770) );
  IV U256 ( .A(B[4019]), .Z(n77) );
  IV U257 ( .A(B[3327]), .Z(n769) );
  IV U258 ( .A(B[3328]), .Z(n768) );
  IV U259 ( .A(B[3329]), .Z(n767) );
  IV U260 ( .A(B[3330]), .Z(n766) );
  IV U261 ( .A(B[3331]), .Z(n765) );
  IV U262 ( .A(B[3332]), .Z(n764) );
  IV U263 ( .A(B[3333]), .Z(n763) );
  IV U264 ( .A(B[3334]), .Z(n762) );
  IV U265 ( .A(B[3335]), .Z(n761) );
  IV U266 ( .A(B[3336]), .Z(n760) );
  IV U267 ( .A(B[4020]), .Z(n76) );
  IV U268 ( .A(B[3337]), .Z(n759) );
  IV U269 ( .A(B[3338]), .Z(n758) );
  IV U270 ( .A(B[3339]), .Z(n757) );
  IV U271 ( .A(B[3340]), .Z(n756) );
  IV U272 ( .A(B[3341]), .Z(n755) );
  IV U273 ( .A(B[3342]), .Z(n754) );
  IV U274 ( .A(B[3343]), .Z(n753) );
  IV U275 ( .A(B[3344]), .Z(n752) );
  IV U276 ( .A(B[3345]), .Z(n751) );
  IV U277 ( .A(B[3346]), .Z(n750) );
  IV U278 ( .A(B[4021]), .Z(n75) );
  IV U279 ( .A(B[3347]), .Z(n749) );
  IV U280 ( .A(B[3348]), .Z(n748) );
  IV U281 ( .A(B[3349]), .Z(n747) );
  IV U282 ( .A(B[3350]), .Z(n746) );
  IV U283 ( .A(B[3351]), .Z(n745) );
  IV U284 ( .A(B[3352]), .Z(n744) );
  IV U285 ( .A(B[3353]), .Z(n743) );
  IV U286 ( .A(B[3354]), .Z(n742) );
  IV U287 ( .A(B[3355]), .Z(n741) );
  IV U288 ( .A(B[3356]), .Z(n740) );
  IV U289 ( .A(B[4022]), .Z(n74) );
  IV U290 ( .A(B[3357]), .Z(n739) );
  IV U291 ( .A(B[3358]), .Z(n738) );
  IV U292 ( .A(B[3359]), .Z(n737) );
  IV U293 ( .A(B[3360]), .Z(n736) );
  IV U294 ( .A(B[3361]), .Z(n735) );
  IV U295 ( .A(B[3362]), .Z(n734) );
  IV U296 ( .A(B[3363]), .Z(n733) );
  IV U297 ( .A(B[3364]), .Z(n732) );
  IV U298 ( .A(B[3365]), .Z(n731) );
  IV U299 ( .A(B[3366]), .Z(n730) );
  IV U300 ( .A(B[4023]), .Z(n73) );
  IV U301 ( .A(B[3367]), .Z(n729) );
  IV U302 ( .A(B[3368]), .Z(n728) );
  IV U303 ( .A(B[3369]), .Z(n727) );
  IV U304 ( .A(B[3370]), .Z(n726) );
  IV U305 ( .A(B[3371]), .Z(n725) );
  IV U306 ( .A(B[3372]), .Z(n724) );
  IV U307 ( .A(B[3373]), .Z(n723) );
  IV U308 ( .A(B[3374]), .Z(n722) );
  IV U309 ( .A(B[3375]), .Z(n721) );
  IV U310 ( .A(B[3376]), .Z(n720) );
  IV U311 ( .A(B[4024]), .Z(n72) );
  IV U312 ( .A(B[3377]), .Z(n719) );
  IV U313 ( .A(B[3378]), .Z(n718) );
  IV U314 ( .A(B[3379]), .Z(n717) );
  IV U315 ( .A(B[3380]), .Z(n716) );
  IV U316 ( .A(B[3381]), .Z(n715) );
  IV U317 ( .A(B[3382]), .Z(n714) );
  IV U318 ( .A(B[3383]), .Z(n713) );
  IV U319 ( .A(B[3384]), .Z(n712) );
  IV U320 ( .A(B[3385]), .Z(n711) );
  IV U321 ( .A(B[3386]), .Z(n710) );
  IV U322 ( .A(B[4025]), .Z(n71) );
  IV U323 ( .A(B[3387]), .Z(n709) );
  IV U324 ( .A(B[3388]), .Z(n708) );
  IV U325 ( .A(B[3389]), .Z(n707) );
  IV U326 ( .A(B[3390]), .Z(n706) );
  IV U327 ( .A(B[3391]), .Z(n705) );
  IV U328 ( .A(B[3392]), .Z(n704) );
  IV U329 ( .A(B[3393]), .Z(n703) );
  IV U330 ( .A(B[3394]), .Z(n702) );
  IV U331 ( .A(B[3395]), .Z(n701) );
  IV U332 ( .A(B[3396]), .Z(n700) );
  IV U333 ( .A(B[4026]), .Z(n70) );
  IV U334 ( .A(B[4089]), .Z(n7) );
  IV U335 ( .A(B[3397]), .Z(n699) );
  IV U336 ( .A(B[3398]), .Z(n698) );
  IV U337 ( .A(B[3399]), .Z(n697) );
  IV U338 ( .A(B[3400]), .Z(n696) );
  IV U339 ( .A(B[3401]), .Z(n695) );
  IV U340 ( .A(B[3402]), .Z(n694) );
  IV U341 ( .A(B[3403]), .Z(n693) );
  IV U342 ( .A(B[3404]), .Z(n692) );
  IV U343 ( .A(B[3405]), .Z(n691) );
  IV U344 ( .A(B[3406]), .Z(n690) );
  IV U345 ( .A(B[4027]), .Z(n69) );
  IV U346 ( .A(B[3407]), .Z(n689) );
  IV U347 ( .A(B[3408]), .Z(n688) );
  IV U348 ( .A(B[3409]), .Z(n687) );
  IV U349 ( .A(B[3410]), .Z(n686) );
  IV U350 ( .A(B[3411]), .Z(n685) );
  IV U351 ( .A(B[3412]), .Z(n684) );
  IV U352 ( .A(B[3413]), .Z(n683) );
  IV U353 ( .A(B[3414]), .Z(n682) );
  IV U354 ( .A(B[3415]), .Z(n681) );
  IV U355 ( .A(B[3416]), .Z(n680) );
  IV U356 ( .A(B[4028]), .Z(n68) );
  IV U357 ( .A(B[3417]), .Z(n679) );
  IV U358 ( .A(B[3418]), .Z(n678) );
  IV U359 ( .A(B[3419]), .Z(n677) );
  IV U360 ( .A(B[3420]), .Z(n676) );
  IV U361 ( .A(B[3421]), .Z(n675) );
  IV U362 ( .A(B[3422]), .Z(n674) );
  IV U363 ( .A(B[3423]), .Z(n673) );
  IV U364 ( .A(B[3424]), .Z(n672) );
  IV U365 ( .A(B[3425]), .Z(n671) );
  IV U366 ( .A(B[3426]), .Z(n670) );
  IV U367 ( .A(B[4029]), .Z(n67) );
  IV U368 ( .A(B[3427]), .Z(n669) );
  IV U369 ( .A(B[3428]), .Z(n668) );
  IV U370 ( .A(B[3429]), .Z(n667) );
  IV U371 ( .A(B[3430]), .Z(n666) );
  IV U372 ( .A(B[3431]), .Z(n665) );
  IV U373 ( .A(B[3432]), .Z(n664) );
  IV U374 ( .A(B[3433]), .Z(n663) );
  IV U375 ( .A(B[3434]), .Z(n662) );
  IV U376 ( .A(B[3435]), .Z(n661) );
  IV U377 ( .A(B[3436]), .Z(n660) );
  IV U378 ( .A(B[4030]), .Z(n66) );
  IV U379 ( .A(B[3437]), .Z(n659) );
  IV U380 ( .A(B[3438]), .Z(n658) );
  IV U381 ( .A(B[3439]), .Z(n657) );
  IV U382 ( .A(B[3440]), .Z(n656) );
  IV U383 ( .A(B[3441]), .Z(n655) );
  IV U384 ( .A(B[3442]), .Z(n654) );
  IV U385 ( .A(B[3443]), .Z(n653) );
  IV U386 ( .A(B[3444]), .Z(n652) );
  IV U387 ( .A(B[3445]), .Z(n651) );
  IV U388 ( .A(B[3446]), .Z(n650) );
  IV U389 ( .A(B[4031]), .Z(n65) );
  IV U390 ( .A(B[3447]), .Z(n649) );
  IV U391 ( .A(B[3448]), .Z(n648) );
  IV U392 ( .A(B[3449]), .Z(n647) );
  IV U393 ( .A(B[3450]), .Z(n646) );
  IV U394 ( .A(B[3451]), .Z(n645) );
  IV U395 ( .A(B[3452]), .Z(n644) );
  IV U396 ( .A(B[3453]), .Z(n643) );
  IV U397 ( .A(B[3454]), .Z(n642) );
  IV U398 ( .A(B[3455]), .Z(n641) );
  IV U399 ( .A(B[3456]), .Z(n640) );
  IV U400 ( .A(B[4032]), .Z(n64) );
  IV U401 ( .A(B[3457]), .Z(n639) );
  IV U402 ( .A(B[3458]), .Z(n638) );
  IV U403 ( .A(B[3459]), .Z(n637) );
  IV U404 ( .A(B[3460]), .Z(n636) );
  IV U405 ( .A(B[3461]), .Z(n635) );
  IV U406 ( .A(B[3462]), .Z(n634) );
  IV U407 ( .A(B[3463]), .Z(n633) );
  IV U408 ( .A(B[3464]), .Z(n632) );
  IV U409 ( .A(B[3465]), .Z(n631) );
  IV U410 ( .A(B[3466]), .Z(n630) );
  IV U411 ( .A(B[4033]), .Z(n63) );
  IV U412 ( .A(B[3467]), .Z(n629) );
  IV U413 ( .A(B[3468]), .Z(n628) );
  IV U414 ( .A(B[3469]), .Z(n627) );
  IV U415 ( .A(B[3470]), .Z(n626) );
  IV U416 ( .A(B[3471]), .Z(n625) );
  IV U417 ( .A(B[3472]), .Z(n624) );
  IV U418 ( .A(B[3473]), .Z(n623) );
  IV U419 ( .A(B[3474]), .Z(n622) );
  IV U420 ( .A(B[3475]), .Z(n621) );
  IV U421 ( .A(B[3476]), .Z(n620) );
  IV U422 ( .A(B[4034]), .Z(n62) );
  IV U423 ( .A(B[3477]), .Z(n619) );
  IV U424 ( .A(B[3478]), .Z(n618) );
  IV U425 ( .A(B[3479]), .Z(n617) );
  IV U426 ( .A(B[3480]), .Z(n616) );
  IV U427 ( .A(B[3481]), .Z(n615) );
  IV U428 ( .A(B[3482]), .Z(n614) );
  IV U429 ( .A(B[3483]), .Z(n613) );
  IV U430 ( .A(B[3484]), .Z(n612) );
  IV U431 ( .A(B[3485]), .Z(n611) );
  IV U432 ( .A(B[3486]), .Z(n610) );
  IV U433 ( .A(B[4035]), .Z(n61) );
  IV U434 ( .A(B[3487]), .Z(n609) );
  IV U435 ( .A(B[3488]), .Z(n608) );
  IV U436 ( .A(B[3489]), .Z(n607) );
  IV U437 ( .A(B[3490]), .Z(n606) );
  IV U438 ( .A(B[3491]), .Z(n605) );
  IV U439 ( .A(B[3492]), .Z(n604) );
  IV U440 ( .A(B[3493]), .Z(n603) );
  IV U441 ( .A(B[3494]), .Z(n602) );
  IV U442 ( .A(B[3495]), .Z(n601) );
  IV U443 ( .A(B[3496]), .Z(n600) );
  IV U444 ( .A(B[4036]), .Z(n60) );
  IV U445 ( .A(B[4090]), .Z(n6) );
  IV U446 ( .A(B[3497]), .Z(n599) );
  IV U447 ( .A(B[3498]), .Z(n598) );
  IV U448 ( .A(B[3499]), .Z(n597) );
  IV U449 ( .A(B[3500]), .Z(n596) );
  IV U450 ( .A(B[3501]), .Z(n595) );
  IV U451 ( .A(B[3502]), .Z(n594) );
  IV U452 ( .A(B[3503]), .Z(n593) );
  IV U453 ( .A(B[3504]), .Z(n592) );
  IV U454 ( .A(B[3505]), .Z(n591) );
  IV U455 ( .A(B[3506]), .Z(n590) );
  IV U456 ( .A(B[4037]), .Z(n59) );
  IV U457 ( .A(B[3507]), .Z(n589) );
  IV U458 ( .A(B[3508]), .Z(n588) );
  IV U459 ( .A(B[3509]), .Z(n587) );
  IV U460 ( .A(B[3510]), .Z(n586) );
  IV U461 ( .A(B[3511]), .Z(n585) );
  IV U462 ( .A(B[3512]), .Z(n584) );
  IV U463 ( .A(B[3513]), .Z(n583) );
  IV U464 ( .A(B[3514]), .Z(n582) );
  IV U465 ( .A(B[3515]), .Z(n581) );
  IV U466 ( .A(B[3516]), .Z(n580) );
  IV U467 ( .A(B[4038]), .Z(n58) );
  IV U468 ( .A(B[3517]), .Z(n579) );
  IV U469 ( .A(B[3518]), .Z(n578) );
  IV U470 ( .A(B[3519]), .Z(n577) );
  IV U471 ( .A(B[3520]), .Z(n576) );
  IV U472 ( .A(B[3521]), .Z(n575) );
  IV U473 ( .A(B[3522]), .Z(n574) );
  IV U474 ( .A(B[3523]), .Z(n573) );
  IV U475 ( .A(B[3524]), .Z(n572) );
  IV U476 ( .A(B[3525]), .Z(n571) );
  IV U477 ( .A(B[3526]), .Z(n570) );
  IV U478 ( .A(B[4039]), .Z(n57) );
  IV U479 ( .A(B[3527]), .Z(n569) );
  IV U480 ( .A(B[3528]), .Z(n568) );
  IV U481 ( .A(B[3529]), .Z(n567) );
  IV U482 ( .A(B[3530]), .Z(n566) );
  IV U483 ( .A(B[3531]), .Z(n565) );
  IV U484 ( .A(B[3532]), .Z(n564) );
  IV U485 ( .A(B[3533]), .Z(n563) );
  IV U486 ( .A(B[3534]), .Z(n562) );
  IV U487 ( .A(B[3535]), .Z(n561) );
  IV U488 ( .A(B[3536]), .Z(n560) );
  IV U489 ( .A(B[4040]), .Z(n56) );
  IV U490 ( .A(B[3537]), .Z(n559) );
  IV U491 ( .A(B[3538]), .Z(n558) );
  IV U492 ( .A(B[3539]), .Z(n557) );
  IV U493 ( .A(B[3540]), .Z(n556) );
  IV U494 ( .A(B[3541]), .Z(n555) );
  IV U495 ( .A(B[3542]), .Z(n554) );
  IV U496 ( .A(B[3543]), .Z(n553) );
  IV U497 ( .A(B[3544]), .Z(n552) );
  IV U498 ( .A(B[3545]), .Z(n551) );
  IV U499 ( .A(B[3546]), .Z(n550) );
  IV U500 ( .A(B[4041]), .Z(n55) );
  IV U501 ( .A(B[3547]), .Z(n549) );
  IV U502 ( .A(B[3548]), .Z(n548) );
  IV U503 ( .A(B[3549]), .Z(n547) );
  IV U504 ( .A(B[3550]), .Z(n546) );
  IV U505 ( .A(B[3551]), .Z(n545) );
  IV U506 ( .A(B[3552]), .Z(n544) );
  IV U507 ( .A(B[3553]), .Z(n543) );
  IV U508 ( .A(B[3554]), .Z(n542) );
  IV U509 ( .A(B[3555]), .Z(n541) );
  IV U510 ( .A(B[3556]), .Z(n540) );
  IV U511 ( .A(B[4042]), .Z(n54) );
  IV U512 ( .A(B[3557]), .Z(n539) );
  IV U513 ( .A(B[3558]), .Z(n538) );
  IV U514 ( .A(B[3559]), .Z(n537) );
  IV U515 ( .A(B[3560]), .Z(n536) );
  IV U516 ( .A(B[3561]), .Z(n535) );
  IV U517 ( .A(B[3562]), .Z(n534) );
  IV U518 ( .A(B[3563]), .Z(n533) );
  IV U519 ( .A(B[3564]), .Z(n532) );
  IV U520 ( .A(B[3565]), .Z(n531) );
  IV U521 ( .A(B[3566]), .Z(n530) );
  IV U522 ( .A(B[4043]), .Z(n53) );
  IV U523 ( .A(B[3567]), .Z(n529) );
  IV U524 ( .A(B[3568]), .Z(n528) );
  IV U525 ( .A(B[3569]), .Z(n527) );
  IV U526 ( .A(B[3570]), .Z(n526) );
  IV U527 ( .A(B[3571]), .Z(n525) );
  IV U528 ( .A(B[3572]), .Z(n524) );
  IV U529 ( .A(B[3573]), .Z(n523) );
  IV U530 ( .A(B[3574]), .Z(n522) );
  IV U531 ( .A(B[3575]), .Z(n521) );
  IV U532 ( .A(B[3576]), .Z(n520) );
  IV U533 ( .A(B[4044]), .Z(n52) );
  IV U534 ( .A(B[3577]), .Z(n519) );
  IV U535 ( .A(B[3578]), .Z(n518) );
  IV U536 ( .A(B[3579]), .Z(n517) );
  IV U537 ( .A(B[3580]), .Z(n516) );
  IV U538 ( .A(B[3581]), .Z(n515) );
  IV U539 ( .A(B[3582]), .Z(n514) );
  IV U540 ( .A(B[3583]), .Z(n513) );
  IV U541 ( .A(B[3584]), .Z(n512) );
  IV U542 ( .A(B[3585]), .Z(n511) );
  IV U543 ( .A(B[3586]), .Z(n510) );
  IV U544 ( .A(B[4045]), .Z(n51) );
  IV U545 ( .A(B[3587]), .Z(n509) );
  IV U546 ( .A(B[3588]), .Z(n508) );
  IV U547 ( .A(B[3589]), .Z(n507) );
  IV U548 ( .A(B[3590]), .Z(n506) );
  IV U549 ( .A(B[3591]), .Z(n505) );
  IV U550 ( .A(B[3592]), .Z(n504) );
  IV U551 ( .A(B[3593]), .Z(n503) );
  IV U552 ( .A(B[3594]), .Z(n502) );
  IV U553 ( .A(B[3595]), .Z(n501) );
  IV U554 ( .A(B[3596]), .Z(n500) );
  IV U555 ( .A(B[4046]), .Z(n50) );
  IV U556 ( .A(B[4091]), .Z(n5) );
  IV U557 ( .A(B[3597]), .Z(n499) );
  IV U558 ( .A(B[3598]), .Z(n498) );
  IV U559 ( .A(B[3599]), .Z(n497) );
  IV U560 ( .A(B[3600]), .Z(n496) );
  IV U561 ( .A(B[3601]), .Z(n495) );
  IV U562 ( .A(B[3602]), .Z(n494) );
  IV U563 ( .A(B[3603]), .Z(n493) );
  IV U564 ( .A(B[3604]), .Z(n492) );
  IV U565 ( .A(B[3605]), .Z(n491) );
  IV U566 ( .A(B[3606]), .Z(n490) );
  IV U567 ( .A(B[4047]), .Z(n49) );
  IV U568 ( .A(B[3607]), .Z(n489) );
  IV U569 ( .A(B[3608]), .Z(n488) );
  IV U570 ( .A(B[3609]), .Z(n487) );
  IV U571 ( .A(B[3610]), .Z(n486) );
  IV U572 ( .A(B[3611]), .Z(n485) );
  IV U573 ( .A(B[3612]), .Z(n484) );
  IV U574 ( .A(B[3613]), .Z(n483) );
  IV U575 ( .A(B[3614]), .Z(n482) );
  IV U576 ( .A(B[3615]), .Z(n481) );
  IV U577 ( .A(B[3616]), .Z(n480) );
  IV U578 ( .A(B[4048]), .Z(n48) );
  IV U579 ( .A(B[3617]), .Z(n479) );
  IV U580 ( .A(B[3618]), .Z(n478) );
  IV U581 ( .A(B[3619]), .Z(n477) );
  IV U582 ( .A(B[3620]), .Z(n476) );
  IV U583 ( .A(B[3621]), .Z(n475) );
  IV U584 ( .A(B[3622]), .Z(n474) );
  IV U585 ( .A(B[3623]), .Z(n473) );
  IV U586 ( .A(B[3624]), .Z(n472) );
  IV U587 ( .A(B[3625]), .Z(n471) );
  IV U588 ( .A(B[3626]), .Z(n470) );
  IV U589 ( .A(B[4049]), .Z(n47) );
  IV U590 ( .A(B[3627]), .Z(n469) );
  IV U591 ( .A(B[3628]), .Z(n468) );
  IV U592 ( .A(B[3629]), .Z(n467) );
  IV U593 ( .A(B[3630]), .Z(n466) );
  IV U594 ( .A(B[3631]), .Z(n465) );
  IV U595 ( .A(B[3632]), .Z(n464) );
  IV U596 ( .A(B[3633]), .Z(n463) );
  IV U597 ( .A(B[3634]), .Z(n462) );
  IV U598 ( .A(B[3635]), .Z(n461) );
  IV U599 ( .A(B[3636]), .Z(n460) );
  IV U600 ( .A(B[4050]), .Z(n46) );
  IV U601 ( .A(B[3637]), .Z(n459) );
  IV U602 ( .A(B[3638]), .Z(n458) );
  IV U603 ( .A(B[3639]), .Z(n457) );
  IV U604 ( .A(B[3640]), .Z(n456) );
  IV U605 ( .A(B[3641]), .Z(n455) );
  IV U606 ( .A(B[3642]), .Z(n454) );
  IV U607 ( .A(B[3643]), .Z(n453) );
  IV U608 ( .A(B[3644]), .Z(n452) );
  IV U609 ( .A(B[3645]), .Z(n451) );
  IV U610 ( .A(B[3646]), .Z(n450) );
  IV U611 ( .A(B[4051]), .Z(n45) );
  IV U612 ( .A(B[3647]), .Z(n449) );
  IV U613 ( .A(B[3648]), .Z(n448) );
  IV U614 ( .A(B[3649]), .Z(n447) );
  IV U615 ( .A(B[3650]), .Z(n446) );
  IV U616 ( .A(B[3651]), .Z(n445) );
  IV U617 ( .A(B[3652]), .Z(n444) );
  IV U618 ( .A(B[3653]), .Z(n443) );
  IV U619 ( .A(B[3654]), .Z(n442) );
  IV U620 ( .A(B[3655]), .Z(n441) );
  IV U621 ( .A(B[3656]), .Z(n440) );
  IV U622 ( .A(B[4052]), .Z(n44) );
  IV U623 ( .A(B[3657]), .Z(n439) );
  IV U624 ( .A(B[3658]), .Z(n438) );
  IV U625 ( .A(B[3659]), .Z(n437) );
  IV U626 ( .A(B[3660]), .Z(n436) );
  IV U627 ( .A(B[3661]), .Z(n435) );
  IV U628 ( .A(B[3662]), .Z(n434) );
  IV U629 ( .A(B[3663]), .Z(n433) );
  IV U630 ( .A(B[3664]), .Z(n432) );
  IV U631 ( .A(B[3665]), .Z(n431) );
  IV U632 ( .A(B[3666]), .Z(n430) );
  IV U633 ( .A(B[4053]), .Z(n43) );
  IV U634 ( .A(B[3667]), .Z(n429) );
  IV U635 ( .A(B[3668]), .Z(n428) );
  IV U636 ( .A(B[3669]), .Z(n427) );
  IV U637 ( .A(B[3670]), .Z(n426) );
  IV U638 ( .A(B[3671]), .Z(n425) );
  IV U639 ( .A(B[3672]), .Z(n424) );
  IV U640 ( .A(B[3673]), .Z(n423) );
  IV U641 ( .A(B[3674]), .Z(n422) );
  IV U642 ( .A(B[3675]), .Z(n421) );
  IV U643 ( .A(B[3676]), .Z(n420) );
  IV U644 ( .A(B[4054]), .Z(n42) );
  IV U645 ( .A(B[3677]), .Z(n419) );
  IV U646 ( .A(B[3678]), .Z(n418) );
  IV U647 ( .A(B[3679]), .Z(n417) );
  IV U648 ( .A(B[3680]), .Z(n416) );
  IV U649 ( .A(B[3681]), .Z(n415) );
  IV U650 ( .A(B[3682]), .Z(n414) );
  IV U651 ( .A(B[3683]), .Z(n413) );
  IV U652 ( .A(B[3684]), .Z(n412) );
  IV U653 ( .A(B[3685]), .Z(n411) );
  IV U654 ( .A(B[3686]), .Z(n410) );
  IV U655 ( .A(B[4055]), .Z(n41) );
  IV U656 ( .A(B[0]), .Z(n4096) );
  IV U657 ( .A(B[1]), .Z(n4095) );
  IV U658 ( .A(B[2]), .Z(n4094) );
  IV U659 ( .A(B[3]), .Z(n4093) );
  IV U660 ( .A(B[4]), .Z(n4092) );
  IV U661 ( .A(B[5]), .Z(n4091) );
  IV U662 ( .A(B[6]), .Z(n4090) );
  IV U663 ( .A(B[3687]), .Z(n409) );
  IV U664 ( .A(B[7]), .Z(n4089) );
  IV U665 ( .A(B[8]), .Z(n4088) );
  IV U666 ( .A(B[9]), .Z(n4087) );
  IV U667 ( .A(B[10]), .Z(n4086) );
  IV U668 ( .A(B[11]), .Z(n4085) );
  IV U669 ( .A(B[12]), .Z(n4084) );
  IV U670 ( .A(B[13]), .Z(n4083) );
  IV U671 ( .A(B[14]), .Z(n4082) );
  IV U672 ( .A(B[15]), .Z(n4081) );
  IV U673 ( .A(B[16]), .Z(n4080) );
  IV U674 ( .A(B[3688]), .Z(n408) );
  IV U675 ( .A(B[17]), .Z(n4079) );
  IV U676 ( .A(B[18]), .Z(n4078) );
  IV U677 ( .A(B[19]), .Z(n4077) );
  IV U678 ( .A(B[20]), .Z(n4076) );
  IV U679 ( .A(B[21]), .Z(n4075) );
  IV U680 ( .A(B[22]), .Z(n4074) );
  IV U681 ( .A(B[23]), .Z(n4073) );
  IV U682 ( .A(B[24]), .Z(n4072) );
  IV U683 ( .A(B[25]), .Z(n4071) );
  IV U684 ( .A(B[26]), .Z(n4070) );
  IV U685 ( .A(B[3689]), .Z(n407) );
  IV U686 ( .A(B[27]), .Z(n4069) );
  IV U687 ( .A(B[28]), .Z(n4068) );
  IV U688 ( .A(B[29]), .Z(n4067) );
  IV U689 ( .A(B[30]), .Z(n4066) );
  IV U690 ( .A(B[31]), .Z(n4065) );
  IV U691 ( .A(B[32]), .Z(n4064) );
  IV U692 ( .A(B[33]), .Z(n4063) );
  IV U693 ( .A(B[34]), .Z(n4062) );
  IV U694 ( .A(B[35]), .Z(n4061) );
  IV U695 ( .A(B[36]), .Z(n4060) );
  IV U696 ( .A(B[3690]), .Z(n406) );
  IV U697 ( .A(B[37]), .Z(n4059) );
  IV U698 ( .A(B[38]), .Z(n4058) );
  IV U699 ( .A(B[39]), .Z(n4057) );
  IV U700 ( .A(B[40]), .Z(n4056) );
  IV U701 ( .A(B[41]), .Z(n4055) );
  IV U702 ( .A(B[42]), .Z(n4054) );
  IV U703 ( .A(B[43]), .Z(n4053) );
  IV U704 ( .A(B[44]), .Z(n4052) );
  IV U705 ( .A(B[45]), .Z(n4051) );
  IV U706 ( .A(B[46]), .Z(n4050) );
  IV U707 ( .A(B[3691]), .Z(n405) );
  IV U708 ( .A(B[47]), .Z(n4049) );
  IV U709 ( .A(B[48]), .Z(n4048) );
  IV U710 ( .A(B[49]), .Z(n4047) );
  IV U711 ( .A(B[50]), .Z(n4046) );
  IV U712 ( .A(B[51]), .Z(n4045) );
  IV U713 ( .A(B[52]), .Z(n4044) );
  IV U714 ( .A(B[53]), .Z(n4043) );
  IV U715 ( .A(B[54]), .Z(n4042) );
  IV U716 ( .A(B[55]), .Z(n4041) );
  IV U717 ( .A(B[56]), .Z(n4040) );
  IV U718 ( .A(B[3692]), .Z(n404) );
  IV U719 ( .A(B[57]), .Z(n4039) );
  IV U720 ( .A(B[58]), .Z(n4038) );
  IV U721 ( .A(B[59]), .Z(n4037) );
  IV U722 ( .A(B[60]), .Z(n4036) );
  IV U723 ( .A(B[61]), .Z(n4035) );
  IV U724 ( .A(B[62]), .Z(n4034) );
  IV U725 ( .A(B[63]), .Z(n4033) );
  IV U726 ( .A(B[64]), .Z(n4032) );
  IV U727 ( .A(B[65]), .Z(n4031) );
  IV U728 ( .A(B[66]), .Z(n4030) );
  IV U729 ( .A(B[3693]), .Z(n403) );
  IV U730 ( .A(B[67]), .Z(n4029) );
  IV U731 ( .A(B[68]), .Z(n4028) );
  IV U732 ( .A(B[69]), .Z(n4027) );
  IV U733 ( .A(B[70]), .Z(n4026) );
  IV U734 ( .A(B[71]), .Z(n4025) );
  IV U735 ( .A(B[72]), .Z(n4024) );
  IV U736 ( .A(B[73]), .Z(n4023) );
  IV U737 ( .A(B[74]), .Z(n4022) );
  IV U738 ( .A(B[75]), .Z(n4021) );
  IV U739 ( .A(B[76]), .Z(n4020) );
  IV U740 ( .A(B[3694]), .Z(n402) );
  IV U741 ( .A(B[77]), .Z(n4019) );
  IV U742 ( .A(B[78]), .Z(n4018) );
  IV U743 ( .A(B[79]), .Z(n4017) );
  IV U744 ( .A(B[80]), .Z(n4016) );
  IV U745 ( .A(B[81]), .Z(n4015) );
  IV U746 ( .A(B[82]), .Z(n4014) );
  IV U747 ( .A(B[83]), .Z(n4013) );
  IV U748 ( .A(B[84]), .Z(n4012) );
  IV U749 ( .A(B[85]), .Z(n4011) );
  IV U750 ( .A(B[86]), .Z(n4010) );
  IV U751 ( .A(B[3695]), .Z(n401) );
  IV U752 ( .A(B[87]), .Z(n4009) );
  IV U753 ( .A(B[88]), .Z(n4008) );
  IV U754 ( .A(B[89]), .Z(n4007) );
  IV U755 ( .A(B[90]), .Z(n4006) );
  IV U756 ( .A(B[91]), .Z(n4005) );
  IV U757 ( .A(B[92]), .Z(n4004) );
  IV U758 ( .A(B[93]), .Z(n4003) );
  IV U759 ( .A(B[94]), .Z(n4002) );
  IV U760 ( .A(B[95]), .Z(n4001) );
  IV U761 ( .A(B[96]), .Z(n4000) );
  IV U762 ( .A(B[3696]), .Z(n400) );
  IV U763 ( .A(B[4056]), .Z(n40) );
  IV U764 ( .A(B[4092]), .Z(n4) );
  IV U765 ( .A(B[97]), .Z(n3999) );
  IV U766 ( .A(B[98]), .Z(n3998) );
  IV U767 ( .A(B[99]), .Z(n3997) );
  IV U768 ( .A(B[100]), .Z(n3996) );
  IV U769 ( .A(B[101]), .Z(n3995) );
  IV U770 ( .A(B[102]), .Z(n3994) );
  IV U771 ( .A(B[103]), .Z(n3993) );
  IV U772 ( .A(B[104]), .Z(n3992) );
  IV U773 ( .A(B[105]), .Z(n3991) );
  IV U774 ( .A(B[106]), .Z(n3990) );
  IV U775 ( .A(B[3697]), .Z(n399) );
  IV U776 ( .A(B[107]), .Z(n3989) );
  IV U777 ( .A(B[108]), .Z(n3988) );
  IV U778 ( .A(B[109]), .Z(n3987) );
  IV U779 ( .A(B[110]), .Z(n3986) );
  IV U780 ( .A(B[111]), .Z(n3985) );
  IV U781 ( .A(B[112]), .Z(n3984) );
  IV U782 ( .A(B[113]), .Z(n3983) );
  IV U783 ( .A(B[114]), .Z(n3982) );
  IV U784 ( .A(B[115]), .Z(n3981) );
  IV U785 ( .A(B[116]), .Z(n3980) );
  IV U786 ( .A(B[3698]), .Z(n398) );
  IV U787 ( .A(B[117]), .Z(n3979) );
  IV U788 ( .A(B[118]), .Z(n3978) );
  IV U789 ( .A(B[119]), .Z(n3977) );
  IV U790 ( .A(B[120]), .Z(n3976) );
  IV U791 ( .A(B[121]), .Z(n3975) );
  IV U792 ( .A(B[122]), .Z(n3974) );
  IV U793 ( .A(B[123]), .Z(n3973) );
  IV U794 ( .A(B[124]), .Z(n3972) );
  IV U795 ( .A(B[125]), .Z(n3971) );
  IV U796 ( .A(B[126]), .Z(n3970) );
  IV U797 ( .A(B[3699]), .Z(n397) );
  IV U798 ( .A(B[127]), .Z(n3969) );
  IV U799 ( .A(B[128]), .Z(n3968) );
  IV U800 ( .A(B[129]), .Z(n3967) );
  IV U801 ( .A(B[130]), .Z(n3966) );
  IV U802 ( .A(B[131]), .Z(n3965) );
  IV U803 ( .A(B[132]), .Z(n3964) );
  IV U804 ( .A(B[133]), .Z(n3963) );
  IV U805 ( .A(B[134]), .Z(n3962) );
  IV U806 ( .A(B[135]), .Z(n3961) );
  IV U807 ( .A(B[136]), .Z(n3960) );
  IV U808 ( .A(B[3700]), .Z(n396) );
  IV U809 ( .A(B[137]), .Z(n3959) );
  IV U810 ( .A(B[138]), .Z(n3958) );
  IV U811 ( .A(B[139]), .Z(n3957) );
  IV U812 ( .A(B[140]), .Z(n3956) );
  IV U813 ( .A(B[141]), .Z(n3955) );
  IV U814 ( .A(B[142]), .Z(n3954) );
  IV U815 ( .A(B[143]), .Z(n3953) );
  IV U816 ( .A(B[144]), .Z(n3952) );
  IV U817 ( .A(B[145]), .Z(n3951) );
  IV U818 ( .A(B[146]), .Z(n3950) );
  IV U819 ( .A(B[3701]), .Z(n395) );
  IV U820 ( .A(B[147]), .Z(n3949) );
  IV U821 ( .A(B[148]), .Z(n3948) );
  IV U822 ( .A(B[149]), .Z(n3947) );
  IV U823 ( .A(B[150]), .Z(n3946) );
  IV U824 ( .A(B[151]), .Z(n3945) );
  IV U825 ( .A(B[152]), .Z(n3944) );
  IV U826 ( .A(B[153]), .Z(n3943) );
  IV U827 ( .A(B[154]), .Z(n3942) );
  IV U828 ( .A(B[155]), .Z(n3941) );
  IV U829 ( .A(B[156]), .Z(n3940) );
  IV U830 ( .A(B[3702]), .Z(n394) );
  IV U831 ( .A(B[157]), .Z(n3939) );
  IV U832 ( .A(B[158]), .Z(n3938) );
  IV U833 ( .A(B[159]), .Z(n3937) );
  IV U834 ( .A(B[160]), .Z(n3936) );
  IV U835 ( .A(B[161]), .Z(n3935) );
  IV U836 ( .A(B[162]), .Z(n3934) );
  IV U837 ( .A(B[163]), .Z(n3933) );
  IV U838 ( .A(B[164]), .Z(n3932) );
  IV U839 ( .A(B[165]), .Z(n3931) );
  IV U840 ( .A(B[166]), .Z(n3930) );
  IV U841 ( .A(B[3703]), .Z(n393) );
  IV U842 ( .A(B[167]), .Z(n3929) );
  IV U843 ( .A(B[168]), .Z(n3928) );
  IV U844 ( .A(B[169]), .Z(n3927) );
  IV U845 ( .A(B[170]), .Z(n3926) );
  IV U846 ( .A(B[171]), .Z(n3925) );
  IV U847 ( .A(B[172]), .Z(n3924) );
  IV U848 ( .A(B[173]), .Z(n3923) );
  IV U849 ( .A(B[174]), .Z(n3922) );
  IV U850 ( .A(B[175]), .Z(n3921) );
  IV U851 ( .A(B[176]), .Z(n3920) );
  IV U852 ( .A(B[3704]), .Z(n392) );
  IV U853 ( .A(B[177]), .Z(n3919) );
  IV U854 ( .A(B[178]), .Z(n3918) );
  IV U855 ( .A(B[179]), .Z(n3917) );
  IV U856 ( .A(B[180]), .Z(n3916) );
  IV U857 ( .A(B[181]), .Z(n3915) );
  IV U858 ( .A(B[182]), .Z(n3914) );
  IV U859 ( .A(B[183]), .Z(n3913) );
  IV U860 ( .A(B[184]), .Z(n3912) );
  IV U861 ( .A(B[185]), .Z(n3911) );
  IV U862 ( .A(B[186]), .Z(n3910) );
  IV U863 ( .A(B[3705]), .Z(n391) );
  IV U864 ( .A(B[187]), .Z(n3909) );
  IV U865 ( .A(B[188]), .Z(n3908) );
  IV U866 ( .A(B[189]), .Z(n3907) );
  IV U867 ( .A(B[190]), .Z(n3906) );
  IV U868 ( .A(B[191]), .Z(n3905) );
  IV U869 ( .A(B[192]), .Z(n3904) );
  IV U870 ( .A(B[193]), .Z(n3903) );
  IV U871 ( .A(B[194]), .Z(n3902) );
  IV U872 ( .A(B[195]), .Z(n3901) );
  IV U873 ( .A(B[196]), .Z(n3900) );
  IV U874 ( .A(B[3706]), .Z(n390) );
  IV U875 ( .A(B[4057]), .Z(n39) );
  IV U876 ( .A(B[197]), .Z(n3899) );
  IV U877 ( .A(B[198]), .Z(n3898) );
  IV U878 ( .A(B[199]), .Z(n3897) );
  IV U879 ( .A(B[200]), .Z(n3896) );
  IV U880 ( .A(B[201]), .Z(n3895) );
  IV U881 ( .A(B[202]), .Z(n3894) );
  IV U882 ( .A(B[203]), .Z(n3893) );
  IV U883 ( .A(B[204]), .Z(n3892) );
  IV U884 ( .A(B[205]), .Z(n3891) );
  IV U885 ( .A(B[206]), .Z(n3890) );
  IV U886 ( .A(B[3707]), .Z(n389) );
  IV U887 ( .A(B[207]), .Z(n3889) );
  IV U888 ( .A(B[208]), .Z(n3888) );
  IV U889 ( .A(B[209]), .Z(n3887) );
  IV U890 ( .A(B[210]), .Z(n3886) );
  IV U891 ( .A(B[211]), .Z(n3885) );
  IV U892 ( .A(B[212]), .Z(n3884) );
  IV U893 ( .A(B[213]), .Z(n3883) );
  IV U894 ( .A(B[214]), .Z(n3882) );
  IV U895 ( .A(B[215]), .Z(n3881) );
  IV U896 ( .A(B[216]), .Z(n3880) );
  IV U897 ( .A(B[3708]), .Z(n388) );
  IV U898 ( .A(B[217]), .Z(n3879) );
  IV U899 ( .A(B[218]), .Z(n3878) );
  IV U900 ( .A(B[219]), .Z(n3877) );
  IV U901 ( .A(B[220]), .Z(n3876) );
  IV U902 ( .A(B[221]), .Z(n3875) );
  IV U903 ( .A(B[222]), .Z(n3874) );
  IV U904 ( .A(B[223]), .Z(n3873) );
  IV U905 ( .A(B[224]), .Z(n3872) );
  IV U906 ( .A(B[225]), .Z(n3871) );
  IV U907 ( .A(B[226]), .Z(n3870) );
  IV U908 ( .A(B[3709]), .Z(n387) );
  IV U909 ( .A(B[227]), .Z(n3869) );
  IV U910 ( .A(B[228]), .Z(n3868) );
  IV U911 ( .A(B[229]), .Z(n3867) );
  IV U912 ( .A(B[230]), .Z(n3866) );
  IV U913 ( .A(B[231]), .Z(n3865) );
  IV U914 ( .A(B[232]), .Z(n3864) );
  IV U915 ( .A(B[233]), .Z(n3863) );
  IV U916 ( .A(B[234]), .Z(n3862) );
  IV U917 ( .A(B[235]), .Z(n3861) );
  IV U918 ( .A(B[236]), .Z(n3860) );
  IV U919 ( .A(B[3710]), .Z(n386) );
  IV U920 ( .A(B[237]), .Z(n3859) );
  IV U921 ( .A(B[238]), .Z(n3858) );
  IV U922 ( .A(B[239]), .Z(n3857) );
  IV U923 ( .A(B[240]), .Z(n3856) );
  IV U924 ( .A(B[241]), .Z(n3855) );
  IV U925 ( .A(B[242]), .Z(n3854) );
  IV U926 ( .A(B[243]), .Z(n3853) );
  IV U927 ( .A(B[244]), .Z(n3852) );
  IV U928 ( .A(B[245]), .Z(n3851) );
  IV U929 ( .A(B[246]), .Z(n3850) );
  IV U930 ( .A(B[3711]), .Z(n385) );
  IV U931 ( .A(B[247]), .Z(n3849) );
  IV U932 ( .A(B[248]), .Z(n3848) );
  IV U933 ( .A(B[249]), .Z(n3847) );
  IV U934 ( .A(B[250]), .Z(n3846) );
  IV U935 ( .A(B[251]), .Z(n3845) );
  IV U936 ( .A(B[252]), .Z(n3844) );
  IV U937 ( .A(B[253]), .Z(n3843) );
  IV U938 ( .A(B[254]), .Z(n3842) );
  IV U939 ( .A(B[255]), .Z(n3841) );
  IV U940 ( .A(B[256]), .Z(n3840) );
  IV U941 ( .A(B[3712]), .Z(n384) );
  IV U942 ( .A(B[257]), .Z(n3839) );
  IV U943 ( .A(B[258]), .Z(n3838) );
  IV U944 ( .A(B[259]), .Z(n3837) );
  IV U945 ( .A(B[260]), .Z(n3836) );
  IV U946 ( .A(B[261]), .Z(n3835) );
  IV U947 ( .A(B[262]), .Z(n3834) );
  IV U948 ( .A(B[263]), .Z(n3833) );
  IV U949 ( .A(B[264]), .Z(n3832) );
  IV U950 ( .A(B[265]), .Z(n3831) );
  IV U951 ( .A(B[266]), .Z(n3830) );
  IV U952 ( .A(B[3713]), .Z(n383) );
  IV U953 ( .A(B[267]), .Z(n3829) );
  IV U954 ( .A(B[268]), .Z(n3828) );
  IV U955 ( .A(B[269]), .Z(n3827) );
  IV U956 ( .A(B[270]), .Z(n3826) );
  IV U957 ( .A(B[271]), .Z(n3825) );
  IV U958 ( .A(B[272]), .Z(n3824) );
  IV U959 ( .A(B[273]), .Z(n3823) );
  IV U960 ( .A(B[274]), .Z(n3822) );
  IV U961 ( .A(B[275]), .Z(n3821) );
  IV U962 ( .A(B[276]), .Z(n3820) );
  IV U963 ( .A(B[3714]), .Z(n382) );
  IV U964 ( .A(B[277]), .Z(n3819) );
  IV U965 ( .A(B[278]), .Z(n3818) );
  IV U966 ( .A(B[279]), .Z(n3817) );
  IV U967 ( .A(B[280]), .Z(n3816) );
  IV U968 ( .A(B[281]), .Z(n3815) );
  IV U969 ( .A(B[282]), .Z(n3814) );
  IV U970 ( .A(B[283]), .Z(n3813) );
  IV U971 ( .A(B[284]), .Z(n3812) );
  IV U972 ( .A(B[285]), .Z(n3811) );
  IV U973 ( .A(B[286]), .Z(n3810) );
  IV U974 ( .A(B[3715]), .Z(n381) );
  IV U975 ( .A(B[287]), .Z(n3809) );
  IV U976 ( .A(B[288]), .Z(n3808) );
  IV U977 ( .A(B[289]), .Z(n3807) );
  IV U978 ( .A(B[290]), .Z(n3806) );
  IV U979 ( .A(B[291]), .Z(n3805) );
  IV U980 ( .A(B[292]), .Z(n3804) );
  IV U981 ( .A(B[293]), .Z(n3803) );
  IV U982 ( .A(B[294]), .Z(n3802) );
  IV U983 ( .A(B[295]), .Z(n3801) );
  IV U984 ( .A(B[296]), .Z(n3800) );
  IV U985 ( .A(B[3716]), .Z(n380) );
  IV U986 ( .A(B[4058]), .Z(n38) );
  IV U987 ( .A(B[297]), .Z(n3799) );
  IV U988 ( .A(B[298]), .Z(n3798) );
  IV U989 ( .A(B[299]), .Z(n3797) );
  IV U990 ( .A(B[300]), .Z(n3796) );
  IV U991 ( .A(B[301]), .Z(n3795) );
  IV U992 ( .A(B[302]), .Z(n3794) );
  IV U993 ( .A(B[303]), .Z(n3793) );
  IV U994 ( .A(B[304]), .Z(n3792) );
  IV U995 ( .A(B[305]), .Z(n3791) );
  IV U996 ( .A(B[306]), .Z(n3790) );
  IV U997 ( .A(B[3717]), .Z(n379) );
  IV U998 ( .A(B[307]), .Z(n3789) );
  IV U999 ( .A(B[308]), .Z(n3788) );
  IV U1000 ( .A(B[309]), .Z(n3787) );
  IV U1001 ( .A(B[310]), .Z(n3786) );
  IV U1002 ( .A(B[311]), .Z(n3785) );
  IV U1003 ( .A(B[312]), .Z(n3784) );
  IV U1004 ( .A(B[313]), .Z(n3783) );
  IV U1005 ( .A(B[314]), .Z(n3782) );
  IV U1006 ( .A(B[315]), .Z(n3781) );
  IV U1007 ( .A(B[316]), .Z(n3780) );
  IV U1008 ( .A(B[3718]), .Z(n378) );
  IV U1009 ( .A(B[317]), .Z(n3779) );
  IV U1010 ( .A(B[318]), .Z(n3778) );
  IV U1011 ( .A(B[319]), .Z(n3777) );
  IV U1012 ( .A(B[320]), .Z(n3776) );
  IV U1013 ( .A(B[321]), .Z(n3775) );
  IV U1014 ( .A(B[322]), .Z(n3774) );
  IV U1015 ( .A(B[323]), .Z(n3773) );
  IV U1016 ( .A(B[324]), .Z(n3772) );
  IV U1017 ( .A(B[325]), .Z(n3771) );
  IV U1018 ( .A(B[326]), .Z(n3770) );
  IV U1019 ( .A(B[3719]), .Z(n377) );
  IV U1020 ( .A(B[327]), .Z(n3769) );
  IV U1021 ( .A(B[328]), .Z(n3768) );
  IV U1022 ( .A(B[329]), .Z(n3767) );
  IV U1023 ( .A(B[330]), .Z(n3766) );
  IV U1024 ( .A(B[331]), .Z(n3765) );
  IV U1025 ( .A(B[332]), .Z(n3764) );
  IV U1026 ( .A(B[333]), .Z(n3763) );
  IV U1027 ( .A(B[334]), .Z(n3762) );
  IV U1028 ( .A(B[335]), .Z(n3761) );
  IV U1029 ( .A(B[336]), .Z(n3760) );
  IV U1030 ( .A(B[3720]), .Z(n376) );
  IV U1031 ( .A(B[337]), .Z(n3759) );
  IV U1032 ( .A(B[338]), .Z(n3758) );
  IV U1033 ( .A(B[339]), .Z(n3757) );
  IV U1034 ( .A(B[340]), .Z(n3756) );
  IV U1035 ( .A(B[341]), .Z(n3755) );
  IV U1036 ( .A(B[342]), .Z(n3754) );
  IV U1037 ( .A(B[343]), .Z(n3753) );
  IV U1038 ( .A(B[344]), .Z(n3752) );
  IV U1039 ( .A(B[345]), .Z(n3751) );
  IV U1040 ( .A(B[346]), .Z(n3750) );
  IV U1041 ( .A(B[3721]), .Z(n375) );
  IV U1042 ( .A(B[347]), .Z(n3749) );
  IV U1043 ( .A(B[348]), .Z(n3748) );
  IV U1044 ( .A(B[349]), .Z(n3747) );
  IV U1045 ( .A(B[350]), .Z(n3746) );
  IV U1046 ( .A(B[351]), .Z(n3745) );
  IV U1047 ( .A(B[352]), .Z(n3744) );
  IV U1048 ( .A(B[353]), .Z(n3743) );
  IV U1049 ( .A(B[354]), .Z(n3742) );
  IV U1050 ( .A(B[355]), .Z(n3741) );
  IV U1051 ( .A(B[356]), .Z(n3740) );
  IV U1052 ( .A(B[3722]), .Z(n374) );
  IV U1053 ( .A(B[357]), .Z(n3739) );
  IV U1054 ( .A(B[358]), .Z(n3738) );
  IV U1055 ( .A(B[359]), .Z(n3737) );
  IV U1056 ( .A(B[360]), .Z(n3736) );
  IV U1057 ( .A(B[361]), .Z(n3735) );
  IV U1058 ( .A(B[362]), .Z(n3734) );
  IV U1059 ( .A(B[363]), .Z(n3733) );
  IV U1060 ( .A(B[364]), .Z(n3732) );
  IV U1061 ( .A(B[365]), .Z(n3731) );
  IV U1062 ( .A(B[366]), .Z(n3730) );
  IV U1063 ( .A(B[3723]), .Z(n373) );
  IV U1064 ( .A(B[367]), .Z(n3729) );
  IV U1065 ( .A(B[368]), .Z(n3728) );
  IV U1066 ( .A(B[369]), .Z(n3727) );
  IV U1067 ( .A(B[370]), .Z(n3726) );
  IV U1068 ( .A(B[371]), .Z(n3725) );
  IV U1069 ( .A(B[372]), .Z(n3724) );
  IV U1070 ( .A(B[373]), .Z(n3723) );
  IV U1071 ( .A(B[374]), .Z(n3722) );
  IV U1072 ( .A(B[375]), .Z(n3721) );
  IV U1073 ( .A(B[376]), .Z(n3720) );
  IV U1074 ( .A(B[3724]), .Z(n372) );
  IV U1075 ( .A(B[377]), .Z(n3719) );
  IV U1076 ( .A(B[378]), .Z(n3718) );
  IV U1077 ( .A(B[379]), .Z(n3717) );
  IV U1078 ( .A(B[380]), .Z(n3716) );
  IV U1079 ( .A(B[381]), .Z(n3715) );
  IV U1080 ( .A(B[382]), .Z(n3714) );
  IV U1081 ( .A(B[383]), .Z(n3713) );
  IV U1082 ( .A(B[384]), .Z(n3712) );
  IV U1083 ( .A(B[385]), .Z(n3711) );
  IV U1084 ( .A(B[386]), .Z(n3710) );
  IV U1085 ( .A(B[3725]), .Z(n371) );
  IV U1086 ( .A(B[387]), .Z(n3709) );
  IV U1087 ( .A(B[388]), .Z(n3708) );
  IV U1088 ( .A(B[389]), .Z(n3707) );
  IV U1089 ( .A(B[390]), .Z(n3706) );
  IV U1090 ( .A(B[391]), .Z(n3705) );
  IV U1091 ( .A(B[392]), .Z(n3704) );
  IV U1092 ( .A(B[393]), .Z(n3703) );
  IV U1093 ( .A(B[394]), .Z(n3702) );
  IV U1094 ( .A(B[395]), .Z(n3701) );
  IV U1095 ( .A(B[396]), .Z(n3700) );
  IV U1096 ( .A(B[3726]), .Z(n370) );
  IV U1097 ( .A(B[4059]), .Z(n37) );
  IV U1098 ( .A(B[397]), .Z(n3699) );
  IV U1099 ( .A(B[398]), .Z(n3698) );
  IV U1100 ( .A(B[399]), .Z(n3697) );
  IV U1101 ( .A(B[400]), .Z(n3696) );
  IV U1102 ( .A(B[401]), .Z(n3695) );
  IV U1103 ( .A(B[402]), .Z(n3694) );
  IV U1104 ( .A(B[403]), .Z(n3693) );
  IV U1105 ( .A(B[404]), .Z(n3692) );
  IV U1106 ( .A(B[405]), .Z(n3691) );
  IV U1107 ( .A(B[406]), .Z(n3690) );
  IV U1108 ( .A(B[3727]), .Z(n369) );
  IV U1109 ( .A(B[407]), .Z(n3689) );
  IV U1110 ( .A(B[408]), .Z(n3688) );
  IV U1111 ( .A(B[409]), .Z(n3687) );
  IV U1112 ( .A(B[410]), .Z(n3686) );
  IV U1113 ( .A(B[411]), .Z(n3685) );
  IV U1114 ( .A(B[412]), .Z(n3684) );
  IV U1115 ( .A(B[413]), .Z(n3683) );
  IV U1116 ( .A(B[414]), .Z(n3682) );
  IV U1117 ( .A(B[415]), .Z(n3681) );
  IV U1118 ( .A(B[416]), .Z(n3680) );
  IV U1119 ( .A(B[3728]), .Z(n368) );
  IV U1120 ( .A(B[417]), .Z(n3679) );
  IV U1121 ( .A(B[418]), .Z(n3678) );
  IV U1122 ( .A(B[419]), .Z(n3677) );
  IV U1123 ( .A(B[420]), .Z(n3676) );
  IV U1124 ( .A(B[421]), .Z(n3675) );
  IV U1125 ( .A(B[422]), .Z(n3674) );
  IV U1126 ( .A(B[423]), .Z(n3673) );
  IV U1127 ( .A(B[424]), .Z(n3672) );
  IV U1128 ( .A(B[425]), .Z(n3671) );
  IV U1129 ( .A(B[426]), .Z(n3670) );
  IV U1130 ( .A(B[3729]), .Z(n367) );
  IV U1131 ( .A(B[427]), .Z(n3669) );
  IV U1132 ( .A(B[428]), .Z(n3668) );
  IV U1133 ( .A(B[429]), .Z(n3667) );
  IV U1134 ( .A(B[430]), .Z(n3666) );
  IV U1135 ( .A(B[431]), .Z(n3665) );
  IV U1136 ( .A(B[432]), .Z(n3664) );
  IV U1137 ( .A(B[433]), .Z(n3663) );
  IV U1138 ( .A(B[434]), .Z(n3662) );
  IV U1139 ( .A(B[435]), .Z(n3661) );
  IV U1140 ( .A(B[436]), .Z(n3660) );
  IV U1141 ( .A(B[3730]), .Z(n366) );
  IV U1142 ( .A(B[437]), .Z(n3659) );
  IV U1143 ( .A(B[438]), .Z(n3658) );
  IV U1144 ( .A(B[439]), .Z(n3657) );
  IV U1145 ( .A(B[440]), .Z(n3656) );
  IV U1146 ( .A(B[441]), .Z(n3655) );
  IV U1147 ( .A(B[442]), .Z(n3654) );
  IV U1148 ( .A(B[443]), .Z(n3653) );
  IV U1149 ( .A(B[444]), .Z(n3652) );
  IV U1150 ( .A(B[445]), .Z(n3651) );
  IV U1151 ( .A(B[446]), .Z(n3650) );
  IV U1152 ( .A(B[3731]), .Z(n365) );
  IV U1153 ( .A(B[447]), .Z(n3649) );
  IV U1154 ( .A(B[448]), .Z(n3648) );
  IV U1155 ( .A(B[449]), .Z(n3647) );
  IV U1156 ( .A(B[450]), .Z(n3646) );
  IV U1157 ( .A(B[451]), .Z(n3645) );
  IV U1158 ( .A(B[452]), .Z(n3644) );
  IV U1159 ( .A(B[453]), .Z(n3643) );
  IV U1160 ( .A(B[454]), .Z(n3642) );
  IV U1161 ( .A(B[455]), .Z(n3641) );
  IV U1162 ( .A(B[456]), .Z(n3640) );
  IV U1163 ( .A(B[3732]), .Z(n364) );
  IV U1164 ( .A(B[457]), .Z(n3639) );
  IV U1165 ( .A(B[458]), .Z(n3638) );
  IV U1166 ( .A(B[459]), .Z(n3637) );
  IV U1167 ( .A(B[460]), .Z(n3636) );
  IV U1168 ( .A(B[461]), .Z(n3635) );
  IV U1169 ( .A(B[462]), .Z(n3634) );
  IV U1170 ( .A(B[463]), .Z(n3633) );
  IV U1171 ( .A(B[464]), .Z(n3632) );
  IV U1172 ( .A(B[465]), .Z(n3631) );
  IV U1173 ( .A(B[466]), .Z(n3630) );
  IV U1174 ( .A(B[3733]), .Z(n363) );
  IV U1175 ( .A(B[467]), .Z(n3629) );
  IV U1176 ( .A(B[468]), .Z(n3628) );
  IV U1177 ( .A(B[469]), .Z(n3627) );
  IV U1178 ( .A(B[470]), .Z(n3626) );
  IV U1179 ( .A(B[471]), .Z(n3625) );
  IV U1180 ( .A(B[472]), .Z(n3624) );
  IV U1181 ( .A(B[473]), .Z(n3623) );
  IV U1182 ( .A(B[474]), .Z(n3622) );
  IV U1183 ( .A(B[475]), .Z(n3621) );
  IV U1184 ( .A(B[476]), .Z(n3620) );
  IV U1185 ( .A(B[3734]), .Z(n362) );
  IV U1186 ( .A(B[477]), .Z(n3619) );
  IV U1187 ( .A(B[478]), .Z(n3618) );
  IV U1188 ( .A(B[479]), .Z(n3617) );
  IV U1189 ( .A(B[480]), .Z(n3616) );
  IV U1190 ( .A(B[481]), .Z(n3615) );
  IV U1191 ( .A(B[482]), .Z(n3614) );
  IV U1192 ( .A(B[483]), .Z(n3613) );
  IV U1193 ( .A(B[484]), .Z(n3612) );
  IV U1194 ( .A(B[485]), .Z(n3611) );
  IV U1195 ( .A(B[486]), .Z(n3610) );
  IV U1196 ( .A(B[3735]), .Z(n361) );
  IV U1197 ( .A(B[487]), .Z(n3609) );
  IV U1198 ( .A(B[488]), .Z(n3608) );
  IV U1199 ( .A(B[489]), .Z(n3607) );
  IV U1200 ( .A(B[490]), .Z(n3606) );
  IV U1201 ( .A(B[491]), .Z(n3605) );
  IV U1202 ( .A(B[492]), .Z(n3604) );
  IV U1203 ( .A(B[493]), .Z(n3603) );
  IV U1204 ( .A(B[494]), .Z(n3602) );
  IV U1205 ( .A(B[495]), .Z(n3601) );
  IV U1206 ( .A(B[496]), .Z(n3600) );
  IV U1207 ( .A(B[3736]), .Z(n360) );
  IV U1208 ( .A(B[4060]), .Z(n36) );
  IV U1209 ( .A(B[497]), .Z(n3599) );
  IV U1210 ( .A(B[498]), .Z(n3598) );
  IV U1211 ( .A(B[499]), .Z(n3597) );
  IV U1212 ( .A(B[500]), .Z(n3596) );
  IV U1213 ( .A(B[501]), .Z(n3595) );
  IV U1214 ( .A(B[502]), .Z(n3594) );
  IV U1215 ( .A(B[503]), .Z(n3593) );
  IV U1216 ( .A(B[504]), .Z(n3592) );
  IV U1217 ( .A(B[505]), .Z(n3591) );
  IV U1218 ( .A(B[506]), .Z(n3590) );
  IV U1219 ( .A(B[3737]), .Z(n359) );
  IV U1220 ( .A(B[507]), .Z(n3589) );
  IV U1221 ( .A(B[508]), .Z(n3588) );
  IV U1222 ( .A(B[509]), .Z(n3587) );
  IV U1223 ( .A(B[510]), .Z(n3586) );
  IV U1224 ( .A(B[511]), .Z(n3585) );
  IV U1225 ( .A(B[512]), .Z(n3584) );
  IV U1226 ( .A(B[513]), .Z(n3583) );
  IV U1227 ( .A(B[514]), .Z(n3582) );
  IV U1228 ( .A(B[515]), .Z(n3581) );
  IV U1229 ( .A(B[516]), .Z(n3580) );
  IV U1230 ( .A(B[3738]), .Z(n358) );
  IV U1231 ( .A(B[517]), .Z(n3579) );
  IV U1232 ( .A(B[518]), .Z(n3578) );
  IV U1233 ( .A(B[519]), .Z(n3577) );
  IV U1234 ( .A(B[520]), .Z(n3576) );
  IV U1235 ( .A(B[521]), .Z(n3575) );
  IV U1236 ( .A(B[522]), .Z(n3574) );
  IV U1237 ( .A(B[523]), .Z(n3573) );
  IV U1238 ( .A(B[524]), .Z(n3572) );
  IV U1239 ( .A(B[525]), .Z(n3571) );
  IV U1240 ( .A(B[526]), .Z(n3570) );
  IV U1241 ( .A(B[3739]), .Z(n357) );
  IV U1242 ( .A(B[527]), .Z(n3569) );
  IV U1243 ( .A(B[528]), .Z(n3568) );
  IV U1244 ( .A(B[529]), .Z(n3567) );
  IV U1245 ( .A(B[530]), .Z(n3566) );
  IV U1246 ( .A(B[531]), .Z(n3565) );
  IV U1247 ( .A(B[532]), .Z(n3564) );
  IV U1248 ( .A(B[533]), .Z(n3563) );
  IV U1249 ( .A(B[534]), .Z(n3562) );
  IV U1250 ( .A(B[535]), .Z(n3561) );
  IV U1251 ( .A(B[536]), .Z(n3560) );
  IV U1252 ( .A(B[3740]), .Z(n356) );
  IV U1253 ( .A(B[537]), .Z(n3559) );
  IV U1254 ( .A(B[538]), .Z(n3558) );
  IV U1255 ( .A(B[539]), .Z(n3557) );
  IV U1256 ( .A(B[540]), .Z(n3556) );
  IV U1257 ( .A(B[541]), .Z(n3555) );
  IV U1258 ( .A(B[542]), .Z(n3554) );
  IV U1259 ( .A(B[543]), .Z(n3553) );
  IV U1260 ( .A(B[544]), .Z(n3552) );
  IV U1261 ( .A(B[545]), .Z(n3551) );
  IV U1262 ( .A(B[546]), .Z(n3550) );
  IV U1263 ( .A(B[3741]), .Z(n355) );
  IV U1264 ( .A(B[547]), .Z(n3549) );
  IV U1265 ( .A(B[548]), .Z(n3548) );
  IV U1266 ( .A(B[549]), .Z(n3547) );
  IV U1267 ( .A(B[550]), .Z(n3546) );
  IV U1268 ( .A(B[551]), .Z(n3545) );
  IV U1269 ( .A(B[552]), .Z(n3544) );
  IV U1270 ( .A(B[553]), .Z(n3543) );
  IV U1271 ( .A(B[554]), .Z(n3542) );
  IV U1272 ( .A(B[555]), .Z(n3541) );
  IV U1273 ( .A(B[556]), .Z(n3540) );
  IV U1274 ( .A(B[3742]), .Z(n354) );
  IV U1275 ( .A(B[557]), .Z(n3539) );
  IV U1276 ( .A(B[558]), .Z(n3538) );
  IV U1277 ( .A(B[559]), .Z(n3537) );
  IV U1278 ( .A(B[560]), .Z(n3536) );
  IV U1279 ( .A(B[561]), .Z(n3535) );
  IV U1280 ( .A(B[562]), .Z(n3534) );
  IV U1281 ( .A(B[563]), .Z(n3533) );
  IV U1282 ( .A(B[564]), .Z(n3532) );
  IV U1283 ( .A(B[565]), .Z(n3531) );
  IV U1284 ( .A(B[566]), .Z(n3530) );
  IV U1285 ( .A(B[3743]), .Z(n353) );
  IV U1286 ( .A(B[567]), .Z(n3529) );
  IV U1287 ( .A(B[568]), .Z(n3528) );
  IV U1288 ( .A(B[569]), .Z(n3527) );
  IV U1289 ( .A(B[570]), .Z(n3526) );
  IV U1290 ( .A(B[571]), .Z(n3525) );
  IV U1291 ( .A(B[572]), .Z(n3524) );
  IV U1292 ( .A(B[573]), .Z(n3523) );
  IV U1293 ( .A(B[574]), .Z(n3522) );
  IV U1294 ( .A(B[575]), .Z(n3521) );
  IV U1295 ( .A(B[576]), .Z(n3520) );
  IV U1296 ( .A(B[3744]), .Z(n352) );
  IV U1297 ( .A(B[577]), .Z(n3519) );
  IV U1298 ( .A(B[578]), .Z(n3518) );
  IV U1299 ( .A(B[579]), .Z(n3517) );
  IV U1300 ( .A(B[580]), .Z(n3516) );
  IV U1301 ( .A(B[581]), .Z(n3515) );
  IV U1302 ( .A(B[582]), .Z(n3514) );
  IV U1303 ( .A(B[583]), .Z(n3513) );
  IV U1304 ( .A(B[584]), .Z(n3512) );
  IV U1305 ( .A(B[585]), .Z(n3511) );
  IV U1306 ( .A(B[586]), .Z(n3510) );
  IV U1307 ( .A(B[3745]), .Z(n351) );
  IV U1308 ( .A(B[587]), .Z(n3509) );
  IV U1309 ( .A(B[588]), .Z(n3508) );
  IV U1310 ( .A(B[589]), .Z(n3507) );
  IV U1311 ( .A(B[590]), .Z(n3506) );
  IV U1312 ( .A(B[591]), .Z(n3505) );
  IV U1313 ( .A(B[592]), .Z(n3504) );
  IV U1314 ( .A(B[593]), .Z(n3503) );
  IV U1315 ( .A(B[594]), .Z(n3502) );
  IV U1316 ( .A(B[595]), .Z(n3501) );
  IV U1317 ( .A(B[596]), .Z(n3500) );
  IV U1318 ( .A(B[3746]), .Z(n350) );
  IV U1319 ( .A(B[4061]), .Z(n35) );
  IV U1320 ( .A(B[597]), .Z(n3499) );
  IV U1321 ( .A(B[598]), .Z(n3498) );
  IV U1322 ( .A(B[599]), .Z(n3497) );
  IV U1323 ( .A(B[600]), .Z(n3496) );
  IV U1324 ( .A(B[601]), .Z(n3495) );
  IV U1325 ( .A(B[602]), .Z(n3494) );
  IV U1326 ( .A(B[603]), .Z(n3493) );
  IV U1327 ( .A(B[604]), .Z(n3492) );
  IV U1328 ( .A(B[605]), .Z(n3491) );
  IV U1329 ( .A(B[606]), .Z(n3490) );
  IV U1330 ( .A(B[3747]), .Z(n349) );
  IV U1331 ( .A(B[607]), .Z(n3489) );
  IV U1332 ( .A(B[608]), .Z(n3488) );
  IV U1333 ( .A(B[609]), .Z(n3487) );
  IV U1334 ( .A(B[610]), .Z(n3486) );
  IV U1335 ( .A(B[611]), .Z(n3485) );
  IV U1336 ( .A(B[612]), .Z(n3484) );
  IV U1337 ( .A(B[613]), .Z(n3483) );
  IV U1338 ( .A(B[614]), .Z(n3482) );
  IV U1339 ( .A(B[615]), .Z(n3481) );
  IV U1340 ( .A(B[616]), .Z(n3480) );
  IV U1341 ( .A(B[3748]), .Z(n348) );
  IV U1342 ( .A(B[617]), .Z(n3479) );
  IV U1343 ( .A(B[618]), .Z(n3478) );
  IV U1344 ( .A(B[619]), .Z(n3477) );
  IV U1345 ( .A(B[620]), .Z(n3476) );
  IV U1346 ( .A(B[621]), .Z(n3475) );
  IV U1347 ( .A(B[622]), .Z(n3474) );
  IV U1348 ( .A(B[623]), .Z(n3473) );
  IV U1349 ( .A(B[624]), .Z(n3472) );
  IV U1350 ( .A(B[625]), .Z(n3471) );
  IV U1351 ( .A(B[626]), .Z(n3470) );
  IV U1352 ( .A(B[3749]), .Z(n347) );
  IV U1353 ( .A(B[627]), .Z(n3469) );
  IV U1354 ( .A(B[628]), .Z(n3468) );
  IV U1355 ( .A(B[629]), .Z(n3467) );
  IV U1356 ( .A(B[630]), .Z(n3466) );
  IV U1357 ( .A(B[631]), .Z(n3465) );
  IV U1358 ( .A(B[632]), .Z(n3464) );
  IV U1359 ( .A(B[633]), .Z(n3463) );
  IV U1360 ( .A(B[634]), .Z(n3462) );
  IV U1361 ( .A(B[635]), .Z(n3461) );
  IV U1362 ( .A(B[636]), .Z(n3460) );
  IV U1363 ( .A(B[3750]), .Z(n346) );
  IV U1364 ( .A(B[637]), .Z(n3459) );
  IV U1365 ( .A(B[638]), .Z(n3458) );
  IV U1366 ( .A(B[639]), .Z(n3457) );
  IV U1367 ( .A(B[640]), .Z(n3456) );
  IV U1368 ( .A(B[641]), .Z(n3455) );
  IV U1369 ( .A(B[642]), .Z(n3454) );
  IV U1370 ( .A(B[643]), .Z(n3453) );
  IV U1371 ( .A(B[644]), .Z(n3452) );
  IV U1372 ( .A(B[645]), .Z(n3451) );
  IV U1373 ( .A(B[646]), .Z(n3450) );
  IV U1374 ( .A(B[3751]), .Z(n345) );
  IV U1375 ( .A(B[647]), .Z(n3449) );
  IV U1376 ( .A(B[648]), .Z(n3448) );
  IV U1377 ( .A(B[649]), .Z(n3447) );
  IV U1378 ( .A(B[650]), .Z(n3446) );
  IV U1379 ( .A(B[651]), .Z(n3445) );
  IV U1380 ( .A(B[652]), .Z(n3444) );
  IV U1381 ( .A(B[653]), .Z(n3443) );
  IV U1382 ( .A(B[654]), .Z(n3442) );
  IV U1383 ( .A(B[655]), .Z(n3441) );
  IV U1384 ( .A(B[656]), .Z(n3440) );
  IV U1385 ( .A(B[3752]), .Z(n344) );
  IV U1386 ( .A(B[657]), .Z(n3439) );
  IV U1387 ( .A(B[658]), .Z(n3438) );
  IV U1388 ( .A(B[659]), .Z(n3437) );
  IV U1389 ( .A(B[660]), .Z(n3436) );
  IV U1390 ( .A(B[661]), .Z(n3435) );
  IV U1391 ( .A(B[662]), .Z(n3434) );
  IV U1392 ( .A(B[663]), .Z(n3433) );
  IV U1393 ( .A(B[664]), .Z(n3432) );
  IV U1394 ( .A(B[665]), .Z(n3431) );
  IV U1395 ( .A(B[666]), .Z(n3430) );
  IV U1396 ( .A(B[3753]), .Z(n343) );
  IV U1397 ( .A(B[667]), .Z(n3429) );
  IV U1398 ( .A(B[668]), .Z(n3428) );
  IV U1399 ( .A(B[669]), .Z(n3427) );
  IV U1400 ( .A(B[670]), .Z(n3426) );
  IV U1401 ( .A(B[671]), .Z(n3425) );
  IV U1402 ( .A(B[672]), .Z(n3424) );
  IV U1403 ( .A(B[673]), .Z(n3423) );
  IV U1404 ( .A(B[674]), .Z(n3422) );
  IV U1405 ( .A(B[675]), .Z(n3421) );
  IV U1406 ( .A(B[676]), .Z(n3420) );
  IV U1407 ( .A(B[3754]), .Z(n342) );
  IV U1408 ( .A(B[677]), .Z(n3419) );
  IV U1409 ( .A(B[678]), .Z(n3418) );
  IV U1410 ( .A(B[679]), .Z(n3417) );
  IV U1411 ( .A(B[680]), .Z(n3416) );
  IV U1412 ( .A(B[681]), .Z(n3415) );
  IV U1413 ( .A(B[682]), .Z(n3414) );
  IV U1414 ( .A(B[683]), .Z(n3413) );
  IV U1415 ( .A(B[684]), .Z(n3412) );
  IV U1416 ( .A(B[685]), .Z(n3411) );
  IV U1417 ( .A(B[686]), .Z(n3410) );
  IV U1418 ( .A(B[3755]), .Z(n341) );
  IV U1419 ( .A(B[687]), .Z(n3409) );
  IV U1420 ( .A(B[688]), .Z(n3408) );
  IV U1421 ( .A(B[689]), .Z(n3407) );
  IV U1422 ( .A(B[690]), .Z(n3406) );
  IV U1423 ( .A(B[691]), .Z(n3405) );
  IV U1424 ( .A(B[692]), .Z(n3404) );
  IV U1425 ( .A(B[693]), .Z(n3403) );
  IV U1426 ( .A(B[694]), .Z(n3402) );
  IV U1427 ( .A(B[695]), .Z(n3401) );
  IV U1428 ( .A(B[696]), .Z(n3400) );
  IV U1429 ( .A(B[3756]), .Z(n340) );
  IV U1430 ( .A(B[4062]), .Z(n34) );
  IV U1431 ( .A(B[697]), .Z(n3399) );
  IV U1432 ( .A(B[698]), .Z(n3398) );
  IV U1433 ( .A(B[699]), .Z(n3397) );
  IV U1434 ( .A(B[700]), .Z(n3396) );
  IV U1435 ( .A(B[701]), .Z(n3395) );
  IV U1436 ( .A(B[702]), .Z(n3394) );
  IV U1437 ( .A(B[703]), .Z(n3393) );
  IV U1438 ( .A(B[704]), .Z(n3392) );
  IV U1439 ( .A(B[705]), .Z(n3391) );
  IV U1440 ( .A(B[706]), .Z(n3390) );
  IV U1441 ( .A(B[3757]), .Z(n339) );
  IV U1442 ( .A(B[707]), .Z(n3389) );
  IV U1443 ( .A(B[708]), .Z(n3388) );
  IV U1444 ( .A(B[709]), .Z(n3387) );
  IV U1445 ( .A(B[710]), .Z(n3386) );
  IV U1446 ( .A(B[711]), .Z(n3385) );
  IV U1447 ( .A(B[712]), .Z(n3384) );
  IV U1448 ( .A(B[713]), .Z(n3383) );
  IV U1449 ( .A(B[714]), .Z(n3382) );
  IV U1450 ( .A(B[715]), .Z(n3381) );
  IV U1451 ( .A(B[716]), .Z(n3380) );
  IV U1452 ( .A(B[3758]), .Z(n338) );
  IV U1453 ( .A(B[717]), .Z(n3379) );
  IV U1454 ( .A(B[718]), .Z(n3378) );
  IV U1455 ( .A(B[719]), .Z(n3377) );
  IV U1456 ( .A(B[720]), .Z(n3376) );
  IV U1457 ( .A(B[721]), .Z(n3375) );
  IV U1458 ( .A(B[722]), .Z(n3374) );
  IV U1459 ( .A(B[723]), .Z(n3373) );
  IV U1460 ( .A(B[724]), .Z(n3372) );
  IV U1461 ( .A(B[725]), .Z(n3371) );
  IV U1462 ( .A(B[726]), .Z(n3370) );
  IV U1463 ( .A(B[3759]), .Z(n337) );
  IV U1464 ( .A(B[727]), .Z(n3369) );
  IV U1465 ( .A(B[728]), .Z(n3368) );
  IV U1466 ( .A(B[729]), .Z(n3367) );
  IV U1467 ( .A(B[730]), .Z(n3366) );
  IV U1468 ( .A(B[731]), .Z(n3365) );
  IV U1469 ( .A(B[732]), .Z(n3364) );
  IV U1470 ( .A(B[733]), .Z(n3363) );
  IV U1471 ( .A(B[734]), .Z(n3362) );
  IV U1472 ( .A(B[735]), .Z(n3361) );
  IV U1473 ( .A(B[736]), .Z(n3360) );
  IV U1474 ( .A(B[3760]), .Z(n336) );
  IV U1475 ( .A(B[737]), .Z(n3359) );
  IV U1476 ( .A(B[738]), .Z(n3358) );
  IV U1477 ( .A(B[739]), .Z(n3357) );
  IV U1478 ( .A(B[740]), .Z(n3356) );
  IV U1479 ( .A(B[741]), .Z(n3355) );
  IV U1480 ( .A(B[742]), .Z(n3354) );
  IV U1481 ( .A(B[743]), .Z(n3353) );
  IV U1482 ( .A(B[744]), .Z(n3352) );
  IV U1483 ( .A(B[745]), .Z(n3351) );
  IV U1484 ( .A(B[746]), .Z(n3350) );
  IV U1485 ( .A(B[3761]), .Z(n335) );
  IV U1486 ( .A(B[747]), .Z(n3349) );
  IV U1487 ( .A(B[748]), .Z(n3348) );
  IV U1488 ( .A(B[749]), .Z(n3347) );
  IV U1489 ( .A(B[750]), .Z(n3346) );
  IV U1490 ( .A(B[751]), .Z(n3345) );
  IV U1491 ( .A(B[752]), .Z(n3344) );
  IV U1492 ( .A(B[753]), .Z(n3343) );
  IV U1493 ( .A(B[754]), .Z(n3342) );
  IV U1494 ( .A(B[755]), .Z(n3341) );
  IV U1495 ( .A(B[756]), .Z(n3340) );
  IV U1496 ( .A(B[3762]), .Z(n334) );
  IV U1497 ( .A(B[757]), .Z(n3339) );
  IV U1498 ( .A(B[758]), .Z(n3338) );
  IV U1499 ( .A(B[759]), .Z(n3337) );
  IV U1500 ( .A(B[760]), .Z(n3336) );
  IV U1501 ( .A(B[761]), .Z(n3335) );
  IV U1502 ( .A(B[762]), .Z(n3334) );
  IV U1503 ( .A(B[763]), .Z(n3333) );
  IV U1504 ( .A(B[764]), .Z(n3332) );
  IV U1505 ( .A(B[765]), .Z(n3331) );
  IV U1506 ( .A(B[766]), .Z(n3330) );
  IV U1507 ( .A(B[3763]), .Z(n333) );
  IV U1508 ( .A(B[767]), .Z(n3329) );
  IV U1509 ( .A(B[768]), .Z(n3328) );
  IV U1510 ( .A(B[769]), .Z(n3327) );
  IV U1511 ( .A(B[770]), .Z(n3326) );
  IV U1512 ( .A(B[771]), .Z(n3325) );
  IV U1513 ( .A(B[772]), .Z(n3324) );
  IV U1514 ( .A(B[773]), .Z(n3323) );
  IV U1515 ( .A(B[774]), .Z(n3322) );
  IV U1516 ( .A(B[775]), .Z(n3321) );
  IV U1517 ( .A(B[776]), .Z(n3320) );
  IV U1518 ( .A(B[3764]), .Z(n332) );
  IV U1519 ( .A(B[777]), .Z(n3319) );
  IV U1520 ( .A(B[778]), .Z(n3318) );
  IV U1521 ( .A(B[779]), .Z(n3317) );
  IV U1522 ( .A(B[780]), .Z(n3316) );
  IV U1523 ( .A(B[781]), .Z(n3315) );
  IV U1524 ( .A(B[782]), .Z(n3314) );
  IV U1525 ( .A(B[783]), .Z(n3313) );
  IV U1526 ( .A(B[784]), .Z(n3312) );
  IV U1527 ( .A(B[785]), .Z(n3311) );
  IV U1528 ( .A(B[786]), .Z(n3310) );
  IV U1529 ( .A(B[3765]), .Z(n331) );
  IV U1530 ( .A(B[787]), .Z(n3309) );
  IV U1531 ( .A(B[788]), .Z(n3308) );
  IV U1532 ( .A(B[789]), .Z(n3307) );
  IV U1533 ( .A(B[790]), .Z(n3306) );
  IV U1534 ( .A(B[791]), .Z(n3305) );
  IV U1535 ( .A(B[792]), .Z(n3304) );
  IV U1536 ( .A(B[793]), .Z(n3303) );
  IV U1537 ( .A(B[794]), .Z(n3302) );
  IV U1538 ( .A(B[795]), .Z(n3301) );
  IV U1539 ( .A(B[796]), .Z(n3300) );
  IV U1540 ( .A(B[3766]), .Z(n330) );
  IV U1541 ( .A(B[4063]), .Z(n33) );
  IV U1542 ( .A(B[797]), .Z(n3299) );
  IV U1543 ( .A(B[798]), .Z(n3298) );
  IV U1544 ( .A(B[799]), .Z(n3297) );
  IV U1545 ( .A(B[800]), .Z(n3296) );
  IV U1546 ( .A(B[801]), .Z(n3295) );
  IV U1547 ( .A(B[802]), .Z(n3294) );
  IV U1548 ( .A(B[803]), .Z(n3293) );
  IV U1549 ( .A(B[804]), .Z(n3292) );
  IV U1550 ( .A(B[805]), .Z(n3291) );
  IV U1551 ( .A(B[806]), .Z(n3290) );
  IV U1552 ( .A(B[3767]), .Z(n329) );
  IV U1553 ( .A(B[807]), .Z(n3289) );
  IV U1554 ( .A(B[808]), .Z(n3288) );
  IV U1555 ( .A(B[809]), .Z(n3287) );
  IV U1556 ( .A(B[810]), .Z(n3286) );
  IV U1557 ( .A(B[811]), .Z(n3285) );
  IV U1558 ( .A(B[812]), .Z(n3284) );
  IV U1559 ( .A(B[813]), .Z(n3283) );
  IV U1560 ( .A(B[814]), .Z(n3282) );
  IV U1561 ( .A(B[815]), .Z(n3281) );
  IV U1562 ( .A(B[816]), .Z(n3280) );
  IV U1563 ( .A(B[3768]), .Z(n328) );
  IV U1564 ( .A(B[817]), .Z(n3279) );
  IV U1565 ( .A(B[818]), .Z(n3278) );
  IV U1566 ( .A(B[819]), .Z(n3277) );
  IV U1567 ( .A(B[820]), .Z(n3276) );
  IV U1568 ( .A(B[821]), .Z(n3275) );
  IV U1569 ( .A(B[822]), .Z(n3274) );
  IV U1570 ( .A(B[823]), .Z(n3273) );
  IV U1571 ( .A(B[824]), .Z(n3272) );
  IV U1572 ( .A(B[825]), .Z(n3271) );
  IV U1573 ( .A(B[826]), .Z(n3270) );
  IV U1574 ( .A(B[3769]), .Z(n327) );
  IV U1575 ( .A(B[827]), .Z(n3269) );
  IV U1576 ( .A(B[828]), .Z(n3268) );
  IV U1577 ( .A(B[829]), .Z(n3267) );
  IV U1578 ( .A(B[830]), .Z(n3266) );
  IV U1579 ( .A(B[831]), .Z(n3265) );
  IV U1580 ( .A(B[832]), .Z(n3264) );
  IV U1581 ( .A(B[833]), .Z(n3263) );
  IV U1582 ( .A(B[834]), .Z(n3262) );
  IV U1583 ( .A(B[835]), .Z(n3261) );
  IV U1584 ( .A(B[836]), .Z(n3260) );
  IV U1585 ( .A(B[3770]), .Z(n326) );
  IV U1586 ( .A(B[837]), .Z(n3259) );
  IV U1587 ( .A(B[838]), .Z(n3258) );
  IV U1588 ( .A(B[839]), .Z(n3257) );
  IV U1589 ( .A(B[840]), .Z(n3256) );
  IV U1590 ( .A(B[841]), .Z(n3255) );
  IV U1591 ( .A(B[842]), .Z(n3254) );
  IV U1592 ( .A(B[843]), .Z(n3253) );
  IV U1593 ( .A(B[844]), .Z(n3252) );
  IV U1594 ( .A(B[845]), .Z(n3251) );
  IV U1595 ( .A(B[846]), .Z(n3250) );
  IV U1596 ( .A(B[3771]), .Z(n325) );
  IV U1597 ( .A(B[847]), .Z(n3249) );
  IV U1598 ( .A(B[848]), .Z(n3248) );
  IV U1599 ( .A(B[849]), .Z(n3247) );
  IV U1600 ( .A(B[850]), .Z(n3246) );
  IV U1601 ( .A(B[851]), .Z(n3245) );
  IV U1602 ( .A(B[852]), .Z(n3244) );
  IV U1603 ( .A(B[853]), .Z(n3243) );
  IV U1604 ( .A(B[854]), .Z(n3242) );
  IV U1605 ( .A(B[855]), .Z(n3241) );
  IV U1606 ( .A(B[856]), .Z(n3240) );
  IV U1607 ( .A(B[3772]), .Z(n324) );
  IV U1608 ( .A(B[857]), .Z(n3239) );
  IV U1609 ( .A(B[858]), .Z(n3238) );
  IV U1610 ( .A(B[859]), .Z(n3237) );
  IV U1611 ( .A(B[860]), .Z(n3236) );
  IV U1612 ( .A(B[861]), .Z(n3235) );
  IV U1613 ( .A(B[862]), .Z(n3234) );
  IV U1614 ( .A(B[863]), .Z(n3233) );
  IV U1615 ( .A(B[864]), .Z(n3232) );
  IV U1616 ( .A(B[865]), .Z(n3231) );
  IV U1617 ( .A(B[866]), .Z(n3230) );
  IV U1618 ( .A(B[3773]), .Z(n323) );
  IV U1619 ( .A(B[867]), .Z(n3229) );
  IV U1620 ( .A(B[868]), .Z(n3228) );
  IV U1621 ( .A(B[869]), .Z(n3227) );
  IV U1622 ( .A(B[870]), .Z(n3226) );
  IV U1623 ( .A(B[871]), .Z(n3225) );
  IV U1624 ( .A(B[872]), .Z(n3224) );
  IV U1625 ( .A(B[873]), .Z(n3223) );
  IV U1626 ( .A(B[874]), .Z(n3222) );
  IV U1627 ( .A(B[875]), .Z(n3221) );
  IV U1628 ( .A(B[876]), .Z(n3220) );
  IV U1629 ( .A(B[3774]), .Z(n322) );
  IV U1630 ( .A(B[877]), .Z(n3219) );
  IV U1631 ( .A(B[878]), .Z(n3218) );
  IV U1632 ( .A(B[879]), .Z(n3217) );
  IV U1633 ( .A(B[880]), .Z(n3216) );
  IV U1634 ( .A(B[881]), .Z(n3215) );
  IV U1635 ( .A(B[882]), .Z(n3214) );
  IV U1636 ( .A(B[883]), .Z(n3213) );
  IV U1637 ( .A(B[884]), .Z(n3212) );
  IV U1638 ( .A(B[885]), .Z(n3211) );
  IV U1639 ( .A(B[886]), .Z(n3210) );
  IV U1640 ( .A(B[3775]), .Z(n321) );
  IV U1641 ( .A(B[887]), .Z(n3209) );
  IV U1642 ( .A(B[888]), .Z(n3208) );
  IV U1643 ( .A(B[889]), .Z(n3207) );
  IV U1644 ( .A(B[890]), .Z(n3206) );
  IV U1645 ( .A(B[891]), .Z(n3205) );
  IV U1646 ( .A(B[892]), .Z(n3204) );
  IV U1647 ( .A(B[893]), .Z(n3203) );
  IV U1648 ( .A(B[894]), .Z(n3202) );
  IV U1649 ( .A(B[895]), .Z(n3201) );
  IV U1650 ( .A(B[896]), .Z(n3200) );
  IV U1651 ( .A(B[3776]), .Z(n320) );
  IV U1652 ( .A(B[4064]), .Z(n32) );
  IV U1653 ( .A(B[897]), .Z(n3199) );
  IV U1654 ( .A(B[898]), .Z(n3198) );
  IV U1655 ( .A(B[899]), .Z(n3197) );
  IV U1656 ( .A(B[900]), .Z(n3196) );
  IV U1657 ( .A(B[901]), .Z(n3195) );
  IV U1658 ( .A(B[902]), .Z(n3194) );
  IV U1659 ( .A(B[903]), .Z(n3193) );
  IV U1660 ( .A(B[904]), .Z(n3192) );
  IV U1661 ( .A(B[905]), .Z(n3191) );
  IV U1662 ( .A(B[906]), .Z(n3190) );
  IV U1663 ( .A(B[3777]), .Z(n319) );
  IV U1664 ( .A(B[907]), .Z(n3189) );
  IV U1665 ( .A(B[908]), .Z(n3188) );
  IV U1666 ( .A(B[909]), .Z(n3187) );
  IV U1667 ( .A(B[910]), .Z(n3186) );
  IV U1668 ( .A(B[911]), .Z(n3185) );
  IV U1669 ( .A(B[912]), .Z(n3184) );
  IV U1670 ( .A(B[913]), .Z(n3183) );
  IV U1671 ( .A(B[914]), .Z(n3182) );
  IV U1672 ( .A(B[915]), .Z(n3181) );
  IV U1673 ( .A(B[916]), .Z(n3180) );
  IV U1674 ( .A(B[3778]), .Z(n318) );
  IV U1675 ( .A(B[917]), .Z(n3179) );
  IV U1676 ( .A(B[918]), .Z(n3178) );
  IV U1677 ( .A(B[919]), .Z(n3177) );
  IV U1678 ( .A(B[920]), .Z(n3176) );
  IV U1679 ( .A(B[921]), .Z(n3175) );
  IV U1680 ( .A(B[922]), .Z(n3174) );
  IV U1681 ( .A(B[923]), .Z(n3173) );
  IV U1682 ( .A(B[924]), .Z(n3172) );
  IV U1683 ( .A(B[925]), .Z(n3171) );
  IV U1684 ( .A(B[926]), .Z(n3170) );
  IV U1685 ( .A(B[3779]), .Z(n317) );
  IV U1686 ( .A(B[927]), .Z(n3169) );
  IV U1687 ( .A(B[928]), .Z(n3168) );
  IV U1688 ( .A(B[929]), .Z(n3167) );
  IV U1689 ( .A(B[930]), .Z(n3166) );
  IV U1690 ( .A(B[931]), .Z(n3165) );
  IV U1691 ( .A(B[932]), .Z(n3164) );
  IV U1692 ( .A(B[933]), .Z(n3163) );
  IV U1693 ( .A(B[934]), .Z(n3162) );
  IV U1694 ( .A(B[935]), .Z(n3161) );
  IV U1695 ( .A(B[936]), .Z(n3160) );
  IV U1696 ( .A(B[3780]), .Z(n316) );
  IV U1697 ( .A(B[937]), .Z(n3159) );
  IV U1698 ( .A(B[938]), .Z(n3158) );
  IV U1699 ( .A(B[939]), .Z(n3157) );
  IV U1700 ( .A(B[940]), .Z(n3156) );
  IV U1701 ( .A(B[941]), .Z(n3155) );
  IV U1702 ( .A(B[942]), .Z(n3154) );
  IV U1703 ( .A(B[943]), .Z(n3153) );
  IV U1704 ( .A(B[944]), .Z(n3152) );
  IV U1705 ( .A(B[945]), .Z(n3151) );
  IV U1706 ( .A(B[946]), .Z(n3150) );
  IV U1707 ( .A(B[3781]), .Z(n315) );
  IV U1708 ( .A(B[947]), .Z(n3149) );
  IV U1709 ( .A(B[948]), .Z(n3148) );
  IV U1710 ( .A(B[949]), .Z(n3147) );
  IV U1711 ( .A(B[950]), .Z(n3146) );
  IV U1712 ( .A(B[951]), .Z(n3145) );
  IV U1713 ( .A(B[952]), .Z(n3144) );
  IV U1714 ( .A(B[953]), .Z(n3143) );
  IV U1715 ( .A(B[954]), .Z(n3142) );
  IV U1716 ( .A(B[955]), .Z(n3141) );
  IV U1717 ( .A(B[956]), .Z(n3140) );
  IV U1718 ( .A(B[3782]), .Z(n314) );
  IV U1719 ( .A(B[957]), .Z(n3139) );
  IV U1720 ( .A(B[958]), .Z(n3138) );
  IV U1721 ( .A(B[959]), .Z(n3137) );
  IV U1722 ( .A(B[960]), .Z(n3136) );
  IV U1723 ( .A(B[961]), .Z(n3135) );
  IV U1724 ( .A(B[962]), .Z(n3134) );
  IV U1725 ( .A(B[963]), .Z(n3133) );
  IV U1726 ( .A(B[964]), .Z(n3132) );
  IV U1727 ( .A(B[965]), .Z(n3131) );
  IV U1728 ( .A(B[966]), .Z(n3130) );
  IV U1729 ( .A(B[3783]), .Z(n313) );
  IV U1730 ( .A(B[967]), .Z(n3129) );
  IV U1731 ( .A(B[968]), .Z(n3128) );
  IV U1732 ( .A(B[969]), .Z(n3127) );
  IV U1733 ( .A(B[970]), .Z(n3126) );
  IV U1734 ( .A(B[971]), .Z(n3125) );
  IV U1735 ( .A(B[972]), .Z(n3124) );
  IV U1736 ( .A(B[973]), .Z(n3123) );
  IV U1737 ( .A(B[974]), .Z(n3122) );
  IV U1738 ( .A(B[975]), .Z(n3121) );
  IV U1739 ( .A(B[976]), .Z(n3120) );
  IV U1740 ( .A(B[3784]), .Z(n312) );
  IV U1741 ( .A(B[977]), .Z(n3119) );
  IV U1742 ( .A(B[978]), .Z(n3118) );
  IV U1743 ( .A(B[979]), .Z(n3117) );
  IV U1744 ( .A(B[980]), .Z(n3116) );
  IV U1745 ( .A(B[981]), .Z(n3115) );
  IV U1746 ( .A(B[982]), .Z(n3114) );
  IV U1747 ( .A(B[983]), .Z(n3113) );
  IV U1748 ( .A(B[984]), .Z(n3112) );
  IV U1749 ( .A(B[985]), .Z(n3111) );
  IV U1750 ( .A(B[986]), .Z(n3110) );
  IV U1751 ( .A(B[3785]), .Z(n311) );
  IV U1752 ( .A(B[987]), .Z(n3109) );
  IV U1753 ( .A(B[988]), .Z(n3108) );
  IV U1754 ( .A(B[989]), .Z(n3107) );
  IV U1755 ( .A(B[990]), .Z(n3106) );
  IV U1756 ( .A(B[991]), .Z(n3105) );
  IV U1757 ( .A(B[992]), .Z(n3104) );
  IV U1758 ( .A(B[993]), .Z(n3103) );
  IV U1759 ( .A(B[994]), .Z(n3102) );
  IV U1760 ( .A(B[995]), .Z(n3101) );
  IV U1761 ( .A(B[996]), .Z(n3100) );
  IV U1762 ( .A(B[3786]), .Z(n310) );
  IV U1763 ( .A(B[4065]), .Z(n31) );
  IV U1764 ( .A(B[997]), .Z(n3099) );
  IV U1765 ( .A(B[998]), .Z(n3098) );
  IV U1766 ( .A(B[999]), .Z(n3097) );
  IV U1767 ( .A(B[1000]), .Z(n3096) );
  IV U1768 ( .A(B[1001]), .Z(n3095) );
  IV U1769 ( .A(B[1002]), .Z(n3094) );
  IV U1770 ( .A(B[1003]), .Z(n3093) );
  IV U1771 ( .A(B[1004]), .Z(n3092) );
  IV U1772 ( .A(B[1005]), .Z(n3091) );
  IV U1773 ( .A(B[1006]), .Z(n3090) );
  IV U1774 ( .A(B[3787]), .Z(n309) );
  IV U1775 ( .A(B[1007]), .Z(n3089) );
  IV U1776 ( .A(B[1008]), .Z(n3088) );
  IV U1777 ( .A(B[1009]), .Z(n3087) );
  IV U1778 ( .A(B[1010]), .Z(n3086) );
  IV U1779 ( .A(B[1011]), .Z(n3085) );
  IV U1780 ( .A(B[1012]), .Z(n3084) );
  IV U1781 ( .A(B[1013]), .Z(n3083) );
  IV U1782 ( .A(B[1014]), .Z(n3082) );
  IV U1783 ( .A(B[1015]), .Z(n3081) );
  IV U1784 ( .A(B[1016]), .Z(n3080) );
  IV U1785 ( .A(B[3788]), .Z(n308) );
  IV U1786 ( .A(B[1017]), .Z(n3079) );
  IV U1787 ( .A(B[1018]), .Z(n3078) );
  IV U1788 ( .A(B[1019]), .Z(n3077) );
  IV U1789 ( .A(B[1020]), .Z(n3076) );
  IV U1790 ( .A(B[1021]), .Z(n3075) );
  IV U1791 ( .A(B[1022]), .Z(n3074) );
  IV U1792 ( .A(B[1023]), .Z(n3073) );
  IV U1793 ( .A(B[1024]), .Z(n3072) );
  IV U1794 ( .A(B[1025]), .Z(n3071) );
  IV U1795 ( .A(B[1026]), .Z(n3070) );
  IV U1796 ( .A(B[3789]), .Z(n307) );
  IV U1797 ( .A(B[1027]), .Z(n3069) );
  IV U1798 ( .A(B[1028]), .Z(n3068) );
  IV U1799 ( .A(B[1029]), .Z(n3067) );
  IV U1800 ( .A(B[1030]), .Z(n3066) );
  IV U1801 ( .A(B[1031]), .Z(n3065) );
  IV U1802 ( .A(B[1032]), .Z(n3064) );
  IV U1803 ( .A(B[1033]), .Z(n3063) );
  IV U1804 ( .A(B[1034]), .Z(n3062) );
  IV U1805 ( .A(B[1035]), .Z(n3061) );
  IV U1806 ( .A(B[1036]), .Z(n3060) );
  IV U1807 ( .A(B[3790]), .Z(n306) );
  IV U1808 ( .A(B[1037]), .Z(n3059) );
  IV U1809 ( .A(B[1038]), .Z(n3058) );
  IV U1810 ( .A(B[1039]), .Z(n3057) );
  IV U1811 ( .A(B[1040]), .Z(n3056) );
  IV U1812 ( .A(B[1041]), .Z(n3055) );
  IV U1813 ( .A(B[1042]), .Z(n3054) );
  IV U1814 ( .A(B[1043]), .Z(n3053) );
  IV U1815 ( .A(B[1044]), .Z(n3052) );
  IV U1816 ( .A(B[1045]), .Z(n3051) );
  IV U1817 ( .A(B[1046]), .Z(n3050) );
  IV U1818 ( .A(B[3791]), .Z(n305) );
  IV U1819 ( .A(B[1047]), .Z(n3049) );
  IV U1820 ( .A(B[1048]), .Z(n3048) );
  IV U1821 ( .A(B[1049]), .Z(n3047) );
  IV U1822 ( .A(B[1050]), .Z(n3046) );
  IV U1823 ( .A(B[1051]), .Z(n3045) );
  IV U1824 ( .A(B[1052]), .Z(n3044) );
  IV U1825 ( .A(B[1053]), .Z(n3043) );
  IV U1826 ( .A(B[1054]), .Z(n3042) );
  IV U1827 ( .A(B[1055]), .Z(n3041) );
  IV U1828 ( .A(B[1056]), .Z(n3040) );
  IV U1829 ( .A(B[3792]), .Z(n304) );
  IV U1830 ( .A(B[1057]), .Z(n3039) );
  IV U1831 ( .A(B[1058]), .Z(n3038) );
  IV U1832 ( .A(B[1059]), .Z(n3037) );
  IV U1833 ( .A(B[1060]), .Z(n3036) );
  IV U1834 ( .A(B[1061]), .Z(n3035) );
  IV U1835 ( .A(B[1062]), .Z(n3034) );
  IV U1836 ( .A(B[1063]), .Z(n3033) );
  IV U1837 ( .A(B[1064]), .Z(n3032) );
  IV U1838 ( .A(B[1065]), .Z(n3031) );
  IV U1839 ( .A(B[1066]), .Z(n3030) );
  IV U1840 ( .A(B[3793]), .Z(n303) );
  IV U1841 ( .A(B[1067]), .Z(n3029) );
  IV U1842 ( .A(B[1068]), .Z(n3028) );
  IV U1843 ( .A(B[1069]), .Z(n3027) );
  IV U1844 ( .A(B[1070]), .Z(n3026) );
  IV U1845 ( .A(B[1071]), .Z(n3025) );
  IV U1846 ( .A(B[1072]), .Z(n3024) );
  IV U1847 ( .A(B[1073]), .Z(n3023) );
  IV U1848 ( .A(B[1074]), .Z(n3022) );
  IV U1849 ( .A(B[1075]), .Z(n3021) );
  IV U1850 ( .A(B[1076]), .Z(n3020) );
  IV U1851 ( .A(B[3794]), .Z(n302) );
  IV U1852 ( .A(B[1077]), .Z(n3019) );
  IV U1853 ( .A(B[1078]), .Z(n3018) );
  IV U1854 ( .A(B[1079]), .Z(n3017) );
  IV U1855 ( .A(B[1080]), .Z(n3016) );
  IV U1856 ( .A(B[1081]), .Z(n3015) );
  IV U1857 ( .A(B[1082]), .Z(n3014) );
  IV U1858 ( .A(B[1083]), .Z(n3013) );
  IV U1859 ( .A(B[1084]), .Z(n3012) );
  IV U1860 ( .A(B[1085]), .Z(n3011) );
  IV U1861 ( .A(B[1086]), .Z(n3010) );
  IV U1862 ( .A(B[3795]), .Z(n301) );
  IV U1863 ( .A(B[1087]), .Z(n3009) );
  IV U1864 ( .A(B[1088]), .Z(n3008) );
  IV U1865 ( .A(B[1089]), .Z(n3007) );
  IV U1866 ( .A(B[1090]), .Z(n3006) );
  IV U1867 ( .A(B[1091]), .Z(n3005) );
  IV U1868 ( .A(B[1092]), .Z(n3004) );
  IV U1869 ( .A(B[1093]), .Z(n3003) );
  IV U1870 ( .A(B[1094]), .Z(n3002) );
  IV U1871 ( .A(B[1095]), .Z(n3001) );
  IV U1872 ( .A(B[1096]), .Z(n3000) );
  IV U1873 ( .A(B[3796]), .Z(n300) );
  IV U1874 ( .A(B[4066]), .Z(n30) );
  IV U1875 ( .A(B[4093]), .Z(n3) );
  IV U1876 ( .A(B[1097]), .Z(n2999) );
  IV U1877 ( .A(B[1098]), .Z(n2998) );
  IV U1878 ( .A(B[1099]), .Z(n2997) );
  IV U1879 ( .A(B[1100]), .Z(n2996) );
  IV U1880 ( .A(B[1101]), .Z(n2995) );
  IV U1881 ( .A(B[1102]), .Z(n2994) );
  IV U1882 ( .A(B[1103]), .Z(n2993) );
  IV U1883 ( .A(B[1104]), .Z(n2992) );
  IV U1884 ( .A(B[1105]), .Z(n2991) );
  IV U1885 ( .A(B[1106]), .Z(n2990) );
  IV U1886 ( .A(B[3797]), .Z(n299) );
  IV U1887 ( .A(B[1107]), .Z(n2989) );
  IV U1888 ( .A(B[1108]), .Z(n2988) );
  IV U1889 ( .A(B[1109]), .Z(n2987) );
  IV U1890 ( .A(B[1110]), .Z(n2986) );
  IV U1891 ( .A(B[1111]), .Z(n2985) );
  IV U1892 ( .A(B[1112]), .Z(n2984) );
  IV U1893 ( .A(B[1113]), .Z(n2983) );
  IV U1894 ( .A(B[1114]), .Z(n2982) );
  IV U1895 ( .A(B[1115]), .Z(n2981) );
  IV U1896 ( .A(B[1116]), .Z(n2980) );
  IV U1897 ( .A(B[3798]), .Z(n298) );
  IV U1898 ( .A(B[1117]), .Z(n2979) );
  IV U1899 ( .A(B[1118]), .Z(n2978) );
  IV U1900 ( .A(B[1119]), .Z(n2977) );
  IV U1901 ( .A(B[1120]), .Z(n2976) );
  IV U1902 ( .A(B[1121]), .Z(n2975) );
  IV U1903 ( .A(B[1122]), .Z(n2974) );
  IV U1904 ( .A(B[1123]), .Z(n2973) );
  IV U1905 ( .A(B[1124]), .Z(n2972) );
  IV U1906 ( .A(B[1125]), .Z(n2971) );
  IV U1907 ( .A(B[1126]), .Z(n2970) );
  IV U1908 ( .A(B[3799]), .Z(n297) );
  IV U1909 ( .A(B[1127]), .Z(n2969) );
  IV U1910 ( .A(B[1128]), .Z(n2968) );
  IV U1911 ( .A(B[1129]), .Z(n2967) );
  IV U1912 ( .A(B[1130]), .Z(n2966) );
  IV U1913 ( .A(B[1131]), .Z(n2965) );
  IV U1914 ( .A(B[1132]), .Z(n2964) );
  IV U1915 ( .A(B[1133]), .Z(n2963) );
  IV U1916 ( .A(B[1134]), .Z(n2962) );
  IV U1917 ( .A(B[1135]), .Z(n2961) );
  IV U1918 ( .A(B[1136]), .Z(n2960) );
  IV U1919 ( .A(B[3800]), .Z(n296) );
  IV U1920 ( .A(B[1137]), .Z(n2959) );
  IV U1921 ( .A(B[1138]), .Z(n2958) );
  IV U1922 ( .A(B[1139]), .Z(n2957) );
  IV U1923 ( .A(B[1140]), .Z(n2956) );
  IV U1924 ( .A(B[1141]), .Z(n2955) );
  IV U1925 ( .A(B[1142]), .Z(n2954) );
  IV U1926 ( .A(B[1143]), .Z(n2953) );
  IV U1927 ( .A(B[1144]), .Z(n2952) );
  IV U1928 ( .A(B[1145]), .Z(n2951) );
  IV U1929 ( .A(B[1146]), .Z(n2950) );
  IV U1930 ( .A(B[3801]), .Z(n295) );
  IV U1931 ( .A(B[1147]), .Z(n2949) );
  IV U1932 ( .A(B[1148]), .Z(n2948) );
  IV U1933 ( .A(B[1149]), .Z(n2947) );
  IV U1934 ( .A(B[1150]), .Z(n2946) );
  IV U1935 ( .A(B[1151]), .Z(n2945) );
  IV U1936 ( .A(B[1152]), .Z(n2944) );
  IV U1937 ( .A(B[1153]), .Z(n2943) );
  IV U1938 ( .A(B[1154]), .Z(n2942) );
  IV U1939 ( .A(B[1155]), .Z(n2941) );
  IV U1940 ( .A(B[1156]), .Z(n2940) );
  IV U1941 ( .A(B[3802]), .Z(n294) );
  IV U1942 ( .A(B[1157]), .Z(n2939) );
  IV U1943 ( .A(B[1158]), .Z(n2938) );
  IV U1944 ( .A(B[1159]), .Z(n2937) );
  IV U1945 ( .A(B[1160]), .Z(n2936) );
  IV U1946 ( .A(B[1161]), .Z(n2935) );
  IV U1947 ( .A(B[1162]), .Z(n2934) );
  IV U1948 ( .A(B[1163]), .Z(n2933) );
  IV U1949 ( .A(B[1164]), .Z(n2932) );
  IV U1950 ( .A(B[1165]), .Z(n2931) );
  IV U1951 ( .A(B[1166]), .Z(n2930) );
  IV U1952 ( .A(B[3803]), .Z(n293) );
  IV U1953 ( .A(B[1167]), .Z(n2929) );
  IV U1954 ( .A(B[1168]), .Z(n2928) );
  IV U1955 ( .A(B[1169]), .Z(n2927) );
  IV U1956 ( .A(B[1170]), .Z(n2926) );
  IV U1957 ( .A(B[1171]), .Z(n2925) );
  IV U1958 ( .A(B[1172]), .Z(n2924) );
  IV U1959 ( .A(B[1173]), .Z(n2923) );
  IV U1960 ( .A(B[1174]), .Z(n2922) );
  IV U1961 ( .A(B[1175]), .Z(n2921) );
  IV U1962 ( .A(B[1176]), .Z(n2920) );
  IV U1963 ( .A(B[3804]), .Z(n292) );
  IV U1964 ( .A(B[1177]), .Z(n2919) );
  IV U1965 ( .A(B[1178]), .Z(n2918) );
  IV U1966 ( .A(B[1179]), .Z(n2917) );
  IV U1967 ( .A(B[1180]), .Z(n2916) );
  IV U1968 ( .A(B[1181]), .Z(n2915) );
  IV U1969 ( .A(B[1182]), .Z(n2914) );
  IV U1970 ( .A(B[1183]), .Z(n2913) );
  IV U1971 ( .A(B[1184]), .Z(n2912) );
  IV U1972 ( .A(B[1185]), .Z(n2911) );
  IV U1973 ( .A(B[1186]), .Z(n2910) );
  IV U1974 ( .A(B[3805]), .Z(n291) );
  IV U1975 ( .A(B[1187]), .Z(n2909) );
  IV U1976 ( .A(B[1188]), .Z(n2908) );
  IV U1977 ( .A(B[1189]), .Z(n2907) );
  IV U1978 ( .A(B[1190]), .Z(n2906) );
  IV U1979 ( .A(B[1191]), .Z(n2905) );
  IV U1980 ( .A(B[1192]), .Z(n2904) );
  IV U1981 ( .A(B[1193]), .Z(n2903) );
  IV U1982 ( .A(B[1194]), .Z(n2902) );
  IV U1983 ( .A(B[1195]), .Z(n2901) );
  IV U1984 ( .A(B[1196]), .Z(n2900) );
  IV U1985 ( .A(B[3806]), .Z(n290) );
  IV U1986 ( .A(B[4067]), .Z(n29) );
  IV U1987 ( .A(B[1197]), .Z(n2899) );
  IV U1988 ( .A(B[1198]), .Z(n2898) );
  IV U1989 ( .A(B[1199]), .Z(n2897) );
  IV U1990 ( .A(B[1200]), .Z(n2896) );
  IV U1991 ( .A(B[1201]), .Z(n2895) );
  IV U1992 ( .A(B[1202]), .Z(n2894) );
  IV U1993 ( .A(B[1203]), .Z(n2893) );
  IV U1994 ( .A(B[1204]), .Z(n2892) );
  IV U1995 ( .A(B[1205]), .Z(n2891) );
  IV U1996 ( .A(B[1206]), .Z(n2890) );
  IV U1997 ( .A(B[3807]), .Z(n289) );
  IV U1998 ( .A(B[1207]), .Z(n2889) );
  IV U1999 ( .A(B[1208]), .Z(n2888) );
  IV U2000 ( .A(B[1209]), .Z(n2887) );
  IV U2001 ( .A(B[1210]), .Z(n2886) );
  IV U2002 ( .A(B[1211]), .Z(n2885) );
  IV U2003 ( .A(B[1212]), .Z(n2884) );
  IV U2004 ( .A(B[1213]), .Z(n2883) );
  IV U2005 ( .A(B[1214]), .Z(n2882) );
  IV U2006 ( .A(B[1215]), .Z(n2881) );
  IV U2007 ( .A(B[1216]), .Z(n2880) );
  IV U2008 ( .A(B[3808]), .Z(n288) );
  IV U2009 ( .A(B[1217]), .Z(n2879) );
  IV U2010 ( .A(B[1218]), .Z(n2878) );
  IV U2011 ( .A(B[1219]), .Z(n2877) );
  IV U2012 ( .A(B[1220]), .Z(n2876) );
  IV U2013 ( .A(B[1221]), .Z(n2875) );
  IV U2014 ( .A(B[1222]), .Z(n2874) );
  IV U2015 ( .A(B[1223]), .Z(n2873) );
  IV U2016 ( .A(B[1224]), .Z(n2872) );
  IV U2017 ( .A(B[1225]), .Z(n2871) );
  IV U2018 ( .A(B[1226]), .Z(n2870) );
  IV U2019 ( .A(B[3809]), .Z(n287) );
  IV U2020 ( .A(B[1227]), .Z(n2869) );
  IV U2021 ( .A(B[1228]), .Z(n2868) );
  IV U2022 ( .A(B[1229]), .Z(n2867) );
  IV U2023 ( .A(B[1230]), .Z(n2866) );
  IV U2024 ( .A(B[1231]), .Z(n2865) );
  IV U2025 ( .A(B[1232]), .Z(n2864) );
  IV U2026 ( .A(B[1233]), .Z(n2863) );
  IV U2027 ( .A(B[1234]), .Z(n2862) );
  IV U2028 ( .A(B[1235]), .Z(n2861) );
  IV U2029 ( .A(B[1236]), .Z(n2860) );
  IV U2030 ( .A(B[3810]), .Z(n286) );
  IV U2031 ( .A(B[1237]), .Z(n2859) );
  IV U2032 ( .A(B[1238]), .Z(n2858) );
  IV U2033 ( .A(B[1239]), .Z(n2857) );
  IV U2034 ( .A(B[1240]), .Z(n2856) );
  IV U2035 ( .A(B[1241]), .Z(n2855) );
  IV U2036 ( .A(B[1242]), .Z(n2854) );
  IV U2037 ( .A(B[1243]), .Z(n2853) );
  IV U2038 ( .A(B[1244]), .Z(n2852) );
  IV U2039 ( .A(B[1245]), .Z(n2851) );
  IV U2040 ( .A(B[1246]), .Z(n2850) );
  IV U2041 ( .A(B[3811]), .Z(n285) );
  IV U2042 ( .A(B[1247]), .Z(n2849) );
  IV U2043 ( .A(B[1248]), .Z(n2848) );
  IV U2044 ( .A(B[1249]), .Z(n2847) );
  IV U2045 ( .A(B[1250]), .Z(n2846) );
  IV U2046 ( .A(B[1251]), .Z(n2845) );
  IV U2047 ( .A(B[1252]), .Z(n2844) );
  IV U2048 ( .A(B[1253]), .Z(n2843) );
  IV U2049 ( .A(B[1254]), .Z(n2842) );
  IV U2050 ( .A(B[1255]), .Z(n2841) );
  IV U2051 ( .A(B[1256]), .Z(n2840) );
  IV U2052 ( .A(B[3812]), .Z(n284) );
  IV U2053 ( .A(B[1257]), .Z(n2839) );
  IV U2054 ( .A(B[1258]), .Z(n2838) );
  IV U2055 ( .A(B[1259]), .Z(n2837) );
  IV U2056 ( .A(B[1260]), .Z(n2836) );
  IV U2057 ( .A(B[1261]), .Z(n2835) );
  IV U2058 ( .A(B[1262]), .Z(n2834) );
  IV U2059 ( .A(B[1263]), .Z(n2833) );
  IV U2060 ( .A(B[1264]), .Z(n2832) );
  IV U2061 ( .A(B[1265]), .Z(n2831) );
  IV U2062 ( .A(B[1266]), .Z(n2830) );
  IV U2063 ( .A(B[3813]), .Z(n283) );
  IV U2064 ( .A(B[1267]), .Z(n2829) );
  IV U2065 ( .A(B[1268]), .Z(n2828) );
  IV U2066 ( .A(B[1269]), .Z(n2827) );
  IV U2067 ( .A(B[1270]), .Z(n2826) );
  IV U2068 ( .A(B[1271]), .Z(n2825) );
  IV U2069 ( .A(B[1272]), .Z(n2824) );
  IV U2070 ( .A(B[1273]), .Z(n2823) );
  IV U2071 ( .A(B[1274]), .Z(n2822) );
  IV U2072 ( .A(B[1275]), .Z(n2821) );
  IV U2073 ( .A(B[1276]), .Z(n2820) );
  IV U2074 ( .A(B[3814]), .Z(n282) );
  IV U2075 ( .A(B[1277]), .Z(n2819) );
  IV U2076 ( .A(B[1278]), .Z(n2818) );
  IV U2077 ( .A(B[1279]), .Z(n2817) );
  IV U2078 ( .A(B[1280]), .Z(n2816) );
  IV U2079 ( .A(B[1281]), .Z(n2815) );
  IV U2080 ( .A(B[1282]), .Z(n2814) );
  IV U2081 ( .A(B[1283]), .Z(n2813) );
  IV U2082 ( .A(B[1284]), .Z(n2812) );
  IV U2083 ( .A(B[1285]), .Z(n2811) );
  IV U2084 ( .A(B[1286]), .Z(n2810) );
  IV U2085 ( .A(B[3815]), .Z(n281) );
  IV U2086 ( .A(B[1287]), .Z(n2809) );
  IV U2087 ( .A(B[1288]), .Z(n2808) );
  IV U2088 ( .A(B[1289]), .Z(n2807) );
  IV U2089 ( .A(B[1290]), .Z(n2806) );
  IV U2090 ( .A(B[1291]), .Z(n2805) );
  IV U2091 ( .A(B[1292]), .Z(n2804) );
  IV U2092 ( .A(B[1293]), .Z(n2803) );
  IV U2093 ( .A(B[1294]), .Z(n2802) );
  IV U2094 ( .A(B[1295]), .Z(n2801) );
  IV U2095 ( .A(B[1296]), .Z(n2800) );
  IV U2096 ( .A(B[3816]), .Z(n280) );
  IV U2097 ( .A(B[4068]), .Z(n28) );
  IV U2098 ( .A(B[1297]), .Z(n2799) );
  IV U2099 ( .A(B[1298]), .Z(n2798) );
  IV U2100 ( .A(B[1299]), .Z(n2797) );
  IV U2101 ( .A(B[1300]), .Z(n2796) );
  IV U2102 ( .A(B[1301]), .Z(n2795) );
  IV U2103 ( .A(B[1302]), .Z(n2794) );
  IV U2104 ( .A(B[1303]), .Z(n2793) );
  IV U2105 ( .A(B[1304]), .Z(n2792) );
  IV U2106 ( .A(B[1305]), .Z(n2791) );
  IV U2107 ( .A(B[1306]), .Z(n2790) );
  IV U2108 ( .A(B[3817]), .Z(n279) );
  IV U2109 ( .A(B[1307]), .Z(n2789) );
  IV U2110 ( .A(B[1308]), .Z(n2788) );
  IV U2111 ( .A(B[1309]), .Z(n2787) );
  IV U2112 ( .A(B[1310]), .Z(n2786) );
  IV U2113 ( .A(B[1311]), .Z(n2785) );
  IV U2114 ( .A(B[1312]), .Z(n2784) );
  IV U2115 ( .A(B[1313]), .Z(n2783) );
  IV U2116 ( .A(B[1314]), .Z(n2782) );
  IV U2117 ( .A(B[1315]), .Z(n2781) );
  IV U2118 ( .A(B[1316]), .Z(n2780) );
  IV U2119 ( .A(B[3818]), .Z(n278) );
  IV U2120 ( .A(B[1317]), .Z(n2779) );
  IV U2121 ( .A(B[1318]), .Z(n2778) );
  IV U2122 ( .A(B[1319]), .Z(n2777) );
  IV U2123 ( .A(B[1320]), .Z(n2776) );
  IV U2124 ( .A(B[1321]), .Z(n2775) );
  IV U2125 ( .A(B[1322]), .Z(n2774) );
  IV U2126 ( .A(B[1323]), .Z(n2773) );
  IV U2127 ( .A(B[1324]), .Z(n2772) );
  IV U2128 ( .A(B[1325]), .Z(n2771) );
  IV U2129 ( .A(B[1326]), .Z(n2770) );
  IV U2130 ( .A(B[3819]), .Z(n277) );
  IV U2131 ( .A(B[1327]), .Z(n2769) );
  IV U2132 ( .A(B[1328]), .Z(n2768) );
  IV U2133 ( .A(B[1329]), .Z(n2767) );
  IV U2134 ( .A(B[1330]), .Z(n2766) );
  IV U2135 ( .A(B[1331]), .Z(n2765) );
  IV U2136 ( .A(B[1332]), .Z(n2764) );
  IV U2137 ( .A(B[1333]), .Z(n2763) );
  IV U2138 ( .A(B[1334]), .Z(n2762) );
  IV U2139 ( .A(B[1335]), .Z(n2761) );
  IV U2140 ( .A(B[1336]), .Z(n2760) );
  IV U2141 ( .A(B[3820]), .Z(n276) );
  IV U2142 ( .A(B[1337]), .Z(n2759) );
  IV U2143 ( .A(B[1338]), .Z(n2758) );
  IV U2144 ( .A(B[1339]), .Z(n2757) );
  IV U2145 ( .A(B[1340]), .Z(n2756) );
  IV U2146 ( .A(B[1341]), .Z(n2755) );
  IV U2147 ( .A(B[1342]), .Z(n2754) );
  IV U2148 ( .A(B[1343]), .Z(n2753) );
  IV U2149 ( .A(B[1344]), .Z(n2752) );
  IV U2150 ( .A(B[1345]), .Z(n2751) );
  IV U2151 ( .A(B[1346]), .Z(n2750) );
  IV U2152 ( .A(B[3821]), .Z(n275) );
  IV U2153 ( .A(B[1347]), .Z(n2749) );
  IV U2154 ( .A(B[1348]), .Z(n2748) );
  IV U2155 ( .A(B[1349]), .Z(n2747) );
  IV U2156 ( .A(B[1350]), .Z(n2746) );
  IV U2157 ( .A(B[1351]), .Z(n2745) );
  IV U2158 ( .A(B[1352]), .Z(n2744) );
  IV U2159 ( .A(B[1353]), .Z(n2743) );
  IV U2160 ( .A(B[1354]), .Z(n2742) );
  IV U2161 ( .A(B[1355]), .Z(n2741) );
  IV U2162 ( .A(B[1356]), .Z(n2740) );
  IV U2163 ( .A(B[3822]), .Z(n274) );
  IV U2164 ( .A(B[1357]), .Z(n2739) );
  IV U2165 ( .A(B[1358]), .Z(n2738) );
  IV U2166 ( .A(B[1359]), .Z(n2737) );
  IV U2167 ( .A(B[1360]), .Z(n2736) );
  IV U2168 ( .A(B[1361]), .Z(n2735) );
  IV U2169 ( .A(B[1362]), .Z(n2734) );
  IV U2170 ( .A(B[1363]), .Z(n2733) );
  IV U2171 ( .A(B[1364]), .Z(n2732) );
  IV U2172 ( .A(B[1365]), .Z(n2731) );
  IV U2173 ( .A(B[1366]), .Z(n2730) );
  IV U2174 ( .A(B[3823]), .Z(n273) );
  IV U2175 ( .A(B[1367]), .Z(n2729) );
  IV U2176 ( .A(B[1368]), .Z(n2728) );
  IV U2177 ( .A(B[1369]), .Z(n2727) );
  IV U2178 ( .A(B[1370]), .Z(n2726) );
  IV U2179 ( .A(B[1371]), .Z(n2725) );
  IV U2180 ( .A(B[1372]), .Z(n2724) );
  IV U2181 ( .A(B[1373]), .Z(n2723) );
  IV U2182 ( .A(B[1374]), .Z(n2722) );
  IV U2183 ( .A(B[1375]), .Z(n2721) );
  IV U2184 ( .A(B[1376]), .Z(n2720) );
  IV U2185 ( .A(B[3824]), .Z(n272) );
  IV U2186 ( .A(B[1377]), .Z(n2719) );
  IV U2187 ( .A(B[1378]), .Z(n2718) );
  IV U2188 ( .A(B[1379]), .Z(n2717) );
  IV U2189 ( .A(B[1380]), .Z(n2716) );
  IV U2190 ( .A(B[1381]), .Z(n2715) );
  IV U2191 ( .A(B[1382]), .Z(n2714) );
  IV U2192 ( .A(B[1383]), .Z(n2713) );
  IV U2193 ( .A(B[1384]), .Z(n2712) );
  IV U2194 ( .A(B[1385]), .Z(n2711) );
  IV U2195 ( .A(B[1386]), .Z(n2710) );
  IV U2196 ( .A(B[3825]), .Z(n271) );
  IV U2197 ( .A(B[1387]), .Z(n2709) );
  IV U2198 ( .A(B[1388]), .Z(n2708) );
  IV U2199 ( .A(B[1389]), .Z(n2707) );
  IV U2200 ( .A(B[1390]), .Z(n2706) );
  IV U2201 ( .A(B[1391]), .Z(n2705) );
  IV U2202 ( .A(B[1392]), .Z(n2704) );
  IV U2203 ( .A(B[1393]), .Z(n2703) );
  IV U2204 ( .A(B[1394]), .Z(n2702) );
  IV U2205 ( .A(B[1395]), .Z(n2701) );
  IV U2206 ( .A(B[1396]), .Z(n2700) );
  IV U2207 ( .A(B[3826]), .Z(n270) );
  IV U2208 ( .A(B[4069]), .Z(n27) );
  IV U2209 ( .A(B[1397]), .Z(n2699) );
  IV U2210 ( .A(B[1398]), .Z(n2698) );
  IV U2211 ( .A(B[1399]), .Z(n2697) );
  IV U2212 ( .A(B[1400]), .Z(n2696) );
  IV U2213 ( .A(B[1401]), .Z(n2695) );
  IV U2214 ( .A(B[1402]), .Z(n2694) );
  IV U2215 ( .A(B[1403]), .Z(n2693) );
  IV U2216 ( .A(B[1404]), .Z(n2692) );
  IV U2217 ( .A(B[1405]), .Z(n2691) );
  IV U2218 ( .A(B[1406]), .Z(n2690) );
  IV U2219 ( .A(B[3827]), .Z(n269) );
  IV U2220 ( .A(B[1407]), .Z(n2689) );
  IV U2221 ( .A(B[1408]), .Z(n2688) );
  IV U2222 ( .A(B[1409]), .Z(n2687) );
  IV U2223 ( .A(B[1410]), .Z(n2686) );
  IV U2224 ( .A(B[1411]), .Z(n2685) );
  IV U2225 ( .A(B[1412]), .Z(n2684) );
  IV U2226 ( .A(B[1413]), .Z(n2683) );
  IV U2227 ( .A(B[1414]), .Z(n2682) );
  IV U2228 ( .A(B[1415]), .Z(n2681) );
  IV U2229 ( .A(B[1416]), .Z(n2680) );
  IV U2230 ( .A(B[3828]), .Z(n268) );
  IV U2231 ( .A(B[1417]), .Z(n2679) );
  IV U2232 ( .A(B[1418]), .Z(n2678) );
  IV U2233 ( .A(B[1419]), .Z(n2677) );
  IV U2234 ( .A(B[1420]), .Z(n2676) );
  IV U2235 ( .A(B[1421]), .Z(n2675) );
  IV U2236 ( .A(B[1422]), .Z(n2674) );
  IV U2237 ( .A(B[1423]), .Z(n2673) );
  IV U2238 ( .A(B[1424]), .Z(n2672) );
  IV U2239 ( .A(B[1425]), .Z(n2671) );
  IV U2240 ( .A(B[1426]), .Z(n2670) );
  IV U2241 ( .A(B[3829]), .Z(n267) );
  IV U2242 ( .A(B[1427]), .Z(n2669) );
  IV U2243 ( .A(B[1428]), .Z(n2668) );
  IV U2244 ( .A(B[1429]), .Z(n2667) );
  IV U2245 ( .A(B[1430]), .Z(n2666) );
  IV U2246 ( .A(B[1431]), .Z(n2665) );
  IV U2247 ( .A(B[1432]), .Z(n2664) );
  IV U2248 ( .A(B[1433]), .Z(n2663) );
  IV U2249 ( .A(B[1434]), .Z(n2662) );
  IV U2250 ( .A(B[1435]), .Z(n2661) );
  IV U2251 ( .A(B[1436]), .Z(n2660) );
  IV U2252 ( .A(B[3830]), .Z(n266) );
  IV U2253 ( .A(B[1437]), .Z(n2659) );
  IV U2254 ( .A(B[1438]), .Z(n2658) );
  IV U2255 ( .A(B[1439]), .Z(n2657) );
  IV U2256 ( .A(B[1440]), .Z(n2656) );
  IV U2257 ( .A(B[1441]), .Z(n2655) );
  IV U2258 ( .A(B[1442]), .Z(n2654) );
  IV U2259 ( .A(B[1443]), .Z(n2653) );
  IV U2260 ( .A(B[1444]), .Z(n2652) );
  IV U2261 ( .A(B[1445]), .Z(n2651) );
  IV U2262 ( .A(B[1446]), .Z(n2650) );
  IV U2263 ( .A(B[3831]), .Z(n265) );
  IV U2264 ( .A(B[1447]), .Z(n2649) );
  IV U2265 ( .A(B[1448]), .Z(n2648) );
  IV U2266 ( .A(B[1449]), .Z(n2647) );
  IV U2267 ( .A(B[1450]), .Z(n2646) );
  IV U2268 ( .A(B[1451]), .Z(n2645) );
  IV U2269 ( .A(B[1452]), .Z(n2644) );
  IV U2270 ( .A(B[1453]), .Z(n2643) );
  IV U2271 ( .A(B[1454]), .Z(n2642) );
  IV U2272 ( .A(B[1455]), .Z(n2641) );
  IV U2273 ( .A(B[1456]), .Z(n2640) );
  IV U2274 ( .A(B[3832]), .Z(n264) );
  IV U2275 ( .A(B[1457]), .Z(n2639) );
  IV U2276 ( .A(B[1458]), .Z(n2638) );
  IV U2277 ( .A(B[1459]), .Z(n2637) );
  IV U2278 ( .A(B[1460]), .Z(n2636) );
  IV U2279 ( .A(B[1461]), .Z(n2635) );
  IV U2280 ( .A(B[1462]), .Z(n2634) );
  IV U2281 ( .A(B[1463]), .Z(n2633) );
  IV U2282 ( .A(B[1464]), .Z(n2632) );
  IV U2283 ( .A(B[1465]), .Z(n2631) );
  IV U2284 ( .A(B[1466]), .Z(n2630) );
  IV U2285 ( .A(B[3833]), .Z(n263) );
  IV U2286 ( .A(B[1467]), .Z(n2629) );
  IV U2287 ( .A(B[1468]), .Z(n2628) );
  IV U2288 ( .A(B[1469]), .Z(n2627) );
  IV U2289 ( .A(B[1470]), .Z(n2626) );
  IV U2290 ( .A(B[1471]), .Z(n2625) );
  IV U2291 ( .A(B[1472]), .Z(n2624) );
  IV U2292 ( .A(B[1473]), .Z(n2623) );
  IV U2293 ( .A(B[1474]), .Z(n2622) );
  IV U2294 ( .A(B[1475]), .Z(n2621) );
  IV U2295 ( .A(B[1476]), .Z(n2620) );
  IV U2296 ( .A(B[3834]), .Z(n262) );
  IV U2297 ( .A(B[1477]), .Z(n2619) );
  IV U2298 ( .A(B[1478]), .Z(n2618) );
  IV U2299 ( .A(B[1479]), .Z(n2617) );
  IV U2300 ( .A(B[1480]), .Z(n2616) );
  IV U2301 ( .A(B[1481]), .Z(n2615) );
  IV U2302 ( .A(B[1482]), .Z(n2614) );
  IV U2303 ( .A(B[1483]), .Z(n2613) );
  IV U2304 ( .A(B[1484]), .Z(n2612) );
  IV U2305 ( .A(B[1485]), .Z(n2611) );
  IV U2306 ( .A(B[1486]), .Z(n2610) );
  IV U2307 ( .A(B[3835]), .Z(n261) );
  IV U2308 ( .A(B[1487]), .Z(n2609) );
  IV U2309 ( .A(B[1488]), .Z(n2608) );
  IV U2310 ( .A(B[1489]), .Z(n2607) );
  IV U2311 ( .A(B[1490]), .Z(n2606) );
  IV U2312 ( .A(B[1491]), .Z(n2605) );
  IV U2313 ( .A(B[1492]), .Z(n2604) );
  IV U2314 ( .A(B[1493]), .Z(n2603) );
  IV U2315 ( .A(B[1494]), .Z(n2602) );
  IV U2316 ( .A(B[1495]), .Z(n2601) );
  IV U2317 ( .A(B[1496]), .Z(n2600) );
  IV U2318 ( .A(B[3836]), .Z(n260) );
  IV U2319 ( .A(B[4070]), .Z(n26) );
  IV U2320 ( .A(B[1497]), .Z(n2599) );
  IV U2321 ( .A(B[1498]), .Z(n2598) );
  IV U2322 ( .A(B[1499]), .Z(n2597) );
  IV U2323 ( .A(B[1500]), .Z(n2596) );
  IV U2324 ( .A(B[1501]), .Z(n2595) );
  IV U2325 ( .A(B[1502]), .Z(n2594) );
  IV U2326 ( .A(B[1503]), .Z(n2593) );
  IV U2327 ( .A(B[1504]), .Z(n2592) );
  IV U2328 ( .A(B[1505]), .Z(n2591) );
  IV U2329 ( .A(B[1506]), .Z(n2590) );
  IV U2330 ( .A(B[3837]), .Z(n259) );
  IV U2331 ( .A(B[1507]), .Z(n2589) );
  IV U2332 ( .A(B[1508]), .Z(n2588) );
  IV U2333 ( .A(B[1509]), .Z(n2587) );
  IV U2334 ( .A(B[1510]), .Z(n2586) );
  IV U2335 ( .A(B[1511]), .Z(n2585) );
  IV U2336 ( .A(B[1512]), .Z(n2584) );
  IV U2337 ( .A(B[1513]), .Z(n2583) );
  IV U2338 ( .A(B[1514]), .Z(n2582) );
  IV U2339 ( .A(B[1515]), .Z(n2581) );
  IV U2340 ( .A(B[1516]), .Z(n2580) );
  IV U2341 ( .A(B[3838]), .Z(n258) );
  IV U2342 ( .A(B[1517]), .Z(n2579) );
  IV U2343 ( .A(B[1518]), .Z(n2578) );
  IV U2344 ( .A(B[1519]), .Z(n2577) );
  IV U2345 ( .A(B[1520]), .Z(n2576) );
  IV U2346 ( .A(B[1521]), .Z(n2575) );
  IV U2347 ( .A(B[1522]), .Z(n2574) );
  IV U2348 ( .A(B[1523]), .Z(n2573) );
  IV U2349 ( .A(B[1524]), .Z(n2572) );
  IV U2350 ( .A(B[1525]), .Z(n2571) );
  IV U2351 ( .A(B[1526]), .Z(n2570) );
  IV U2352 ( .A(B[3839]), .Z(n257) );
  IV U2353 ( .A(B[1527]), .Z(n2569) );
  IV U2354 ( .A(B[1528]), .Z(n2568) );
  IV U2355 ( .A(B[1529]), .Z(n2567) );
  IV U2356 ( .A(B[1530]), .Z(n2566) );
  IV U2357 ( .A(B[1531]), .Z(n2565) );
  IV U2358 ( .A(B[1532]), .Z(n2564) );
  IV U2359 ( .A(B[1533]), .Z(n2563) );
  IV U2360 ( .A(B[1534]), .Z(n2562) );
  IV U2361 ( .A(B[1535]), .Z(n2561) );
  IV U2362 ( .A(B[1536]), .Z(n2560) );
  IV U2363 ( .A(B[3840]), .Z(n256) );
  IV U2364 ( .A(B[1537]), .Z(n2559) );
  IV U2365 ( .A(B[1538]), .Z(n2558) );
  IV U2366 ( .A(B[1539]), .Z(n2557) );
  IV U2367 ( .A(B[1540]), .Z(n2556) );
  IV U2368 ( .A(B[1541]), .Z(n2555) );
  IV U2369 ( .A(B[1542]), .Z(n2554) );
  IV U2370 ( .A(B[1543]), .Z(n2553) );
  IV U2371 ( .A(B[1544]), .Z(n2552) );
  IV U2372 ( .A(B[1545]), .Z(n2551) );
  IV U2373 ( .A(B[1546]), .Z(n2550) );
  IV U2374 ( .A(B[3841]), .Z(n255) );
  IV U2375 ( .A(B[1547]), .Z(n2549) );
  IV U2376 ( .A(B[1548]), .Z(n2548) );
  IV U2377 ( .A(B[1549]), .Z(n2547) );
  IV U2378 ( .A(B[1550]), .Z(n2546) );
  IV U2379 ( .A(B[1551]), .Z(n2545) );
  IV U2380 ( .A(B[1552]), .Z(n2544) );
  IV U2381 ( .A(B[1553]), .Z(n2543) );
  IV U2382 ( .A(B[1554]), .Z(n2542) );
  IV U2383 ( .A(B[1555]), .Z(n2541) );
  IV U2384 ( .A(B[1556]), .Z(n2540) );
  IV U2385 ( .A(B[3842]), .Z(n254) );
  IV U2386 ( .A(B[1557]), .Z(n2539) );
  IV U2387 ( .A(B[1558]), .Z(n2538) );
  IV U2388 ( .A(B[1559]), .Z(n2537) );
  IV U2389 ( .A(B[1560]), .Z(n2536) );
  IV U2390 ( .A(B[1561]), .Z(n2535) );
  IV U2391 ( .A(B[1562]), .Z(n2534) );
  IV U2392 ( .A(B[1563]), .Z(n2533) );
  IV U2393 ( .A(B[1564]), .Z(n2532) );
  IV U2394 ( .A(B[1565]), .Z(n2531) );
  IV U2395 ( .A(B[1566]), .Z(n2530) );
  IV U2396 ( .A(B[3843]), .Z(n253) );
  IV U2397 ( .A(B[1567]), .Z(n2529) );
  IV U2398 ( .A(B[1568]), .Z(n2528) );
  IV U2399 ( .A(B[1569]), .Z(n2527) );
  IV U2400 ( .A(B[1570]), .Z(n2526) );
  IV U2401 ( .A(B[1571]), .Z(n2525) );
  IV U2402 ( .A(B[1572]), .Z(n2524) );
  IV U2403 ( .A(B[1573]), .Z(n2523) );
  IV U2404 ( .A(B[1574]), .Z(n2522) );
  IV U2405 ( .A(B[1575]), .Z(n2521) );
  IV U2406 ( .A(B[1576]), .Z(n2520) );
  IV U2407 ( .A(B[3844]), .Z(n252) );
  IV U2408 ( .A(B[1577]), .Z(n2519) );
  IV U2409 ( .A(B[1578]), .Z(n2518) );
  IV U2410 ( .A(B[1579]), .Z(n2517) );
  IV U2411 ( .A(B[1580]), .Z(n2516) );
  IV U2412 ( .A(B[1581]), .Z(n2515) );
  IV U2413 ( .A(B[1582]), .Z(n2514) );
  IV U2414 ( .A(B[1583]), .Z(n2513) );
  IV U2415 ( .A(B[1584]), .Z(n2512) );
  IV U2416 ( .A(B[1585]), .Z(n2511) );
  IV U2417 ( .A(B[1586]), .Z(n2510) );
  IV U2418 ( .A(B[3845]), .Z(n251) );
  IV U2419 ( .A(B[1587]), .Z(n2509) );
  IV U2420 ( .A(B[1588]), .Z(n2508) );
  IV U2421 ( .A(B[1589]), .Z(n2507) );
  IV U2422 ( .A(B[1590]), .Z(n2506) );
  IV U2423 ( .A(B[1591]), .Z(n2505) );
  IV U2424 ( .A(B[1592]), .Z(n2504) );
  IV U2425 ( .A(B[1593]), .Z(n2503) );
  IV U2426 ( .A(B[1594]), .Z(n2502) );
  IV U2427 ( .A(B[1595]), .Z(n2501) );
  IV U2428 ( .A(B[1596]), .Z(n2500) );
  IV U2429 ( .A(B[3846]), .Z(n250) );
  IV U2430 ( .A(B[4071]), .Z(n25) );
  IV U2431 ( .A(B[1597]), .Z(n2499) );
  IV U2432 ( .A(B[1598]), .Z(n2498) );
  IV U2433 ( .A(B[1599]), .Z(n2497) );
  IV U2434 ( .A(B[1600]), .Z(n2496) );
  IV U2435 ( .A(B[1601]), .Z(n2495) );
  IV U2436 ( .A(B[1602]), .Z(n2494) );
  IV U2437 ( .A(B[1603]), .Z(n2493) );
  IV U2438 ( .A(B[1604]), .Z(n2492) );
  IV U2439 ( .A(B[1605]), .Z(n2491) );
  IV U2440 ( .A(B[1606]), .Z(n2490) );
  IV U2441 ( .A(B[3847]), .Z(n249) );
  IV U2442 ( .A(B[1607]), .Z(n2489) );
  IV U2443 ( .A(B[1608]), .Z(n2488) );
  IV U2444 ( .A(B[1609]), .Z(n2487) );
  IV U2445 ( .A(B[1610]), .Z(n2486) );
  IV U2446 ( .A(B[1611]), .Z(n2485) );
  IV U2447 ( .A(B[1612]), .Z(n2484) );
  IV U2448 ( .A(B[1613]), .Z(n2483) );
  IV U2449 ( .A(B[1614]), .Z(n2482) );
  IV U2450 ( .A(B[1615]), .Z(n2481) );
  IV U2451 ( .A(B[1616]), .Z(n2480) );
  IV U2452 ( .A(B[3848]), .Z(n248) );
  IV U2453 ( .A(B[1617]), .Z(n2479) );
  IV U2454 ( .A(B[1618]), .Z(n2478) );
  IV U2455 ( .A(B[1619]), .Z(n2477) );
  IV U2456 ( .A(B[1620]), .Z(n2476) );
  IV U2457 ( .A(B[1621]), .Z(n2475) );
  IV U2458 ( .A(B[1622]), .Z(n2474) );
  IV U2459 ( .A(B[1623]), .Z(n2473) );
  IV U2460 ( .A(B[1624]), .Z(n2472) );
  IV U2461 ( .A(B[1625]), .Z(n2471) );
  IV U2462 ( .A(B[1626]), .Z(n2470) );
  IV U2463 ( .A(B[3849]), .Z(n247) );
  IV U2464 ( .A(B[1627]), .Z(n2469) );
  IV U2465 ( .A(B[1628]), .Z(n2468) );
  IV U2466 ( .A(B[1629]), .Z(n2467) );
  IV U2467 ( .A(B[1630]), .Z(n2466) );
  IV U2468 ( .A(B[1631]), .Z(n2465) );
  IV U2469 ( .A(B[1632]), .Z(n2464) );
  IV U2470 ( .A(B[1633]), .Z(n2463) );
  IV U2471 ( .A(B[1634]), .Z(n2462) );
  IV U2472 ( .A(B[1635]), .Z(n2461) );
  IV U2473 ( .A(B[1636]), .Z(n2460) );
  IV U2474 ( .A(B[3850]), .Z(n246) );
  IV U2475 ( .A(B[1637]), .Z(n2459) );
  IV U2476 ( .A(B[1638]), .Z(n2458) );
  IV U2477 ( .A(B[1639]), .Z(n2457) );
  IV U2478 ( .A(B[1640]), .Z(n2456) );
  IV U2479 ( .A(B[1641]), .Z(n2455) );
  IV U2480 ( .A(B[1642]), .Z(n2454) );
  IV U2481 ( .A(B[1643]), .Z(n2453) );
  IV U2482 ( .A(B[1644]), .Z(n2452) );
  IV U2483 ( .A(B[1645]), .Z(n2451) );
  IV U2484 ( .A(B[1646]), .Z(n2450) );
  IV U2485 ( .A(B[3851]), .Z(n245) );
  IV U2486 ( .A(B[1647]), .Z(n2449) );
  IV U2487 ( .A(B[1648]), .Z(n2448) );
  IV U2488 ( .A(B[1649]), .Z(n2447) );
  IV U2489 ( .A(B[1650]), .Z(n2446) );
  IV U2490 ( .A(B[1651]), .Z(n2445) );
  IV U2491 ( .A(B[1652]), .Z(n2444) );
  IV U2492 ( .A(B[1653]), .Z(n2443) );
  IV U2493 ( .A(B[1654]), .Z(n2442) );
  IV U2494 ( .A(B[1655]), .Z(n2441) );
  IV U2495 ( .A(B[1656]), .Z(n2440) );
  IV U2496 ( .A(B[3852]), .Z(n244) );
  IV U2497 ( .A(B[1657]), .Z(n2439) );
  IV U2498 ( .A(B[1658]), .Z(n2438) );
  IV U2499 ( .A(B[1659]), .Z(n2437) );
  IV U2500 ( .A(B[1660]), .Z(n2436) );
  IV U2501 ( .A(B[1661]), .Z(n2435) );
  IV U2502 ( .A(B[1662]), .Z(n2434) );
  IV U2503 ( .A(B[1663]), .Z(n2433) );
  IV U2504 ( .A(B[1664]), .Z(n2432) );
  IV U2505 ( .A(B[1665]), .Z(n2431) );
  IV U2506 ( .A(B[1666]), .Z(n2430) );
  IV U2507 ( .A(B[3853]), .Z(n243) );
  IV U2508 ( .A(B[1667]), .Z(n2429) );
  IV U2509 ( .A(B[1668]), .Z(n2428) );
  IV U2510 ( .A(B[1669]), .Z(n2427) );
  IV U2511 ( .A(B[1670]), .Z(n2426) );
  IV U2512 ( .A(B[1671]), .Z(n2425) );
  IV U2513 ( .A(B[1672]), .Z(n2424) );
  IV U2514 ( .A(B[1673]), .Z(n2423) );
  IV U2515 ( .A(B[1674]), .Z(n2422) );
  IV U2516 ( .A(B[1675]), .Z(n2421) );
  IV U2517 ( .A(B[1676]), .Z(n2420) );
  IV U2518 ( .A(B[3854]), .Z(n242) );
  IV U2519 ( .A(B[1677]), .Z(n2419) );
  IV U2520 ( .A(B[1678]), .Z(n2418) );
  IV U2521 ( .A(B[1679]), .Z(n2417) );
  IV U2522 ( .A(B[1680]), .Z(n2416) );
  IV U2523 ( .A(B[1681]), .Z(n2415) );
  IV U2524 ( .A(B[1682]), .Z(n2414) );
  IV U2525 ( .A(B[1683]), .Z(n2413) );
  IV U2526 ( .A(B[1684]), .Z(n2412) );
  IV U2527 ( .A(B[1685]), .Z(n2411) );
  IV U2528 ( .A(B[1686]), .Z(n2410) );
  IV U2529 ( .A(B[3855]), .Z(n241) );
  IV U2530 ( .A(B[1687]), .Z(n2409) );
  IV U2531 ( .A(B[1688]), .Z(n2408) );
  IV U2532 ( .A(B[1689]), .Z(n2407) );
  IV U2533 ( .A(B[1690]), .Z(n2406) );
  IV U2534 ( .A(B[1691]), .Z(n2405) );
  IV U2535 ( .A(B[1692]), .Z(n2404) );
  IV U2536 ( .A(B[1693]), .Z(n2403) );
  IV U2537 ( .A(B[1694]), .Z(n2402) );
  IV U2538 ( .A(B[1695]), .Z(n2401) );
  IV U2539 ( .A(B[1696]), .Z(n2400) );
  IV U2540 ( .A(B[3856]), .Z(n240) );
  IV U2541 ( .A(B[4072]), .Z(n24) );
  IV U2542 ( .A(B[1697]), .Z(n2399) );
  IV U2543 ( .A(B[1698]), .Z(n2398) );
  IV U2544 ( .A(B[1699]), .Z(n2397) );
  IV U2545 ( .A(B[1700]), .Z(n2396) );
  IV U2546 ( .A(B[1701]), .Z(n2395) );
  IV U2547 ( .A(B[1702]), .Z(n2394) );
  IV U2548 ( .A(B[1703]), .Z(n2393) );
  IV U2549 ( .A(B[1704]), .Z(n2392) );
  IV U2550 ( .A(B[1705]), .Z(n2391) );
  IV U2551 ( .A(B[1706]), .Z(n2390) );
  IV U2552 ( .A(B[3857]), .Z(n239) );
  IV U2553 ( .A(B[1707]), .Z(n2389) );
  IV U2554 ( .A(B[1708]), .Z(n2388) );
  IV U2555 ( .A(B[1709]), .Z(n2387) );
  IV U2556 ( .A(B[1710]), .Z(n2386) );
  IV U2557 ( .A(B[1711]), .Z(n2385) );
  IV U2558 ( .A(B[1712]), .Z(n2384) );
  IV U2559 ( .A(B[1713]), .Z(n2383) );
  IV U2560 ( .A(B[1714]), .Z(n2382) );
  IV U2561 ( .A(B[1715]), .Z(n2381) );
  IV U2562 ( .A(B[1716]), .Z(n2380) );
  IV U2563 ( .A(B[3858]), .Z(n238) );
  IV U2564 ( .A(B[1717]), .Z(n2379) );
  IV U2565 ( .A(B[1718]), .Z(n2378) );
  IV U2566 ( .A(B[1719]), .Z(n2377) );
  IV U2567 ( .A(B[1720]), .Z(n2376) );
  IV U2568 ( .A(B[1721]), .Z(n2375) );
  IV U2569 ( .A(B[1722]), .Z(n2374) );
  IV U2570 ( .A(B[1723]), .Z(n2373) );
  IV U2571 ( .A(B[1724]), .Z(n2372) );
  IV U2572 ( .A(B[1725]), .Z(n2371) );
  IV U2573 ( .A(B[1726]), .Z(n2370) );
  IV U2574 ( .A(B[3859]), .Z(n237) );
  IV U2575 ( .A(B[1727]), .Z(n2369) );
  IV U2576 ( .A(B[1728]), .Z(n2368) );
  IV U2577 ( .A(B[1729]), .Z(n2367) );
  IV U2578 ( .A(B[1730]), .Z(n2366) );
  IV U2579 ( .A(B[1731]), .Z(n2365) );
  IV U2580 ( .A(B[1732]), .Z(n2364) );
  IV U2581 ( .A(B[1733]), .Z(n2363) );
  IV U2582 ( .A(B[1734]), .Z(n2362) );
  IV U2583 ( .A(B[1735]), .Z(n2361) );
  IV U2584 ( .A(B[1736]), .Z(n2360) );
  IV U2585 ( .A(B[3860]), .Z(n236) );
  IV U2586 ( .A(B[1737]), .Z(n2359) );
  IV U2587 ( .A(B[1738]), .Z(n2358) );
  IV U2588 ( .A(B[1739]), .Z(n2357) );
  IV U2589 ( .A(B[1740]), .Z(n2356) );
  IV U2590 ( .A(B[1741]), .Z(n2355) );
  IV U2591 ( .A(B[1742]), .Z(n2354) );
  IV U2592 ( .A(B[1743]), .Z(n2353) );
  IV U2593 ( .A(B[1744]), .Z(n2352) );
  IV U2594 ( .A(B[1745]), .Z(n2351) );
  IV U2595 ( .A(B[1746]), .Z(n2350) );
  IV U2596 ( .A(B[3861]), .Z(n235) );
  IV U2597 ( .A(B[1747]), .Z(n2349) );
  IV U2598 ( .A(B[1748]), .Z(n2348) );
  IV U2599 ( .A(B[1749]), .Z(n2347) );
  IV U2600 ( .A(B[1750]), .Z(n2346) );
  IV U2601 ( .A(B[1751]), .Z(n2345) );
  IV U2602 ( .A(B[1752]), .Z(n2344) );
  IV U2603 ( .A(B[1753]), .Z(n2343) );
  IV U2604 ( .A(B[1754]), .Z(n2342) );
  IV U2605 ( .A(B[1755]), .Z(n2341) );
  IV U2606 ( .A(B[1756]), .Z(n2340) );
  IV U2607 ( .A(B[3862]), .Z(n234) );
  IV U2608 ( .A(B[1757]), .Z(n2339) );
  IV U2609 ( .A(B[1758]), .Z(n2338) );
  IV U2610 ( .A(B[1759]), .Z(n2337) );
  IV U2611 ( .A(B[1760]), .Z(n2336) );
  IV U2612 ( .A(B[1761]), .Z(n2335) );
  IV U2613 ( .A(B[1762]), .Z(n2334) );
  IV U2614 ( .A(B[1763]), .Z(n2333) );
  IV U2615 ( .A(B[1764]), .Z(n2332) );
  IV U2616 ( .A(B[1765]), .Z(n2331) );
  IV U2617 ( .A(B[1766]), .Z(n2330) );
  IV U2618 ( .A(B[3863]), .Z(n233) );
  IV U2619 ( .A(B[1767]), .Z(n2329) );
  IV U2620 ( .A(B[1768]), .Z(n2328) );
  IV U2621 ( .A(B[1769]), .Z(n2327) );
  IV U2622 ( .A(B[1770]), .Z(n2326) );
  IV U2623 ( .A(B[1771]), .Z(n2325) );
  IV U2624 ( .A(B[1772]), .Z(n2324) );
  IV U2625 ( .A(B[1773]), .Z(n2323) );
  IV U2626 ( .A(B[1774]), .Z(n2322) );
  IV U2627 ( .A(B[1775]), .Z(n2321) );
  IV U2628 ( .A(B[1776]), .Z(n2320) );
  IV U2629 ( .A(B[3864]), .Z(n232) );
  IV U2630 ( .A(B[1777]), .Z(n2319) );
  IV U2631 ( .A(B[1778]), .Z(n2318) );
  IV U2632 ( .A(B[1779]), .Z(n2317) );
  IV U2633 ( .A(B[1780]), .Z(n2316) );
  IV U2634 ( .A(B[1781]), .Z(n2315) );
  IV U2635 ( .A(B[1782]), .Z(n2314) );
  IV U2636 ( .A(B[1783]), .Z(n2313) );
  IV U2637 ( .A(B[1784]), .Z(n2312) );
  IV U2638 ( .A(B[1785]), .Z(n2311) );
  IV U2639 ( .A(B[1786]), .Z(n2310) );
  IV U2640 ( .A(B[3865]), .Z(n231) );
  IV U2641 ( .A(B[1787]), .Z(n2309) );
  IV U2642 ( .A(B[1788]), .Z(n2308) );
  IV U2643 ( .A(B[1789]), .Z(n2307) );
  IV U2644 ( .A(B[1790]), .Z(n2306) );
  IV U2645 ( .A(B[1791]), .Z(n2305) );
  IV U2646 ( .A(B[1792]), .Z(n2304) );
  IV U2647 ( .A(B[1793]), .Z(n2303) );
  IV U2648 ( .A(B[1794]), .Z(n2302) );
  IV U2649 ( .A(B[1795]), .Z(n2301) );
  IV U2650 ( .A(B[1796]), .Z(n2300) );
  IV U2651 ( .A(B[3866]), .Z(n230) );
  IV U2652 ( .A(B[4073]), .Z(n23) );
  IV U2653 ( .A(B[1797]), .Z(n2299) );
  IV U2654 ( .A(B[1798]), .Z(n2298) );
  IV U2655 ( .A(B[1799]), .Z(n2297) );
  IV U2656 ( .A(B[1800]), .Z(n2296) );
  IV U2657 ( .A(B[1801]), .Z(n2295) );
  IV U2658 ( .A(B[1802]), .Z(n2294) );
  IV U2659 ( .A(B[1803]), .Z(n2293) );
  IV U2660 ( .A(B[1804]), .Z(n2292) );
  IV U2661 ( .A(B[1805]), .Z(n2291) );
  IV U2662 ( .A(B[1806]), .Z(n2290) );
  IV U2663 ( .A(B[3867]), .Z(n229) );
  IV U2664 ( .A(B[1807]), .Z(n2289) );
  IV U2665 ( .A(B[1808]), .Z(n2288) );
  IV U2666 ( .A(B[1809]), .Z(n2287) );
  IV U2667 ( .A(B[1810]), .Z(n2286) );
  IV U2668 ( .A(B[1811]), .Z(n2285) );
  IV U2669 ( .A(B[1812]), .Z(n2284) );
  IV U2670 ( .A(B[1813]), .Z(n2283) );
  IV U2671 ( .A(B[1814]), .Z(n2282) );
  IV U2672 ( .A(B[1815]), .Z(n2281) );
  IV U2673 ( .A(B[1816]), .Z(n2280) );
  IV U2674 ( .A(B[3868]), .Z(n228) );
  IV U2675 ( .A(B[1817]), .Z(n2279) );
  IV U2676 ( .A(B[1818]), .Z(n2278) );
  IV U2677 ( .A(B[1819]), .Z(n2277) );
  IV U2678 ( .A(B[1820]), .Z(n2276) );
  IV U2679 ( .A(B[1821]), .Z(n2275) );
  IV U2680 ( .A(B[1822]), .Z(n2274) );
  IV U2681 ( .A(B[1823]), .Z(n2273) );
  IV U2682 ( .A(B[1824]), .Z(n2272) );
  IV U2683 ( .A(B[1825]), .Z(n2271) );
  IV U2684 ( .A(B[1826]), .Z(n2270) );
  IV U2685 ( .A(B[3869]), .Z(n227) );
  IV U2686 ( .A(B[1827]), .Z(n2269) );
  IV U2687 ( .A(B[1828]), .Z(n2268) );
  IV U2688 ( .A(B[1829]), .Z(n2267) );
  IV U2689 ( .A(B[1830]), .Z(n2266) );
  IV U2690 ( .A(B[1831]), .Z(n2265) );
  IV U2691 ( .A(B[1832]), .Z(n2264) );
  IV U2692 ( .A(B[1833]), .Z(n2263) );
  IV U2693 ( .A(B[1834]), .Z(n2262) );
  IV U2694 ( .A(B[1835]), .Z(n2261) );
  IV U2695 ( .A(B[1836]), .Z(n2260) );
  IV U2696 ( .A(B[3870]), .Z(n226) );
  IV U2697 ( .A(B[1837]), .Z(n2259) );
  IV U2698 ( .A(B[1838]), .Z(n2258) );
  IV U2699 ( .A(B[1839]), .Z(n2257) );
  IV U2700 ( .A(B[1840]), .Z(n2256) );
  IV U2701 ( .A(B[1841]), .Z(n2255) );
  IV U2702 ( .A(B[1842]), .Z(n2254) );
  IV U2703 ( .A(B[1843]), .Z(n2253) );
  IV U2704 ( .A(B[1844]), .Z(n2252) );
  IV U2705 ( .A(B[1845]), .Z(n2251) );
  IV U2706 ( .A(B[1846]), .Z(n2250) );
  IV U2707 ( .A(B[3871]), .Z(n225) );
  IV U2708 ( .A(B[1847]), .Z(n2249) );
  IV U2709 ( .A(B[1848]), .Z(n2248) );
  IV U2710 ( .A(B[1849]), .Z(n2247) );
  IV U2711 ( .A(B[1850]), .Z(n2246) );
  IV U2712 ( .A(B[1851]), .Z(n2245) );
  IV U2713 ( .A(B[1852]), .Z(n2244) );
  IV U2714 ( .A(B[1853]), .Z(n2243) );
  IV U2715 ( .A(B[1854]), .Z(n2242) );
  IV U2716 ( .A(B[1855]), .Z(n2241) );
  IV U2717 ( .A(B[1856]), .Z(n2240) );
  IV U2718 ( .A(B[3872]), .Z(n224) );
  IV U2719 ( .A(B[1857]), .Z(n2239) );
  IV U2720 ( .A(B[1858]), .Z(n2238) );
  IV U2721 ( .A(B[1859]), .Z(n2237) );
  IV U2722 ( .A(B[1860]), .Z(n2236) );
  IV U2723 ( .A(B[1861]), .Z(n2235) );
  IV U2724 ( .A(B[1862]), .Z(n2234) );
  IV U2725 ( .A(B[1863]), .Z(n2233) );
  IV U2726 ( .A(B[1864]), .Z(n2232) );
  IV U2727 ( .A(B[1865]), .Z(n2231) );
  IV U2728 ( .A(B[1866]), .Z(n2230) );
  IV U2729 ( .A(B[3873]), .Z(n223) );
  IV U2730 ( .A(B[1867]), .Z(n2229) );
  IV U2731 ( .A(B[1868]), .Z(n2228) );
  IV U2732 ( .A(B[1869]), .Z(n2227) );
  IV U2733 ( .A(B[1870]), .Z(n2226) );
  IV U2734 ( .A(B[1871]), .Z(n2225) );
  IV U2735 ( .A(B[1872]), .Z(n2224) );
  IV U2736 ( .A(B[1873]), .Z(n2223) );
  IV U2737 ( .A(B[1874]), .Z(n2222) );
  IV U2738 ( .A(B[1875]), .Z(n2221) );
  IV U2739 ( .A(B[1876]), .Z(n2220) );
  IV U2740 ( .A(B[3874]), .Z(n222) );
  IV U2741 ( .A(B[1877]), .Z(n2219) );
  IV U2742 ( .A(B[1878]), .Z(n2218) );
  IV U2743 ( .A(B[1879]), .Z(n2217) );
  IV U2744 ( .A(B[1880]), .Z(n2216) );
  IV U2745 ( .A(B[1881]), .Z(n2215) );
  IV U2746 ( .A(B[1882]), .Z(n2214) );
  IV U2747 ( .A(B[1883]), .Z(n2213) );
  IV U2748 ( .A(B[1884]), .Z(n2212) );
  IV U2749 ( .A(B[1885]), .Z(n2211) );
  IV U2750 ( .A(B[1886]), .Z(n2210) );
  IV U2751 ( .A(B[3875]), .Z(n221) );
  IV U2752 ( .A(B[1887]), .Z(n2209) );
  IV U2753 ( .A(B[1888]), .Z(n2208) );
  IV U2754 ( .A(B[1889]), .Z(n2207) );
  IV U2755 ( .A(B[1890]), .Z(n2206) );
  IV U2756 ( .A(B[1891]), .Z(n2205) );
  IV U2757 ( .A(B[1892]), .Z(n2204) );
  IV U2758 ( .A(B[1893]), .Z(n2203) );
  IV U2759 ( .A(B[1894]), .Z(n2202) );
  IV U2760 ( .A(B[1895]), .Z(n2201) );
  IV U2761 ( .A(B[1896]), .Z(n2200) );
  IV U2762 ( .A(B[3876]), .Z(n220) );
  IV U2763 ( .A(B[4074]), .Z(n22) );
  IV U2764 ( .A(B[1897]), .Z(n2199) );
  IV U2765 ( .A(B[1898]), .Z(n2198) );
  IV U2766 ( .A(B[1899]), .Z(n2197) );
  IV U2767 ( .A(B[1900]), .Z(n2196) );
  IV U2768 ( .A(B[1901]), .Z(n2195) );
  IV U2769 ( .A(B[1902]), .Z(n2194) );
  IV U2770 ( .A(B[1903]), .Z(n2193) );
  IV U2771 ( .A(B[1904]), .Z(n2192) );
  IV U2772 ( .A(B[1905]), .Z(n2191) );
  IV U2773 ( .A(B[1906]), .Z(n2190) );
  IV U2774 ( .A(B[3877]), .Z(n219) );
  IV U2775 ( .A(B[1907]), .Z(n2189) );
  IV U2776 ( .A(B[1908]), .Z(n2188) );
  IV U2777 ( .A(B[1909]), .Z(n2187) );
  IV U2778 ( .A(B[1910]), .Z(n2186) );
  IV U2779 ( .A(B[1911]), .Z(n2185) );
  IV U2780 ( .A(B[1912]), .Z(n2184) );
  IV U2781 ( .A(B[1913]), .Z(n2183) );
  IV U2782 ( .A(B[1914]), .Z(n2182) );
  IV U2783 ( .A(B[1915]), .Z(n2181) );
  IV U2784 ( .A(B[1916]), .Z(n2180) );
  IV U2785 ( .A(B[3878]), .Z(n218) );
  IV U2786 ( .A(B[1917]), .Z(n2179) );
  IV U2787 ( .A(B[1918]), .Z(n2178) );
  IV U2788 ( .A(B[1919]), .Z(n2177) );
  IV U2789 ( .A(B[1920]), .Z(n2176) );
  IV U2790 ( .A(B[1921]), .Z(n2175) );
  IV U2791 ( .A(B[1922]), .Z(n2174) );
  IV U2792 ( .A(B[1923]), .Z(n2173) );
  IV U2793 ( .A(B[1924]), .Z(n2172) );
  IV U2794 ( .A(B[1925]), .Z(n2171) );
  IV U2795 ( .A(B[1926]), .Z(n2170) );
  IV U2796 ( .A(B[3879]), .Z(n217) );
  IV U2797 ( .A(B[1927]), .Z(n2169) );
  IV U2798 ( .A(B[1928]), .Z(n2168) );
  IV U2799 ( .A(B[1929]), .Z(n2167) );
  IV U2800 ( .A(B[1930]), .Z(n2166) );
  IV U2801 ( .A(B[1931]), .Z(n2165) );
  IV U2802 ( .A(B[1932]), .Z(n2164) );
  IV U2803 ( .A(B[1933]), .Z(n2163) );
  IV U2804 ( .A(B[1934]), .Z(n2162) );
  IV U2805 ( .A(B[1935]), .Z(n2161) );
  IV U2806 ( .A(B[1936]), .Z(n2160) );
  IV U2807 ( .A(B[3880]), .Z(n216) );
  IV U2808 ( .A(B[1937]), .Z(n2159) );
  IV U2809 ( .A(B[1938]), .Z(n2158) );
  IV U2810 ( .A(B[1939]), .Z(n2157) );
  IV U2811 ( .A(B[1940]), .Z(n2156) );
  IV U2812 ( .A(B[1941]), .Z(n2155) );
  IV U2813 ( .A(B[1942]), .Z(n2154) );
  IV U2814 ( .A(B[1943]), .Z(n2153) );
  IV U2815 ( .A(B[1944]), .Z(n2152) );
  IV U2816 ( .A(B[1945]), .Z(n2151) );
  IV U2817 ( .A(B[1946]), .Z(n2150) );
  IV U2818 ( .A(B[3881]), .Z(n215) );
  IV U2819 ( .A(B[1947]), .Z(n2149) );
  IV U2820 ( .A(B[1948]), .Z(n2148) );
  IV U2821 ( .A(B[1949]), .Z(n2147) );
  IV U2822 ( .A(B[1950]), .Z(n2146) );
  IV U2823 ( .A(B[1951]), .Z(n2145) );
  IV U2824 ( .A(B[1952]), .Z(n2144) );
  IV U2825 ( .A(B[1953]), .Z(n2143) );
  IV U2826 ( .A(B[1954]), .Z(n2142) );
  IV U2827 ( .A(B[1955]), .Z(n2141) );
  IV U2828 ( .A(B[1956]), .Z(n2140) );
  IV U2829 ( .A(B[3882]), .Z(n214) );
  IV U2830 ( .A(B[1957]), .Z(n2139) );
  IV U2831 ( .A(B[1958]), .Z(n2138) );
  IV U2832 ( .A(B[1959]), .Z(n2137) );
  IV U2833 ( .A(B[1960]), .Z(n2136) );
  IV U2834 ( .A(B[1961]), .Z(n2135) );
  IV U2835 ( .A(B[1962]), .Z(n2134) );
  IV U2836 ( .A(B[1963]), .Z(n2133) );
  IV U2837 ( .A(B[1964]), .Z(n2132) );
  IV U2838 ( .A(B[1965]), .Z(n2131) );
  IV U2839 ( .A(B[1966]), .Z(n2130) );
  IV U2840 ( .A(B[3883]), .Z(n213) );
  IV U2841 ( .A(B[1967]), .Z(n2129) );
  IV U2842 ( .A(B[1968]), .Z(n2128) );
  IV U2843 ( .A(B[1969]), .Z(n2127) );
  IV U2844 ( .A(B[1970]), .Z(n2126) );
  IV U2845 ( .A(B[1971]), .Z(n2125) );
  IV U2846 ( .A(B[1972]), .Z(n2124) );
  IV U2847 ( .A(B[1973]), .Z(n2123) );
  IV U2848 ( .A(B[1974]), .Z(n2122) );
  IV U2849 ( .A(B[1975]), .Z(n2121) );
  IV U2850 ( .A(B[1976]), .Z(n2120) );
  IV U2851 ( .A(B[3884]), .Z(n212) );
  IV U2852 ( .A(B[1977]), .Z(n2119) );
  IV U2853 ( .A(B[1978]), .Z(n2118) );
  IV U2854 ( .A(B[1979]), .Z(n2117) );
  IV U2855 ( .A(B[1980]), .Z(n2116) );
  IV U2856 ( .A(B[1981]), .Z(n2115) );
  IV U2857 ( .A(B[1982]), .Z(n2114) );
  IV U2858 ( .A(B[1983]), .Z(n2113) );
  IV U2859 ( .A(B[1984]), .Z(n2112) );
  IV U2860 ( .A(B[1985]), .Z(n2111) );
  IV U2861 ( .A(B[1986]), .Z(n2110) );
  IV U2862 ( .A(B[3885]), .Z(n211) );
  IV U2863 ( .A(B[1987]), .Z(n2109) );
  IV U2864 ( .A(B[1988]), .Z(n2108) );
  IV U2865 ( .A(B[1989]), .Z(n2107) );
  IV U2866 ( .A(B[1990]), .Z(n2106) );
  IV U2867 ( .A(B[1991]), .Z(n2105) );
  IV U2868 ( .A(B[1992]), .Z(n2104) );
  IV U2869 ( .A(B[1993]), .Z(n2103) );
  IV U2870 ( .A(B[1994]), .Z(n2102) );
  IV U2871 ( .A(B[1995]), .Z(n2101) );
  IV U2872 ( .A(B[1996]), .Z(n2100) );
  IV U2873 ( .A(B[3886]), .Z(n210) );
  IV U2874 ( .A(B[4075]), .Z(n21) );
  IV U2875 ( .A(B[1997]), .Z(n2099) );
  IV U2876 ( .A(B[1998]), .Z(n2098) );
  IV U2877 ( .A(B[1999]), .Z(n2097) );
  IV U2878 ( .A(B[2000]), .Z(n2096) );
  IV U2879 ( .A(B[2001]), .Z(n2095) );
  IV U2880 ( .A(B[2002]), .Z(n2094) );
  IV U2881 ( .A(B[2003]), .Z(n2093) );
  IV U2882 ( .A(B[2004]), .Z(n2092) );
  IV U2883 ( .A(B[2005]), .Z(n2091) );
  IV U2884 ( .A(B[2006]), .Z(n2090) );
  IV U2885 ( .A(B[3887]), .Z(n209) );
  IV U2886 ( .A(B[2007]), .Z(n2089) );
  IV U2887 ( .A(B[2008]), .Z(n2088) );
  IV U2888 ( .A(B[2009]), .Z(n2087) );
  IV U2889 ( .A(B[2010]), .Z(n2086) );
  IV U2890 ( .A(B[2011]), .Z(n2085) );
  IV U2891 ( .A(B[2012]), .Z(n2084) );
  IV U2892 ( .A(B[2013]), .Z(n2083) );
  IV U2893 ( .A(B[2014]), .Z(n2082) );
  IV U2894 ( .A(B[2015]), .Z(n2081) );
  IV U2895 ( .A(B[2016]), .Z(n2080) );
  IV U2896 ( .A(B[3888]), .Z(n208) );
  IV U2897 ( .A(B[2017]), .Z(n2079) );
  IV U2898 ( .A(B[2018]), .Z(n2078) );
  IV U2899 ( .A(B[2019]), .Z(n2077) );
  IV U2900 ( .A(B[2020]), .Z(n2076) );
  IV U2901 ( .A(B[2021]), .Z(n2075) );
  IV U2902 ( .A(B[2022]), .Z(n2074) );
  IV U2903 ( .A(B[2023]), .Z(n2073) );
  IV U2904 ( .A(B[2024]), .Z(n2072) );
  IV U2905 ( .A(B[2025]), .Z(n2071) );
  IV U2906 ( .A(B[2026]), .Z(n2070) );
  IV U2907 ( .A(B[3889]), .Z(n207) );
  IV U2908 ( .A(B[2027]), .Z(n2069) );
  IV U2909 ( .A(B[2028]), .Z(n2068) );
  IV U2910 ( .A(B[2029]), .Z(n2067) );
  IV U2911 ( .A(B[2030]), .Z(n2066) );
  IV U2912 ( .A(B[2031]), .Z(n2065) );
  IV U2913 ( .A(B[2032]), .Z(n2064) );
  IV U2914 ( .A(B[2033]), .Z(n2063) );
  IV U2915 ( .A(B[2034]), .Z(n2062) );
  IV U2916 ( .A(B[2035]), .Z(n2061) );
  IV U2917 ( .A(B[2036]), .Z(n2060) );
  IV U2918 ( .A(B[3890]), .Z(n206) );
  IV U2919 ( .A(B[2037]), .Z(n2059) );
  IV U2920 ( .A(B[2038]), .Z(n2058) );
  IV U2921 ( .A(B[2039]), .Z(n2057) );
  IV U2922 ( .A(B[2040]), .Z(n2056) );
  IV U2923 ( .A(B[2041]), .Z(n2055) );
  IV U2924 ( .A(B[2042]), .Z(n2054) );
  IV U2925 ( .A(B[2043]), .Z(n2053) );
  IV U2926 ( .A(B[2044]), .Z(n2052) );
  IV U2927 ( .A(B[2045]), .Z(n2051) );
  IV U2928 ( .A(B[2046]), .Z(n2050) );
  IV U2929 ( .A(B[3891]), .Z(n205) );
  IV U2930 ( .A(B[2047]), .Z(n2049) );
  IV U2931 ( .A(B[2048]), .Z(n2048) );
  IV U2932 ( .A(B[2049]), .Z(n2047) );
  IV U2933 ( .A(B[2050]), .Z(n2046) );
  IV U2934 ( .A(B[2051]), .Z(n2045) );
  IV U2935 ( .A(B[2052]), .Z(n2044) );
  IV U2936 ( .A(B[2053]), .Z(n2043) );
  IV U2937 ( .A(B[2054]), .Z(n2042) );
  IV U2938 ( .A(B[2055]), .Z(n2041) );
  IV U2939 ( .A(B[2056]), .Z(n2040) );
  IV U2940 ( .A(B[3892]), .Z(n204) );
  IV U2941 ( .A(B[2057]), .Z(n2039) );
  IV U2942 ( .A(B[2058]), .Z(n2038) );
  IV U2943 ( .A(B[2059]), .Z(n2037) );
  IV U2944 ( .A(B[2060]), .Z(n2036) );
  IV U2945 ( .A(B[2061]), .Z(n2035) );
  IV U2946 ( .A(B[2062]), .Z(n2034) );
  IV U2947 ( .A(B[2063]), .Z(n2033) );
  IV U2948 ( .A(B[2064]), .Z(n2032) );
  IV U2949 ( .A(B[2065]), .Z(n2031) );
  IV U2950 ( .A(B[2066]), .Z(n2030) );
  IV U2951 ( .A(B[3893]), .Z(n203) );
  IV U2952 ( .A(B[2067]), .Z(n2029) );
  IV U2953 ( .A(B[2068]), .Z(n2028) );
  IV U2954 ( .A(B[2069]), .Z(n2027) );
  IV U2955 ( .A(B[2070]), .Z(n2026) );
  IV U2956 ( .A(B[2071]), .Z(n2025) );
  IV U2957 ( .A(B[2072]), .Z(n2024) );
  IV U2958 ( .A(B[2073]), .Z(n2023) );
  IV U2959 ( .A(B[2074]), .Z(n2022) );
  IV U2960 ( .A(B[2075]), .Z(n2021) );
  IV U2961 ( .A(B[2076]), .Z(n2020) );
  IV U2962 ( .A(B[3894]), .Z(n202) );
  IV U2963 ( .A(B[2077]), .Z(n2019) );
  IV U2964 ( .A(B[2078]), .Z(n2018) );
  IV U2965 ( .A(B[2079]), .Z(n2017) );
  IV U2966 ( .A(B[2080]), .Z(n2016) );
  IV U2967 ( .A(B[2081]), .Z(n2015) );
  IV U2968 ( .A(B[2082]), .Z(n2014) );
  IV U2969 ( .A(B[2083]), .Z(n2013) );
  IV U2970 ( .A(B[2084]), .Z(n2012) );
  IV U2971 ( .A(B[2085]), .Z(n2011) );
  IV U2972 ( .A(B[2086]), .Z(n2010) );
  IV U2973 ( .A(B[3895]), .Z(n201) );
  IV U2974 ( .A(B[2087]), .Z(n2009) );
  IV U2975 ( .A(B[2088]), .Z(n2008) );
  IV U2976 ( .A(B[2089]), .Z(n2007) );
  IV U2977 ( .A(B[2090]), .Z(n2006) );
  IV U2978 ( .A(B[2091]), .Z(n2005) );
  IV U2979 ( .A(B[2092]), .Z(n2004) );
  IV U2980 ( .A(B[2093]), .Z(n2003) );
  IV U2981 ( .A(B[2094]), .Z(n2002) );
  IV U2982 ( .A(B[2095]), .Z(n2001) );
  IV U2983 ( .A(B[2096]), .Z(n2000) );
  IV U2984 ( .A(B[3896]), .Z(n200) );
  IV U2985 ( .A(B[4076]), .Z(n20) );
  IV U2986 ( .A(B[4094]), .Z(n2) );
  IV U2987 ( .A(B[2097]), .Z(n1999) );
  IV U2988 ( .A(B[2098]), .Z(n1998) );
  IV U2989 ( .A(B[2099]), .Z(n1997) );
  IV U2990 ( .A(B[2100]), .Z(n1996) );
  IV U2991 ( .A(B[2101]), .Z(n1995) );
  IV U2992 ( .A(B[2102]), .Z(n1994) );
  IV U2993 ( .A(B[2103]), .Z(n1993) );
  IV U2994 ( .A(B[2104]), .Z(n1992) );
  IV U2995 ( .A(B[2105]), .Z(n1991) );
  IV U2996 ( .A(B[2106]), .Z(n1990) );
  IV U2997 ( .A(B[3897]), .Z(n199) );
  IV U2998 ( .A(B[2107]), .Z(n1989) );
  IV U2999 ( .A(B[2108]), .Z(n1988) );
  IV U3000 ( .A(B[2109]), .Z(n1987) );
  IV U3001 ( .A(B[2110]), .Z(n1986) );
  IV U3002 ( .A(B[2111]), .Z(n1985) );
  IV U3003 ( .A(B[2112]), .Z(n1984) );
  IV U3004 ( .A(B[2113]), .Z(n1983) );
  IV U3005 ( .A(B[2114]), .Z(n1982) );
  IV U3006 ( .A(B[2115]), .Z(n1981) );
  IV U3007 ( .A(B[2116]), .Z(n1980) );
  IV U3008 ( .A(B[3898]), .Z(n198) );
  IV U3009 ( .A(B[2117]), .Z(n1979) );
  IV U3010 ( .A(B[2118]), .Z(n1978) );
  IV U3011 ( .A(B[2119]), .Z(n1977) );
  IV U3012 ( .A(B[2120]), .Z(n1976) );
  IV U3013 ( .A(B[2121]), .Z(n1975) );
  IV U3014 ( .A(B[2122]), .Z(n1974) );
  IV U3015 ( .A(B[2123]), .Z(n1973) );
  IV U3016 ( .A(B[2124]), .Z(n1972) );
  IV U3017 ( .A(B[2125]), .Z(n1971) );
  IV U3018 ( .A(B[2126]), .Z(n1970) );
  IV U3019 ( .A(B[3899]), .Z(n197) );
  IV U3020 ( .A(B[2127]), .Z(n1969) );
  IV U3021 ( .A(B[2128]), .Z(n1968) );
  IV U3022 ( .A(B[2129]), .Z(n1967) );
  IV U3023 ( .A(B[2130]), .Z(n1966) );
  IV U3024 ( .A(B[2131]), .Z(n1965) );
  IV U3025 ( .A(B[2132]), .Z(n1964) );
  IV U3026 ( .A(B[2133]), .Z(n1963) );
  IV U3027 ( .A(B[2134]), .Z(n1962) );
  IV U3028 ( .A(B[2135]), .Z(n1961) );
  IV U3029 ( .A(B[2136]), .Z(n1960) );
  IV U3030 ( .A(B[3900]), .Z(n196) );
  IV U3031 ( .A(B[2137]), .Z(n1959) );
  IV U3032 ( .A(B[2138]), .Z(n1958) );
  IV U3033 ( .A(B[2139]), .Z(n1957) );
  IV U3034 ( .A(B[2140]), .Z(n1956) );
  IV U3035 ( .A(B[2141]), .Z(n1955) );
  IV U3036 ( .A(B[2142]), .Z(n1954) );
  IV U3037 ( .A(B[2143]), .Z(n1953) );
  IV U3038 ( .A(B[2144]), .Z(n1952) );
  IV U3039 ( .A(B[2145]), .Z(n1951) );
  IV U3040 ( .A(B[2146]), .Z(n1950) );
  IV U3041 ( .A(B[3901]), .Z(n195) );
  IV U3042 ( .A(B[2147]), .Z(n1949) );
  IV U3043 ( .A(B[2148]), .Z(n1948) );
  IV U3044 ( .A(B[2149]), .Z(n1947) );
  IV U3045 ( .A(B[2150]), .Z(n1946) );
  IV U3046 ( .A(B[2151]), .Z(n1945) );
  IV U3047 ( .A(B[2152]), .Z(n1944) );
  IV U3048 ( .A(B[2153]), .Z(n1943) );
  IV U3049 ( .A(B[2154]), .Z(n1942) );
  IV U3050 ( .A(B[2155]), .Z(n1941) );
  IV U3051 ( .A(B[2156]), .Z(n1940) );
  IV U3052 ( .A(B[3902]), .Z(n194) );
  IV U3053 ( .A(B[2157]), .Z(n1939) );
  IV U3054 ( .A(B[2158]), .Z(n1938) );
  IV U3055 ( .A(B[2159]), .Z(n1937) );
  IV U3056 ( .A(B[2160]), .Z(n1936) );
  IV U3057 ( .A(B[2161]), .Z(n1935) );
  IV U3058 ( .A(B[2162]), .Z(n1934) );
  IV U3059 ( .A(B[2163]), .Z(n1933) );
  IV U3060 ( .A(B[2164]), .Z(n1932) );
  IV U3061 ( .A(B[2165]), .Z(n1931) );
  IV U3062 ( .A(B[2166]), .Z(n1930) );
  IV U3063 ( .A(B[3903]), .Z(n193) );
  IV U3064 ( .A(B[2167]), .Z(n1929) );
  IV U3065 ( .A(B[2168]), .Z(n1928) );
  IV U3066 ( .A(B[2169]), .Z(n1927) );
  IV U3067 ( .A(B[2170]), .Z(n1926) );
  IV U3068 ( .A(B[2171]), .Z(n1925) );
  IV U3069 ( .A(B[2172]), .Z(n1924) );
  IV U3070 ( .A(B[2173]), .Z(n1923) );
  IV U3071 ( .A(B[2174]), .Z(n1922) );
  IV U3072 ( .A(B[2175]), .Z(n1921) );
  IV U3073 ( .A(B[2176]), .Z(n1920) );
  IV U3074 ( .A(B[3904]), .Z(n192) );
  IV U3075 ( .A(B[2177]), .Z(n1919) );
  IV U3076 ( .A(B[2178]), .Z(n1918) );
  IV U3077 ( .A(B[2179]), .Z(n1917) );
  IV U3078 ( .A(B[2180]), .Z(n1916) );
  IV U3079 ( .A(B[2181]), .Z(n1915) );
  IV U3080 ( .A(B[2182]), .Z(n1914) );
  IV U3081 ( .A(B[2183]), .Z(n1913) );
  IV U3082 ( .A(B[2184]), .Z(n1912) );
  IV U3083 ( .A(B[2185]), .Z(n1911) );
  IV U3084 ( .A(B[2186]), .Z(n1910) );
  IV U3085 ( .A(B[3905]), .Z(n191) );
  IV U3086 ( .A(B[2187]), .Z(n1909) );
  IV U3087 ( .A(B[2188]), .Z(n1908) );
  IV U3088 ( .A(B[2189]), .Z(n1907) );
  IV U3089 ( .A(B[2190]), .Z(n1906) );
  IV U3090 ( .A(B[2191]), .Z(n1905) );
  IV U3091 ( .A(B[2192]), .Z(n1904) );
  IV U3092 ( .A(B[2193]), .Z(n1903) );
  IV U3093 ( .A(B[2194]), .Z(n1902) );
  IV U3094 ( .A(B[2195]), .Z(n1901) );
  IV U3095 ( .A(B[2196]), .Z(n1900) );
  IV U3096 ( .A(B[3906]), .Z(n190) );
  IV U3097 ( .A(B[4077]), .Z(n19) );
  IV U3098 ( .A(B[2197]), .Z(n1899) );
  IV U3099 ( .A(B[2198]), .Z(n1898) );
  IV U3100 ( .A(B[2199]), .Z(n1897) );
  IV U3101 ( .A(B[2200]), .Z(n1896) );
  IV U3102 ( .A(B[2201]), .Z(n1895) );
  IV U3103 ( .A(B[2202]), .Z(n1894) );
  IV U3104 ( .A(B[2203]), .Z(n1893) );
  IV U3105 ( .A(B[2204]), .Z(n1892) );
  IV U3106 ( .A(B[2205]), .Z(n1891) );
  IV U3107 ( .A(B[2206]), .Z(n1890) );
  IV U3108 ( .A(B[3907]), .Z(n189) );
  IV U3109 ( .A(B[2207]), .Z(n1889) );
  IV U3110 ( .A(B[2208]), .Z(n1888) );
  IV U3111 ( .A(B[2209]), .Z(n1887) );
  IV U3112 ( .A(B[2210]), .Z(n1886) );
  IV U3113 ( .A(B[2211]), .Z(n1885) );
  IV U3114 ( .A(B[2212]), .Z(n1884) );
  IV U3115 ( .A(B[2213]), .Z(n1883) );
  IV U3116 ( .A(B[2214]), .Z(n1882) );
  IV U3117 ( .A(B[2215]), .Z(n1881) );
  IV U3118 ( .A(B[2216]), .Z(n1880) );
  IV U3119 ( .A(B[3908]), .Z(n188) );
  IV U3120 ( .A(B[2217]), .Z(n1879) );
  IV U3121 ( .A(B[2218]), .Z(n1878) );
  IV U3122 ( .A(B[2219]), .Z(n1877) );
  IV U3123 ( .A(B[2220]), .Z(n1876) );
  IV U3124 ( .A(B[2221]), .Z(n1875) );
  IV U3125 ( .A(B[2222]), .Z(n1874) );
  IV U3126 ( .A(B[2223]), .Z(n1873) );
  IV U3127 ( .A(B[2224]), .Z(n1872) );
  IV U3128 ( .A(B[2225]), .Z(n1871) );
  IV U3129 ( .A(B[2226]), .Z(n1870) );
  IV U3130 ( .A(B[3909]), .Z(n187) );
  IV U3131 ( .A(B[2227]), .Z(n1869) );
  IV U3132 ( .A(B[2228]), .Z(n1868) );
  IV U3133 ( .A(B[2229]), .Z(n1867) );
  IV U3134 ( .A(B[2230]), .Z(n1866) );
  IV U3135 ( .A(B[2231]), .Z(n1865) );
  IV U3136 ( .A(B[2232]), .Z(n1864) );
  IV U3137 ( .A(B[2233]), .Z(n1863) );
  IV U3138 ( .A(B[2234]), .Z(n1862) );
  IV U3139 ( .A(B[2235]), .Z(n1861) );
  IV U3140 ( .A(B[2236]), .Z(n1860) );
  IV U3141 ( .A(B[3910]), .Z(n186) );
  IV U3142 ( .A(B[2237]), .Z(n1859) );
  IV U3143 ( .A(B[2238]), .Z(n1858) );
  IV U3144 ( .A(B[2239]), .Z(n1857) );
  IV U3145 ( .A(B[2240]), .Z(n1856) );
  IV U3146 ( .A(B[2241]), .Z(n1855) );
  IV U3147 ( .A(B[2242]), .Z(n1854) );
  IV U3148 ( .A(B[2243]), .Z(n1853) );
  IV U3149 ( .A(B[2244]), .Z(n1852) );
  IV U3150 ( .A(B[2245]), .Z(n1851) );
  IV U3151 ( .A(B[2246]), .Z(n1850) );
  IV U3152 ( .A(B[3911]), .Z(n185) );
  IV U3153 ( .A(B[2247]), .Z(n1849) );
  IV U3154 ( .A(B[2248]), .Z(n1848) );
  IV U3155 ( .A(B[2249]), .Z(n1847) );
  IV U3156 ( .A(B[2250]), .Z(n1846) );
  IV U3157 ( .A(B[2251]), .Z(n1845) );
  IV U3158 ( .A(B[2252]), .Z(n1844) );
  IV U3159 ( .A(B[2253]), .Z(n1843) );
  IV U3160 ( .A(B[2254]), .Z(n1842) );
  IV U3161 ( .A(B[2255]), .Z(n1841) );
  IV U3162 ( .A(B[2256]), .Z(n1840) );
  IV U3163 ( .A(B[3912]), .Z(n184) );
  IV U3164 ( .A(B[2257]), .Z(n1839) );
  IV U3165 ( .A(B[2258]), .Z(n1838) );
  IV U3166 ( .A(B[2259]), .Z(n1837) );
  IV U3167 ( .A(B[2260]), .Z(n1836) );
  IV U3168 ( .A(B[2261]), .Z(n1835) );
  IV U3169 ( .A(B[2262]), .Z(n1834) );
  IV U3170 ( .A(B[2263]), .Z(n1833) );
  IV U3171 ( .A(B[2264]), .Z(n1832) );
  IV U3172 ( .A(B[2265]), .Z(n1831) );
  IV U3173 ( .A(B[2266]), .Z(n1830) );
  IV U3174 ( .A(B[3913]), .Z(n183) );
  IV U3175 ( .A(B[2267]), .Z(n1829) );
  IV U3176 ( .A(B[2268]), .Z(n1828) );
  IV U3177 ( .A(B[2269]), .Z(n1827) );
  IV U3178 ( .A(B[2270]), .Z(n1826) );
  IV U3179 ( .A(B[2271]), .Z(n1825) );
  IV U3180 ( .A(B[2272]), .Z(n1824) );
  IV U3181 ( .A(B[2273]), .Z(n1823) );
  IV U3182 ( .A(B[2274]), .Z(n1822) );
  IV U3183 ( .A(B[2275]), .Z(n1821) );
  IV U3184 ( .A(B[2276]), .Z(n1820) );
  IV U3185 ( .A(B[3914]), .Z(n182) );
  IV U3186 ( .A(B[2277]), .Z(n1819) );
  IV U3187 ( .A(B[2278]), .Z(n1818) );
  IV U3188 ( .A(B[2279]), .Z(n1817) );
  IV U3189 ( .A(B[2280]), .Z(n1816) );
  IV U3190 ( .A(B[2281]), .Z(n1815) );
  IV U3191 ( .A(B[2282]), .Z(n1814) );
  IV U3192 ( .A(B[2283]), .Z(n1813) );
  IV U3193 ( .A(B[2284]), .Z(n1812) );
  IV U3194 ( .A(B[2285]), .Z(n1811) );
  IV U3195 ( .A(B[2286]), .Z(n1810) );
  IV U3196 ( .A(B[3915]), .Z(n181) );
  IV U3197 ( .A(B[2287]), .Z(n1809) );
  IV U3198 ( .A(B[2288]), .Z(n1808) );
  IV U3199 ( .A(B[2289]), .Z(n1807) );
  IV U3200 ( .A(B[2290]), .Z(n1806) );
  IV U3201 ( .A(B[2291]), .Z(n1805) );
  IV U3202 ( .A(B[2292]), .Z(n1804) );
  IV U3203 ( .A(B[2293]), .Z(n1803) );
  IV U3204 ( .A(B[2294]), .Z(n1802) );
  IV U3205 ( .A(B[2295]), .Z(n1801) );
  IV U3206 ( .A(B[2296]), .Z(n1800) );
  IV U3207 ( .A(B[3916]), .Z(n180) );
  IV U3208 ( .A(B[4078]), .Z(n18) );
  IV U3209 ( .A(B[2297]), .Z(n1799) );
  IV U3210 ( .A(B[2298]), .Z(n1798) );
  IV U3211 ( .A(B[2299]), .Z(n1797) );
  IV U3212 ( .A(B[2300]), .Z(n1796) );
  IV U3213 ( .A(B[2301]), .Z(n1795) );
  IV U3214 ( .A(B[2302]), .Z(n1794) );
  IV U3215 ( .A(B[2303]), .Z(n1793) );
  IV U3216 ( .A(B[2304]), .Z(n1792) );
  IV U3217 ( .A(B[2305]), .Z(n1791) );
  IV U3218 ( .A(B[2306]), .Z(n1790) );
  IV U3219 ( .A(B[3917]), .Z(n179) );
  IV U3220 ( .A(B[2307]), .Z(n1789) );
  IV U3221 ( .A(B[2308]), .Z(n1788) );
  IV U3222 ( .A(B[2309]), .Z(n1787) );
  IV U3223 ( .A(B[2310]), .Z(n1786) );
  IV U3224 ( .A(B[2311]), .Z(n1785) );
  IV U3225 ( .A(B[2312]), .Z(n1784) );
  IV U3226 ( .A(B[2313]), .Z(n1783) );
  IV U3227 ( .A(B[2314]), .Z(n1782) );
  IV U3228 ( .A(B[2315]), .Z(n1781) );
  IV U3229 ( .A(B[2316]), .Z(n1780) );
  IV U3230 ( .A(B[3918]), .Z(n178) );
  IV U3231 ( .A(B[2317]), .Z(n1779) );
  IV U3232 ( .A(B[2318]), .Z(n1778) );
  IV U3233 ( .A(B[2319]), .Z(n1777) );
  IV U3234 ( .A(B[2320]), .Z(n1776) );
  IV U3235 ( .A(B[2321]), .Z(n1775) );
  IV U3236 ( .A(B[2322]), .Z(n1774) );
  IV U3237 ( .A(B[2323]), .Z(n1773) );
  IV U3238 ( .A(B[2324]), .Z(n1772) );
  IV U3239 ( .A(B[2325]), .Z(n1771) );
  IV U3240 ( .A(B[2326]), .Z(n1770) );
  IV U3241 ( .A(B[3919]), .Z(n177) );
  IV U3242 ( .A(B[2327]), .Z(n1769) );
  IV U3243 ( .A(B[2328]), .Z(n1768) );
  IV U3244 ( .A(B[2329]), .Z(n1767) );
  IV U3245 ( .A(B[2330]), .Z(n1766) );
  IV U3246 ( .A(B[2331]), .Z(n1765) );
  IV U3247 ( .A(B[2332]), .Z(n1764) );
  IV U3248 ( .A(B[2333]), .Z(n1763) );
  IV U3249 ( .A(B[2334]), .Z(n1762) );
  IV U3250 ( .A(B[2335]), .Z(n1761) );
  IV U3251 ( .A(B[2336]), .Z(n1760) );
  IV U3252 ( .A(B[3920]), .Z(n176) );
  IV U3253 ( .A(B[2337]), .Z(n1759) );
  IV U3254 ( .A(B[2338]), .Z(n1758) );
  IV U3255 ( .A(B[2339]), .Z(n1757) );
  IV U3256 ( .A(B[2340]), .Z(n1756) );
  IV U3257 ( .A(B[2341]), .Z(n1755) );
  IV U3258 ( .A(B[2342]), .Z(n1754) );
  IV U3259 ( .A(B[2343]), .Z(n1753) );
  IV U3260 ( .A(B[2344]), .Z(n1752) );
  IV U3261 ( .A(B[2345]), .Z(n1751) );
  IV U3262 ( .A(B[2346]), .Z(n1750) );
  IV U3263 ( .A(B[3921]), .Z(n175) );
  IV U3264 ( .A(B[2347]), .Z(n1749) );
  IV U3265 ( .A(B[2348]), .Z(n1748) );
  IV U3266 ( .A(B[2349]), .Z(n1747) );
  IV U3267 ( .A(B[2350]), .Z(n1746) );
  IV U3268 ( .A(B[2351]), .Z(n1745) );
  IV U3269 ( .A(B[2352]), .Z(n1744) );
  IV U3270 ( .A(B[2353]), .Z(n1743) );
  IV U3271 ( .A(B[2354]), .Z(n1742) );
  IV U3272 ( .A(B[2355]), .Z(n1741) );
  IV U3273 ( .A(B[2356]), .Z(n1740) );
  IV U3274 ( .A(B[3922]), .Z(n174) );
  IV U3275 ( .A(B[2357]), .Z(n1739) );
  IV U3276 ( .A(B[2358]), .Z(n1738) );
  IV U3277 ( .A(B[2359]), .Z(n1737) );
  IV U3278 ( .A(B[2360]), .Z(n1736) );
  IV U3279 ( .A(B[2361]), .Z(n1735) );
  IV U3280 ( .A(B[2362]), .Z(n1734) );
  IV U3281 ( .A(B[2363]), .Z(n1733) );
  IV U3282 ( .A(B[2364]), .Z(n1732) );
  IV U3283 ( .A(B[2365]), .Z(n1731) );
  IV U3284 ( .A(B[2366]), .Z(n1730) );
  IV U3285 ( .A(B[3923]), .Z(n173) );
  IV U3286 ( .A(B[2367]), .Z(n1729) );
  IV U3287 ( .A(B[2368]), .Z(n1728) );
  IV U3288 ( .A(B[2369]), .Z(n1727) );
  IV U3289 ( .A(B[2370]), .Z(n1726) );
  IV U3290 ( .A(B[2371]), .Z(n1725) );
  IV U3291 ( .A(B[2372]), .Z(n1724) );
  IV U3292 ( .A(B[2373]), .Z(n1723) );
  IV U3293 ( .A(B[2374]), .Z(n1722) );
  IV U3294 ( .A(B[2375]), .Z(n1721) );
  IV U3295 ( .A(B[2376]), .Z(n1720) );
  IV U3296 ( .A(B[3924]), .Z(n172) );
  IV U3297 ( .A(B[2377]), .Z(n1719) );
  IV U3298 ( .A(B[2378]), .Z(n1718) );
  IV U3299 ( .A(B[2379]), .Z(n1717) );
  IV U3300 ( .A(B[2380]), .Z(n1716) );
  IV U3301 ( .A(B[2381]), .Z(n1715) );
  IV U3302 ( .A(B[2382]), .Z(n1714) );
  IV U3303 ( .A(B[2383]), .Z(n1713) );
  IV U3304 ( .A(B[2384]), .Z(n1712) );
  IV U3305 ( .A(B[2385]), .Z(n1711) );
  IV U3306 ( .A(B[2386]), .Z(n1710) );
  IV U3307 ( .A(B[3925]), .Z(n171) );
  IV U3308 ( .A(B[2387]), .Z(n1709) );
  IV U3309 ( .A(B[2388]), .Z(n1708) );
  IV U3310 ( .A(B[2389]), .Z(n1707) );
  IV U3311 ( .A(B[2390]), .Z(n1706) );
  IV U3312 ( .A(B[2391]), .Z(n1705) );
  IV U3313 ( .A(B[2392]), .Z(n1704) );
  IV U3314 ( .A(B[2393]), .Z(n1703) );
  IV U3315 ( .A(B[2394]), .Z(n1702) );
  IV U3316 ( .A(B[2395]), .Z(n1701) );
  IV U3317 ( .A(B[2396]), .Z(n1700) );
  IV U3318 ( .A(B[3926]), .Z(n170) );
  IV U3319 ( .A(B[4079]), .Z(n17) );
  IV U3320 ( .A(B[2397]), .Z(n1699) );
  IV U3321 ( .A(B[2398]), .Z(n1698) );
  IV U3322 ( .A(B[2399]), .Z(n1697) );
  IV U3323 ( .A(B[2400]), .Z(n1696) );
  IV U3324 ( .A(B[2401]), .Z(n1695) );
  IV U3325 ( .A(B[2402]), .Z(n1694) );
  IV U3326 ( .A(B[2403]), .Z(n1693) );
  IV U3327 ( .A(B[2404]), .Z(n1692) );
  IV U3328 ( .A(B[2405]), .Z(n1691) );
  IV U3329 ( .A(B[2406]), .Z(n1690) );
  IV U3330 ( .A(B[3927]), .Z(n169) );
  IV U3331 ( .A(B[2407]), .Z(n1689) );
  IV U3332 ( .A(B[2408]), .Z(n1688) );
  IV U3333 ( .A(B[2409]), .Z(n1687) );
  IV U3334 ( .A(B[2410]), .Z(n1686) );
  IV U3335 ( .A(B[2411]), .Z(n1685) );
  IV U3336 ( .A(B[2412]), .Z(n1684) );
  IV U3337 ( .A(B[2413]), .Z(n1683) );
  IV U3338 ( .A(B[2414]), .Z(n1682) );
  IV U3339 ( .A(B[2415]), .Z(n1681) );
  IV U3340 ( .A(B[2416]), .Z(n1680) );
  IV U3341 ( .A(B[3928]), .Z(n168) );
  IV U3342 ( .A(B[2417]), .Z(n1679) );
  IV U3343 ( .A(B[2418]), .Z(n1678) );
  IV U3344 ( .A(B[2419]), .Z(n1677) );
  IV U3345 ( .A(B[2420]), .Z(n1676) );
  IV U3346 ( .A(B[2421]), .Z(n1675) );
  IV U3347 ( .A(B[2422]), .Z(n1674) );
  IV U3348 ( .A(B[2423]), .Z(n1673) );
  IV U3349 ( .A(B[2424]), .Z(n1672) );
  IV U3350 ( .A(B[2425]), .Z(n1671) );
  IV U3351 ( .A(B[2426]), .Z(n1670) );
  IV U3352 ( .A(B[3929]), .Z(n167) );
  IV U3353 ( .A(B[2427]), .Z(n1669) );
  IV U3354 ( .A(B[2428]), .Z(n1668) );
  IV U3355 ( .A(B[2429]), .Z(n1667) );
  IV U3356 ( .A(B[2430]), .Z(n1666) );
  IV U3357 ( .A(B[2431]), .Z(n1665) );
  IV U3358 ( .A(B[2432]), .Z(n1664) );
  IV U3359 ( .A(B[2433]), .Z(n1663) );
  IV U3360 ( .A(B[2434]), .Z(n1662) );
  IV U3361 ( .A(B[2435]), .Z(n1661) );
  IV U3362 ( .A(B[2436]), .Z(n1660) );
  IV U3363 ( .A(B[3930]), .Z(n166) );
  IV U3364 ( .A(B[2437]), .Z(n1659) );
  IV U3365 ( .A(B[2438]), .Z(n1658) );
  IV U3366 ( .A(B[2439]), .Z(n1657) );
  IV U3367 ( .A(B[2440]), .Z(n1656) );
  IV U3368 ( .A(B[2441]), .Z(n1655) );
  IV U3369 ( .A(B[2442]), .Z(n1654) );
  IV U3370 ( .A(B[2443]), .Z(n1653) );
  IV U3371 ( .A(B[2444]), .Z(n1652) );
  IV U3372 ( .A(B[2445]), .Z(n1651) );
  IV U3373 ( .A(B[2446]), .Z(n1650) );
  IV U3374 ( .A(B[3931]), .Z(n165) );
  IV U3375 ( .A(B[2447]), .Z(n1649) );
  IV U3376 ( .A(B[2448]), .Z(n1648) );
  IV U3377 ( .A(B[2449]), .Z(n1647) );
  IV U3378 ( .A(B[2450]), .Z(n1646) );
  IV U3379 ( .A(B[2451]), .Z(n1645) );
  IV U3380 ( .A(B[2452]), .Z(n1644) );
  IV U3381 ( .A(B[2453]), .Z(n1643) );
  IV U3382 ( .A(B[2454]), .Z(n1642) );
  IV U3383 ( .A(B[2455]), .Z(n1641) );
  IV U3384 ( .A(B[2456]), .Z(n1640) );
  IV U3385 ( .A(B[3932]), .Z(n164) );
  IV U3386 ( .A(B[2457]), .Z(n1639) );
  IV U3387 ( .A(B[2458]), .Z(n1638) );
  IV U3388 ( .A(B[2459]), .Z(n1637) );
  IV U3389 ( .A(B[2460]), .Z(n1636) );
  IV U3390 ( .A(B[2461]), .Z(n1635) );
  IV U3391 ( .A(B[2462]), .Z(n1634) );
  IV U3392 ( .A(B[2463]), .Z(n1633) );
  IV U3393 ( .A(B[2464]), .Z(n1632) );
  IV U3394 ( .A(B[2465]), .Z(n1631) );
  IV U3395 ( .A(B[2466]), .Z(n1630) );
  IV U3396 ( .A(B[3933]), .Z(n163) );
  IV U3397 ( .A(B[2467]), .Z(n1629) );
  IV U3398 ( .A(B[2468]), .Z(n1628) );
  IV U3399 ( .A(B[2469]), .Z(n1627) );
  IV U3400 ( .A(B[2470]), .Z(n1626) );
  IV U3401 ( .A(B[2471]), .Z(n1625) );
  IV U3402 ( .A(B[2472]), .Z(n1624) );
  IV U3403 ( .A(B[2473]), .Z(n1623) );
  IV U3404 ( .A(B[2474]), .Z(n1622) );
  IV U3405 ( .A(B[2475]), .Z(n1621) );
  IV U3406 ( .A(B[2476]), .Z(n1620) );
  IV U3407 ( .A(B[3934]), .Z(n162) );
  IV U3408 ( .A(B[2477]), .Z(n1619) );
  IV U3409 ( .A(B[2478]), .Z(n1618) );
  IV U3410 ( .A(B[2479]), .Z(n1617) );
  IV U3411 ( .A(B[2480]), .Z(n1616) );
  IV U3412 ( .A(B[2481]), .Z(n1615) );
  IV U3413 ( .A(B[2482]), .Z(n1614) );
  IV U3414 ( .A(B[2483]), .Z(n1613) );
  IV U3415 ( .A(B[2484]), .Z(n1612) );
  IV U3416 ( .A(B[2485]), .Z(n1611) );
  IV U3417 ( .A(B[2486]), .Z(n1610) );
  IV U3418 ( .A(B[3935]), .Z(n161) );
  IV U3419 ( .A(B[2487]), .Z(n1609) );
  IV U3420 ( .A(B[2488]), .Z(n1608) );
  IV U3421 ( .A(B[2489]), .Z(n1607) );
  IV U3422 ( .A(B[2490]), .Z(n1606) );
  IV U3423 ( .A(B[2491]), .Z(n1605) );
  IV U3424 ( .A(B[2492]), .Z(n1604) );
  IV U3425 ( .A(B[2493]), .Z(n1603) );
  IV U3426 ( .A(B[2494]), .Z(n1602) );
  IV U3427 ( .A(B[2495]), .Z(n1601) );
  IV U3428 ( .A(B[2496]), .Z(n1600) );
  IV U3429 ( .A(B[3936]), .Z(n160) );
  IV U3430 ( .A(B[4080]), .Z(n16) );
  IV U3431 ( .A(B[2497]), .Z(n1599) );
  IV U3432 ( .A(B[2498]), .Z(n1598) );
  IV U3433 ( .A(B[2499]), .Z(n1597) );
  IV U3434 ( .A(B[2500]), .Z(n1596) );
  IV U3435 ( .A(B[2501]), .Z(n1595) );
  IV U3436 ( .A(B[2502]), .Z(n1594) );
  IV U3437 ( .A(B[2503]), .Z(n1593) );
  IV U3438 ( .A(B[2504]), .Z(n1592) );
  IV U3439 ( .A(B[2505]), .Z(n1591) );
  IV U3440 ( .A(B[2506]), .Z(n1590) );
  IV U3441 ( .A(B[3937]), .Z(n159) );
  IV U3442 ( .A(B[2507]), .Z(n1589) );
  IV U3443 ( .A(B[2508]), .Z(n1588) );
  IV U3444 ( .A(B[2509]), .Z(n1587) );
  IV U3445 ( .A(B[2510]), .Z(n1586) );
  IV U3446 ( .A(B[2511]), .Z(n1585) );
  IV U3447 ( .A(B[2512]), .Z(n1584) );
  IV U3448 ( .A(B[2513]), .Z(n1583) );
  IV U3449 ( .A(B[2514]), .Z(n1582) );
  IV U3450 ( .A(B[2515]), .Z(n1581) );
  IV U3451 ( .A(B[2516]), .Z(n1580) );
  IV U3452 ( .A(B[3938]), .Z(n158) );
  IV U3453 ( .A(B[2517]), .Z(n1579) );
  IV U3454 ( .A(B[2518]), .Z(n1578) );
  IV U3455 ( .A(B[2519]), .Z(n1577) );
  IV U3456 ( .A(B[2520]), .Z(n1576) );
  IV U3457 ( .A(B[2521]), .Z(n1575) );
  IV U3458 ( .A(B[2522]), .Z(n1574) );
  IV U3459 ( .A(B[2523]), .Z(n1573) );
  IV U3460 ( .A(B[2524]), .Z(n1572) );
  IV U3461 ( .A(B[2525]), .Z(n1571) );
  IV U3462 ( .A(B[2526]), .Z(n1570) );
  IV U3463 ( .A(B[3939]), .Z(n157) );
  IV U3464 ( .A(B[2527]), .Z(n1569) );
  IV U3465 ( .A(B[2528]), .Z(n1568) );
  IV U3466 ( .A(B[2529]), .Z(n1567) );
  IV U3467 ( .A(B[2530]), .Z(n1566) );
  IV U3468 ( .A(B[2531]), .Z(n1565) );
  IV U3469 ( .A(B[2532]), .Z(n1564) );
  IV U3470 ( .A(B[2533]), .Z(n1563) );
  IV U3471 ( .A(B[2534]), .Z(n1562) );
  IV U3472 ( .A(B[2535]), .Z(n1561) );
  IV U3473 ( .A(B[2536]), .Z(n1560) );
  IV U3474 ( .A(B[3940]), .Z(n156) );
  IV U3475 ( .A(B[2537]), .Z(n1559) );
  IV U3476 ( .A(B[2538]), .Z(n1558) );
  IV U3477 ( .A(B[2539]), .Z(n1557) );
  IV U3478 ( .A(B[2540]), .Z(n1556) );
  IV U3479 ( .A(B[2541]), .Z(n1555) );
  IV U3480 ( .A(B[2542]), .Z(n1554) );
  IV U3481 ( .A(B[2543]), .Z(n1553) );
  IV U3482 ( .A(B[2544]), .Z(n1552) );
  IV U3483 ( .A(B[2545]), .Z(n1551) );
  IV U3484 ( .A(B[2546]), .Z(n1550) );
  IV U3485 ( .A(B[3941]), .Z(n155) );
  IV U3486 ( .A(B[2547]), .Z(n1549) );
  IV U3487 ( .A(B[2548]), .Z(n1548) );
  IV U3488 ( .A(B[2549]), .Z(n1547) );
  IV U3489 ( .A(B[2550]), .Z(n1546) );
  IV U3490 ( .A(B[2551]), .Z(n1545) );
  IV U3491 ( .A(B[2552]), .Z(n1544) );
  IV U3492 ( .A(B[2553]), .Z(n1543) );
  IV U3493 ( .A(B[2554]), .Z(n1542) );
  IV U3494 ( .A(B[2555]), .Z(n1541) );
  IV U3495 ( .A(B[2556]), .Z(n1540) );
  IV U3496 ( .A(B[3942]), .Z(n154) );
  IV U3497 ( .A(B[2557]), .Z(n1539) );
  IV U3498 ( .A(B[2558]), .Z(n1538) );
  IV U3499 ( .A(B[2559]), .Z(n1537) );
  IV U3500 ( .A(B[2560]), .Z(n1536) );
  IV U3501 ( .A(B[2561]), .Z(n1535) );
  IV U3502 ( .A(B[2562]), .Z(n1534) );
  IV U3503 ( .A(B[2563]), .Z(n1533) );
  IV U3504 ( .A(B[2564]), .Z(n1532) );
  IV U3505 ( .A(B[2565]), .Z(n1531) );
  IV U3506 ( .A(B[2566]), .Z(n1530) );
  IV U3507 ( .A(B[3943]), .Z(n153) );
  IV U3508 ( .A(B[2567]), .Z(n1529) );
  IV U3509 ( .A(B[2568]), .Z(n1528) );
  IV U3510 ( .A(B[2569]), .Z(n1527) );
  IV U3511 ( .A(B[2570]), .Z(n1526) );
  IV U3512 ( .A(B[2571]), .Z(n1525) );
  IV U3513 ( .A(B[2572]), .Z(n1524) );
  IV U3514 ( .A(B[2573]), .Z(n1523) );
  IV U3515 ( .A(B[2574]), .Z(n1522) );
  IV U3516 ( .A(B[2575]), .Z(n1521) );
  IV U3517 ( .A(B[2576]), .Z(n1520) );
  IV U3518 ( .A(B[3944]), .Z(n152) );
  IV U3519 ( .A(B[2577]), .Z(n1519) );
  IV U3520 ( .A(B[2578]), .Z(n1518) );
  IV U3521 ( .A(B[2579]), .Z(n1517) );
  IV U3522 ( .A(B[2580]), .Z(n1516) );
  IV U3523 ( .A(B[2581]), .Z(n1515) );
  IV U3524 ( .A(B[2582]), .Z(n1514) );
  IV U3525 ( .A(B[2583]), .Z(n1513) );
  IV U3526 ( .A(B[2584]), .Z(n1512) );
  IV U3527 ( .A(B[2585]), .Z(n1511) );
  IV U3528 ( .A(B[2586]), .Z(n1510) );
  IV U3529 ( .A(B[3945]), .Z(n151) );
  IV U3530 ( .A(B[2587]), .Z(n1509) );
  IV U3531 ( .A(B[2588]), .Z(n1508) );
  IV U3532 ( .A(B[2589]), .Z(n1507) );
  IV U3533 ( .A(B[2590]), .Z(n1506) );
  IV U3534 ( .A(B[2591]), .Z(n1505) );
  IV U3535 ( .A(B[2592]), .Z(n1504) );
  IV U3536 ( .A(B[2593]), .Z(n1503) );
  IV U3537 ( .A(B[2594]), .Z(n1502) );
  IV U3538 ( .A(B[2595]), .Z(n1501) );
  IV U3539 ( .A(B[2596]), .Z(n1500) );
  IV U3540 ( .A(B[3946]), .Z(n150) );
  IV U3541 ( .A(B[4081]), .Z(n15) );
  IV U3542 ( .A(B[2597]), .Z(n1499) );
  IV U3543 ( .A(B[2598]), .Z(n1498) );
  IV U3544 ( .A(B[2599]), .Z(n1497) );
  IV U3545 ( .A(B[2600]), .Z(n1496) );
  IV U3546 ( .A(B[2601]), .Z(n1495) );
  IV U3547 ( .A(B[2602]), .Z(n1494) );
  IV U3548 ( .A(B[2603]), .Z(n1493) );
  IV U3549 ( .A(B[2604]), .Z(n1492) );
  IV U3550 ( .A(B[2605]), .Z(n1491) );
  IV U3551 ( .A(B[2606]), .Z(n1490) );
  IV U3552 ( .A(B[3947]), .Z(n149) );
  IV U3553 ( .A(B[2607]), .Z(n1489) );
  IV U3554 ( .A(B[2608]), .Z(n1488) );
  IV U3555 ( .A(B[2609]), .Z(n1487) );
  IV U3556 ( .A(B[2610]), .Z(n1486) );
  IV U3557 ( .A(B[2611]), .Z(n1485) );
  IV U3558 ( .A(B[2612]), .Z(n1484) );
  IV U3559 ( .A(B[2613]), .Z(n1483) );
  IV U3560 ( .A(B[2614]), .Z(n1482) );
  IV U3561 ( .A(B[2615]), .Z(n1481) );
  IV U3562 ( .A(B[2616]), .Z(n1480) );
  IV U3563 ( .A(B[3948]), .Z(n148) );
  IV U3564 ( .A(B[2617]), .Z(n1479) );
  IV U3565 ( .A(B[2618]), .Z(n1478) );
  IV U3566 ( .A(B[2619]), .Z(n1477) );
  IV U3567 ( .A(B[2620]), .Z(n1476) );
  IV U3568 ( .A(B[2621]), .Z(n1475) );
  IV U3569 ( .A(B[2622]), .Z(n1474) );
  IV U3570 ( .A(B[2623]), .Z(n1473) );
  IV U3571 ( .A(B[2624]), .Z(n1472) );
  IV U3572 ( .A(B[2625]), .Z(n1471) );
  IV U3573 ( .A(B[2626]), .Z(n1470) );
  IV U3574 ( .A(B[3949]), .Z(n147) );
  IV U3575 ( .A(B[2627]), .Z(n1469) );
  IV U3576 ( .A(B[2628]), .Z(n1468) );
  IV U3577 ( .A(B[2629]), .Z(n1467) );
  IV U3578 ( .A(B[2630]), .Z(n1466) );
  IV U3579 ( .A(B[2631]), .Z(n1465) );
  IV U3580 ( .A(B[2632]), .Z(n1464) );
  IV U3581 ( .A(B[2633]), .Z(n1463) );
  IV U3582 ( .A(B[2634]), .Z(n1462) );
  IV U3583 ( .A(B[2635]), .Z(n1461) );
  IV U3584 ( .A(B[2636]), .Z(n1460) );
  IV U3585 ( .A(B[3950]), .Z(n146) );
  IV U3586 ( .A(B[2637]), .Z(n1459) );
  IV U3587 ( .A(B[2638]), .Z(n1458) );
  IV U3588 ( .A(B[2639]), .Z(n1457) );
  IV U3589 ( .A(B[2640]), .Z(n1456) );
  IV U3590 ( .A(B[2641]), .Z(n1455) );
  IV U3591 ( .A(B[2642]), .Z(n1454) );
  IV U3592 ( .A(B[2643]), .Z(n1453) );
  IV U3593 ( .A(B[2644]), .Z(n1452) );
  IV U3594 ( .A(B[2645]), .Z(n1451) );
  IV U3595 ( .A(B[2646]), .Z(n1450) );
  IV U3596 ( .A(B[3951]), .Z(n145) );
  IV U3597 ( .A(B[2647]), .Z(n1449) );
  IV U3598 ( .A(B[2648]), .Z(n1448) );
  IV U3599 ( .A(B[2649]), .Z(n1447) );
  IV U3600 ( .A(B[2650]), .Z(n1446) );
  IV U3601 ( .A(B[2651]), .Z(n1445) );
  IV U3602 ( .A(B[2652]), .Z(n1444) );
  IV U3603 ( .A(B[2653]), .Z(n1443) );
  IV U3604 ( .A(B[2654]), .Z(n1442) );
  IV U3605 ( .A(B[2655]), .Z(n1441) );
  IV U3606 ( .A(B[2656]), .Z(n1440) );
  IV U3607 ( .A(B[3952]), .Z(n144) );
  IV U3608 ( .A(B[2657]), .Z(n1439) );
  IV U3609 ( .A(B[2658]), .Z(n1438) );
  IV U3610 ( .A(B[2659]), .Z(n1437) );
  IV U3611 ( .A(B[2660]), .Z(n1436) );
  IV U3612 ( .A(B[2661]), .Z(n1435) );
  IV U3613 ( .A(B[2662]), .Z(n1434) );
  IV U3614 ( .A(B[2663]), .Z(n1433) );
  IV U3615 ( .A(B[2664]), .Z(n1432) );
  IV U3616 ( .A(B[2665]), .Z(n1431) );
  IV U3617 ( .A(B[2666]), .Z(n1430) );
  IV U3618 ( .A(B[3953]), .Z(n143) );
  IV U3619 ( .A(B[2667]), .Z(n1429) );
  IV U3620 ( .A(B[2668]), .Z(n1428) );
  IV U3621 ( .A(B[2669]), .Z(n1427) );
  IV U3622 ( .A(B[2670]), .Z(n1426) );
  IV U3623 ( .A(B[2671]), .Z(n1425) );
  IV U3624 ( .A(B[2672]), .Z(n1424) );
  IV U3625 ( .A(B[2673]), .Z(n1423) );
  IV U3626 ( .A(B[2674]), .Z(n1422) );
  IV U3627 ( .A(B[2675]), .Z(n1421) );
  IV U3628 ( .A(B[2676]), .Z(n1420) );
  IV U3629 ( .A(B[3954]), .Z(n142) );
  IV U3630 ( .A(B[2677]), .Z(n1419) );
  IV U3631 ( .A(B[2678]), .Z(n1418) );
  IV U3632 ( .A(B[2679]), .Z(n1417) );
  IV U3633 ( .A(B[2680]), .Z(n1416) );
  IV U3634 ( .A(B[2681]), .Z(n1415) );
  IV U3635 ( .A(B[2682]), .Z(n1414) );
  IV U3636 ( .A(B[2683]), .Z(n1413) );
  IV U3637 ( .A(B[2684]), .Z(n1412) );
  IV U3638 ( .A(B[2685]), .Z(n1411) );
  IV U3639 ( .A(B[2686]), .Z(n1410) );
  IV U3640 ( .A(B[3955]), .Z(n141) );
  IV U3641 ( .A(B[2687]), .Z(n1409) );
  IV U3642 ( .A(B[2688]), .Z(n1408) );
  IV U3643 ( .A(B[2689]), .Z(n1407) );
  IV U3644 ( .A(B[2690]), .Z(n1406) );
  IV U3645 ( .A(B[2691]), .Z(n1405) );
  IV U3646 ( .A(B[2692]), .Z(n1404) );
  IV U3647 ( .A(B[2693]), .Z(n1403) );
  IV U3648 ( .A(B[2694]), .Z(n1402) );
  IV U3649 ( .A(B[2695]), .Z(n1401) );
  IV U3650 ( .A(B[2696]), .Z(n1400) );
  IV U3651 ( .A(B[3956]), .Z(n140) );
  IV U3652 ( .A(B[4082]), .Z(n14) );
  IV U3653 ( .A(B[2697]), .Z(n1399) );
  IV U3654 ( .A(B[2698]), .Z(n1398) );
  IV U3655 ( .A(B[2699]), .Z(n1397) );
  IV U3656 ( .A(B[2700]), .Z(n1396) );
  IV U3657 ( .A(B[2701]), .Z(n1395) );
  IV U3658 ( .A(B[2702]), .Z(n1394) );
  IV U3659 ( .A(B[2703]), .Z(n1393) );
  IV U3660 ( .A(B[2704]), .Z(n1392) );
  IV U3661 ( .A(B[2705]), .Z(n1391) );
  IV U3662 ( .A(B[2706]), .Z(n1390) );
  IV U3663 ( .A(B[3957]), .Z(n139) );
  IV U3664 ( .A(B[2707]), .Z(n1389) );
  IV U3665 ( .A(B[2708]), .Z(n1388) );
  IV U3666 ( .A(B[2709]), .Z(n1387) );
  IV U3667 ( .A(B[2710]), .Z(n1386) );
  IV U3668 ( .A(B[2711]), .Z(n1385) );
  IV U3669 ( .A(B[2712]), .Z(n1384) );
  IV U3670 ( .A(B[2713]), .Z(n1383) );
  IV U3671 ( .A(B[2714]), .Z(n1382) );
  IV U3672 ( .A(B[2715]), .Z(n1381) );
  IV U3673 ( .A(B[2716]), .Z(n1380) );
  IV U3674 ( .A(B[3958]), .Z(n138) );
  IV U3675 ( .A(B[2717]), .Z(n1379) );
  IV U3676 ( .A(B[2718]), .Z(n1378) );
  IV U3677 ( .A(B[2719]), .Z(n1377) );
  IV U3678 ( .A(B[2720]), .Z(n1376) );
  IV U3679 ( .A(B[2721]), .Z(n1375) );
  IV U3680 ( .A(B[2722]), .Z(n1374) );
  IV U3681 ( .A(B[2723]), .Z(n1373) );
  IV U3682 ( .A(B[2724]), .Z(n1372) );
  IV U3683 ( .A(B[2725]), .Z(n1371) );
  IV U3684 ( .A(B[2726]), .Z(n1370) );
  IV U3685 ( .A(B[3959]), .Z(n137) );
  IV U3686 ( .A(B[2727]), .Z(n1369) );
  IV U3687 ( .A(B[2728]), .Z(n1368) );
  IV U3688 ( .A(B[2729]), .Z(n1367) );
  IV U3689 ( .A(B[2730]), .Z(n1366) );
  IV U3690 ( .A(B[2731]), .Z(n1365) );
  IV U3691 ( .A(B[2732]), .Z(n1364) );
  IV U3692 ( .A(B[2733]), .Z(n1363) );
  IV U3693 ( .A(B[2734]), .Z(n1362) );
  IV U3694 ( .A(B[2735]), .Z(n1361) );
  IV U3695 ( .A(B[2736]), .Z(n1360) );
  IV U3696 ( .A(B[3960]), .Z(n136) );
  IV U3697 ( .A(B[2737]), .Z(n1359) );
  IV U3698 ( .A(B[2738]), .Z(n1358) );
  IV U3699 ( .A(B[2739]), .Z(n1357) );
  IV U3700 ( .A(B[2740]), .Z(n1356) );
  IV U3701 ( .A(B[2741]), .Z(n1355) );
  IV U3702 ( .A(B[2742]), .Z(n1354) );
  IV U3703 ( .A(B[2743]), .Z(n1353) );
  IV U3704 ( .A(B[2744]), .Z(n1352) );
  IV U3705 ( .A(B[2745]), .Z(n1351) );
  IV U3706 ( .A(B[2746]), .Z(n1350) );
  IV U3707 ( .A(B[3961]), .Z(n135) );
  IV U3708 ( .A(B[2747]), .Z(n1349) );
  IV U3709 ( .A(B[2748]), .Z(n1348) );
  IV U3710 ( .A(B[2749]), .Z(n1347) );
  IV U3711 ( .A(B[2750]), .Z(n1346) );
  IV U3712 ( .A(B[2751]), .Z(n1345) );
  IV U3713 ( .A(B[2752]), .Z(n1344) );
  IV U3714 ( .A(B[2753]), .Z(n1343) );
  IV U3715 ( .A(B[2754]), .Z(n1342) );
  IV U3716 ( .A(B[2755]), .Z(n1341) );
  IV U3717 ( .A(B[2756]), .Z(n1340) );
  IV U3718 ( .A(B[3962]), .Z(n134) );
  IV U3719 ( .A(B[2757]), .Z(n1339) );
  IV U3720 ( .A(B[2758]), .Z(n1338) );
  IV U3721 ( .A(B[2759]), .Z(n1337) );
  IV U3722 ( .A(B[2760]), .Z(n1336) );
  IV U3723 ( .A(B[2761]), .Z(n1335) );
  IV U3724 ( .A(B[2762]), .Z(n1334) );
  IV U3725 ( .A(B[2763]), .Z(n1333) );
  IV U3726 ( .A(B[2764]), .Z(n1332) );
  IV U3727 ( .A(B[2765]), .Z(n1331) );
  IV U3728 ( .A(B[2766]), .Z(n1330) );
  IV U3729 ( .A(B[3963]), .Z(n133) );
  IV U3730 ( .A(B[2767]), .Z(n1329) );
  IV U3731 ( .A(B[2768]), .Z(n1328) );
  IV U3732 ( .A(B[2769]), .Z(n1327) );
  IV U3733 ( .A(B[2770]), .Z(n1326) );
  IV U3734 ( .A(B[2771]), .Z(n1325) );
  IV U3735 ( .A(B[2772]), .Z(n1324) );
  IV U3736 ( .A(B[2773]), .Z(n1323) );
  IV U3737 ( .A(B[2774]), .Z(n1322) );
  IV U3738 ( .A(B[2775]), .Z(n1321) );
  IV U3739 ( .A(B[2776]), .Z(n1320) );
  IV U3740 ( .A(B[3964]), .Z(n132) );
  IV U3741 ( .A(B[2777]), .Z(n1319) );
  IV U3742 ( .A(B[2778]), .Z(n1318) );
  IV U3743 ( .A(B[2779]), .Z(n1317) );
  IV U3744 ( .A(B[2780]), .Z(n1316) );
  IV U3745 ( .A(B[2781]), .Z(n1315) );
  IV U3746 ( .A(B[2782]), .Z(n1314) );
  IV U3747 ( .A(B[2783]), .Z(n1313) );
  IV U3748 ( .A(B[2784]), .Z(n1312) );
  IV U3749 ( .A(B[2785]), .Z(n1311) );
  IV U3750 ( .A(B[2786]), .Z(n1310) );
  IV U3751 ( .A(B[3965]), .Z(n131) );
  IV U3752 ( .A(B[2787]), .Z(n1309) );
  IV U3753 ( .A(B[2788]), .Z(n1308) );
  IV U3754 ( .A(B[2789]), .Z(n1307) );
  IV U3755 ( .A(B[2790]), .Z(n1306) );
  IV U3756 ( .A(B[2791]), .Z(n1305) );
  IV U3757 ( .A(B[2792]), .Z(n1304) );
  IV U3758 ( .A(B[2793]), .Z(n1303) );
  IV U3759 ( .A(B[2794]), .Z(n1302) );
  IV U3760 ( .A(B[2795]), .Z(n1301) );
  IV U3761 ( .A(B[2796]), .Z(n1300) );
  IV U3762 ( .A(B[3966]), .Z(n130) );
  IV U3763 ( .A(B[4083]), .Z(n13) );
  IV U3764 ( .A(B[2797]), .Z(n1299) );
  IV U3765 ( .A(B[2798]), .Z(n1298) );
  IV U3766 ( .A(B[2799]), .Z(n1297) );
  IV U3767 ( .A(B[2800]), .Z(n1296) );
  IV U3768 ( .A(B[2801]), .Z(n1295) );
  IV U3769 ( .A(B[2802]), .Z(n1294) );
  IV U3770 ( .A(B[2803]), .Z(n1293) );
  IV U3771 ( .A(B[2804]), .Z(n1292) );
  IV U3772 ( .A(B[2805]), .Z(n1291) );
  IV U3773 ( .A(B[2806]), .Z(n1290) );
  IV U3774 ( .A(B[3967]), .Z(n129) );
  IV U3775 ( .A(B[2807]), .Z(n1289) );
  IV U3776 ( .A(B[2808]), .Z(n1288) );
  IV U3777 ( .A(B[2809]), .Z(n1287) );
  IV U3778 ( .A(B[2810]), .Z(n1286) );
  IV U3779 ( .A(B[2811]), .Z(n1285) );
  IV U3780 ( .A(B[2812]), .Z(n1284) );
  IV U3781 ( .A(B[2813]), .Z(n1283) );
  IV U3782 ( .A(B[2814]), .Z(n1282) );
  IV U3783 ( .A(B[2815]), .Z(n1281) );
  IV U3784 ( .A(B[2816]), .Z(n1280) );
  IV U3785 ( .A(B[3968]), .Z(n128) );
  IV U3786 ( .A(B[2817]), .Z(n1279) );
  IV U3787 ( .A(B[2818]), .Z(n1278) );
  IV U3788 ( .A(B[2819]), .Z(n1277) );
  IV U3789 ( .A(B[2820]), .Z(n1276) );
  IV U3790 ( .A(B[2821]), .Z(n1275) );
  IV U3791 ( .A(B[2822]), .Z(n1274) );
  IV U3792 ( .A(B[2823]), .Z(n1273) );
  IV U3793 ( .A(B[2824]), .Z(n1272) );
  IV U3794 ( .A(B[2825]), .Z(n1271) );
  IV U3795 ( .A(B[2826]), .Z(n1270) );
  IV U3796 ( .A(B[3969]), .Z(n127) );
  IV U3797 ( .A(B[2827]), .Z(n1269) );
  IV U3798 ( .A(B[2828]), .Z(n1268) );
  IV U3799 ( .A(B[2829]), .Z(n1267) );
  IV U3800 ( .A(B[2830]), .Z(n1266) );
  IV U3801 ( .A(B[2831]), .Z(n1265) );
  IV U3802 ( .A(B[2832]), .Z(n1264) );
  IV U3803 ( .A(B[2833]), .Z(n1263) );
  IV U3804 ( .A(B[2834]), .Z(n1262) );
  IV U3805 ( .A(B[2835]), .Z(n1261) );
  IV U3806 ( .A(B[2836]), .Z(n1260) );
  IV U3807 ( .A(B[3970]), .Z(n126) );
  IV U3808 ( .A(B[2837]), .Z(n1259) );
  IV U3809 ( .A(B[2838]), .Z(n1258) );
  IV U3810 ( .A(B[2839]), .Z(n1257) );
  IV U3811 ( .A(B[2840]), .Z(n1256) );
  IV U3812 ( .A(B[2841]), .Z(n1255) );
  IV U3813 ( .A(B[2842]), .Z(n1254) );
  IV U3814 ( .A(B[2843]), .Z(n1253) );
  IV U3815 ( .A(B[2844]), .Z(n1252) );
  IV U3816 ( .A(B[2845]), .Z(n1251) );
  IV U3817 ( .A(B[2846]), .Z(n1250) );
  IV U3818 ( .A(B[3971]), .Z(n125) );
  IV U3819 ( .A(B[2847]), .Z(n1249) );
  IV U3820 ( .A(B[2848]), .Z(n1248) );
  IV U3821 ( .A(B[2849]), .Z(n1247) );
  IV U3822 ( .A(B[2850]), .Z(n1246) );
  IV U3823 ( .A(B[2851]), .Z(n1245) );
  IV U3824 ( .A(B[2852]), .Z(n1244) );
  IV U3825 ( .A(B[2853]), .Z(n1243) );
  IV U3826 ( .A(B[2854]), .Z(n1242) );
  IV U3827 ( .A(B[2855]), .Z(n1241) );
  IV U3828 ( .A(B[2856]), .Z(n1240) );
  IV U3829 ( .A(B[3972]), .Z(n124) );
  IV U3830 ( .A(B[2857]), .Z(n1239) );
  IV U3831 ( .A(B[2858]), .Z(n1238) );
  IV U3832 ( .A(B[2859]), .Z(n1237) );
  IV U3833 ( .A(B[2860]), .Z(n1236) );
  IV U3834 ( .A(B[2861]), .Z(n1235) );
  IV U3835 ( .A(B[2862]), .Z(n1234) );
  IV U3836 ( .A(B[2863]), .Z(n1233) );
  IV U3837 ( .A(B[2864]), .Z(n1232) );
  IV U3838 ( .A(B[2865]), .Z(n1231) );
  IV U3839 ( .A(B[2866]), .Z(n1230) );
  IV U3840 ( .A(B[3973]), .Z(n123) );
  IV U3841 ( .A(B[2867]), .Z(n1229) );
  IV U3842 ( .A(B[2868]), .Z(n1228) );
  IV U3843 ( .A(B[2869]), .Z(n1227) );
  IV U3844 ( .A(B[2870]), .Z(n1226) );
  IV U3845 ( .A(B[2871]), .Z(n1225) );
  IV U3846 ( .A(B[2872]), .Z(n1224) );
  IV U3847 ( .A(B[2873]), .Z(n1223) );
  IV U3848 ( .A(B[2874]), .Z(n1222) );
  IV U3849 ( .A(B[2875]), .Z(n1221) );
  IV U3850 ( .A(B[2876]), .Z(n1220) );
  IV U3851 ( .A(B[3974]), .Z(n122) );
  IV U3852 ( .A(B[2877]), .Z(n1219) );
  IV U3853 ( .A(B[2878]), .Z(n1218) );
  IV U3854 ( .A(B[2879]), .Z(n1217) );
  IV U3855 ( .A(B[2880]), .Z(n1216) );
  IV U3856 ( .A(B[2881]), .Z(n1215) );
  IV U3857 ( .A(B[2882]), .Z(n1214) );
  IV U3858 ( .A(B[2883]), .Z(n1213) );
  IV U3859 ( .A(B[2884]), .Z(n1212) );
  IV U3860 ( .A(B[2885]), .Z(n1211) );
  IV U3861 ( .A(B[2886]), .Z(n1210) );
  IV U3862 ( .A(B[3975]), .Z(n121) );
  IV U3863 ( .A(B[2887]), .Z(n1209) );
  IV U3864 ( .A(B[2888]), .Z(n1208) );
  IV U3865 ( .A(B[2889]), .Z(n1207) );
  IV U3866 ( .A(B[2890]), .Z(n1206) );
  IV U3867 ( .A(B[2891]), .Z(n1205) );
  IV U3868 ( .A(B[2892]), .Z(n1204) );
  IV U3869 ( .A(B[2893]), .Z(n1203) );
  IV U3870 ( .A(B[2894]), .Z(n1202) );
  IV U3871 ( .A(B[2895]), .Z(n1201) );
  IV U3872 ( .A(B[2896]), .Z(n1200) );
  IV U3873 ( .A(B[3976]), .Z(n120) );
  IV U3874 ( .A(B[4084]), .Z(n12) );
  IV U3875 ( .A(B[2897]), .Z(n1199) );
  IV U3876 ( .A(B[2898]), .Z(n1198) );
  IV U3877 ( .A(B[2899]), .Z(n1197) );
  IV U3878 ( .A(B[2900]), .Z(n1196) );
  IV U3879 ( .A(B[2901]), .Z(n1195) );
  IV U3880 ( .A(B[2902]), .Z(n1194) );
  IV U3881 ( .A(B[2903]), .Z(n1193) );
  IV U3882 ( .A(B[2904]), .Z(n1192) );
  IV U3883 ( .A(B[2905]), .Z(n1191) );
  IV U3884 ( .A(B[2906]), .Z(n1190) );
  IV U3885 ( .A(B[3977]), .Z(n119) );
  IV U3886 ( .A(B[2907]), .Z(n1189) );
  IV U3887 ( .A(B[2908]), .Z(n1188) );
  IV U3888 ( .A(B[2909]), .Z(n1187) );
  IV U3889 ( .A(B[2910]), .Z(n1186) );
  IV U3890 ( .A(B[2911]), .Z(n1185) );
  IV U3891 ( .A(B[2912]), .Z(n1184) );
  IV U3892 ( .A(B[2913]), .Z(n1183) );
  IV U3893 ( .A(B[2914]), .Z(n1182) );
  IV U3894 ( .A(B[2915]), .Z(n1181) );
  IV U3895 ( .A(B[2916]), .Z(n1180) );
  IV U3896 ( .A(B[3978]), .Z(n118) );
  IV U3897 ( .A(B[2917]), .Z(n1179) );
  IV U3898 ( .A(B[2918]), .Z(n1178) );
  IV U3899 ( .A(B[2919]), .Z(n1177) );
  IV U3900 ( .A(B[2920]), .Z(n1176) );
  IV U3901 ( .A(B[2921]), .Z(n1175) );
  IV U3902 ( .A(B[2922]), .Z(n1174) );
  IV U3903 ( .A(B[2923]), .Z(n1173) );
  IV U3904 ( .A(B[2924]), .Z(n1172) );
  IV U3905 ( .A(B[2925]), .Z(n1171) );
  IV U3906 ( .A(B[2926]), .Z(n1170) );
  IV U3907 ( .A(B[3979]), .Z(n117) );
  IV U3908 ( .A(B[2927]), .Z(n1169) );
  IV U3909 ( .A(B[2928]), .Z(n1168) );
  IV U3910 ( .A(B[2929]), .Z(n1167) );
  IV U3911 ( .A(B[2930]), .Z(n1166) );
  IV U3912 ( .A(B[2931]), .Z(n1165) );
  IV U3913 ( .A(B[2932]), .Z(n1164) );
  IV U3914 ( .A(B[2933]), .Z(n1163) );
  IV U3915 ( .A(B[2934]), .Z(n1162) );
  IV U3916 ( .A(B[2935]), .Z(n1161) );
  IV U3917 ( .A(B[2936]), .Z(n1160) );
  IV U3918 ( .A(B[3980]), .Z(n116) );
  IV U3919 ( .A(B[2937]), .Z(n1159) );
  IV U3920 ( .A(B[2938]), .Z(n1158) );
  IV U3921 ( .A(B[2939]), .Z(n1157) );
  IV U3922 ( .A(B[2940]), .Z(n1156) );
  IV U3923 ( .A(B[2941]), .Z(n1155) );
  IV U3924 ( .A(B[2942]), .Z(n1154) );
  IV U3925 ( .A(B[2943]), .Z(n1153) );
  IV U3926 ( .A(B[2944]), .Z(n1152) );
  IV U3927 ( .A(B[2945]), .Z(n1151) );
  IV U3928 ( .A(B[2946]), .Z(n1150) );
  IV U3929 ( .A(B[3981]), .Z(n115) );
  IV U3930 ( .A(B[2947]), .Z(n1149) );
  IV U3931 ( .A(B[2948]), .Z(n1148) );
  IV U3932 ( .A(B[2949]), .Z(n1147) );
  IV U3933 ( .A(B[2950]), .Z(n1146) );
  IV U3934 ( .A(B[2951]), .Z(n1145) );
  IV U3935 ( .A(B[2952]), .Z(n1144) );
  IV U3936 ( .A(B[2953]), .Z(n1143) );
  IV U3937 ( .A(B[2954]), .Z(n1142) );
  IV U3938 ( .A(B[2955]), .Z(n1141) );
  IV U3939 ( .A(B[2956]), .Z(n1140) );
  IV U3940 ( .A(B[3982]), .Z(n114) );
  IV U3941 ( .A(B[2957]), .Z(n1139) );
  IV U3942 ( .A(B[2958]), .Z(n1138) );
  IV U3943 ( .A(B[2959]), .Z(n1137) );
  IV U3944 ( .A(B[2960]), .Z(n1136) );
  IV U3945 ( .A(B[2961]), .Z(n1135) );
  IV U3946 ( .A(B[2962]), .Z(n1134) );
  IV U3947 ( .A(B[2963]), .Z(n1133) );
  IV U3948 ( .A(B[2964]), .Z(n1132) );
  IV U3949 ( .A(B[2965]), .Z(n1131) );
  IV U3950 ( .A(B[2966]), .Z(n1130) );
  IV U3951 ( .A(B[3983]), .Z(n113) );
  IV U3952 ( .A(B[2967]), .Z(n1129) );
  IV U3953 ( .A(B[2968]), .Z(n1128) );
  IV U3954 ( .A(B[2969]), .Z(n1127) );
  IV U3955 ( .A(B[2970]), .Z(n1126) );
  IV U3956 ( .A(B[2971]), .Z(n1125) );
  IV U3957 ( .A(B[2972]), .Z(n1124) );
  IV U3958 ( .A(B[2973]), .Z(n1123) );
  IV U3959 ( .A(B[2974]), .Z(n1122) );
  IV U3960 ( .A(B[2975]), .Z(n1121) );
  IV U3961 ( .A(B[2976]), .Z(n1120) );
  IV U3962 ( .A(B[3984]), .Z(n112) );
  IV U3963 ( .A(B[2977]), .Z(n1119) );
  IV U3964 ( .A(B[2978]), .Z(n1118) );
  IV U3965 ( .A(B[2979]), .Z(n1117) );
  IV U3966 ( .A(B[2980]), .Z(n1116) );
  IV U3967 ( .A(B[2981]), .Z(n1115) );
  IV U3968 ( .A(B[2982]), .Z(n1114) );
  IV U3969 ( .A(B[2983]), .Z(n1113) );
  IV U3970 ( .A(B[2984]), .Z(n1112) );
  IV U3971 ( .A(B[2985]), .Z(n1111) );
  IV U3972 ( .A(B[2986]), .Z(n1110) );
  IV U3973 ( .A(B[3985]), .Z(n111) );
  IV U3974 ( .A(B[2987]), .Z(n1109) );
  IV U3975 ( .A(B[2988]), .Z(n1108) );
  IV U3976 ( .A(B[2989]), .Z(n1107) );
  IV U3977 ( .A(B[2990]), .Z(n1106) );
  IV U3978 ( .A(B[2991]), .Z(n1105) );
  IV U3979 ( .A(B[2992]), .Z(n1104) );
  IV U3980 ( .A(B[2993]), .Z(n1103) );
  IV U3981 ( .A(B[2994]), .Z(n1102) );
  IV U3982 ( .A(B[2995]), .Z(n1101) );
  IV U3983 ( .A(B[2996]), .Z(n1100) );
  IV U3984 ( .A(B[3986]), .Z(n110) );
  IV U3985 ( .A(B[4085]), .Z(n11) );
  IV U3986 ( .A(B[2997]), .Z(n1099) );
  IV U3987 ( .A(B[2998]), .Z(n1098) );
  IV U3988 ( .A(B[2999]), .Z(n1097) );
  IV U3989 ( .A(B[3000]), .Z(n1096) );
  IV U3990 ( .A(B[3001]), .Z(n1095) );
  IV U3991 ( .A(B[3002]), .Z(n1094) );
  IV U3992 ( .A(B[3003]), .Z(n1093) );
  IV U3993 ( .A(B[3004]), .Z(n1092) );
  IV U3994 ( .A(B[3005]), .Z(n1091) );
  IV U3995 ( .A(B[3006]), .Z(n1090) );
  IV U3996 ( .A(B[3987]), .Z(n109) );
  IV U3997 ( .A(B[3007]), .Z(n1089) );
  IV U3998 ( .A(B[3008]), .Z(n1088) );
  IV U3999 ( .A(B[3009]), .Z(n1087) );
  IV U4000 ( .A(B[3010]), .Z(n1086) );
  IV U4001 ( .A(B[3011]), .Z(n1085) );
  IV U4002 ( .A(B[3012]), .Z(n1084) );
  IV U4003 ( .A(B[3013]), .Z(n1083) );
  IV U4004 ( .A(B[3014]), .Z(n1082) );
  IV U4005 ( .A(B[3015]), .Z(n1081) );
  IV U4006 ( .A(B[3016]), .Z(n1080) );
  IV U4007 ( .A(B[3988]), .Z(n108) );
  IV U4008 ( .A(B[3017]), .Z(n1079) );
  IV U4009 ( .A(B[3018]), .Z(n1078) );
  IV U4010 ( .A(B[3019]), .Z(n1077) );
  IV U4011 ( .A(B[3020]), .Z(n1076) );
  IV U4012 ( .A(B[3021]), .Z(n1075) );
  IV U4013 ( .A(B[3022]), .Z(n1074) );
  IV U4014 ( .A(B[3023]), .Z(n1073) );
  IV U4015 ( .A(B[3024]), .Z(n1072) );
  IV U4016 ( .A(B[3025]), .Z(n1071) );
  IV U4017 ( .A(B[3026]), .Z(n1070) );
  IV U4018 ( .A(B[3989]), .Z(n107) );
  IV U4019 ( .A(B[3027]), .Z(n1069) );
  IV U4020 ( .A(B[3028]), .Z(n1068) );
  IV U4021 ( .A(B[3029]), .Z(n1067) );
  IV U4022 ( .A(B[3030]), .Z(n1066) );
  IV U4023 ( .A(B[3031]), .Z(n1065) );
  IV U4024 ( .A(B[3032]), .Z(n1064) );
  IV U4025 ( .A(B[3033]), .Z(n1063) );
  IV U4026 ( .A(B[3034]), .Z(n1062) );
  IV U4027 ( .A(B[3035]), .Z(n1061) );
  IV U4028 ( .A(B[3036]), .Z(n1060) );
  IV U4029 ( .A(B[3990]), .Z(n106) );
  IV U4030 ( .A(B[3037]), .Z(n1059) );
  IV U4031 ( .A(B[3038]), .Z(n1058) );
  IV U4032 ( .A(B[3039]), .Z(n1057) );
  IV U4033 ( .A(B[3040]), .Z(n1056) );
  IV U4034 ( .A(B[3041]), .Z(n1055) );
  IV U4035 ( .A(B[3042]), .Z(n1054) );
  IV U4036 ( .A(B[3043]), .Z(n1053) );
  IV U4037 ( .A(B[3044]), .Z(n1052) );
  IV U4038 ( .A(B[3045]), .Z(n1051) );
  IV U4039 ( .A(B[3046]), .Z(n1050) );
  IV U4040 ( .A(B[3991]), .Z(n105) );
  IV U4041 ( .A(B[3047]), .Z(n1049) );
  IV U4042 ( .A(B[3048]), .Z(n1048) );
  IV U4043 ( .A(B[3049]), .Z(n1047) );
  IV U4044 ( .A(B[3050]), .Z(n1046) );
  IV U4045 ( .A(B[3051]), .Z(n1045) );
  IV U4046 ( .A(B[3052]), .Z(n1044) );
  IV U4047 ( .A(B[3053]), .Z(n1043) );
  IV U4048 ( .A(B[3054]), .Z(n1042) );
  IV U4049 ( .A(B[3055]), .Z(n1041) );
  IV U4050 ( .A(B[3056]), .Z(n1040) );
  IV U4051 ( .A(B[3992]), .Z(n104) );
  IV U4052 ( .A(B[3057]), .Z(n1039) );
  IV U4053 ( .A(B[3058]), .Z(n1038) );
  IV U4054 ( .A(B[3059]), .Z(n1037) );
  IV U4055 ( .A(B[3060]), .Z(n1036) );
  IV U4056 ( .A(B[3061]), .Z(n1035) );
  IV U4057 ( .A(B[3062]), .Z(n1034) );
  IV U4058 ( .A(B[3063]), .Z(n1033) );
  IV U4059 ( .A(B[3064]), .Z(n1032) );
  IV U4060 ( .A(B[3065]), .Z(n1031) );
  IV U4061 ( .A(B[3066]), .Z(n1030) );
  IV U4062 ( .A(B[3993]), .Z(n103) );
  IV U4063 ( .A(B[3067]), .Z(n1029) );
  IV U4064 ( .A(B[3068]), .Z(n1028) );
  IV U4065 ( .A(B[3069]), .Z(n1027) );
  IV U4066 ( .A(B[3070]), .Z(n1026) );
  IV U4067 ( .A(B[3071]), .Z(n1025) );
  IV U4068 ( .A(B[3072]), .Z(n1024) );
  IV U4069 ( .A(B[3073]), .Z(n1023) );
  IV U4070 ( .A(B[3074]), .Z(n1022) );
  IV U4071 ( .A(B[3075]), .Z(n1021) );
  IV U4072 ( .A(B[3076]), .Z(n1020) );
  IV U4073 ( .A(B[3994]), .Z(n102) );
  IV U4074 ( .A(B[3077]), .Z(n1019) );
  IV U4075 ( .A(B[3078]), .Z(n1018) );
  IV U4076 ( .A(B[3079]), .Z(n1017) );
  IV U4077 ( .A(B[3080]), .Z(n1016) );
  IV U4078 ( .A(B[3081]), .Z(n1015) );
  IV U4079 ( .A(B[3082]), .Z(n1014) );
  IV U4080 ( .A(B[3083]), .Z(n1013) );
  IV U4081 ( .A(B[3084]), .Z(n1012) );
  IV U4082 ( .A(B[3085]), .Z(n1011) );
  IV U4083 ( .A(B[3086]), .Z(n1010) );
  IV U4084 ( .A(B[3995]), .Z(n101) );
  IV U4085 ( .A(B[3087]), .Z(n1009) );
  IV U4086 ( .A(B[3088]), .Z(n1008) );
  IV U4087 ( .A(B[3089]), .Z(n1007) );
  IV U4088 ( .A(B[3090]), .Z(n1006) );
  IV U4089 ( .A(B[3091]), .Z(n1005) );
  IV U4090 ( .A(B[3092]), .Z(n1004) );
  IV U4091 ( .A(B[3093]), .Z(n1003) );
  IV U4092 ( .A(B[3094]), .Z(n1002) );
  IV U4093 ( .A(B[3095]), .Z(n1001) );
  IV U4094 ( .A(B[3096]), .Z(n1000) );
  IV U4095 ( .A(B[3996]), .Z(n100) );
  IV U4096 ( .A(B[4086]), .Z(n10) );
  IV U4097 ( .A(B[4095]), .Z(n1) );
endmodule


module compare_N16384_CC4 ( clk, rst, x, y, g, e );
  input [4095:0] x;
  input [4095:0] y;
  input clk, rst;
  output g, e;
  wire   xly, ebreg, ebnew, gnew, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389;

  COMP_N4096 UCOMP ( .A(x), .B(y), .O(xly) );
  DFF ebreg_reg ( .D(ebnew), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(gnew), .CLK(clk), .RST(rst), .Q(g) );
  XOR U8200 ( .A(g), .B(n8196), .Z(gnew) );
  AND U8201 ( .A(n8197), .B(n8198), .Z(n8196) );
  XOR U8202 ( .A(xly), .B(g), .Z(n8198) );
  OR U8203 ( .A(n8197), .B(ebreg), .Z(ebnew) );
  AND U8204 ( .A(n8199), .B(e), .Z(n8197) );
  NAND U8205 ( .A(n8200), .B(n8201), .Z(n8199) );
  AND U8206 ( .A(n8202), .B(n8203), .Z(n8201) );
  AND U8207 ( .A(n8204), .B(n8205), .Z(n8203) );
  AND U8208 ( .A(n8206), .B(n8207), .Z(n8205) );
  AND U8209 ( .A(n8208), .B(n8209), .Z(n8207) );
  AND U8210 ( .A(n8210), .B(n8211), .Z(n8209) );
  AND U8211 ( .A(n8212), .B(n8213), .Z(n8211) );
  AND U8212 ( .A(n8214), .B(n8215), .Z(n8213) );
  AND U8213 ( .A(n8216), .B(n8217), .Z(n8215) );
  AND U8214 ( .A(n8218), .B(n8219), .Z(n8217) );
  AND U8215 ( .A(n8220), .B(n8221), .Z(n8219) );
  AND U8216 ( .A(n8222), .B(n8223), .Z(n8221) );
  AND U8217 ( .A(n8224), .B(n8225), .Z(n8223) );
  AND U8218 ( .A(n8226), .B(n8227), .Z(n8225) );
  AND U8219 ( .A(n8228), .B(n8229), .Z(n8227) );
  AND U8220 ( .A(n8230), .B(n8231), .Z(n8229) );
  AND U8221 ( .A(n8232), .B(n8233), .Z(n8231) );
  XNOR U8222 ( .A(y[0]), .B(x[0]), .Z(n8233) );
  XNOR U8223 ( .A(y[1]), .B(x[1]), .Z(n8232) );
  AND U8224 ( .A(n8234), .B(n8235), .Z(n8230) );
  XNOR U8225 ( .A(y[2]), .B(x[2]), .Z(n8235) );
  XNOR U8226 ( .A(y[3]), .B(x[3]), .Z(n8234) );
  AND U8227 ( .A(n8236), .B(n8237), .Z(n8228) );
  XNOR U8228 ( .A(y[5]), .B(x[5]), .Z(n8237) );
  AND U8229 ( .A(n8238), .B(n8239), .Z(n8236) );
  XNOR U8230 ( .A(y[6]), .B(x[6]), .Z(n8239) );
  XNOR U8231 ( .A(y[4]), .B(x[4]), .Z(n8238) );
  AND U8232 ( .A(n8240), .B(n8241), .Z(n8226) );
  AND U8233 ( .A(n8242), .B(n8243), .Z(n8241) );
  XNOR U8234 ( .A(y[8]), .B(x[8]), .Z(n8243) );
  AND U8235 ( .A(n8244), .B(n8245), .Z(n8242) );
  XNOR U8236 ( .A(y[9]), .B(x[9]), .Z(n8245) );
  XNOR U8237 ( .A(y[7]), .B(x[7]), .Z(n8244) );
  AND U8238 ( .A(n8246), .B(n8247), .Z(n8240) );
  XNOR U8239 ( .A(y[11]), .B(x[11]), .Z(n8247) );
  AND U8240 ( .A(n8248), .B(n8249), .Z(n8246) );
  XNOR U8241 ( .A(y[12]), .B(x[12]), .Z(n8249) );
  XNOR U8242 ( .A(y[10]), .B(x[10]), .Z(n8248) );
  AND U8243 ( .A(n8250), .B(n8251), .Z(n8224) );
  AND U8244 ( .A(n8252), .B(n8253), .Z(n8251) );
  AND U8245 ( .A(n8254), .B(n8255), .Z(n8253) );
  XNOR U8246 ( .A(y[14]), .B(x[14]), .Z(n8255) );
  AND U8247 ( .A(n8256), .B(n8257), .Z(n8254) );
  XNOR U8248 ( .A(y[17]), .B(x[17]), .Z(n8257) );
  XNOR U8249 ( .A(y[13]), .B(x[13]), .Z(n8256) );
  AND U8250 ( .A(n8258), .B(n8259), .Z(n8252) );
  XNOR U8251 ( .A(y[16]), .B(x[16]), .Z(n8259) );
  AND U8252 ( .A(n8260), .B(n8261), .Z(n8258) );
  XNOR U8253 ( .A(y[18]), .B(x[18]), .Z(n8261) );
  XNOR U8254 ( .A(y[15]), .B(x[15]), .Z(n8260) );
  AND U8255 ( .A(n8262), .B(n8263), .Z(n8250) );
  AND U8256 ( .A(n8264), .B(n8265), .Z(n8263) );
  XNOR U8257 ( .A(y[20]), .B(x[20]), .Z(n8265) );
  AND U8258 ( .A(n8266), .B(n8267), .Z(n8264) );
  XNOR U8259 ( .A(y[21]), .B(x[21]), .Z(n8267) );
  XNOR U8260 ( .A(y[19]), .B(x[19]), .Z(n8266) );
  AND U8261 ( .A(n8268), .B(n8269), .Z(n8262) );
  XNOR U8262 ( .A(y[23]), .B(x[23]), .Z(n8269) );
  AND U8263 ( .A(n8270), .B(n8271), .Z(n8268) );
  XNOR U8264 ( .A(y[24]), .B(x[24]), .Z(n8271) );
  XNOR U8265 ( .A(y[22]), .B(x[22]), .Z(n8270) );
  AND U8266 ( .A(n8272), .B(n8273), .Z(n8222) );
  AND U8267 ( .A(n8274), .B(n8275), .Z(n8273) );
  AND U8268 ( .A(n8276), .B(n8277), .Z(n8275) );
  AND U8269 ( .A(n8278), .B(n8279), .Z(n8277) );
  AND U8270 ( .A(n8280), .B(n8281), .Z(n8279) );
  XNOR U8271 ( .A(y[25]), .B(x[25]), .Z(n8281) );
  XNOR U8272 ( .A(y[26]), .B(x[26]), .Z(n8280) );
  AND U8273 ( .A(n8282), .B(n8283), .Z(n8278) );
  XNOR U8274 ( .A(y[27]), .B(x[27]), .Z(n8283) );
  XNOR U8275 ( .A(y[28]), .B(x[28]), .Z(n8282) );
  AND U8276 ( .A(n8284), .B(n8285), .Z(n8276) );
  XNOR U8277 ( .A(y[30]), .B(x[30]), .Z(n8285) );
  AND U8278 ( .A(n8286), .B(n8287), .Z(n8284) );
  XNOR U8279 ( .A(y[31]), .B(x[31]), .Z(n8287) );
  XNOR U8280 ( .A(y[29]), .B(x[29]), .Z(n8286) );
  AND U8281 ( .A(n8288), .B(n8289), .Z(n8274) );
  AND U8282 ( .A(n8290), .B(n8291), .Z(n8289) );
  XNOR U8283 ( .A(y[33]), .B(x[33]), .Z(n8291) );
  AND U8284 ( .A(n8292), .B(n8293), .Z(n8290) );
  XNOR U8285 ( .A(y[34]), .B(x[34]), .Z(n8293) );
  XNOR U8286 ( .A(y[32]), .B(x[32]), .Z(n8292) );
  AND U8287 ( .A(n8294), .B(n8295), .Z(n8288) );
  XNOR U8288 ( .A(y[36]), .B(x[36]), .Z(n8295) );
  AND U8289 ( .A(n8296), .B(n8297), .Z(n8294) );
  XNOR U8290 ( .A(y[37]), .B(x[37]), .Z(n8297) );
  XNOR U8291 ( .A(y[35]), .B(x[35]), .Z(n8296) );
  AND U8292 ( .A(n8298), .B(n8299), .Z(n8272) );
  AND U8293 ( .A(n8300), .B(n8301), .Z(n8299) );
  AND U8294 ( .A(n8302), .B(n8303), .Z(n8301) );
  XNOR U8295 ( .A(y[39]), .B(x[39]), .Z(n8303) );
  AND U8296 ( .A(n8304), .B(n8305), .Z(n8302) );
  XNOR U8297 ( .A(y[40]), .B(x[40]), .Z(n8305) );
  XNOR U8298 ( .A(y[38]), .B(x[38]), .Z(n8304) );
  AND U8299 ( .A(n8306), .B(n8307), .Z(n8300) );
  XNOR U8300 ( .A(y[42]), .B(x[42]), .Z(n8307) );
  AND U8301 ( .A(n8308), .B(n8309), .Z(n8306) );
  XNOR U8302 ( .A(y[43]), .B(x[43]), .Z(n8309) );
  XNOR U8303 ( .A(y[41]), .B(x[41]), .Z(n8308) );
  AND U8304 ( .A(n8310), .B(n8311), .Z(n8298) );
  AND U8305 ( .A(n8312), .B(n8313), .Z(n8311) );
  XNOR U8306 ( .A(y[45]), .B(x[45]), .Z(n8313) );
  AND U8307 ( .A(n8314), .B(n8315), .Z(n8312) );
  XNOR U8308 ( .A(y[46]), .B(x[46]), .Z(n8315) );
  XNOR U8309 ( .A(y[44]), .B(x[44]), .Z(n8314) );
  AND U8310 ( .A(n8316), .B(n8317), .Z(n8310) );
  XNOR U8311 ( .A(y[48]), .B(x[48]), .Z(n8317) );
  AND U8312 ( .A(n8318), .B(n8319), .Z(n8316) );
  XNOR U8313 ( .A(y[49]), .B(x[49]), .Z(n8319) );
  XNOR U8314 ( .A(y[47]), .B(x[47]), .Z(n8318) );
  AND U8315 ( .A(n8320), .B(n8321), .Z(n8220) );
  AND U8316 ( .A(n8322), .B(n8323), .Z(n8321) );
  AND U8317 ( .A(n8324), .B(n8325), .Z(n8323) );
  AND U8318 ( .A(n8326), .B(n8327), .Z(n8325) );
  AND U8319 ( .A(n8328), .B(n8329), .Z(n8327) );
  AND U8320 ( .A(n8330), .B(n8331), .Z(n8329) );
  XNOR U8321 ( .A(y[50]), .B(x[50]), .Z(n8331) );
  XNOR U8322 ( .A(y[51]), .B(x[51]), .Z(n8330) );
  AND U8323 ( .A(n8332), .B(n8333), .Z(n8328) );
  XNOR U8324 ( .A(y[52]), .B(x[52]), .Z(n8333) );
  XNOR U8325 ( .A(y[53]), .B(x[53]), .Z(n8332) );
  AND U8326 ( .A(n8334), .B(n8335), .Z(n8326) );
  XNOR U8327 ( .A(y[55]), .B(x[55]), .Z(n8335) );
  AND U8328 ( .A(n8336), .B(n8337), .Z(n8334) );
  XNOR U8329 ( .A(y[56]), .B(x[56]), .Z(n8337) );
  XNOR U8330 ( .A(y[54]), .B(x[54]), .Z(n8336) );
  AND U8331 ( .A(n8338), .B(n8339), .Z(n8324) );
  AND U8332 ( .A(n8340), .B(n8341), .Z(n8339) );
  XNOR U8333 ( .A(y[58]), .B(x[58]), .Z(n8341) );
  AND U8334 ( .A(n8342), .B(n8343), .Z(n8340) );
  XNOR U8335 ( .A(y[59]), .B(x[59]), .Z(n8343) );
  XNOR U8336 ( .A(y[57]), .B(x[57]), .Z(n8342) );
  AND U8337 ( .A(n8344), .B(n8345), .Z(n8338) );
  XNOR U8338 ( .A(y[61]), .B(x[61]), .Z(n8345) );
  AND U8339 ( .A(n8346), .B(n8347), .Z(n8344) );
  XNOR U8340 ( .A(y[62]), .B(x[62]), .Z(n8347) );
  XNOR U8341 ( .A(y[60]), .B(x[60]), .Z(n8346) );
  AND U8342 ( .A(n8348), .B(n8349), .Z(n8322) );
  AND U8343 ( .A(n8350), .B(n8351), .Z(n8349) );
  AND U8344 ( .A(n8352), .B(n8353), .Z(n8351) );
  XNOR U8345 ( .A(y[64]), .B(x[64]), .Z(n8353) );
  AND U8346 ( .A(n8354), .B(n8355), .Z(n8352) );
  XNOR U8347 ( .A(y[65]), .B(x[65]), .Z(n8355) );
  XNOR U8348 ( .A(y[63]), .B(x[63]), .Z(n8354) );
  AND U8349 ( .A(n8356), .B(n8357), .Z(n8350) );
  XNOR U8350 ( .A(y[67]), .B(x[67]), .Z(n8357) );
  AND U8351 ( .A(n8358), .B(n8359), .Z(n8356) );
  XNOR U8352 ( .A(y[68]), .B(x[68]), .Z(n8359) );
  XNOR U8353 ( .A(y[66]), .B(x[66]), .Z(n8358) );
  AND U8354 ( .A(n8360), .B(n8361), .Z(n8348) );
  AND U8355 ( .A(n8362), .B(n8363), .Z(n8361) );
  XNOR U8356 ( .A(y[70]), .B(x[70]), .Z(n8363) );
  AND U8357 ( .A(n8364), .B(n8365), .Z(n8362) );
  XNOR U8358 ( .A(y[71]), .B(x[71]), .Z(n8365) );
  XNOR U8359 ( .A(y[69]), .B(x[69]), .Z(n8364) );
  AND U8360 ( .A(n8366), .B(n8367), .Z(n8360) );
  XNOR U8361 ( .A(y[73]), .B(x[73]), .Z(n8367) );
  AND U8362 ( .A(n8368), .B(n8369), .Z(n8366) );
  XNOR U8363 ( .A(y[74]), .B(x[74]), .Z(n8369) );
  XNOR U8364 ( .A(y[72]), .B(x[72]), .Z(n8368) );
  AND U8365 ( .A(n8370), .B(n8371), .Z(n8320) );
  AND U8366 ( .A(n8372), .B(n8373), .Z(n8371) );
  AND U8367 ( .A(n8374), .B(n8375), .Z(n8373) );
  AND U8368 ( .A(n8376), .B(n8377), .Z(n8375) );
  AND U8369 ( .A(n8378), .B(n8379), .Z(n8377) );
  XNOR U8370 ( .A(y[75]), .B(x[75]), .Z(n8379) );
  XNOR U8371 ( .A(y[76]), .B(x[76]), .Z(n8378) );
  AND U8372 ( .A(n8380), .B(n8381), .Z(n8376) );
  XNOR U8373 ( .A(y[77]), .B(x[77]), .Z(n8381) );
  XNOR U8374 ( .A(y[78]), .B(x[78]), .Z(n8380) );
  AND U8375 ( .A(n8382), .B(n8383), .Z(n8374) );
  XNOR U8376 ( .A(y[80]), .B(x[80]), .Z(n8383) );
  AND U8377 ( .A(n8384), .B(n8385), .Z(n8382) );
  XNOR U8378 ( .A(y[81]), .B(x[81]), .Z(n8385) );
  XNOR U8379 ( .A(y[79]), .B(x[79]), .Z(n8384) );
  AND U8380 ( .A(n8386), .B(n8387), .Z(n8372) );
  AND U8381 ( .A(n8388), .B(n8389), .Z(n8387) );
  XNOR U8382 ( .A(y[83]), .B(x[83]), .Z(n8389) );
  AND U8383 ( .A(n8390), .B(n8391), .Z(n8388) );
  XNOR U8384 ( .A(y[84]), .B(x[84]), .Z(n8391) );
  XNOR U8385 ( .A(y[82]), .B(x[82]), .Z(n8390) );
  AND U8386 ( .A(n8392), .B(n8393), .Z(n8386) );
  XNOR U8387 ( .A(y[86]), .B(x[86]), .Z(n8393) );
  AND U8388 ( .A(n8394), .B(n8395), .Z(n8392) );
  XNOR U8389 ( .A(y[87]), .B(x[87]), .Z(n8395) );
  XNOR U8390 ( .A(y[85]), .B(x[85]), .Z(n8394) );
  AND U8391 ( .A(n8396), .B(n8397), .Z(n8370) );
  AND U8392 ( .A(n8398), .B(n8399), .Z(n8397) );
  AND U8393 ( .A(n8400), .B(n8401), .Z(n8399) );
  XNOR U8394 ( .A(y[89]), .B(x[89]), .Z(n8401) );
  AND U8395 ( .A(n8402), .B(n8403), .Z(n8400) );
  XNOR U8396 ( .A(y[90]), .B(x[90]), .Z(n8403) );
  XNOR U8397 ( .A(y[88]), .B(x[88]), .Z(n8402) );
  AND U8398 ( .A(n8404), .B(n8405), .Z(n8398) );
  XNOR U8399 ( .A(y[92]), .B(x[92]), .Z(n8405) );
  AND U8400 ( .A(n8406), .B(n8407), .Z(n8404) );
  XNOR U8401 ( .A(y[93]), .B(x[93]), .Z(n8407) );
  XNOR U8402 ( .A(y[91]), .B(x[91]), .Z(n8406) );
  AND U8403 ( .A(n8408), .B(n8409), .Z(n8396) );
  AND U8404 ( .A(n8410), .B(n8411), .Z(n8409) );
  XNOR U8405 ( .A(y[95]), .B(x[95]), .Z(n8411) );
  AND U8406 ( .A(n8412), .B(n8413), .Z(n8410) );
  XNOR U8407 ( .A(y[96]), .B(x[96]), .Z(n8413) );
  XNOR U8408 ( .A(y[94]), .B(x[94]), .Z(n8412) );
  AND U8409 ( .A(n8414), .B(n8415), .Z(n8408) );
  XNOR U8410 ( .A(y[98]), .B(x[98]), .Z(n8415) );
  AND U8411 ( .A(n8416), .B(n8417), .Z(n8414) );
  XNOR U8412 ( .A(y[99]), .B(x[99]), .Z(n8417) );
  XNOR U8413 ( .A(y[97]), .B(x[97]), .Z(n8416) );
  AND U8414 ( .A(n8418), .B(n8419), .Z(n8218) );
  AND U8415 ( .A(n8420), .B(n8421), .Z(n8419) );
  AND U8416 ( .A(n8422), .B(n8423), .Z(n8421) );
  AND U8417 ( .A(n8424), .B(n8425), .Z(n8423) );
  AND U8418 ( .A(n8426), .B(n8427), .Z(n8425) );
  AND U8419 ( .A(n8428), .B(n8429), .Z(n8427) );
  AND U8420 ( .A(n8430), .B(n8431), .Z(n8429) );
  XNOR U8421 ( .A(y[100]), .B(x[100]), .Z(n8431) );
  XNOR U8422 ( .A(y[101]), .B(x[101]), .Z(n8430) );
  AND U8423 ( .A(n8432), .B(n8433), .Z(n8428) );
  XNOR U8424 ( .A(y[102]), .B(x[102]), .Z(n8433) );
  XNOR U8425 ( .A(y[103]), .B(x[103]), .Z(n8432) );
  AND U8426 ( .A(n8434), .B(n8435), .Z(n8426) );
  XNOR U8427 ( .A(y[105]), .B(x[105]), .Z(n8435) );
  AND U8428 ( .A(n8436), .B(n8437), .Z(n8434) );
  XNOR U8429 ( .A(y[106]), .B(x[106]), .Z(n8437) );
  XNOR U8430 ( .A(y[104]), .B(x[104]), .Z(n8436) );
  AND U8431 ( .A(n8438), .B(n8439), .Z(n8424) );
  AND U8432 ( .A(n8440), .B(n8441), .Z(n8439) );
  XNOR U8433 ( .A(y[108]), .B(x[108]), .Z(n8441) );
  AND U8434 ( .A(n8442), .B(n8443), .Z(n8440) );
  XNOR U8435 ( .A(y[109]), .B(x[109]), .Z(n8443) );
  XNOR U8436 ( .A(y[107]), .B(x[107]), .Z(n8442) );
  AND U8437 ( .A(n8444), .B(n8445), .Z(n8438) );
  XNOR U8438 ( .A(y[111]), .B(x[111]), .Z(n8445) );
  AND U8439 ( .A(n8446), .B(n8447), .Z(n8444) );
  XNOR U8440 ( .A(y[112]), .B(x[112]), .Z(n8447) );
  XNOR U8441 ( .A(y[110]), .B(x[110]), .Z(n8446) );
  AND U8442 ( .A(n8448), .B(n8449), .Z(n8422) );
  AND U8443 ( .A(n8450), .B(n8451), .Z(n8449) );
  AND U8444 ( .A(n8452), .B(n8453), .Z(n8451) );
  XNOR U8445 ( .A(y[114]), .B(x[114]), .Z(n8453) );
  AND U8446 ( .A(n8454), .B(n8455), .Z(n8452) );
  XNOR U8447 ( .A(y[115]), .B(x[115]), .Z(n8455) );
  XNOR U8448 ( .A(y[113]), .B(x[113]), .Z(n8454) );
  AND U8449 ( .A(n8456), .B(n8457), .Z(n8450) );
  XNOR U8450 ( .A(y[117]), .B(x[117]), .Z(n8457) );
  AND U8451 ( .A(n8458), .B(n8459), .Z(n8456) );
  XNOR U8452 ( .A(y[118]), .B(x[118]), .Z(n8459) );
  XNOR U8453 ( .A(y[116]), .B(x[116]), .Z(n8458) );
  AND U8454 ( .A(n8460), .B(n8461), .Z(n8448) );
  AND U8455 ( .A(n8462), .B(n8463), .Z(n8461) );
  XNOR U8456 ( .A(y[120]), .B(x[120]), .Z(n8463) );
  AND U8457 ( .A(n8464), .B(n8465), .Z(n8462) );
  XNOR U8458 ( .A(y[121]), .B(x[121]), .Z(n8465) );
  XNOR U8459 ( .A(y[119]), .B(x[119]), .Z(n8464) );
  AND U8460 ( .A(n8466), .B(n8467), .Z(n8460) );
  XNOR U8461 ( .A(y[123]), .B(x[123]), .Z(n8467) );
  AND U8462 ( .A(n8468), .B(n8469), .Z(n8466) );
  XNOR U8463 ( .A(y[124]), .B(x[124]), .Z(n8469) );
  XNOR U8464 ( .A(y[122]), .B(x[122]), .Z(n8468) );
  AND U8465 ( .A(n8470), .B(n8471), .Z(n8420) );
  AND U8466 ( .A(n8472), .B(n8473), .Z(n8471) );
  AND U8467 ( .A(n8474), .B(n8475), .Z(n8473) );
  AND U8468 ( .A(n8476), .B(n8477), .Z(n8475) );
  AND U8469 ( .A(n8478), .B(n8479), .Z(n8477) );
  XNOR U8470 ( .A(y[125]), .B(x[125]), .Z(n8479) );
  XNOR U8471 ( .A(y[126]), .B(x[126]), .Z(n8478) );
  AND U8472 ( .A(n8480), .B(n8481), .Z(n8476) );
  XNOR U8473 ( .A(y[127]), .B(x[127]), .Z(n8481) );
  XNOR U8474 ( .A(y[128]), .B(x[128]), .Z(n8480) );
  AND U8475 ( .A(n8482), .B(n8483), .Z(n8474) );
  XNOR U8476 ( .A(y[130]), .B(x[130]), .Z(n8483) );
  AND U8477 ( .A(n8484), .B(n8485), .Z(n8482) );
  XNOR U8478 ( .A(y[131]), .B(x[131]), .Z(n8485) );
  XNOR U8479 ( .A(y[129]), .B(x[129]), .Z(n8484) );
  AND U8480 ( .A(n8486), .B(n8487), .Z(n8472) );
  AND U8481 ( .A(n8488), .B(n8489), .Z(n8487) );
  XNOR U8482 ( .A(y[133]), .B(x[133]), .Z(n8489) );
  AND U8483 ( .A(n8490), .B(n8491), .Z(n8488) );
  XNOR U8484 ( .A(y[134]), .B(x[134]), .Z(n8491) );
  XNOR U8485 ( .A(y[132]), .B(x[132]), .Z(n8490) );
  AND U8486 ( .A(n8492), .B(n8493), .Z(n8486) );
  XNOR U8487 ( .A(y[136]), .B(x[136]), .Z(n8493) );
  AND U8488 ( .A(n8494), .B(n8495), .Z(n8492) );
  XNOR U8489 ( .A(y[137]), .B(x[137]), .Z(n8495) );
  XNOR U8490 ( .A(y[135]), .B(x[135]), .Z(n8494) );
  AND U8491 ( .A(n8496), .B(n8497), .Z(n8470) );
  AND U8492 ( .A(n8498), .B(n8499), .Z(n8497) );
  AND U8493 ( .A(n8500), .B(n8501), .Z(n8499) );
  XNOR U8494 ( .A(y[139]), .B(x[139]), .Z(n8501) );
  AND U8495 ( .A(n8502), .B(n8503), .Z(n8500) );
  XNOR U8496 ( .A(y[140]), .B(x[140]), .Z(n8503) );
  XNOR U8497 ( .A(y[138]), .B(x[138]), .Z(n8502) );
  AND U8498 ( .A(n8504), .B(n8505), .Z(n8498) );
  XNOR U8499 ( .A(y[142]), .B(x[142]), .Z(n8505) );
  AND U8500 ( .A(n8506), .B(n8507), .Z(n8504) );
  XNOR U8501 ( .A(y[143]), .B(x[143]), .Z(n8507) );
  XNOR U8502 ( .A(y[141]), .B(x[141]), .Z(n8506) );
  AND U8503 ( .A(n8508), .B(n8509), .Z(n8496) );
  AND U8504 ( .A(n8510), .B(n8511), .Z(n8509) );
  XNOR U8505 ( .A(y[145]), .B(x[145]), .Z(n8511) );
  AND U8506 ( .A(n8512), .B(n8513), .Z(n8510) );
  XNOR U8507 ( .A(y[146]), .B(x[146]), .Z(n8513) );
  XNOR U8508 ( .A(y[144]), .B(x[144]), .Z(n8512) );
  AND U8509 ( .A(n8514), .B(n8515), .Z(n8508) );
  XNOR U8510 ( .A(y[148]), .B(x[148]), .Z(n8515) );
  AND U8511 ( .A(n8516), .B(n8517), .Z(n8514) );
  XNOR U8512 ( .A(y[149]), .B(x[149]), .Z(n8517) );
  XNOR U8513 ( .A(y[147]), .B(x[147]), .Z(n8516) );
  AND U8514 ( .A(n8518), .B(n8519), .Z(n8418) );
  AND U8515 ( .A(n8520), .B(n8521), .Z(n8519) );
  AND U8516 ( .A(n8522), .B(n8523), .Z(n8521) );
  AND U8517 ( .A(n8524), .B(n8525), .Z(n8523) );
  AND U8518 ( .A(n8526), .B(n8527), .Z(n8525) );
  AND U8519 ( .A(n8528), .B(n8529), .Z(n8527) );
  XNOR U8520 ( .A(y[150]), .B(x[150]), .Z(n8529) );
  XNOR U8521 ( .A(y[151]), .B(x[151]), .Z(n8528) );
  AND U8522 ( .A(n8530), .B(n8531), .Z(n8526) );
  XNOR U8523 ( .A(y[152]), .B(x[152]), .Z(n8531) );
  XNOR U8524 ( .A(y[153]), .B(x[153]), .Z(n8530) );
  AND U8525 ( .A(n8532), .B(n8533), .Z(n8524) );
  XNOR U8526 ( .A(y[155]), .B(x[155]), .Z(n8533) );
  AND U8527 ( .A(n8534), .B(n8535), .Z(n8532) );
  XNOR U8528 ( .A(y[156]), .B(x[156]), .Z(n8535) );
  XNOR U8529 ( .A(y[154]), .B(x[154]), .Z(n8534) );
  AND U8530 ( .A(n8536), .B(n8537), .Z(n8522) );
  AND U8531 ( .A(n8538), .B(n8539), .Z(n8537) );
  XNOR U8532 ( .A(y[158]), .B(x[158]), .Z(n8539) );
  AND U8533 ( .A(n8540), .B(n8541), .Z(n8538) );
  XNOR U8534 ( .A(y[159]), .B(x[159]), .Z(n8541) );
  XNOR U8535 ( .A(y[157]), .B(x[157]), .Z(n8540) );
  AND U8536 ( .A(n8542), .B(n8543), .Z(n8536) );
  XNOR U8537 ( .A(y[161]), .B(x[161]), .Z(n8543) );
  AND U8538 ( .A(n8544), .B(n8545), .Z(n8542) );
  XNOR U8539 ( .A(y[162]), .B(x[162]), .Z(n8545) );
  XNOR U8540 ( .A(y[160]), .B(x[160]), .Z(n8544) );
  AND U8541 ( .A(n8546), .B(n8547), .Z(n8520) );
  AND U8542 ( .A(n8548), .B(n8549), .Z(n8547) );
  AND U8543 ( .A(n8550), .B(n8551), .Z(n8549) );
  XNOR U8544 ( .A(y[164]), .B(x[164]), .Z(n8551) );
  AND U8545 ( .A(n8552), .B(n8553), .Z(n8550) );
  XNOR U8546 ( .A(y[165]), .B(x[165]), .Z(n8553) );
  XNOR U8547 ( .A(y[163]), .B(x[163]), .Z(n8552) );
  AND U8548 ( .A(n8554), .B(n8555), .Z(n8548) );
  XNOR U8549 ( .A(y[167]), .B(x[167]), .Z(n8555) );
  AND U8550 ( .A(n8556), .B(n8557), .Z(n8554) );
  XNOR U8551 ( .A(y[168]), .B(x[168]), .Z(n8557) );
  XNOR U8552 ( .A(y[166]), .B(x[166]), .Z(n8556) );
  AND U8553 ( .A(n8558), .B(n8559), .Z(n8546) );
  AND U8554 ( .A(n8560), .B(n8561), .Z(n8559) );
  XNOR U8555 ( .A(y[170]), .B(x[170]), .Z(n8561) );
  AND U8556 ( .A(n8562), .B(n8563), .Z(n8560) );
  XNOR U8557 ( .A(y[171]), .B(x[171]), .Z(n8563) );
  XNOR U8558 ( .A(y[169]), .B(x[169]), .Z(n8562) );
  AND U8559 ( .A(n8564), .B(n8565), .Z(n8558) );
  XNOR U8560 ( .A(y[173]), .B(x[173]), .Z(n8565) );
  AND U8561 ( .A(n8566), .B(n8567), .Z(n8564) );
  XNOR U8562 ( .A(y[174]), .B(x[174]), .Z(n8567) );
  XNOR U8563 ( .A(y[172]), .B(x[172]), .Z(n8566) );
  AND U8564 ( .A(n8568), .B(n8569), .Z(n8518) );
  AND U8565 ( .A(n8570), .B(n8571), .Z(n8569) );
  AND U8566 ( .A(n8572), .B(n8573), .Z(n8571) );
  AND U8567 ( .A(n8574), .B(n8575), .Z(n8573) );
  AND U8568 ( .A(n8576), .B(n8577), .Z(n8575) );
  XNOR U8569 ( .A(y[175]), .B(x[175]), .Z(n8577) );
  XNOR U8570 ( .A(y[176]), .B(x[176]), .Z(n8576) );
  AND U8571 ( .A(n8578), .B(n8579), .Z(n8574) );
  XNOR U8572 ( .A(y[177]), .B(x[177]), .Z(n8579) );
  XNOR U8573 ( .A(y[178]), .B(x[178]), .Z(n8578) );
  AND U8574 ( .A(n8580), .B(n8581), .Z(n8572) );
  XNOR U8575 ( .A(y[180]), .B(x[180]), .Z(n8581) );
  AND U8576 ( .A(n8582), .B(n8583), .Z(n8580) );
  XNOR U8577 ( .A(y[181]), .B(x[181]), .Z(n8583) );
  XNOR U8578 ( .A(y[179]), .B(x[179]), .Z(n8582) );
  AND U8579 ( .A(n8584), .B(n8585), .Z(n8570) );
  AND U8580 ( .A(n8586), .B(n8587), .Z(n8585) );
  XNOR U8581 ( .A(y[183]), .B(x[183]), .Z(n8587) );
  AND U8582 ( .A(n8588), .B(n8589), .Z(n8586) );
  XNOR U8583 ( .A(y[184]), .B(x[184]), .Z(n8589) );
  XNOR U8584 ( .A(y[182]), .B(x[182]), .Z(n8588) );
  AND U8585 ( .A(n8590), .B(n8591), .Z(n8584) );
  XNOR U8586 ( .A(y[186]), .B(x[186]), .Z(n8591) );
  AND U8587 ( .A(n8592), .B(n8593), .Z(n8590) );
  XNOR U8588 ( .A(y[187]), .B(x[187]), .Z(n8593) );
  XNOR U8589 ( .A(y[185]), .B(x[185]), .Z(n8592) );
  AND U8590 ( .A(n8594), .B(n8595), .Z(n8568) );
  AND U8591 ( .A(n8596), .B(n8597), .Z(n8595) );
  AND U8592 ( .A(n8598), .B(n8599), .Z(n8597) );
  XNOR U8593 ( .A(y[189]), .B(x[189]), .Z(n8599) );
  AND U8594 ( .A(n8600), .B(n8601), .Z(n8598) );
  XNOR U8595 ( .A(y[190]), .B(x[190]), .Z(n8601) );
  XNOR U8596 ( .A(y[188]), .B(x[188]), .Z(n8600) );
  AND U8597 ( .A(n8602), .B(n8603), .Z(n8596) );
  XNOR U8598 ( .A(y[192]), .B(x[192]), .Z(n8603) );
  AND U8599 ( .A(n8604), .B(n8605), .Z(n8602) );
  XNOR U8600 ( .A(y[193]), .B(x[193]), .Z(n8605) );
  XNOR U8601 ( .A(y[191]), .B(x[191]), .Z(n8604) );
  AND U8602 ( .A(n8606), .B(n8607), .Z(n8594) );
  AND U8603 ( .A(n8608), .B(n8609), .Z(n8607) );
  XNOR U8604 ( .A(y[195]), .B(x[195]), .Z(n8609) );
  AND U8605 ( .A(n8610), .B(n8611), .Z(n8608) );
  XNOR U8606 ( .A(y[196]), .B(x[196]), .Z(n8611) );
  XNOR U8607 ( .A(y[194]), .B(x[194]), .Z(n8610) );
  AND U8608 ( .A(n8612), .B(n8613), .Z(n8606) );
  XNOR U8609 ( .A(y[198]), .B(x[198]), .Z(n8613) );
  AND U8610 ( .A(n8614), .B(n8615), .Z(n8612) );
  XNOR U8611 ( .A(y[199]), .B(x[199]), .Z(n8615) );
  XNOR U8612 ( .A(y[197]), .B(x[197]), .Z(n8614) );
  AND U8613 ( .A(n8616), .B(n8617), .Z(n8216) );
  AND U8614 ( .A(n8618), .B(n8619), .Z(n8617) );
  AND U8615 ( .A(n8620), .B(n8621), .Z(n8619) );
  AND U8616 ( .A(n8622), .B(n8623), .Z(n8621) );
  AND U8617 ( .A(n8624), .B(n8625), .Z(n8623) );
  AND U8618 ( .A(n8626), .B(n8627), .Z(n8625) );
  AND U8619 ( .A(n8628), .B(n8629), .Z(n8627) );
  AND U8620 ( .A(n8630), .B(n8631), .Z(n8629) );
  XNOR U8621 ( .A(y[942]), .B(x[942]), .Z(n8631) );
  AND U8622 ( .A(n8632), .B(n8633), .Z(n8630) );
  AND U8623 ( .A(n8634), .B(n8635), .Z(n8633) );
  AND U8624 ( .A(n8636), .B(n8637), .Z(n8635) );
  AND U8625 ( .A(n8638), .B(n8639), .Z(n8637) );
  AND U8626 ( .A(n8640), .B(n8641), .Z(n8639) );
  AND U8627 ( .A(n8642), .B(n8643), .Z(n8641) );
  AND U8628 ( .A(n8644), .B(n8645), .Z(n8643) );
  AND U8629 ( .A(n8646), .B(n8647), .Z(n8645) );
  AND U8630 ( .A(n8648), .B(n8649), .Z(n8647) );
  XNOR U8631 ( .A(y[1500]), .B(x[1500]), .Z(n8649) );
  AND U8632 ( .A(n8650), .B(n8651), .Z(n8648) );
  AND U8633 ( .A(n8652), .B(n8653), .Z(n8651) );
  AND U8634 ( .A(n8654), .B(n8655), .Z(n8653) );
  AND U8635 ( .A(n8656), .B(n8657), .Z(n8655) );
  AND U8636 ( .A(n8658), .B(n8659), .Z(n8657) );
  AND U8637 ( .A(n8660), .B(n8661), .Z(n8659) );
  AND U8638 ( .A(n8662), .B(n8663), .Z(n8661) );
  AND U8639 ( .A(n8664), .B(n8665), .Z(n8663) );
  AND U8640 ( .A(n8666), .B(n8667), .Z(n8665) );
  AND U8641 ( .A(n8668), .B(n8669), .Z(n8667) );
  AND U8642 ( .A(n8670), .B(n8671), .Z(n8669) );
  AND U8643 ( .A(n8672), .B(n8673), .Z(n8671) );
  AND U8644 ( .A(n8674), .B(n8675), .Z(n8673) );
  AND U8645 ( .A(n8676), .B(n8677), .Z(n8675) );
  AND U8646 ( .A(n8678), .B(n8679), .Z(n8677) );
  AND U8647 ( .A(n8680), .B(n8681), .Z(n8679) );
  AND U8648 ( .A(n8682), .B(n8683), .Z(n8681) );
  AND U8649 ( .A(n8684), .B(n8685), .Z(n8683) );
  XNOR U8650 ( .A(y[2048]), .B(x[2048]), .Z(n8685) );
  XNOR U8651 ( .A(y[2049]), .B(x[2049]), .Z(n8684) );
  AND U8652 ( .A(n8686), .B(n8687), .Z(n8682) );
  XNOR U8653 ( .A(y[2050]), .B(x[2050]), .Z(n8687) );
  XNOR U8654 ( .A(y[2051]), .B(x[2051]), .Z(n8686) );
  AND U8655 ( .A(n8688), .B(n8689), .Z(n8680) );
  AND U8656 ( .A(n8690), .B(n8691), .Z(n8689) );
  XNOR U8657 ( .A(y[2052]), .B(x[2052]), .Z(n8691) );
  XNOR U8658 ( .A(y[2053]), .B(x[2053]), .Z(n8690) );
  AND U8659 ( .A(n8692), .B(n8693), .Z(n8688) );
  XNOR U8660 ( .A(y[2054]), .B(x[2054]), .Z(n8693) );
  XNOR U8661 ( .A(y[2057]), .B(x[2057]), .Z(n8692) );
  AND U8662 ( .A(n8694), .B(n8695), .Z(n8678) );
  AND U8663 ( .A(n8696), .B(n8697), .Z(n8695) );
  AND U8664 ( .A(n8698), .B(n8699), .Z(n8697) );
  XNOR U8665 ( .A(y[2055]), .B(x[2055]), .Z(n8699) );
  XNOR U8666 ( .A(y[2056]), .B(x[2056]), .Z(n8698) );
  AND U8667 ( .A(n8700), .B(n8701), .Z(n8696) );
  XNOR U8668 ( .A(y[2058]), .B(x[2058]), .Z(n8701) );
  XNOR U8669 ( .A(y[2059]), .B(x[2059]), .Z(n8700) );
  AND U8670 ( .A(n8702), .B(n8703), .Z(n8694) );
  AND U8671 ( .A(n8704), .B(n8705), .Z(n8703) );
  XNOR U8672 ( .A(y[2060]), .B(x[2060]), .Z(n8705) );
  XNOR U8673 ( .A(y[2061]), .B(x[2061]), .Z(n8704) );
  AND U8674 ( .A(n8706), .B(n8707), .Z(n8702) );
  XNOR U8675 ( .A(y[2062]), .B(x[2062]), .Z(n8707) );
  XNOR U8676 ( .A(y[2063]), .B(x[2063]), .Z(n8706) );
  AND U8677 ( .A(n8708), .B(n8709), .Z(n8676) );
  AND U8678 ( .A(n8710), .B(n8711), .Z(n8709) );
  AND U8679 ( .A(n8712), .B(n8713), .Z(n8711) );
  AND U8680 ( .A(n8714), .B(n8715), .Z(n8713) );
  XNOR U8681 ( .A(y[2064]), .B(x[2064]), .Z(n8715) );
  XNOR U8682 ( .A(y[2065]), .B(x[2065]), .Z(n8714) );
  AND U8683 ( .A(n8716), .B(n8717), .Z(n8712) );
  XNOR U8684 ( .A(y[2066]), .B(x[2066]), .Z(n8717) );
  XNOR U8685 ( .A(y[2067]), .B(x[2067]), .Z(n8716) );
  AND U8686 ( .A(n8718), .B(n8719), .Z(n8710) );
  AND U8687 ( .A(n8720), .B(n8721), .Z(n8719) );
  XNOR U8688 ( .A(y[2068]), .B(x[2068]), .Z(n8721) );
  XNOR U8689 ( .A(y[2069]), .B(x[2069]), .Z(n8720) );
  AND U8690 ( .A(n8722), .B(n8723), .Z(n8718) );
  XNOR U8691 ( .A(y[2070]), .B(x[2070]), .Z(n8723) );
  XNOR U8692 ( .A(y[2071]), .B(x[2071]), .Z(n8722) );
  AND U8693 ( .A(n8724), .B(n8725), .Z(n8708) );
  AND U8694 ( .A(n8726), .B(n8727), .Z(n8725) );
  AND U8695 ( .A(n8728), .B(n8729), .Z(n8727) );
  XNOR U8696 ( .A(y[2072]), .B(x[2072]), .Z(n8729) );
  XNOR U8697 ( .A(y[2073]), .B(x[2073]), .Z(n8728) );
  AND U8698 ( .A(n8730), .B(n8731), .Z(n8726) );
  XNOR U8699 ( .A(y[2074]), .B(x[2074]), .Z(n8731) );
  XNOR U8700 ( .A(y[2075]), .B(x[2075]), .Z(n8730) );
  AND U8701 ( .A(n8732), .B(n8733), .Z(n8724) );
  AND U8702 ( .A(n8734), .B(n8735), .Z(n8733) );
  XNOR U8703 ( .A(y[2076]), .B(x[2076]), .Z(n8735) );
  XNOR U8704 ( .A(y[2077]), .B(x[2077]), .Z(n8734) );
  AND U8705 ( .A(n8736), .B(n8737), .Z(n8732) );
  XNOR U8706 ( .A(y[2078]), .B(x[2078]), .Z(n8737) );
  XNOR U8707 ( .A(y[2079]), .B(x[2079]), .Z(n8736) );
  AND U8708 ( .A(n8738), .B(n8739), .Z(n8674) );
  AND U8709 ( .A(n8740), .B(n8741), .Z(n8739) );
  AND U8710 ( .A(n8742), .B(n8743), .Z(n8741) );
  AND U8711 ( .A(n8744), .B(n8745), .Z(n8743) );
  AND U8712 ( .A(n8746), .B(n8747), .Z(n8745) );
  XNOR U8713 ( .A(y[2080]), .B(x[2080]), .Z(n8747) );
  XNOR U8714 ( .A(y[2081]), .B(x[2081]), .Z(n8746) );
  AND U8715 ( .A(n8748), .B(n8749), .Z(n8744) );
  XNOR U8716 ( .A(y[2082]), .B(x[2082]), .Z(n8749) );
  XNOR U8717 ( .A(y[2083]), .B(x[2083]), .Z(n8748) );
  AND U8718 ( .A(n8750), .B(n8751), .Z(n8742) );
  AND U8719 ( .A(n8752), .B(n8753), .Z(n8751) );
  XNOR U8720 ( .A(y[2084]), .B(x[2084]), .Z(n8753) );
  XNOR U8721 ( .A(y[2085]), .B(x[2085]), .Z(n8752) );
  AND U8722 ( .A(n8754), .B(n8755), .Z(n8750) );
  XNOR U8723 ( .A(y[2086]), .B(x[2086]), .Z(n8755) );
  XNOR U8724 ( .A(y[2087]), .B(x[2087]), .Z(n8754) );
  AND U8725 ( .A(n8756), .B(n8757), .Z(n8740) );
  AND U8726 ( .A(n8758), .B(n8759), .Z(n8757) );
  AND U8727 ( .A(n8760), .B(n8761), .Z(n8759) );
  XNOR U8728 ( .A(y[2088]), .B(x[2088]), .Z(n8761) );
  XNOR U8729 ( .A(y[2089]), .B(x[2089]), .Z(n8760) );
  AND U8730 ( .A(n8762), .B(n8763), .Z(n8758) );
  XNOR U8731 ( .A(y[2090]), .B(x[2090]), .Z(n8763) );
  XNOR U8732 ( .A(y[2091]), .B(x[2091]), .Z(n8762) );
  AND U8733 ( .A(n8764), .B(n8765), .Z(n8756) );
  AND U8734 ( .A(n8766), .B(n8767), .Z(n8765) );
  XNOR U8735 ( .A(y[2092]), .B(x[2092]), .Z(n8767) );
  XNOR U8736 ( .A(y[2093]), .B(x[2093]), .Z(n8766) );
  AND U8737 ( .A(n8768), .B(n8769), .Z(n8764) );
  XNOR U8738 ( .A(y[2094]), .B(x[2094]), .Z(n8769) );
  XNOR U8739 ( .A(y[2095]), .B(x[2095]), .Z(n8768) );
  AND U8740 ( .A(n8770), .B(n8771), .Z(n8738) );
  AND U8741 ( .A(n8772), .B(n8773), .Z(n8771) );
  AND U8742 ( .A(n8774), .B(n8775), .Z(n8773) );
  AND U8743 ( .A(n8776), .B(n8777), .Z(n8775) );
  XNOR U8744 ( .A(y[2096]), .B(x[2096]), .Z(n8777) );
  XNOR U8745 ( .A(y[2097]), .B(x[2097]), .Z(n8776) );
  AND U8746 ( .A(n8778), .B(n8779), .Z(n8774) );
  XNOR U8747 ( .A(y[2098]), .B(x[2098]), .Z(n8779) );
  XNOR U8748 ( .A(y[2099]), .B(x[2099]), .Z(n8778) );
  AND U8749 ( .A(n8780), .B(n8781), .Z(n8772) );
  AND U8750 ( .A(n8782), .B(n8783), .Z(n8781) );
  XNOR U8751 ( .A(y[2100]), .B(x[2100]), .Z(n8783) );
  XNOR U8752 ( .A(y[2101]), .B(x[2101]), .Z(n8782) );
  AND U8753 ( .A(n8784), .B(n8785), .Z(n8780) );
  XNOR U8754 ( .A(y[2102]), .B(x[2102]), .Z(n8785) );
  XNOR U8755 ( .A(y[2103]), .B(x[2103]), .Z(n8784) );
  AND U8756 ( .A(n8786), .B(n8787), .Z(n8770) );
  AND U8757 ( .A(n8788), .B(n8789), .Z(n8787) );
  AND U8758 ( .A(n8790), .B(n8791), .Z(n8789) );
  XNOR U8759 ( .A(y[2104]), .B(x[2104]), .Z(n8791) );
  XNOR U8760 ( .A(y[2105]), .B(x[2105]), .Z(n8790) );
  AND U8761 ( .A(n8792), .B(n8793), .Z(n8788) );
  XNOR U8762 ( .A(y[2106]), .B(x[2106]), .Z(n8793) );
  XNOR U8763 ( .A(y[2107]), .B(x[2107]), .Z(n8792) );
  AND U8764 ( .A(n8794), .B(n8795), .Z(n8786) );
  AND U8765 ( .A(n8796), .B(n8797), .Z(n8795) );
  XNOR U8766 ( .A(y[2108]), .B(x[2108]), .Z(n8797) );
  XNOR U8767 ( .A(y[2109]), .B(x[2109]), .Z(n8796) );
  AND U8768 ( .A(n8798), .B(n8799), .Z(n8794) );
  XNOR U8769 ( .A(y[2110]), .B(x[2110]), .Z(n8799) );
  XNOR U8770 ( .A(y[2111]), .B(x[2111]), .Z(n8798) );
  AND U8771 ( .A(n8800), .B(n8801), .Z(n8672) );
  AND U8772 ( .A(n8802), .B(n8803), .Z(n8801) );
  AND U8773 ( .A(n8804), .B(n8805), .Z(n8803) );
  AND U8774 ( .A(n8806), .B(n8807), .Z(n8805) );
  AND U8775 ( .A(n8808), .B(n8809), .Z(n8807) );
  AND U8776 ( .A(n8810), .B(n8811), .Z(n8809) );
  XNOR U8777 ( .A(y[2112]), .B(x[2112]), .Z(n8811) );
  XNOR U8778 ( .A(y[2113]), .B(x[2113]), .Z(n8810) );
  AND U8779 ( .A(n8812), .B(n8813), .Z(n8808) );
  XNOR U8780 ( .A(y[2114]), .B(x[2114]), .Z(n8813) );
  XNOR U8781 ( .A(y[2115]), .B(x[2115]), .Z(n8812) );
  AND U8782 ( .A(n8814), .B(n8815), .Z(n8806) );
  AND U8783 ( .A(n8816), .B(n8817), .Z(n8815) );
  XNOR U8784 ( .A(y[2116]), .B(x[2116]), .Z(n8817) );
  XNOR U8785 ( .A(y[2117]), .B(x[2117]), .Z(n8816) );
  AND U8786 ( .A(n8818), .B(n8819), .Z(n8814) );
  XNOR U8787 ( .A(y[2118]), .B(x[2118]), .Z(n8819) );
  XNOR U8788 ( .A(y[2119]), .B(x[2119]), .Z(n8818) );
  AND U8789 ( .A(n8820), .B(n8821), .Z(n8804) );
  AND U8790 ( .A(n8822), .B(n8823), .Z(n8821) );
  AND U8791 ( .A(n8824), .B(n8825), .Z(n8823) );
  XNOR U8792 ( .A(y[2120]), .B(x[2120]), .Z(n8825) );
  XNOR U8793 ( .A(y[2121]), .B(x[2121]), .Z(n8824) );
  AND U8794 ( .A(n8826), .B(n8827), .Z(n8822) );
  XNOR U8795 ( .A(y[2122]), .B(x[2122]), .Z(n8827) );
  XNOR U8796 ( .A(y[2123]), .B(x[2123]), .Z(n8826) );
  AND U8797 ( .A(n8828), .B(n8829), .Z(n8820) );
  AND U8798 ( .A(n8830), .B(n8831), .Z(n8829) );
  XNOR U8799 ( .A(y[2124]), .B(x[2124]), .Z(n8831) );
  XNOR U8800 ( .A(y[2125]), .B(x[2125]), .Z(n8830) );
  AND U8801 ( .A(n8832), .B(n8833), .Z(n8828) );
  XNOR U8802 ( .A(y[2126]), .B(x[2126]), .Z(n8833) );
  XNOR U8803 ( .A(y[2127]), .B(x[2127]), .Z(n8832) );
  AND U8804 ( .A(n8834), .B(n8835), .Z(n8802) );
  AND U8805 ( .A(n8836), .B(n8837), .Z(n8835) );
  AND U8806 ( .A(n8838), .B(n8839), .Z(n8837) );
  AND U8807 ( .A(n8840), .B(n8841), .Z(n8839) );
  XNOR U8808 ( .A(y[2128]), .B(x[2128]), .Z(n8841) );
  XNOR U8809 ( .A(y[2129]), .B(x[2129]), .Z(n8840) );
  AND U8810 ( .A(n8842), .B(n8843), .Z(n8838) );
  XNOR U8811 ( .A(y[2130]), .B(x[2130]), .Z(n8843) );
  XNOR U8812 ( .A(y[2131]), .B(x[2131]), .Z(n8842) );
  AND U8813 ( .A(n8844), .B(n8845), .Z(n8836) );
  AND U8814 ( .A(n8846), .B(n8847), .Z(n8845) );
  XNOR U8815 ( .A(y[2132]), .B(x[2132]), .Z(n8847) );
  XNOR U8816 ( .A(y[2133]), .B(x[2133]), .Z(n8846) );
  AND U8817 ( .A(n8848), .B(n8849), .Z(n8844) );
  XNOR U8818 ( .A(y[2134]), .B(x[2134]), .Z(n8849) );
  XNOR U8819 ( .A(y[2135]), .B(x[2135]), .Z(n8848) );
  AND U8820 ( .A(n8850), .B(n8851), .Z(n8834) );
  AND U8821 ( .A(n8852), .B(n8853), .Z(n8851) );
  AND U8822 ( .A(n8854), .B(n8855), .Z(n8853) );
  XNOR U8823 ( .A(y[2136]), .B(x[2136]), .Z(n8855) );
  XNOR U8824 ( .A(y[2137]), .B(x[2137]), .Z(n8854) );
  AND U8825 ( .A(n8856), .B(n8857), .Z(n8852) );
  XNOR U8826 ( .A(y[2138]), .B(x[2138]), .Z(n8857) );
  XNOR U8827 ( .A(y[2139]), .B(x[2139]), .Z(n8856) );
  AND U8828 ( .A(n8858), .B(n8859), .Z(n8850) );
  AND U8829 ( .A(n8860), .B(n8861), .Z(n8859) );
  XNOR U8830 ( .A(y[2140]), .B(x[2140]), .Z(n8861) );
  XNOR U8831 ( .A(y[2141]), .B(x[2141]), .Z(n8860) );
  AND U8832 ( .A(n8862), .B(n8863), .Z(n8858) );
  XNOR U8833 ( .A(y[2142]), .B(x[2142]), .Z(n8863) );
  XNOR U8834 ( .A(y[2143]), .B(x[2143]), .Z(n8862) );
  AND U8835 ( .A(n8864), .B(n8865), .Z(n8800) );
  AND U8836 ( .A(n8866), .B(n8867), .Z(n8865) );
  AND U8837 ( .A(n8868), .B(n8869), .Z(n8867) );
  AND U8838 ( .A(n8870), .B(n8871), .Z(n8869) );
  AND U8839 ( .A(n8872), .B(n8873), .Z(n8871) );
  XNOR U8840 ( .A(y[2144]), .B(x[2144]), .Z(n8873) );
  XNOR U8841 ( .A(y[2145]), .B(x[2145]), .Z(n8872) );
  AND U8842 ( .A(n8874), .B(n8875), .Z(n8870) );
  XNOR U8843 ( .A(y[2146]), .B(x[2146]), .Z(n8875) );
  XNOR U8844 ( .A(y[2147]), .B(x[2147]), .Z(n8874) );
  AND U8845 ( .A(n8876), .B(n8877), .Z(n8868) );
  AND U8846 ( .A(n8878), .B(n8879), .Z(n8877) );
  XNOR U8847 ( .A(y[2148]), .B(x[2148]), .Z(n8879) );
  XNOR U8848 ( .A(y[2149]), .B(x[2149]), .Z(n8878) );
  AND U8849 ( .A(n8880), .B(n8881), .Z(n8876) );
  XNOR U8850 ( .A(y[2150]), .B(x[2150]), .Z(n8881) );
  XNOR U8851 ( .A(y[2151]), .B(x[2151]), .Z(n8880) );
  AND U8852 ( .A(n8882), .B(n8883), .Z(n8866) );
  AND U8853 ( .A(n8884), .B(n8885), .Z(n8883) );
  AND U8854 ( .A(n8886), .B(n8887), .Z(n8885) );
  XNOR U8855 ( .A(y[2152]), .B(x[2152]), .Z(n8887) );
  XNOR U8856 ( .A(y[2153]), .B(x[2153]), .Z(n8886) );
  AND U8857 ( .A(n8888), .B(n8889), .Z(n8884) );
  XNOR U8858 ( .A(y[2154]), .B(x[2154]), .Z(n8889) );
  XNOR U8859 ( .A(y[2155]), .B(x[2155]), .Z(n8888) );
  AND U8860 ( .A(n8890), .B(n8891), .Z(n8882) );
  AND U8861 ( .A(n8892), .B(n8893), .Z(n8891) );
  XNOR U8862 ( .A(y[2156]), .B(x[2156]), .Z(n8893) );
  XNOR U8863 ( .A(y[2157]), .B(x[2157]), .Z(n8892) );
  AND U8864 ( .A(n8894), .B(n8895), .Z(n8890) );
  XNOR U8865 ( .A(y[2158]), .B(x[2158]), .Z(n8895) );
  XNOR U8866 ( .A(y[2159]), .B(x[2159]), .Z(n8894) );
  AND U8867 ( .A(n8896), .B(n8897), .Z(n8864) );
  AND U8868 ( .A(n8898), .B(n8899), .Z(n8897) );
  AND U8869 ( .A(n8900), .B(n8901), .Z(n8899) );
  AND U8870 ( .A(n8902), .B(n8903), .Z(n8901) );
  XNOR U8871 ( .A(y[2160]), .B(x[2160]), .Z(n8903) );
  XNOR U8872 ( .A(y[2161]), .B(x[2161]), .Z(n8902) );
  AND U8873 ( .A(n8904), .B(n8905), .Z(n8900) );
  XNOR U8874 ( .A(y[2162]), .B(x[2162]), .Z(n8905) );
  XNOR U8875 ( .A(y[2163]), .B(x[2163]), .Z(n8904) );
  AND U8876 ( .A(n8906), .B(n8907), .Z(n8898) );
  AND U8877 ( .A(n8908), .B(n8909), .Z(n8907) );
  XNOR U8878 ( .A(y[2164]), .B(x[2164]), .Z(n8909) );
  XNOR U8879 ( .A(y[2165]), .B(x[2165]), .Z(n8908) );
  AND U8880 ( .A(n8910), .B(n8911), .Z(n8906) );
  XNOR U8881 ( .A(y[2166]), .B(x[2166]), .Z(n8911) );
  XNOR U8882 ( .A(y[2167]), .B(x[2167]), .Z(n8910) );
  AND U8883 ( .A(n8912), .B(n8913), .Z(n8896) );
  AND U8884 ( .A(n8914), .B(n8915), .Z(n8913) );
  AND U8885 ( .A(n8916), .B(n8917), .Z(n8915) );
  XNOR U8886 ( .A(y[2168]), .B(x[2168]), .Z(n8917) );
  XNOR U8887 ( .A(y[2169]), .B(x[2169]), .Z(n8916) );
  AND U8888 ( .A(n8918), .B(n8919), .Z(n8914) );
  XNOR U8889 ( .A(y[2170]), .B(x[2170]), .Z(n8919) );
  XNOR U8890 ( .A(y[2171]), .B(x[2171]), .Z(n8918) );
  AND U8891 ( .A(n8920), .B(n8921), .Z(n8912) );
  AND U8892 ( .A(n8922), .B(n8923), .Z(n8921) );
  XNOR U8893 ( .A(y[2172]), .B(x[2172]), .Z(n8923) );
  XNOR U8894 ( .A(y[2173]), .B(x[2173]), .Z(n8922) );
  AND U8895 ( .A(n8924), .B(n8925), .Z(n8920) );
  XNOR U8896 ( .A(y[2174]), .B(x[2174]), .Z(n8925) );
  XNOR U8897 ( .A(y[2175]), .B(x[2175]), .Z(n8924) );
  AND U8898 ( .A(n8926), .B(n8927), .Z(n8670) );
  AND U8899 ( .A(n8928), .B(n8929), .Z(n8927) );
  AND U8900 ( .A(n8930), .B(n8931), .Z(n8929) );
  AND U8901 ( .A(n8932), .B(n8933), .Z(n8931) );
  AND U8902 ( .A(n8934), .B(n8935), .Z(n8933) );
  AND U8903 ( .A(n8936), .B(n8937), .Z(n8935) );
  AND U8904 ( .A(n8938), .B(n8939), .Z(n8937) );
  XNOR U8905 ( .A(y[2176]), .B(x[2176]), .Z(n8939) );
  XNOR U8906 ( .A(y[2177]), .B(x[2177]), .Z(n8938) );
  AND U8907 ( .A(n8940), .B(n8941), .Z(n8936) );
  XNOR U8908 ( .A(y[2178]), .B(x[2178]), .Z(n8941) );
  XNOR U8909 ( .A(y[2179]), .B(x[2179]), .Z(n8940) );
  AND U8910 ( .A(n8942), .B(n8943), .Z(n8934) );
  AND U8911 ( .A(n8944), .B(n8945), .Z(n8943) );
  XNOR U8912 ( .A(y[2180]), .B(x[2180]), .Z(n8945) );
  XNOR U8913 ( .A(y[2181]), .B(x[2181]), .Z(n8944) );
  AND U8914 ( .A(n8946), .B(n8947), .Z(n8942) );
  XNOR U8915 ( .A(y[2182]), .B(x[2182]), .Z(n8947) );
  XNOR U8916 ( .A(y[2183]), .B(x[2183]), .Z(n8946) );
  AND U8917 ( .A(n8948), .B(n8949), .Z(n8932) );
  AND U8918 ( .A(n8950), .B(n8951), .Z(n8949) );
  AND U8919 ( .A(n8952), .B(n8953), .Z(n8951) );
  XNOR U8920 ( .A(y[2184]), .B(x[2184]), .Z(n8953) );
  XNOR U8921 ( .A(y[2185]), .B(x[2185]), .Z(n8952) );
  AND U8922 ( .A(n8954), .B(n8955), .Z(n8950) );
  XNOR U8923 ( .A(y[2186]), .B(x[2186]), .Z(n8955) );
  XNOR U8924 ( .A(y[2187]), .B(x[2187]), .Z(n8954) );
  AND U8925 ( .A(n8956), .B(n8957), .Z(n8948) );
  AND U8926 ( .A(n8958), .B(n8959), .Z(n8957) );
  XNOR U8927 ( .A(y[2188]), .B(x[2188]), .Z(n8959) );
  XNOR U8928 ( .A(y[2189]), .B(x[2189]), .Z(n8958) );
  AND U8929 ( .A(n8960), .B(n8961), .Z(n8956) );
  XNOR U8930 ( .A(y[2190]), .B(x[2190]), .Z(n8961) );
  XNOR U8931 ( .A(y[2191]), .B(x[2191]), .Z(n8960) );
  AND U8932 ( .A(n8962), .B(n8963), .Z(n8930) );
  AND U8933 ( .A(n8964), .B(n8965), .Z(n8963) );
  AND U8934 ( .A(n8966), .B(n8967), .Z(n8965) );
  AND U8935 ( .A(n8968), .B(n8969), .Z(n8967) );
  XNOR U8936 ( .A(y[2192]), .B(x[2192]), .Z(n8969) );
  XNOR U8937 ( .A(y[2193]), .B(x[2193]), .Z(n8968) );
  AND U8938 ( .A(n8970), .B(n8971), .Z(n8966) );
  XNOR U8939 ( .A(y[2194]), .B(x[2194]), .Z(n8971) );
  XNOR U8940 ( .A(y[2195]), .B(x[2195]), .Z(n8970) );
  AND U8941 ( .A(n8972), .B(n8973), .Z(n8964) );
  AND U8942 ( .A(n8974), .B(n8975), .Z(n8973) );
  XNOR U8943 ( .A(y[2196]), .B(x[2196]), .Z(n8975) );
  XNOR U8944 ( .A(y[2197]), .B(x[2197]), .Z(n8974) );
  AND U8945 ( .A(n8976), .B(n8977), .Z(n8972) );
  XNOR U8946 ( .A(y[2198]), .B(x[2198]), .Z(n8977) );
  XNOR U8947 ( .A(y[2199]), .B(x[2199]), .Z(n8976) );
  AND U8948 ( .A(n8978), .B(n8979), .Z(n8962) );
  AND U8949 ( .A(n8980), .B(n8981), .Z(n8979) );
  AND U8950 ( .A(n8982), .B(n8983), .Z(n8981) );
  XNOR U8951 ( .A(y[2200]), .B(x[2200]), .Z(n8983) );
  XNOR U8952 ( .A(y[2201]), .B(x[2201]), .Z(n8982) );
  AND U8953 ( .A(n8984), .B(n8985), .Z(n8980) );
  XNOR U8954 ( .A(y[2202]), .B(x[2202]), .Z(n8985) );
  XNOR U8955 ( .A(y[2203]), .B(x[2203]), .Z(n8984) );
  AND U8956 ( .A(n8986), .B(n8987), .Z(n8978) );
  AND U8957 ( .A(n8988), .B(n8989), .Z(n8987) );
  XNOR U8958 ( .A(y[2204]), .B(x[2204]), .Z(n8989) );
  XNOR U8959 ( .A(y[2205]), .B(x[2205]), .Z(n8988) );
  AND U8960 ( .A(n8990), .B(n8991), .Z(n8986) );
  XNOR U8961 ( .A(y[2206]), .B(x[2206]), .Z(n8991) );
  XNOR U8962 ( .A(y[2207]), .B(x[2207]), .Z(n8990) );
  AND U8963 ( .A(n8992), .B(n8993), .Z(n8928) );
  AND U8964 ( .A(n8994), .B(n8995), .Z(n8993) );
  AND U8965 ( .A(n8996), .B(n8997), .Z(n8995) );
  AND U8966 ( .A(n8998), .B(n8999), .Z(n8997) );
  AND U8967 ( .A(n9000), .B(n9001), .Z(n8999) );
  XNOR U8968 ( .A(y[2208]), .B(x[2208]), .Z(n9001) );
  XNOR U8969 ( .A(y[2209]), .B(x[2209]), .Z(n9000) );
  AND U8970 ( .A(n9002), .B(n9003), .Z(n8998) );
  XNOR U8971 ( .A(y[2210]), .B(x[2210]), .Z(n9003) );
  XNOR U8972 ( .A(y[2211]), .B(x[2211]), .Z(n9002) );
  AND U8973 ( .A(n9004), .B(n9005), .Z(n8996) );
  AND U8974 ( .A(n9006), .B(n9007), .Z(n9005) );
  XNOR U8975 ( .A(y[2212]), .B(x[2212]), .Z(n9007) );
  XNOR U8976 ( .A(y[2213]), .B(x[2213]), .Z(n9006) );
  AND U8977 ( .A(n9008), .B(n9009), .Z(n9004) );
  XNOR U8978 ( .A(y[2214]), .B(x[2214]), .Z(n9009) );
  XNOR U8979 ( .A(y[2215]), .B(x[2215]), .Z(n9008) );
  AND U8980 ( .A(n9010), .B(n9011), .Z(n8994) );
  AND U8981 ( .A(n9012), .B(n9013), .Z(n9011) );
  AND U8982 ( .A(n9014), .B(n9015), .Z(n9013) );
  XNOR U8983 ( .A(y[2216]), .B(x[2216]), .Z(n9015) );
  XNOR U8984 ( .A(y[2217]), .B(x[2217]), .Z(n9014) );
  AND U8985 ( .A(n9016), .B(n9017), .Z(n9012) );
  XNOR U8986 ( .A(y[2218]), .B(x[2218]), .Z(n9017) );
  XNOR U8987 ( .A(y[2219]), .B(x[2219]), .Z(n9016) );
  AND U8988 ( .A(n9018), .B(n9019), .Z(n9010) );
  AND U8989 ( .A(n9020), .B(n9021), .Z(n9019) );
  XNOR U8990 ( .A(y[2220]), .B(x[2220]), .Z(n9021) );
  XNOR U8991 ( .A(y[2221]), .B(x[2221]), .Z(n9020) );
  AND U8992 ( .A(n9022), .B(n9023), .Z(n9018) );
  XNOR U8993 ( .A(y[2222]), .B(x[2222]), .Z(n9023) );
  XNOR U8994 ( .A(y[2223]), .B(x[2223]), .Z(n9022) );
  AND U8995 ( .A(n9024), .B(n9025), .Z(n8992) );
  AND U8996 ( .A(n9026), .B(n9027), .Z(n9025) );
  AND U8997 ( .A(n9028), .B(n9029), .Z(n9027) );
  AND U8998 ( .A(n9030), .B(n9031), .Z(n9029) );
  XNOR U8999 ( .A(y[2224]), .B(x[2224]), .Z(n9031) );
  XNOR U9000 ( .A(y[2225]), .B(x[2225]), .Z(n9030) );
  AND U9001 ( .A(n9032), .B(n9033), .Z(n9028) );
  XNOR U9002 ( .A(y[2226]), .B(x[2226]), .Z(n9033) );
  XNOR U9003 ( .A(y[2227]), .B(x[2227]), .Z(n9032) );
  AND U9004 ( .A(n9034), .B(n9035), .Z(n9026) );
  AND U9005 ( .A(n9036), .B(n9037), .Z(n9035) );
  XNOR U9006 ( .A(y[2228]), .B(x[2228]), .Z(n9037) );
  XNOR U9007 ( .A(y[2229]), .B(x[2229]), .Z(n9036) );
  AND U9008 ( .A(n9038), .B(n9039), .Z(n9034) );
  XNOR U9009 ( .A(y[2230]), .B(x[2230]), .Z(n9039) );
  XNOR U9010 ( .A(y[2231]), .B(x[2231]), .Z(n9038) );
  AND U9011 ( .A(n9040), .B(n9041), .Z(n9024) );
  AND U9012 ( .A(n9042), .B(n9043), .Z(n9041) );
  AND U9013 ( .A(n9044), .B(n9045), .Z(n9043) );
  XNOR U9014 ( .A(y[2232]), .B(x[2232]), .Z(n9045) );
  XNOR U9015 ( .A(y[2233]), .B(x[2233]), .Z(n9044) );
  AND U9016 ( .A(n9046), .B(n9047), .Z(n9042) );
  XNOR U9017 ( .A(y[2234]), .B(x[2234]), .Z(n9047) );
  XNOR U9018 ( .A(y[2235]), .B(x[2235]), .Z(n9046) );
  AND U9019 ( .A(n9048), .B(n9049), .Z(n9040) );
  AND U9020 ( .A(n9050), .B(n9051), .Z(n9049) );
  XNOR U9021 ( .A(y[2236]), .B(x[2236]), .Z(n9051) );
  XNOR U9022 ( .A(y[2237]), .B(x[2237]), .Z(n9050) );
  AND U9023 ( .A(n9052), .B(n9053), .Z(n9048) );
  XNOR U9024 ( .A(y[2238]), .B(x[2238]), .Z(n9053) );
  XNOR U9025 ( .A(y[2239]), .B(x[2239]), .Z(n9052) );
  AND U9026 ( .A(n9054), .B(n9055), .Z(n8926) );
  AND U9027 ( .A(n9056), .B(n9057), .Z(n9055) );
  AND U9028 ( .A(n9058), .B(n9059), .Z(n9057) );
  AND U9029 ( .A(n9060), .B(n9061), .Z(n9059) );
  AND U9030 ( .A(n9062), .B(n9063), .Z(n9061) );
  AND U9031 ( .A(n9064), .B(n9065), .Z(n9063) );
  XNOR U9032 ( .A(y[2240]), .B(x[2240]), .Z(n9065) );
  XNOR U9033 ( .A(y[2241]), .B(x[2241]), .Z(n9064) );
  AND U9034 ( .A(n9066), .B(n9067), .Z(n9062) );
  XNOR U9035 ( .A(y[2242]), .B(x[2242]), .Z(n9067) );
  XNOR U9036 ( .A(y[2243]), .B(x[2243]), .Z(n9066) );
  AND U9037 ( .A(n9068), .B(n9069), .Z(n9060) );
  AND U9038 ( .A(n9070), .B(n9071), .Z(n9069) );
  XNOR U9039 ( .A(y[2244]), .B(x[2244]), .Z(n9071) );
  XNOR U9040 ( .A(y[2245]), .B(x[2245]), .Z(n9070) );
  AND U9041 ( .A(n9072), .B(n9073), .Z(n9068) );
  XNOR U9042 ( .A(y[2246]), .B(x[2246]), .Z(n9073) );
  XNOR U9043 ( .A(y[2247]), .B(x[2247]), .Z(n9072) );
  AND U9044 ( .A(n9074), .B(n9075), .Z(n9058) );
  AND U9045 ( .A(n9076), .B(n9077), .Z(n9075) );
  AND U9046 ( .A(n9078), .B(n9079), .Z(n9077) );
  XNOR U9047 ( .A(y[2248]), .B(x[2248]), .Z(n9079) );
  XNOR U9048 ( .A(y[2249]), .B(x[2249]), .Z(n9078) );
  AND U9049 ( .A(n9080), .B(n9081), .Z(n9076) );
  XNOR U9050 ( .A(y[2250]), .B(x[2250]), .Z(n9081) );
  XNOR U9051 ( .A(y[2251]), .B(x[2251]), .Z(n9080) );
  AND U9052 ( .A(n9082), .B(n9083), .Z(n9074) );
  AND U9053 ( .A(n9084), .B(n9085), .Z(n9083) );
  XNOR U9054 ( .A(y[2252]), .B(x[2252]), .Z(n9085) );
  XNOR U9055 ( .A(y[2253]), .B(x[2253]), .Z(n9084) );
  AND U9056 ( .A(n9086), .B(n9087), .Z(n9082) );
  XNOR U9057 ( .A(y[2254]), .B(x[2254]), .Z(n9087) );
  XNOR U9058 ( .A(y[2255]), .B(x[2255]), .Z(n9086) );
  AND U9059 ( .A(n9088), .B(n9089), .Z(n9056) );
  AND U9060 ( .A(n9090), .B(n9091), .Z(n9089) );
  AND U9061 ( .A(n9092), .B(n9093), .Z(n9091) );
  AND U9062 ( .A(n9094), .B(n9095), .Z(n9093) );
  XNOR U9063 ( .A(y[2256]), .B(x[2256]), .Z(n9095) );
  XNOR U9064 ( .A(y[2257]), .B(x[2257]), .Z(n9094) );
  AND U9065 ( .A(n9096), .B(n9097), .Z(n9092) );
  XNOR U9066 ( .A(y[2258]), .B(x[2258]), .Z(n9097) );
  XNOR U9067 ( .A(y[2259]), .B(x[2259]), .Z(n9096) );
  AND U9068 ( .A(n9098), .B(n9099), .Z(n9090) );
  AND U9069 ( .A(n9100), .B(n9101), .Z(n9099) );
  XNOR U9070 ( .A(y[2260]), .B(x[2260]), .Z(n9101) );
  XNOR U9071 ( .A(y[2261]), .B(x[2261]), .Z(n9100) );
  AND U9072 ( .A(n9102), .B(n9103), .Z(n9098) );
  XNOR U9073 ( .A(y[2262]), .B(x[2262]), .Z(n9103) );
  XNOR U9074 ( .A(y[2263]), .B(x[2263]), .Z(n9102) );
  AND U9075 ( .A(n9104), .B(n9105), .Z(n9088) );
  AND U9076 ( .A(n9106), .B(n9107), .Z(n9105) );
  AND U9077 ( .A(n9108), .B(n9109), .Z(n9107) );
  XNOR U9078 ( .A(y[2264]), .B(x[2264]), .Z(n9109) );
  XNOR U9079 ( .A(y[2265]), .B(x[2265]), .Z(n9108) );
  AND U9080 ( .A(n9110), .B(n9111), .Z(n9106) );
  XNOR U9081 ( .A(y[2266]), .B(x[2266]), .Z(n9111) );
  XNOR U9082 ( .A(y[2267]), .B(x[2267]), .Z(n9110) );
  AND U9083 ( .A(n9112), .B(n9113), .Z(n9104) );
  AND U9084 ( .A(n9114), .B(n9115), .Z(n9113) );
  XNOR U9085 ( .A(y[2268]), .B(x[2268]), .Z(n9115) );
  XNOR U9086 ( .A(y[2269]), .B(x[2269]), .Z(n9114) );
  AND U9087 ( .A(n9116), .B(n9117), .Z(n9112) );
  XNOR U9088 ( .A(y[2270]), .B(x[2270]), .Z(n9117) );
  XNOR U9089 ( .A(y[2271]), .B(x[2271]), .Z(n9116) );
  AND U9090 ( .A(n9118), .B(n9119), .Z(n9054) );
  AND U9091 ( .A(n9120), .B(n9121), .Z(n9119) );
  AND U9092 ( .A(n9122), .B(n9123), .Z(n9121) );
  AND U9093 ( .A(n9124), .B(n9125), .Z(n9123) );
  AND U9094 ( .A(n9126), .B(n9127), .Z(n9125) );
  XNOR U9095 ( .A(y[2272]), .B(x[2272]), .Z(n9127) );
  XNOR U9096 ( .A(y[2273]), .B(x[2273]), .Z(n9126) );
  AND U9097 ( .A(n9128), .B(n9129), .Z(n9124) );
  XNOR U9098 ( .A(y[2274]), .B(x[2274]), .Z(n9129) );
  XNOR U9099 ( .A(y[2275]), .B(x[2275]), .Z(n9128) );
  AND U9100 ( .A(n9130), .B(n9131), .Z(n9122) );
  AND U9101 ( .A(n9132), .B(n9133), .Z(n9131) );
  XNOR U9102 ( .A(y[2276]), .B(x[2276]), .Z(n9133) );
  XNOR U9103 ( .A(y[2277]), .B(x[2277]), .Z(n9132) );
  AND U9104 ( .A(n9134), .B(n9135), .Z(n9130) );
  XNOR U9105 ( .A(y[2278]), .B(x[2278]), .Z(n9135) );
  XNOR U9106 ( .A(y[2279]), .B(x[2279]), .Z(n9134) );
  AND U9107 ( .A(n9136), .B(n9137), .Z(n9120) );
  AND U9108 ( .A(n9138), .B(n9139), .Z(n9137) );
  AND U9109 ( .A(n9140), .B(n9141), .Z(n9139) );
  XNOR U9110 ( .A(y[2280]), .B(x[2280]), .Z(n9141) );
  XNOR U9111 ( .A(y[2281]), .B(x[2281]), .Z(n9140) );
  AND U9112 ( .A(n9142), .B(n9143), .Z(n9138) );
  XNOR U9113 ( .A(y[2282]), .B(x[2282]), .Z(n9143) );
  XNOR U9114 ( .A(y[2283]), .B(x[2283]), .Z(n9142) );
  AND U9115 ( .A(n9144), .B(n9145), .Z(n9136) );
  AND U9116 ( .A(n9146), .B(n9147), .Z(n9145) );
  XNOR U9117 ( .A(y[2284]), .B(x[2284]), .Z(n9147) );
  XNOR U9118 ( .A(y[2285]), .B(x[2285]), .Z(n9146) );
  AND U9119 ( .A(n9148), .B(n9149), .Z(n9144) );
  XNOR U9120 ( .A(y[2286]), .B(x[2286]), .Z(n9149) );
  XNOR U9121 ( .A(y[2287]), .B(x[2287]), .Z(n9148) );
  AND U9122 ( .A(n9150), .B(n9151), .Z(n9118) );
  AND U9123 ( .A(n9152), .B(n9153), .Z(n9151) );
  AND U9124 ( .A(n9154), .B(n9155), .Z(n9153) );
  AND U9125 ( .A(n9156), .B(n9157), .Z(n9155) );
  XNOR U9126 ( .A(y[2288]), .B(x[2288]), .Z(n9157) );
  XNOR U9127 ( .A(y[2289]), .B(x[2289]), .Z(n9156) );
  AND U9128 ( .A(n9158), .B(n9159), .Z(n9154) );
  XNOR U9129 ( .A(y[2290]), .B(x[2290]), .Z(n9159) );
  XNOR U9130 ( .A(y[2291]), .B(x[2291]), .Z(n9158) );
  AND U9131 ( .A(n9160), .B(n9161), .Z(n9152) );
  AND U9132 ( .A(n9162), .B(n9163), .Z(n9161) );
  XNOR U9133 ( .A(y[2292]), .B(x[2292]), .Z(n9163) );
  XNOR U9134 ( .A(y[2293]), .B(x[2293]), .Z(n9162) );
  AND U9135 ( .A(n9164), .B(n9165), .Z(n9160) );
  XNOR U9136 ( .A(y[2294]), .B(x[2294]), .Z(n9165) );
  XNOR U9137 ( .A(y[2295]), .B(x[2295]), .Z(n9164) );
  AND U9138 ( .A(n9166), .B(n9167), .Z(n9150) );
  AND U9139 ( .A(n9168), .B(n9169), .Z(n9167) );
  AND U9140 ( .A(n9170), .B(n9171), .Z(n9169) );
  XNOR U9141 ( .A(y[2296]), .B(x[2296]), .Z(n9171) );
  XNOR U9142 ( .A(y[2297]), .B(x[2297]), .Z(n9170) );
  AND U9143 ( .A(n9172), .B(n9173), .Z(n9168) );
  XNOR U9144 ( .A(y[2298]), .B(x[2298]), .Z(n9173) );
  XNOR U9145 ( .A(y[2299]), .B(x[2299]), .Z(n9172) );
  AND U9146 ( .A(n9174), .B(n9175), .Z(n9166) );
  AND U9147 ( .A(n9176), .B(n9177), .Z(n9175) );
  XNOR U9148 ( .A(y[2300]), .B(x[2300]), .Z(n9177) );
  XNOR U9149 ( .A(y[2301]), .B(x[2301]), .Z(n9176) );
  AND U9150 ( .A(n9178), .B(n9179), .Z(n9174) );
  XNOR U9151 ( .A(y[2302]), .B(x[2302]), .Z(n9179) );
  XNOR U9152 ( .A(y[2303]), .B(x[2303]), .Z(n9178) );
  AND U9153 ( .A(n9180), .B(n9181), .Z(n8668) );
  AND U9154 ( .A(n9182), .B(n9183), .Z(n9181) );
  AND U9155 ( .A(n9184), .B(n9185), .Z(n9183) );
  AND U9156 ( .A(n9186), .B(n9187), .Z(n9185) );
  AND U9157 ( .A(n9188), .B(n9189), .Z(n9187) );
  AND U9158 ( .A(n9190), .B(n9191), .Z(n9189) );
  XNOR U9159 ( .A(y[2946]), .B(x[2946]), .Z(n9191) );
  XNOR U9160 ( .A(y[2947]), .B(x[2947]), .Z(n9190) );
  AND U9161 ( .A(n9192), .B(n9193), .Z(n9188) );
  XNOR U9162 ( .A(y[2948]), .B(x[2948]), .Z(n9193) );
  XNOR U9163 ( .A(y[2949]), .B(x[2949]), .Z(n9192) );
  AND U9164 ( .A(n9194), .B(n9195), .Z(n9186) );
  AND U9165 ( .A(n9196), .B(n9197), .Z(n9195) );
  XNOR U9166 ( .A(y[2950]), .B(x[2950]), .Z(n9197) );
  XNOR U9167 ( .A(y[2951]), .B(x[2951]), .Z(n9196) );
  AND U9168 ( .A(n9198), .B(n9199), .Z(n9194) );
  XNOR U9169 ( .A(y[2952]), .B(x[2952]), .Z(n9199) );
  XNOR U9170 ( .A(y[2953]), .B(x[2953]), .Z(n9198) );
  AND U9171 ( .A(n9200), .B(n9201), .Z(n9184) );
  AND U9172 ( .A(n9202), .B(n9203), .Z(n9201) );
  AND U9173 ( .A(n9204), .B(n9205), .Z(n9203) );
  XNOR U9174 ( .A(y[2954]), .B(x[2954]), .Z(n9205) );
  XNOR U9175 ( .A(y[2955]), .B(x[2955]), .Z(n9204) );
  AND U9176 ( .A(n9206), .B(n9207), .Z(n9202) );
  XNOR U9177 ( .A(y[2956]), .B(x[2956]), .Z(n9207) );
  XNOR U9178 ( .A(y[2957]), .B(x[2957]), .Z(n9206) );
  AND U9179 ( .A(n9208), .B(n9209), .Z(n9200) );
  AND U9180 ( .A(n9210), .B(n9211), .Z(n9209) );
  XNOR U9181 ( .A(y[2958]), .B(x[2958]), .Z(n9211) );
  XNOR U9182 ( .A(y[2959]), .B(x[2959]), .Z(n9210) );
  AND U9183 ( .A(n9212), .B(n9213), .Z(n9208) );
  XNOR U9184 ( .A(y[2960]), .B(x[2960]), .Z(n9213) );
  XNOR U9185 ( .A(y[2961]), .B(x[2961]), .Z(n9212) );
  AND U9186 ( .A(n9214), .B(n9215), .Z(n9182) );
  AND U9187 ( .A(n9216), .B(n9217), .Z(n9215) );
  AND U9188 ( .A(n9218), .B(n9219), .Z(n9217) );
  AND U9189 ( .A(n9220), .B(n9221), .Z(n9219) );
  XNOR U9190 ( .A(y[2962]), .B(x[2962]), .Z(n9221) );
  XNOR U9191 ( .A(y[2963]), .B(x[2963]), .Z(n9220) );
  AND U9192 ( .A(n9222), .B(n9223), .Z(n9218) );
  XNOR U9193 ( .A(y[2964]), .B(x[2964]), .Z(n9223) );
  XNOR U9194 ( .A(y[2965]), .B(x[2965]), .Z(n9222) );
  AND U9195 ( .A(n9224), .B(n9225), .Z(n9216) );
  AND U9196 ( .A(n9226), .B(n9227), .Z(n9225) );
  XNOR U9197 ( .A(y[2966]), .B(x[2966]), .Z(n9227) );
  XNOR U9198 ( .A(y[2967]), .B(x[2967]), .Z(n9226) );
  AND U9199 ( .A(n9228), .B(n9229), .Z(n9224) );
  XNOR U9200 ( .A(y[2968]), .B(x[2968]), .Z(n9229) );
  XNOR U9201 ( .A(y[2969]), .B(x[2969]), .Z(n9228) );
  AND U9202 ( .A(n9230), .B(n9231), .Z(n9214) );
  AND U9203 ( .A(n9232), .B(n9233), .Z(n9231) );
  AND U9204 ( .A(n9234), .B(n9235), .Z(n9233) );
  XNOR U9205 ( .A(y[2970]), .B(x[2970]), .Z(n9235) );
  XNOR U9206 ( .A(y[2971]), .B(x[2971]), .Z(n9234) );
  AND U9207 ( .A(n9236), .B(n9237), .Z(n9232) );
  XNOR U9208 ( .A(y[2972]), .B(x[2972]), .Z(n9237) );
  XNOR U9209 ( .A(y[2973]), .B(x[2973]), .Z(n9236) );
  AND U9210 ( .A(n9238), .B(n9239), .Z(n9230) );
  AND U9211 ( .A(n9240), .B(n9241), .Z(n9239) );
  XNOR U9212 ( .A(y[2974]), .B(x[2974]), .Z(n9241) );
  XNOR U9213 ( .A(y[2975]), .B(x[2975]), .Z(n9240) );
  AND U9214 ( .A(n9242), .B(n9243), .Z(n9238) );
  XNOR U9215 ( .A(y[2976]), .B(x[2976]), .Z(n9243) );
  XNOR U9216 ( .A(y[2977]), .B(x[2977]), .Z(n9242) );
  AND U9217 ( .A(n9244), .B(n9245), .Z(n9180) );
  AND U9218 ( .A(n9246), .B(n9247), .Z(n9245) );
  AND U9219 ( .A(n9248), .B(n9249), .Z(n9247) );
  AND U9220 ( .A(n9250), .B(n9251), .Z(n9249) );
  AND U9221 ( .A(n9252), .B(n9253), .Z(n9251) );
  XNOR U9222 ( .A(y[2978]), .B(x[2978]), .Z(n9253) );
  XNOR U9223 ( .A(y[2979]), .B(x[2979]), .Z(n9252) );
  AND U9224 ( .A(n9254), .B(n9255), .Z(n9250) );
  XNOR U9225 ( .A(y[2980]), .B(x[2980]), .Z(n9255) );
  XNOR U9226 ( .A(y[2981]), .B(x[2981]), .Z(n9254) );
  AND U9227 ( .A(n9256), .B(n9257), .Z(n9248) );
  AND U9228 ( .A(n9258), .B(n9259), .Z(n9257) );
  XNOR U9229 ( .A(y[2982]), .B(x[2982]), .Z(n9259) );
  XNOR U9230 ( .A(y[2983]), .B(x[2983]), .Z(n9258) );
  AND U9231 ( .A(n9260), .B(n9261), .Z(n9256) );
  XNOR U9232 ( .A(y[2984]), .B(x[2984]), .Z(n9261) );
  XNOR U9233 ( .A(y[2985]), .B(x[2985]), .Z(n9260) );
  AND U9234 ( .A(n9262), .B(n9263), .Z(n9246) );
  AND U9235 ( .A(n9264), .B(n9265), .Z(n9263) );
  AND U9236 ( .A(n9266), .B(n9267), .Z(n9265) );
  XNOR U9237 ( .A(y[2986]), .B(x[2986]), .Z(n9267) );
  XNOR U9238 ( .A(y[2987]), .B(x[2987]), .Z(n9266) );
  AND U9239 ( .A(n9268), .B(n9269), .Z(n9264) );
  XNOR U9240 ( .A(y[2988]), .B(x[2988]), .Z(n9269) );
  XNOR U9241 ( .A(y[2989]), .B(x[2989]), .Z(n9268) );
  AND U9242 ( .A(n9270), .B(n9271), .Z(n9262) );
  AND U9243 ( .A(n9272), .B(n9273), .Z(n9271) );
  XNOR U9244 ( .A(y[2990]), .B(x[2990]), .Z(n9273) );
  XNOR U9245 ( .A(y[2991]), .B(x[2991]), .Z(n9272) );
  AND U9246 ( .A(n9274), .B(n9275), .Z(n9270) );
  XNOR U9247 ( .A(y[2992]), .B(x[2992]), .Z(n9275) );
  XNOR U9248 ( .A(y[2993]), .B(x[2993]), .Z(n9274) );
  AND U9249 ( .A(n9276), .B(n9277), .Z(n9244) );
  AND U9250 ( .A(n9278), .B(n9279), .Z(n9277) );
  AND U9251 ( .A(n9280), .B(n9281), .Z(n9279) );
  AND U9252 ( .A(n9282), .B(n9283), .Z(n9281) );
  XNOR U9253 ( .A(y[2994]), .B(x[2994]), .Z(n9283) );
  XNOR U9254 ( .A(y[2995]), .B(x[2995]), .Z(n9282) );
  AND U9255 ( .A(n9284), .B(n9285), .Z(n9280) );
  XNOR U9256 ( .A(y[2996]), .B(x[2996]), .Z(n9285) );
  XNOR U9257 ( .A(y[2997]), .B(x[2997]), .Z(n9284) );
  AND U9258 ( .A(n9286), .B(n9287), .Z(n9278) );
  AND U9259 ( .A(n9288), .B(n9289), .Z(n9287) );
  XNOR U9260 ( .A(y[2998]), .B(x[2998]), .Z(n9289) );
  XNOR U9261 ( .A(y[2999]), .B(x[2999]), .Z(n9288) );
  AND U9262 ( .A(n9290), .B(n9291), .Z(n9286) );
  XNOR U9263 ( .A(y[3000]), .B(x[3000]), .Z(n9291) );
  XNOR U9264 ( .A(y[3001]), .B(x[3001]), .Z(n9290) );
  AND U9265 ( .A(n9292), .B(n9293), .Z(n9276) );
  AND U9266 ( .A(n9294), .B(n9295), .Z(n9293) );
  AND U9267 ( .A(n9296), .B(n9297), .Z(n9295) );
  XNOR U9268 ( .A(y[3002]), .B(x[3002]), .Z(n9297) );
  XNOR U9269 ( .A(y[3003]), .B(x[3003]), .Z(n9296) );
  AND U9270 ( .A(n9298), .B(n9299), .Z(n9294) );
  XNOR U9271 ( .A(y[3004]), .B(x[3004]), .Z(n9299) );
  XNOR U9272 ( .A(y[3005]), .B(x[3005]), .Z(n9298) );
  AND U9273 ( .A(n9300), .B(n9301), .Z(n9292) );
  AND U9274 ( .A(n9302), .B(n9303), .Z(n9301) );
  XNOR U9275 ( .A(y[3006]), .B(x[3006]), .Z(n9303) );
  XNOR U9276 ( .A(y[3007]), .B(x[3007]), .Z(n9302) );
  AND U9277 ( .A(n9304), .B(n9305), .Z(n9300) );
  XNOR U9278 ( .A(y[3008]), .B(x[3008]), .Z(n9305) );
  XNOR U9279 ( .A(y[3009]), .B(x[3009]), .Z(n9304) );
  AND U9280 ( .A(n9306), .B(n9307), .Z(n8666) );
  AND U9281 ( .A(n9308), .B(n9309), .Z(n9307) );
  AND U9282 ( .A(n9310), .B(n9311), .Z(n9309) );
  AND U9283 ( .A(n9312), .B(n9313), .Z(n9311) );
  AND U9284 ( .A(n9314), .B(n9315), .Z(n9313) );
  AND U9285 ( .A(n9316), .B(n9317), .Z(n9315) );
  AND U9286 ( .A(n9318), .B(n9319), .Z(n9317) );
  AND U9287 ( .A(n9320), .B(n9321), .Z(n9319) );
  XNOR U9288 ( .A(y[2818]), .B(x[2818]), .Z(n9321) );
  XNOR U9289 ( .A(y[2819]), .B(x[2819]), .Z(n9320) );
  AND U9290 ( .A(n9322), .B(n9323), .Z(n9318) );
  XNOR U9291 ( .A(y[2820]), .B(x[2820]), .Z(n9323) );
  XNOR U9292 ( .A(y[2821]), .B(x[2821]), .Z(n9322) );
  AND U9293 ( .A(n9324), .B(n9325), .Z(n9316) );
  AND U9294 ( .A(n9326), .B(n9327), .Z(n9325) );
  XNOR U9295 ( .A(y[2822]), .B(x[2822]), .Z(n9327) );
  XNOR U9296 ( .A(y[2823]), .B(x[2823]), .Z(n9326) );
  AND U9297 ( .A(n9328), .B(n9329), .Z(n9324) );
  XNOR U9298 ( .A(y[2824]), .B(x[2824]), .Z(n9329) );
  XNOR U9299 ( .A(y[2825]), .B(x[2825]), .Z(n9328) );
  AND U9300 ( .A(n9330), .B(n9331), .Z(n9314) );
  AND U9301 ( .A(n9332), .B(n9333), .Z(n9331) );
  AND U9302 ( .A(n9334), .B(n9335), .Z(n9333) );
  XNOR U9303 ( .A(y[2826]), .B(x[2826]), .Z(n9335) );
  XNOR U9304 ( .A(y[2827]), .B(x[2827]), .Z(n9334) );
  AND U9305 ( .A(n9336), .B(n9337), .Z(n9332) );
  XNOR U9306 ( .A(y[2828]), .B(x[2828]), .Z(n9337) );
  XNOR U9307 ( .A(y[2829]), .B(x[2829]), .Z(n9336) );
  AND U9308 ( .A(n9338), .B(n9339), .Z(n9330) );
  AND U9309 ( .A(n9340), .B(n9341), .Z(n9339) );
  XNOR U9310 ( .A(y[2830]), .B(x[2830]), .Z(n9341) );
  XNOR U9311 ( .A(y[2831]), .B(x[2831]), .Z(n9340) );
  AND U9312 ( .A(n9342), .B(n9343), .Z(n9338) );
  XNOR U9313 ( .A(y[2832]), .B(x[2832]), .Z(n9343) );
  XNOR U9314 ( .A(y[2833]), .B(x[2833]), .Z(n9342) );
  AND U9315 ( .A(n9344), .B(n9345), .Z(n9312) );
  AND U9316 ( .A(n9346), .B(n9347), .Z(n9345) );
  AND U9317 ( .A(n9348), .B(n9349), .Z(n9347) );
  AND U9318 ( .A(n9350), .B(n9351), .Z(n9349) );
  XNOR U9319 ( .A(y[2834]), .B(x[2834]), .Z(n9351) );
  XNOR U9320 ( .A(y[2835]), .B(x[2835]), .Z(n9350) );
  AND U9321 ( .A(n9352), .B(n9353), .Z(n9348) );
  XNOR U9322 ( .A(y[2836]), .B(x[2836]), .Z(n9353) );
  XNOR U9323 ( .A(y[2837]), .B(x[2837]), .Z(n9352) );
  AND U9324 ( .A(n9354), .B(n9355), .Z(n9346) );
  AND U9325 ( .A(n9356), .B(n9357), .Z(n9355) );
  XNOR U9326 ( .A(y[2838]), .B(x[2838]), .Z(n9357) );
  XNOR U9327 ( .A(y[2839]), .B(x[2839]), .Z(n9356) );
  AND U9328 ( .A(n9358), .B(n9359), .Z(n9354) );
  XNOR U9329 ( .A(y[2840]), .B(x[2840]), .Z(n9359) );
  XNOR U9330 ( .A(y[2841]), .B(x[2841]), .Z(n9358) );
  AND U9331 ( .A(n9360), .B(n9361), .Z(n9344) );
  AND U9332 ( .A(n9362), .B(n9363), .Z(n9361) );
  AND U9333 ( .A(n9364), .B(n9365), .Z(n9363) );
  XNOR U9334 ( .A(y[2842]), .B(x[2842]), .Z(n9365) );
  XNOR U9335 ( .A(y[2843]), .B(x[2843]), .Z(n9364) );
  AND U9336 ( .A(n9366), .B(n9367), .Z(n9362) );
  XNOR U9337 ( .A(y[2844]), .B(x[2844]), .Z(n9367) );
  XNOR U9338 ( .A(y[2845]), .B(x[2845]), .Z(n9366) );
  AND U9339 ( .A(n9368), .B(n9369), .Z(n9360) );
  AND U9340 ( .A(n9370), .B(n9371), .Z(n9369) );
  XNOR U9341 ( .A(y[2846]), .B(x[2846]), .Z(n9371) );
  XNOR U9342 ( .A(y[2847]), .B(x[2847]), .Z(n9370) );
  AND U9343 ( .A(n9372), .B(n9373), .Z(n9368) );
  XNOR U9344 ( .A(y[2848]), .B(x[2848]), .Z(n9373) );
  XNOR U9345 ( .A(y[2849]), .B(x[2849]), .Z(n9372) );
  AND U9346 ( .A(n9374), .B(n9375), .Z(n9310) );
  AND U9347 ( .A(n9376), .B(n9377), .Z(n9375) );
  AND U9348 ( .A(n9378), .B(n9379), .Z(n9377) );
  AND U9349 ( .A(n9380), .B(n9381), .Z(n9379) );
  AND U9350 ( .A(n9382), .B(n9383), .Z(n9381) );
  XNOR U9351 ( .A(y[2850]), .B(x[2850]), .Z(n9383) );
  XNOR U9352 ( .A(y[2851]), .B(x[2851]), .Z(n9382) );
  AND U9353 ( .A(n9384), .B(n9385), .Z(n9380) );
  XNOR U9354 ( .A(y[2852]), .B(x[2852]), .Z(n9385) );
  XNOR U9355 ( .A(y[2853]), .B(x[2853]), .Z(n9384) );
  AND U9356 ( .A(n9386), .B(n9387), .Z(n9378) );
  AND U9357 ( .A(n9388), .B(n9389), .Z(n9387) );
  XNOR U9358 ( .A(y[2854]), .B(x[2854]), .Z(n9389) );
  XNOR U9359 ( .A(y[2855]), .B(x[2855]), .Z(n9388) );
  AND U9360 ( .A(n9390), .B(n9391), .Z(n9386) );
  XNOR U9361 ( .A(y[2856]), .B(x[2856]), .Z(n9391) );
  XNOR U9362 ( .A(y[2857]), .B(x[2857]), .Z(n9390) );
  AND U9363 ( .A(n9392), .B(n9393), .Z(n9376) );
  AND U9364 ( .A(n9394), .B(n9395), .Z(n9393) );
  AND U9365 ( .A(n9396), .B(n9397), .Z(n9395) );
  XNOR U9366 ( .A(y[2858]), .B(x[2858]), .Z(n9397) );
  XNOR U9367 ( .A(y[2859]), .B(x[2859]), .Z(n9396) );
  AND U9368 ( .A(n9398), .B(n9399), .Z(n9394) );
  XNOR U9369 ( .A(y[2860]), .B(x[2860]), .Z(n9399) );
  XNOR U9370 ( .A(y[2861]), .B(x[2861]), .Z(n9398) );
  AND U9371 ( .A(n9400), .B(n9401), .Z(n9392) );
  AND U9372 ( .A(n9402), .B(n9403), .Z(n9401) );
  XNOR U9373 ( .A(y[2862]), .B(x[2862]), .Z(n9403) );
  XNOR U9374 ( .A(y[2863]), .B(x[2863]), .Z(n9402) );
  AND U9375 ( .A(n9404), .B(n9405), .Z(n9400) );
  XNOR U9376 ( .A(y[2864]), .B(x[2864]), .Z(n9405) );
  XNOR U9377 ( .A(y[2865]), .B(x[2865]), .Z(n9404) );
  AND U9378 ( .A(n9406), .B(n9407), .Z(n9374) );
  AND U9379 ( .A(n9408), .B(n9409), .Z(n9407) );
  AND U9380 ( .A(n9410), .B(n9411), .Z(n9409) );
  AND U9381 ( .A(n9412), .B(n9413), .Z(n9411) );
  XNOR U9382 ( .A(y[2866]), .B(x[2866]), .Z(n9413) );
  XNOR U9383 ( .A(y[2867]), .B(x[2867]), .Z(n9412) );
  AND U9384 ( .A(n9414), .B(n9415), .Z(n9410) );
  XNOR U9385 ( .A(y[2868]), .B(x[2868]), .Z(n9415) );
  XNOR U9386 ( .A(y[2869]), .B(x[2869]), .Z(n9414) );
  AND U9387 ( .A(n9416), .B(n9417), .Z(n9408) );
  AND U9388 ( .A(n9418), .B(n9419), .Z(n9417) );
  XNOR U9389 ( .A(y[2870]), .B(x[2870]), .Z(n9419) );
  XNOR U9390 ( .A(y[2871]), .B(x[2871]), .Z(n9418) );
  AND U9391 ( .A(n9420), .B(n9421), .Z(n9416) );
  XNOR U9392 ( .A(y[2872]), .B(x[2872]), .Z(n9421) );
  XNOR U9393 ( .A(y[2873]), .B(x[2873]), .Z(n9420) );
  AND U9394 ( .A(n9422), .B(n9423), .Z(n9406) );
  AND U9395 ( .A(n9424), .B(n9425), .Z(n9423) );
  AND U9396 ( .A(n9426), .B(n9427), .Z(n9425) );
  XNOR U9397 ( .A(y[2874]), .B(x[2874]), .Z(n9427) );
  XNOR U9398 ( .A(y[2875]), .B(x[2875]), .Z(n9426) );
  AND U9399 ( .A(n9428), .B(n9429), .Z(n9424) );
  XNOR U9400 ( .A(y[2876]), .B(x[2876]), .Z(n9429) );
  XNOR U9401 ( .A(y[2877]), .B(x[2877]), .Z(n9428) );
  AND U9402 ( .A(n9430), .B(n9431), .Z(n9422) );
  AND U9403 ( .A(n9432), .B(n9433), .Z(n9431) );
  XNOR U9404 ( .A(y[2878]), .B(x[2878]), .Z(n9433) );
  XNOR U9405 ( .A(y[2879]), .B(x[2879]), .Z(n9432) );
  AND U9406 ( .A(n9434), .B(n9435), .Z(n9430) );
  XNOR U9407 ( .A(y[2880]), .B(x[2880]), .Z(n9435) );
  XNOR U9408 ( .A(y[2881]), .B(x[2881]), .Z(n9434) );
  AND U9409 ( .A(n9436), .B(n9437), .Z(n9308) );
  AND U9410 ( .A(n9438), .B(n9439), .Z(n9437) );
  AND U9411 ( .A(n9440), .B(n9441), .Z(n9439) );
  AND U9412 ( .A(n9442), .B(n9443), .Z(n9441) );
  AND U9413 ( .A(n9444), .B(n9445), .Z(n9443) );
  AND U9414 ( .A(n9446), .B(n9447), .Z(n9445) );
  XNOR U9415 ( .A(y[2882]), .B(x[2882]), .Z(n9447) );
  XNOR U9416 ( .A(y[2883]), .B(x[2883]), .Z(n9446) );
  AND U9417 ( .A(n9448), .B(n9449), .Z(n9444) );
  XNOR U9418 ( .A(y[2884]), .B(x[2884]), .Z(n9449) );
  XNOR U9419 ( .A(y[2885]), .B(x[2885]), .Z(n9448) );
  AND U9420 ( .A(n9450), .B(n9451), .Z(n9442) );
  AND U9421 ( .A(n9452), .B(n9453), .Z(n9451) );
  XNOR U9422 ( .A(y[2886]), .B(x[2886]), .Z(n9453) );
  XNOR U9423 ( .A(y[2887]), .B(x[2887]), .Z(n9452) );
  AND U9424 ( .A(n9454), .B(n9455), .Z(n9450) );
  XNOR U9425 ( .A(y[2888]), .B(x[2888]), .Z(n9455) );
  XNOR U9426 ( .A(y[2889]), .B(x[2889]), .Z(n9454) );
  AND U9427 ( .A(n9456), .B(n9457), .Z(n9440) );
  AND U9428 ( .A(n9458), .B(n9459), .Z(n9457) );
  AND U9429 ( .A(n9460), .B(n9461), .Z(n9459) );
  XNOR U9430 ( .A(y[2890]), .B(x[2890]), .Z(n9461) );
  XNOR U9431 ( .A(y[2891]), .B(x[2891]), .Z(n9460) );
  AND U9432 ( .A(n9462), .B(n9463), .Z(n9458) );
  XNOR U9433 ( .A(y[2892]), .B(x[2892]), .Z(n9463) );
  XNOR U9434 ( .A(y[2893]), .B(x[2893]), .Z(n9462) );
  AND U9435 ( .A(n9464), .B(n9465), .Z(n9456) );
  AND U9436 ( .A(n9466), .B(n9467), .Z(n9465) );
  XNOR U9437 ( .A(y[2894]), .B(x[2894]), .Z(n9467) );
  XNOR U9438 ( .A(y[2895]), .B(x[2895]), .Z(n9466) );
  AND U9439 ( .A(n9468), .B(n9469), .Z(n9464) );
  XNOR U9440 ( .A(y[2896]), .B(x[2896]), .Z(n9469) );
  XNOR U9441 ( .A(y[2897]), .B(x[2897]), .Z(n9468) );
  AND U9442 ( .A(n9470), .B(n9471), .Z(n9438) );
  AND U9443 ( .A(n9472), .B(n9473), .Z(n9471) );
  AND U9444 ( .A(n9474), .B(n9475), .Z(n9473) );
  AND U9445 ( .A(n9476), .B(n9477), .Z(n9475) );
  XNOR U9446 ( .A(y[2898]), .B(x[2898]), .Z(n9477) );
  XNOR U9447 ( .A(y[2899]), .B(x[2899]), .Z(n9476) );
  AND U9448 ( .A(n9478), .B(n9479), .Z(n9474) );
  XNOR U9449 ( .A(y[2900]), .B(x[2900]), .Z(n9479) );
  XNOR U9450 ( .A(y[2901]), .B(x[2901]), .Z(n9478) );
  AND U9451 ( .A(n9480), .B(n9481), .Z(n9472) );
  AND U9452 ( .A(n9482), .B(n9483), .Z(n9481) );
  XNOR U9453 ( .A(y[2902]), .B(x[2902]), .Z(n9483) );
  XNOR U9454 ( .A(y[2903]), .B(x[2903]), .Z(n9482) );
  AND U9455 ( .A(n9484), .B(n9485), .Z(n9480) );
  XNOR U9456 ( .A(y[2904]), .B(x[2904]), .Z(n9485) );
  XNOR U9457 ( .A(y[2905]), .B(x[2905]), .Z(n9484) );
  AND U9458 ( .A(n9486), .B(n9487), .Z(n9470) );
  AND U9459 ( .A(n9488), .B(n9489), .Z(n9487) );
  AND U9460 ( .A(n9490), .B(n9491), .Z(n9489) );
  XNOR U9461 ( .A(y[2906]), .B(x[2906]), .Z(n9491) );
  XNOR U9462 ( .A(y[2907]), .B(x[2907]), .Z(n9490) );
  AND U9463 ( .A(n9492), .B(n9493), .Z(n9488) );
  XNOR U9464 ( .A(y[2908]), .B(x[2908]), .Z(n9493) );
  XNOR U9465 ( .A(y[2909]), .B(x[2909]), .Z(n9492) );
  AND U9466 ( .A(n9494), .B(n9495), .Z(n9486) );
  AND U9467 ( .A(n9496), .B(n9497), .Z(n9495) );
  XNOR U9468 ( .A(y[2910]), .B(x[2910]), .Z(n9497) );
  XNOR U9469 ( .A(y[2911]), .B(x[2911]), .Z(n9496) );
  AND U9470 ( .A(n9498), .B(n9499), .Z(n9494) );
  XNOR U9471 ( .A(y[2912]), .B(x[2912]), .Z(n9499) );
  XNOR U9472 ( .A(y[2913]), .B(x[2913]), .Z(n9498) );
  AND U9473 ( .A(n9500), .B(n9501), .Z(n9436) );
  AND U9474 ( .A(n9502), .B(n9503), .Z(n9501) );
  AND U9475 ( .A(n9504), .B(n9505), .Z(n9503) );
  AND U9476 ( .A(n9506), .B(n9507), .Z(n9505) );
  AND U9477 ( .A(n9508), .B(n9509), .Z(n9507) );
  XNOR U9478 ( .A(y[2914]), .B(x[2914]), .Z(n9509) );
  XNOR U9479 ( .A(y[2915]), .B(x[2915]), .Z(n9508) );
  AND U9480 ( .A(n9510), .B(n9511), .Z(n9506) );
  XNOR U9481 ( .A(y[2916]), .B(x[2916]), .Z(n9511) );
  XNOR U9482 ( .A(y[2917]), .B(x[2917]), .Z(n9510) );
  AND U9483 ( .A(n9512), .B(n9513), .Z(n9504) );
  AND U9484 ( .A(n9514), .B(n9515), .Z(n9513) );
  XNOR U9485 ( .A(y[2918]), .B(x[2918]), .Z(n9515) );
  XNOR U9486 ( .A(y[2919]), .B(x[2919]), .Z(n9514) );
  AND U9487 ( .A(n9516), .B(n9517), .Z(n9512) );
  XNOR U9488 ( .A(y[2920]), .B(x[2920]), .Z(n9517) );
  XNOR U9489 ( .A(y[2921]), .B(x[2921]), .Z(n9516) );
  AND U9490 ( .A(n9518), .B(n9519), .Z(n9502) );
  AND U9491 ( .A(n9520), .B(n9521), .Z(n9519) );
  AND U9492 ( .A(n9522), .B(n9523), .Z(n9521) );
  XNOR U9493 ( .A(y[2922]), .B(x[2922]), .Z(n9523) );
  XNOR U9494 ( .A(y[2923]), .B(x[2923]), .Z(n9522) );
  AND U9495 ( .A(n9524), .B(n9525), .Z(n9520) );
  XNOR U9496 ( .A(y[2924]), .B(x[2924]), .Z(n9525) );
  XNOR U9497 ( .A(y[2925]), .B(x[2925]), .Z(n9524) );
  AND U9498 ( .A(n9526), .B(n9527), .Z(n9518) );
  AND U9499 ( .A(n9528), .B(n9529), .Z(n9527) );
  XNOR U9500 ( .A(y[2926]), .B(x[2926]), .Z(n9529) );
  XNOR U9501 ( .A(y[2927]), .B(x[2927]), .Z(n9528) );
  AND U9502 ( .A(n9530), .B(n9531), .Z(n9526) );
  XNOR U9503 ( .A(y[2928]), .B(x[2928]), .Z(n9531) );
  XNOR U9504 ( .A(y[2929]), .B(x[2929]), .Z(n9530) );
  AND U9505 ( .A(n9532), .B(n9533), .Z(n9500) );
  AND U9506 ( .A(n9534), .B(n9535), .Z(n9533) );
  AND U9507 ( .A(n9536), .B(n9537), .Z(n9535) );
  AND U9508 ( .A(n9538), .B(n9539), .Z(n9537) );
  XNOR U9509 ( .A(y[2930]), .B(x[2930]), .Z(n9539) );
  XNOR U9510 ( .A(y[2931]), .B(x[2931]), .Z(n9538) );
  AND U9511 ( .A(n9540), .B(n9541), .Z(n9536) );
  XNOR U9512 ( .A(y[2932]), .B(x[2932]), .Z(n9541) );
  XNOR U9513 ( .A(y[2933]), .B(x[2933]), .Z(n9540) );
  AND U9514 ( .A(n9542), .B(n9543), .Z(n9534) );
  AND U9515 ( .A(n9544), .B(n9545), .Z(n9543) );
  XNOR U9516 ( .A(y[2934]), .B(x[2934]), .Z(n9545) );
  XNOR U9517 ( .A(y[2935]), .B(x[2935]), .Z(n9544) );
  AND U9518 ( .A(n9546), .B(n9547), .Z(n9542) );
  XNOR U9519 ( .A(y[2936]), .B(x[2936]), .Z(n9547) );
  XNOR U9520 ( .A(y[2937]), .B(x[2937]), .Z(n9546) );
  AND U9521 ( .A(n9548), .B(n9549), .Z(n9532) );
  AND U9522 ( .A(n9550), .B(n9551), .Z(n9549) );
  AND U9523 ( .A(n9552), .B(n9553), .Z(n9551) );
  XNOR U9524 ( .A(y[2938]), .B(x[2938]), .Z(n9553) );
  XNOR U9525 ( .A(y[2939]), .B(x[2939]), .Z(n9552) );
  AND U9526 ( .A(n9554), .B(n9555), .Z(n9550) );
  XNOR U9527 ( .A(y[2940]), .B(x[2940]), .Z(n9555) );
  XNOR U9528 ( .A(y[2941]), .B(x[2941]), .Z(n9554) );
  AND U9529 ( .A(n9556), .B(n9557), .Z(n9548) );
  AND U9530 ( .A(n9558), .B(n9559), .Z(n9557) );
  XNOR U9531 ( .A(y[2942]), .B(x[2942]), .Z(n9559) );
  XNOR U9532 ( .A(y[2943]), .B(x[2943]), .Z(n9558) );
  AND U9533 ( .A(n9560), .B(n9561), .Z(n9556) );
  XNOR U9534 ( .A(y[2944]), .B(x[2944]), .Z(n9561) );
  XNOR U9535 ( .A(y[2945]), .B(x[2945]), .Z(n9560) );
  AND U9536 ( .A(n9562), .B(n9563), .Z(n9306) );
  AND U9537 ( .A(n9564), .B(n9565), .Z(n9563) );
  AND U9538 ( .A(n9566), .B(n9567), .Z(n9565) );
  AND U9539 ( .A(n9568), .B(n9569), .Z(n9567) );
  AND U9540 ( .A(n9570), .B(n9571), .Z(n9569) );
  AND U9541 ( .A(n9572), .B(n9573), .Z(n9571) );
  AND U9542 ( .A(n9574), .B(n9575), .Z(n9573) );
  AND U9543 ( .A(n9576), .B(n9577), .Z(n9575) );
  XNOR U9544 ( .A(y[2562]), .B(x[2562]), .Z(n9577) );
  XNOR U9545 ( .A(y[2563]), .B(x[2563]), .Z(n9576) );
  AND U9546 ( .A(n9578), .B(n9579), .Z(n9574) );
  XNOR U9547 ( .A(y[2564]), .B(x[2564]), .Z(n9579) );
  XNOR U9548 ( .A(y[2567]), .B(x[2567]), .Z(n9578) );
  AND U9549 ( .A(n9580), .B(n9581), .Z(n9572) );
  AND U9550 ( .A(n9582), .B(n9583), .Z(n9581) );
  XNOR U9551 ( .A(y[2565]), .B(x[2565]), .Z(n9583) );
  XNOR U9552 ( .A(y[2566]), .B(x[2566]), .Z(n9582) );
  AND U9553 ( .A(n9584), .B(n9585), .Z(n9580) );
  XNOR U9554 ( .A(y[2568]), .B(x[2568]), .Z(n9585) );
  XNOR U9555 ( .A(y[2569]), .B(x[2569]), .Z(n9584) );
  AND U9556 ( .A(n9586), .B(n9587), .Z(n9570) );
  AND U9557 ( .A(n9588), .B(n9589), .Z(n9587) );
  AND U9558 ( .A(n9590), .B(n9591), .Z(n9589) );
  XNOR U9559 ( .A(y[2570]), .B(x[2570]), .Z(n9591) );
  XNOR U9560 ( .A(y[2571]), .B(x[2571]), .Z(n9590) );
  AND U9561 ( .A(n9592), .B(n9593), .Z(n9588) );
  XNOR U9562 ( .A(y[2572]), .B(x[2572]), .Z(n9593) );
  XNOR U9563 ( .A(y[2573]), .B(x[2573]), .Z(n9592) );
  AND U9564 ( .A(n9594), .B(n9595), .Z(n9586) );
  AND U9565 ( .A(n9596), .B(n9597), .Z(n9595) );
  XNOR U9566 ( .A(y[2574]), .B(x[2574]), .Z(n9597) );
  XNOR U9567 ( .A(y[2575]), .B(x[2575]), .Z(n9596) );
  AND U9568 ( .A(n9598), .B(n9599), .Z(n9594) );
  XNOR U9569 ( .A(y[2576]), .B(x[2576]), .Z(n9599) );
  XNOR U9570 ( .A(y[2577]), .B(x[2577]), .Z(n9598) );
  AND U9571 ( .A(n9600), .B(n9601), .Z(n9568) );
  AND U9572 ( .A(n9602), .B(n9603), .Z(n9601) );
  AND U9573 ( .A(n9604), .B(n9605), .Z(n9603) );
  AND U9574 ( .A(n9606), .B(n9607), .Z(n9605) );
  XNOR U9575 ( .A(y[2578]), .B(x[2578]), .Z(n9607) );
  XNOR U9576 ( .A(y[2579]), .B(x[2579]), .Z(n9606) );
  AND U9577 ( .A(n9608), .B(n9609), .Z(n9604) );
  XNOR U9578 ( .A(y[2580]), .B(x[2580]), .Z(n9609) );
  XNOR U9579 ( .A(y[2581]), .B(x[2581]), .Z(n9608) );
  AND U9580 ( .A(n9610), .B(n9611), .Z(n9602) );
  AND U9581 ( .A(n9612), .B(n9613), .Z(n9611) );
  XNOR U9582 ( .A(y[2582]), .B(x[2582]), .Z(n9613) );
  XNOR U9583 ( .A(y[2583]), .B(x[2583]), .Z(n9612) );
  AND U9584 ( .A(n9614), .B(n9615), .Z(n9610) );
  XNOR U9585 ( .A(y[2584]), .B(x[2584]), .Z(n9615) );
  XNOR U9586 ( .A(y[2585]), .B(x[2585]), .Z(n9614) );
  AND U9587 ( .A(n9616), .B(n9617), .Z(n9600) );
  AND U9588 ( .A(n9618), .B(n9619), .Z(n9617) );
  AND U9589 ( .A(n9620), .B(n9621), .Z(n9619) );
  XNOR U9590 ( .A(y[2586]), .B(x[2586]), .Z(n9621) );
  XNOR U9591 ( .A(y[2587]), .B(x[2587]), .Z(n9620) );
  AND U9592 ( .A(n9622), .B(n9623), .Z(n9618) );
  XNOR U9593 ( .A(y[2588]), .B(x[2588]), .Z(n9623) );
  XNOR U9594 ( .A(y[2589]), .B(x[2589]), .Z(n9622) );
  AND U9595 ( .A(n9624), .B(n9625), .Z(n9616) );
  AND U9596 ( .A(n9626), .B(n9627), .Z(n9625) );
  XNOR U9597 ( .A(y[2590]), .B(x[2590]), .Z(n9627) );
  XNOR U9598 ( .A(y[2591]), .B(x[2591]), .Z(n9626) );
  AND U9599 ( .A(n9628), .B(n9629), .Z(n9624) );
  XNOR U9600 ( .A(y[2592]), .B(x[2592]), .Z(n9629) );
  XNOR U9601 ( .A(y[2593]), .B(x[2593]), .Z(n9628) );
  AND U9602 ( .A(n9630), .B(n9631), .Z(n9566) );
  AND U9603 ( .A(n9632), .B(n9633), .Z(n9631) );
  AND U9604 ( .A(n9634), .B(n9635), .Z(n9633) );
  AND U9605 ( .A(n9636), .B(n9637), .Z(n9635) );
  AND U9606 ( .A(n9638), .B(n9639), .Z(n9637) );
  XNOR U9607 ( .A(y[2594]), .B(x[2594]), .Z(n9639) );
  XNOR U9608 ( .A(y[2595]), .B(x[2595]), .Z(n9638) );
  AND U9609 ( .A(n9640), .B(n9641), .Z(n9636) );
  XNOR U9610 ( .A(y[2596]), .B(x[2596]), .Z(n9641) );
  XNOR U9611 ( .A(y[2597]), .B(x[2597]), .Z(n9640) );
  AND U9612 ( .A(n9642), .B(n9643), .Z(n9634) );
  AND U9613 ( .A(n9644), .B(n9645), .Z(n9643) );
  XNOR U9614 ( .A(y[2598]), .B(x[2598]), .Z(n9645) );
  XNOR U9615 ( .A(y[2599]), .B(x[2599]), .Z(n9644) );
  AND U9616 ( .A(n9646), .B(n9647), .Z(n9642) );
  XNOR U9617 ( .A(y[2600]), .B(x[2600]), .Z(n9647) );
  XNOR U9618 ( .A(y[2601]), .B(x[2601]), .Z(n9646) );
  AND U9619 ( .A(n9648), .B(n9649), .Z(n9632) );
  AND U9620 ( .A(n9650), .B(n9651), .Z(n9649) );
  AND U9621 ( .A(n9652), .B(n9653), .Z(n9651) );
  XNOR U9622 ( .A(y[2602]), .B(x[2602]), .Z(n9653) );
  XNOR U9623 ( .A(y[2603]), .B(x[2603]), .Z(n9652) );
  AND U9624 ( .A(n9654), .B(n9655), .Z(n9650) );
  XNOR U9625 ( .A(y[2604]), .B(x[2604]), .Z(n9655) );
  XNOR U9626 ( .A(y[2605]), .B(x[2605]), .Z(n9654) );
  AND U9627 ( .A(n9656), .B(n9657), .Z(n9648) );
  AND U9628 ( .A(n9658), .B(n9659), .Z(n9657) );
  XNOR U9629 ( .A(y[2606]), .B(x[2606]), .Z(n9659) );
  XNOR U9630 ( .A(y[2607]), .B(x[2607]), .Z(n9658) );
  AND U9631 ( .A(n9660), .B(n9661), .Z(n9656) );
  XNOR U9632 ( .A(y[2608]), .B(x[2608]), .Z(n9661) );
  XNOR U9633 ( .A(y[2609]), .B(x[2609]), .Z(n9660) );
  AND U9634 ( .A(n9662), .B(n9663), .Z(n9630) );
  AND U9635 ( .A(n9664), .B(n9665), .Z(n9663) );
  AND U9636 ( .A(n9666), .B(n9667), .Z(n9665) );
  AND U9637 ( .A(n9668), .B(n9669), .Z(n9667) );
  XNOR U9638 ( .A(y[2610]), .B(x[2610]), .Z(n9669) );
  XNOR U9639 ( .A(y[2611]), .B(x[2611]), .Z(n9668) );
  AND U9640 ( .A(n9670), .B(n9671), .Z(n9666) );
  XNOR U9641 ( .A(y[2612]), .B(x[2612]), .Z(n9671) );
  XNOR U9642 ( .A(y[2613]), .B(x[2613]), .Z(n9670) );
  AND U9643 ( .A(n9672), .B(n9673), .Z(n9664) );
  AND U9644 ( .A(n9674), .B(n9675), .Z(n9673) );
  XNOR U9645 ( .A(y[2614]), .B(x[2614]), .Z(n9675) );
  XNOR U9646 ( .A(y[2615]), .B(x[2615]), .Z(n9674) );
  AND U9647 ( .A(n9676), .B(n9677), .Z(n9672) );
  XNOR U9648 ( .A(y[2616]), .B(x[2616]), .Z(n9677) );
  XNOR U9649 ( .A(y[2617]), .B(x[2617]), .Z(n9676) );
  AND U9650 ( .A(n9678), .B(n9679), .Z(n9662) );
  AND U9651 ( .A(n9680), .B(n9681), .Z(n9679) );
  AND U9652 ( .A(n9682), .B(n9683), .Z(n9681) );
  XNOR U9653 ( .A(y[2618]), .B(x[2618]), .Z(n9683) );
  XNOR U9654 ( .A(y[2619]), .B(x[2619]), .Z(n9682) );
  AND U9655 ( .A(n9684), .B(n9685), .Z(n9680) );
  XNOR U9656 ( .A(y[2620]), .B(x[2620]), .Z(n9685) );
  XNOR U9657 ( .A(y[2621]), .B(x[2621]), .Z(n9684) );
  AND U9658 ( .A(n9686), .B(n9687), .Z(n9678) );
  AND U9659 ( .A(n9688), .B(n9689), .Z(n9687) );
  XNOR U9660 ( .A(y[2622]), .B(x[2622]), .Z(n9689) );
  XNOR U9661 ( .A(y[2623]), .B(x[2623]), .Z(n9688) );
  AND U9662 ( .A(n9690), .B(n9691), .Z(n9686) );
  XNOR U9663 ( .A(y[2624]), .B(x[2624]), .Z(n9691) );
  XNOR U9664 ( .A(y[2625]), .B(x[2625]), .Z(n9690) );
  AND U9665 ( .A(n9692), .B(n9693), .Z(n9564) );
  AND U9666 ( .A(n9694), .B(n9695), .Z(n9693) );
  AND U9667 ( .A(n9696), .B(n9697), .Z(n9695) );
  AND U9668 ( .A(n9698), .B(n9699), .Z(n9697) );
  AND U9669 ( .A(n9700), .B(n9701), .Z(n9699) );
  AND U9670 ( .A(n9702), .B(n9703), .Z(n9701) );
  XNOR U9671 ( .A(y[2626]), .B(x[2626]), .Z(n9703) );
  XNOR U9672 ( .A(y[2627]), .B(x[2627]), .Z(n9702) );
  AND U9673 ( .A(n9704), .B(n9705), .Z(n9700) );
  XNOR U9674 ( .A(y[2628]), .B(x[2628]), .Z(n9705) );
  XNOR U9675 ( .A(y[2629]), .B(x[2629]), .Z(n9704) );
  AND U9676 ( .A(n9706), .B(n9707), .Z(n9698) );
  AND U9677 ( .A(n9708), .B(n9709), .Z(n9707) );
  XNOR U9678 ( .A(y[2630]), .B(x[2630]), .Z(n9709) );
  XNOR U9679 ( .A(y[2631]), .B(x[2631]), .Z(n9708) );
  AND U9680 ( .A(n9710), .B(n9711), .Z(n9706) );
  XNOR U9681 ( .A(y[2632]), .B(x[2632]), .Z(n9711) );
  XNOR U9682 ( .A(y[2633]), .B(x[2633]), .Z(n9710) );
  AND U9683 ( .A(n9712), .B(n9713), .Z(n9696) );
  AND U9684 ( .A(n9714), .B(n9715), .Z(n9713) );
  AND U9685 ( .A(n9716), .B(n9717), .Z(n9715) );
  XNOR U9686 ( .A(y[2634]), .B(x[2634]), .Z(n9717) );
  XNOR U9687 ( .A(y[2635]), .B(x[2635]), .Z(n9716) );
  AND U9688 ( .A(n9718), .B(n9719), .Z(n9714) );
  XNOR U9689 ( .A(y[2636]), .B(x[2636]), .Z(n9719) );
  XNOR U9690 ( .A(y[2637]), .B(x[2637]), .Z(n9718) );
  AND U9691 ( .A(n9720), .B(n9721), .Z(n9712) );
  AND U9692 ( .A(n9722), .B(n9723), .Z(n9721) );
  XNOR U9693 ( .A(y[2638]), .B(x[2638]), .Z(n9723) );
  XNOR U9694 ( .A(y[2639]), .B(x[2639]), .Z(n9722) );
  AND U9695 ( .A(n9724), .B(n9725), .Z(n9720) );
  XNOR U9696 ( .A(y[2640]), .B(x[2640]), .Z(n9725) );
  XNOR U9697 ( .A(y[2641]), .B(x[2641]), .Z(n9724) );
  AND U9698 ( .A(n9726), .B(n9727), .Z(n9694) );
  AND U9699 ( .A(n9728), .B(n9729), .Z(n9727) );
  AND U9700 ( .A(n9730), .B(n9731), .Z(n9729) );
  AND U9701 ( .A(n9732), .B(n9733), .Z(n9731) );
  XNOR U9702 ( .A(y[2642]), .B(x[2642]), .Z(n9733) );
  XNOR U9703 ( .A(y[2643]), .B(x[2643]), .Z(n9732) );
  AND U9704 ( .A(n9734), .B(n9735), .Z(n9730) );
  XNOR U9705 ( .A(y[2644]), .B(x[2644]), .Z(n9735) );
  XNOR U9706 ( .A(y[2645]), .B(x[2645]), .Z(n9734) );
  AND U9707 ( .A(n9736), .B(n9737), .Z(n9728) );
  AND U9708 ( .A(n9738), .B(n9739), .Z(n9737) );
  XNOR U9709 ( .A(y[2646]), .B(x[2646]), .Z(n9739) );
  XNOR U9710 ( .A(y[2647]), .B(x[2647]), .Z(n9738) );
  AND U9711 ( .A(n9740), .B(n9741), .Z(n9736) );
  XNOR U9712 ( .A(y[2648]), .B(x[2648]), .Z(n9741) );
  XNOR U9713 ( .A(y[2649]), .B(x[2649]), .Z(n9740) );
  AND U9714 ( .A(n9742), .B(n9743), .Z(n9726) );
  AND U9715 ( .A(n9744), .B(n9745), .Z(n9743) );
  AND U9716 ( .A(n9746), .B(n9747), .Z(n9745) );
  XNOR U9717 ( .A(y[2650]), .B(x[2650]), .Z(n9747) );
  XNOR U9718 ( .A(y[2651]), .B(x[2651]), .Z(n9746) );
  AND U9719 ( .A(n9748), .B(n9749), .Z(n9744) );
  XNOR U9720 ( .A(y[2652]), .B(x[2652]), .Z(n9749) );
  XNOR U9721 ( .A(y[2653]), .B(x[2653]), .Z(n9748) );
  AND U9722 ( .A(n9750), .B(n9751), .Z(n9742) );
  AND U9723 ( .A(n9752), .B(n9753), .Z(n9751) );
  XNOR U9724 ( .A(y[2654]), .B(x[2654]), .Z(n9753) );
  XNOR U9725 ( .A(y[2655]), .B(x[2655]), .Z(n9752) );
  AND U9726 ( .A(n9754), .B(n9755), .Z(n9750) );
  XNOR U9727 ( .A(y[2656]), .B(x[2656]), .Z(n9755) );
  XNOR U9728 ( .A(y[2657]), .B(x[2657]), .Z(n9754) );
  AND U9729 ( .A(n9756), .B(n9757), .Z(n9692) );
  AND U9730 ( .A(n9758), .B(n9759), .Z(n9757) );
  AND U9731 ( .A(n9760), .B(n9761), .Z(n9759) );
  AND U9732 ( .A(n9762), .B(n9763), .Z(n9761) );
  AND U9733 ( .A(n9764), .B(n9765), .Z(n9763) );
  XNOR U9734 ( .A(y[2658]), .B(x[2658]), .Z(n9765) );
  XNOR U9735 ( .A(y[2659]), .B(x[2659]), .Z(n9764) );
  AND U9736 ( .A(n9766), .B(n9767), .Z(n9762) );
  XNOR U9737 ( .A(y[2660]), .B(x[2660]), .Z(n9767) );
  XNOR U9738 ( .A(y[2661]), .B(x[2661]), .Z(n9766) );
  AND U9739 ( .A(n9768), .B(n9769), .Z(n9760) );
  AND U9740 ( .A(n9770), .B(n9771), .Z(n9769) );
  XNOR U9741 ( .A(y[2662]), .B(x[2662]), .Z(n9771) );
  XNOR U9742 ( .A(y[2663]), .B(x[2663]), .Z(n9770) );
  AND U9743 ( .A(n9772), .B(n9773), .Z(n9768) );
  XNOR U9744 ( .A(y[2664]), .B(x[2664]), .Z(n9773) );
  XNOR U9745 ( .A(y[2665]), .B(x[2665]), .Z(n9772) );
  AND U9746 ( .A(n9774), .B(n9775), .Z(n9758) );
  AND U9747 ( .A(n9776), .B(n9777), .Z(n9775) );
  AND U9748 ( .A(n9778), .B(n9779), .Z(n9777) );
  XNOR U9749 ( .A(y[2666]), .B(x[2666]), .Z(n9779) );
  XNOR U9750 ( .A(y[2667]), .B(x[2667]), .Z(n9778) );
  AND U9751 ( .A(n9780), .B(n9781), .Z(n9776) );
  XNOR U9752 ( .A(y[2668]), .B(x[2668]), .Z(n9781) );
  XNOR U9753 ( .A(y[2669]), .B(x[2669]), .Z(n9780) );
  AND U9754 ( .A(n9782), .B(n9783), .Z(n9774) );
  AND U9755 ( .A(n9784), .B(n9785), .Z(n9783) );
  XNOR U9756 ( .A(y[2670]), .B(x[2670]), .Z(n9785) );
  XNOR U9757 ( .A(y[2671]), .B(x[2671]), .Z(n9784) );
  AND U9758 ( .A(n9786), .B(n9787), .Z(n9782) );
  XNOR U9759 ( .A(y[2672]), .B(x[2672]), .Z(n9787) );
  XNOR U9760 ( .A(y[2673]), .B(x[2673]), .Z(n9786) );
  AND U9761 ( .A(n9788), .B(n9789), .Z(n9756) );
  AND U9762 ( .A(n9790), .B(n9791), .Z(n9789) );
  AND U9763 ( .A(n9792), .B(n9793), .Z(n9791) );
  AND U9764 ( .A(n9794), .B(n9795), .Z(n9793) );
  XNOR U9765 ( .A(y[2674]), .B(x[2674]), .Z(n9795) );
  XNOR U9766 ( .A(y[2675]), .B(x[2675]), .Z(n9794) );
  AND U9767 ( .A(n9796), .B(n9797), .Z(n9792) );
  XNOR U9768 ( .A(y[2676]), .B(x[2676]), .Z(n9797) );
  XNOR U9769 ( .A(y[2677]), .B(x[2677]), .Z(n9796) );
  AND U9770 ( .A(n9798), .B(n9799), .Z(n9790) );
  AND U9771 ( .A(n9800), .B(n9801), .Z(n9799) );
  XNOR U9772 ( .A(y[2678]), .B(x[2678]), .Z(n9801) );
  XNOR U9773 ( .A(y[2679]), .B(x[2679]), .Z(n9800) );
  AND U9774 ( .A(n9802), .B(n9803), .Z(n9798) );
  XNOR U9775 ( .A(y[2680]), .B(x[2680]), .Z(n9803) );
  XNOR U9776 ( .A(y[2681]), .B(x[2681]), .Z(n9802) );
  AND U9777 ( .A(n9804), .B(n9805), .Z(n9788) );
  AND U9778 ( .A(n9806), .B(n9807), .Z(n9805) );
  AND U9779 ( .A(n9808), .B(n9809), .Z(n9807) );
  XNOR U9780 ( .A(y[2682]), .B(x[2682]), .Z(n9809) );
  XNOR U9781 ( .A(y[2683]), .B(x[2683]), .Z(n9808) );
  AND U9782 ( .A(n9810), .B(n9811), .Z(n9806) );
  XNOR U9783 ( .A(y[2684]), .B(x[2684]), .Z(n9811) );
  XNOR U9784 ( .A(y[2685]), .B(x[2685]), .Z(n9810) );
  AND U9785 ( .A(n9812), .B(n9813), .Z(n9804) );
  AND U9786 ( .A(n9814), .B(n9815), .Z(n9813) );
  XNOR U9787 ( .A(y[2686]), .B(x[2686]), .Z(n9815) );
  XNOR U9788 ( .A(y[2687]), .B(x[2687]), .Z(n9814) );
  AND U9789 ( .A(n9816), .B(n9817), .Z(n9812) );
  XNOR U9790 ( .A(y[2688]), .B(x[2688]), .Z(n9817) );
  XNOR U9791 ( .A(y[2689]), .B(x[2689]), .Z(n9816) );
  AND U9792 ( .A(n9818), .B(n9819), .Z(n9562) );
  AND U9793 ( .A(n9820), .B(n9821), .Z(n9819) );
  AND U9794 ( .A(n9822), .B(n9823), .Z(n9821) );
  AND U9795 ( .A(n9824), .B(n9825), .Z(n9823) );
  AND U9796 ( .A(n9826), .B(n9827), .Z(n9825) );
  AND U9797 ( .A(n9828), .B(n9829), .Z(n9827) );
  AND U9798 ( .A(n9830), .B(n9831), .Z(n9829) );
  XNOR U9799 ( .A(y[2690]), .B(x[2690]), .Z(n9831) );
  XNOR U9800 ( .A(y[2691]), .B(x[2691]), .Z(n9830) );
  AND U9801 ( .A(n9832), .B(n9833), .Z(n9828) );
  XNOR U9802 ( .A(y[2692]), .B(x[2692]), .Z(n9833) );
  XNOR U9803 ( .A(y[2693]), .B(x[2693]), .Z(n9832) );
  AND U9804 ( .A(n9834), .B(n9835), .Z(n9826) );
  AND U9805 ( .A(n9836), .B(n9837), .Z(n9835) );
  XNOR U9806 ( .A(y[2694]), .B(x[2694]), .Z(n9837) );
  XNOR U9807 ( .A(y[2695]), .B(x[2695]), .Z(n9836) );
  AND U9808 ( .A(n9838), .B(n9839), .Z(n9834) );
  XNOR U9809 ( .A(y[2696]), .B(x[2696]), .Z(n9839) );
  XNOR U9810 ( .A(y[2697]), .B(x[2697]), .Z(n9838) );
  AND U9811 ( .A(n9840), .B(n9841), .Z(n9824) );
  AND U9812 ( .A(n9842), .B(n9843), .Z(n9841) );
  AND U9813 ( .A(n9844), .B(n9845), .Z(n9843) );
  XNOR U9814 ( .A(y[2698]), .B(x[2698]), .Z(n9845) );
  XNOR U9815 ( .A(y[2699]), .B(x[2699]), .Z(n9844) );
  AND U9816 ( .A(n9846), .B(n9847), .Z(n9842) );
  XNOR U9817 ( .A(y[2700]), .B(x[2700]), .Z(n9847) );
  XNOR U9818 ( .A(y[2701]), .B(x[2701]), .Z(n9846) );
  AND U9819 ( .A(n9848), .B(n9849), .Z(n9840) );
  AND U9820 ( .A(n9850), .B(n9851), .Z(n9849) );
  XNOR U9821 ( .A(y[2702]), .B(x[2702]), .Z(n9851) );
  XNOR U9822 ( .A(y[2703]), .B(x[2703]), .Z(n9850) );
  AND U9823 ( .A(n9852), .B(n9853), .Z(n9848) );
  XNOR U9824 ( .A(y[2704]), .B(x[2704]), .Z(n9853) );
  XNOR U9825 ( .A(y[2705]), .B(x[2705]), .Z(n9852) );
  AND U9826 ( .A(n9854), .B(n9855), .Z(n9822) );
  AND U9827 ( .A(n9856), .B(n9857), .Z(n9855) );
  AND U9828 ( .A(n9858), .B(n9859), .Z(n9857) );
  AND U9829 ( .A(n9860), .B(n9861), .Z(n9859) );
  XNOR U9830 ( .A(y[2706]), .B(x[2706]), .Z(n9861) );
  XNOR U9831 ( .A(y[2707]), .B(x[2707]), .Z(n9860) );
  AND U9832 ( .A(n9862), .B(n9863), .Z(n9858) );
  XNOR U9833 ( .A(y[2708]), .B(x[2708]), .Z(n9863) );
  XNOR U9834 ( .A(y[2709]), .B(x[2709]), .Z(n9862) );
  AND U9835 ( .A(n9864), .B(n9865), .Z(n9856) );
  AND U9836 ( .A(n9866), .B(n9867), .Z(n9865) );
  XNOR U9837 ( .A(y[2710]), .B(x[2710]), .Z(n9867) );
  XNOR U9838 ( .A(y[2711]), .B(x[2711]), .Z(n9866) );
  AND U9839 ( .A(n9868), .B(n9869), .Z(n9864) );
  XNOR U9840 ( .A(y[2712]), .B(x[2712]), .Z(n9869) );
  XNOR U9841 ( .A(y[2713]), .B(x[2713]), .Z(n9868) );
  AND U9842 ( .A(n9870), .B(n9871), .Z(n9854) );
  AND U9843 ( .A(n9872), .B(n9873), .Z(n9871) );
  AND U9844 ( .A(n9874), .B(n9875), .Z(n9873) );
  XNOR U9845 ( .A(y[2714]), .B(x[2714]), .Z(n9875) );
  XNOR U9846 ( .A(y[2715]), .B(x[2715]), .Z(n9874) );
  AND U9847 ( .A(n9876), .B(n9877), .Z(n9872) );
  XNOR U9848 ( .A(y[2716]), .B(x[2716]), .Z(n9877) );
  XNOR U9849 ( .A(y[2717]), .B(x[2717]), .Z(n9876) );
  AND U9850 ( .A(n9878), .B(n9879), .Z(n9870) );
  AND U9851 ( .A(n9880), .B(n9881), .Z(n9879) );
  XNOR U9852 ( .A(y[2718]), .B(x[2718]), .Z(n9881) );
  XNOR U9853 ( .A(y[2719]), .B(x[2719]), .Z(n9880) );
  AND U9854 ( .A(n9882), .B(n9883), .Z(n9878) );
  XNOR U9855 ( .A(y[2720]), .B(x[2720]), .Z(n9883) );
  XNOR U9856 ( .A(y[2721]), .B(x[2721]), .Z(n9882) );
  AND U9857 ( .A(n9884), .B(n9885), .Z(n9820) );
  AND U9858 ( .A(n9886), .B(n9887), .Z(n9885) );
  AND U9859 ( .A(n9888), .B(n9889), .Z(n9887) );
  AND U9860 ( .A(n9890), .B(n9891), .Z(n9889) );
  AND U9861 ( .A(n9892), .B(n9893), .Z(n9891) );
  XNOR U9862 ( .A(y[2722]), .B(x[2722]), .Z(n9893) );
  XNOR U9863 ( .A(y[2723]), .B(x[2723]), .Z(n9892) );
  AND U9864 ( .A(n9894), .B(n9895), .Z(n9890) );
  XNOR U9865 ( .A(y[2724]), .B(x[2724]), .Z(n9895) );
  XNOR U9866 ( .A(y[2725]), .B(x[2725]), .Z(n9894) );
  AND U9867 ( .A(n9896), .B(n9897), .Z(n9888) );
  AND U9868 ( .A(n9898), .B(n9899), .Z(n9897) );
  XNOR U9869 ( .A(y[2726]), .B(x[2726]), .Z(n9899) );
  XNOR U9870 ( .A(y[2727]), .B(x[2727]), .Z(n9898) );
  AND U9871 ( .A(n9900), .B(n9901), .Z(n9896) );
  XNOR U9872 ( .A(y[2728]), .B(x[2728]), .Z(n9901) );
  XNOR U9873 ( .A(y[2729]), .B(x[2729]), .Z(n9900) );
  AND U9874 ( .A(n9902), .B(n9903), .Z(n9886) );
  AND U9875 ( .A(n9904), .B(n9905), .Z(n9903) );
  AND U9876 ( .A(n9906), .B(n9907), .Z(n9905) );
  XNOR U9877 ( .A(y[2730]), .B(x[2730]), .Z(n9907) );
  XNOR U9878 ( .A(y[2731]), .B(x[2731]), .Z(n9906) );
  AND U9879 ( .A(n9908), .B(n9909), .Z(n9904) );
  XNOR U9880 ( .A(y[2732]), .B(x[2732]), .Z(n9909) );
  XNOR U9881 ( .A(y[2733]), .B(x[2733]), .Z(n9908) );
  AND U9882 ( .A(n9910), .B(n9911), .Z(n9902) );
  AND U9883 ( .A(n9912), .B(n9913), .Z(n9911) );
  XNOR U9884 ( .A(y[2734]), .B(x[2734]), .Z(n9913) );
  XNOR U9885 ( .A(y[2735]), .B(x[2735]), .Z(n9912) );
  AND U9886 ( .A(n9914), .B(n9915), .Z(n9910) );
  XNOR U9887 ( .A(y[2736]), .B(x[2736]), .Z(n9915) );
  XNOR U9888 ( .A(y[2737]), .B(x[2737]), .Z(n9914) );
  AND U9889 ( .A(n9916), .B(n9917), .Z(n9884) );
  AND U9890 ( .A(n9918), .B(n9919), .Z(n9917) );
  AND U9891 ( .A(n9920), .B(n9921), .Z(n9919) );
  AND U9892 ( .A(n9922), .B(n9923), .Z(n9921) );
  XNOR U9893 ( .A(y[2738]), .B(x[2738]), .Z(n9923) );
  XNOR U9894 ( .A(y[2739]), .B(x[2739]), .Z(n9922) );
  AND U9895 ( .A(n9924), .B(n9925), .Z(n9920) );
  XNOR U9896 ( .A(y[2740]), .B(x[2740]), .Z(n9925) );
  XNOR U9897 ( .A(y[2741]), .B(x[2741]), .Z(n9924) );
  AND U9898 ( .A(n9926), .B(n9927), .Z(n9918) );
  AND U9899 ( .A(n9928), .B(n9929), .Z(n9927) );
  XNOR U9900 ( .A(y[2742]), .B(x[2742]), .Z(n9929) );
  XNOR U9901 ( .A(y[2743]), .B(x[2743]), .Z(n9928) );
  AND U9902 ( .A(n9930), .B(n9931), .Z(n9926) );
  XNOR U9903 ( .A(y[2744]), .B(x[2744]), .Z(n9931) );
  XNOR U9904 ( .A(y[2745]), .B(x[2745]), .Z(n9930) );
  AND U9905 ( .A(n9932), .B(n9933), .Z(n9916) );
  AND U9906 ( .A(n9934), .B(n9935), .Z(n9933) );
  AND U9907 ( .A(n9936), .B(n9937), .Z(n9935) );
  XNOR U9908 ( .A(y[2746]), .B(x[2746]), .Z(n9937) );
  XNOR U9909 ( .A(y[2747]), .B(x[2747]), .Z(n9936) );
  AND U9910 ( .A(n9938), .B(n9939), .Z(n9934) );
  XNOR U9911 ( .A(y[2748]), .B(x[2748]), .Z(n9939) );
  XNOR U9912 ( .A(y[2749]), .B(x[2749]), .Z(n9938) );
  AND U9913 ( .A(n9940), .B(n9941), .Z(n9932) );
  AND U9914 ( .A(n9942), .B(n9943), .Z(n9941) );
  XNOR U9915 ( .A(y[2750]), .B(x[2750]), .Z(n9943) );
  XNOR U9916 ( .A(y[2751]), .B(x[2751]), .Z(n9942) );
  AND U9917 ( .A(n9944), .B(n9945), .Z(n9940) );
  XNOR U9918 ( .A(y[2752]), .B(x[2752]), .Z(n9945) );
  XNOR U9919 ( .A(y[2753]), .B(x[2753]), .Z(n9944) );
  AND U9920 ( .A(n9946), .B(n9947), .Z(n9818) );
  AND U9921 ( .A(n9948), .B(n9949), .Z(n9947) );
  AND U9922 ( .A(n9950), .B(n9951), .Z(n9949) );
  AND U9923 ( .A(n9952), .B(n9953), .Z(n9951) );
  AND U9924 ( .A(n9954), .B(n9955), .Z(n9953) );
  AND U9925 ( .A(n9956), .B(n9957), .Z(n9955) );
  XNOR U9926 ( .A(y[2754]), .B(x[2754]), .Z(n9957) );
  XNOR U9927 ( .A(y[2755]), .B(x[2755]), .Z(n9956) );
  AND U9928 ( .A(n9958), .B(n9959), .Z(n9954) );
  XNOR U9929 ( .A(y[2756]), .B(x[2756]), .Z(n9959) );
  XNOR U9930 ( .A(y[2757]), .B(x[2757]), .Z(n9958) );
  AND U9931 ( .A(n9960), .B(n9961), .Z(n9952) );
  AND U9932 ( .A(n9962), .B(n9963), .Z(n9961) );
  XNOR U9933 ( .A(y[2758]), .B(x[2758]), .Z(n9963) );
  XNOR U9934 ( .A(y[2759]), .B(x[2759]), .Z(n9962) );
  AND U9935 ( .A(n9964), .B(n9965), .Z(n9960) );
  XNOR U9936 ( .A(y[2760]), .B(x[2760]), .Z(n9965) );
  XNOR U9937 ( .A(y[2761]), .B(x[2761]), .Z(n9964) );
  AND U9938 ( .A(n9966), .B(n9967), .Z(n9950) );
  AND U9939 ( .A(n9968), .B(n9969), .Z(n9967) );
  AND U9940 ( .A(n9970), .B(n9971), .Z(n9969) );
  XNOR U9941 ( .A(y[2762]), .B(x[2762]), .Z(n9971) );
  XNOR U9942 ( .A(y[2763]), .B(x[2763]), .Z(n9970) );
  AND U9943 ( .A(n9972), .B(n9973), .Z(n9968) );
  XNOR U9944 ( .A(y[2764]), .B(x[2764]), .Z(n9973) );
  XNOR U9945 ( .A(y[2765]), .B(x[2765]), .Z(n9972) );
  AND U9946 ( .A(n9974), .B(n9975), .Z(n9966) );
  AND U9947 ( .A(n9976), .B(n9977), .Z(n9975) );
  XNOR U9948 ( .A(y[2766]), .B(x[2766]), .Z(n9977) );
  XNOR U9949 ( .A(y[2767]), .B(x[2767]), .Z(n9976) );
  AND U9950 ( .A(n9978), .B(n9979), .Z(n9974) );
  XNOR U9951 ( .A(y[2768]), .B(x[2768]), .Z(n9979) );
  XNOR U9952 ( .A(y[2769]), .B(x[2769]), .Z(n9978) );
  AND U9953 ( .A(n9980), .B(n9981), .Z(n9948) );
  AND U9954 ( .A(n9982), .B(n9983), .Z(n9981) );
  AND U9955 ( .A(n9984), .B(n9985), .Z(n9983) );
  AND U9956 ( .A(n9986), .B(n9987), .Z(n9985) );
  XNOR U9957 ( .A(y[2770]), .B(x[2770]), .Z(n9987) );
  XNOR U9958 ( .A(y[2771]), .B(x[2771]), .Z(n9986) );
  AND U9959 ( .A(n9988), .B(n9989), .Z(n9984) );
  XNOR U9960 ( .A(y[2772]), .B(x[2772]), .Z(n9989) );
  XNOR U9961 ( .A(y[2773]), .B(x[2773]), .Z(n9988) );
  AND U9962 ( .A(n9990), .B(n9991), .Z(n9982) );
  AND U9963 ( .A(n9992), .B(n9993), .Z(n9991) );
  XNOR U9964 ( .A(y[2774]), .B(x[2774]), .Z(n9993) );
  XNOR U9965 ( .A(y[2775]), .B(x[2775]), .Z(n9992) );
  AND U9966 ( .A(n9994), .B(n9995), .Z(n9990) );
  XNOR U9967 ( .A(y[2776]), .B(x[2776]), .Z(n9995) );
  XNOR U9968 ( .A(y[2777]), .B(x[2777]), .Z(n9994) );
  AND U9969 ( .A(n9996), .B(n9997), .Z(n9980) );
  AND U9970 ( .A(n9998), .B(n9999), .Z(n9997) );
  AND U9971 ( .A(n10000), .B(n10001), .Z(n9999) );
  XNOR U9972 ( .A(y[2778]), .B(x[2778]), .Z(n10001) );
  XNOR U9973 ( .A(y[2779]), .B(x[2779]), .Z(n10000) );
  AND U9974 ( .A(n10002), .B(n10003), .Z(n9998) );
  XNOR U9975 ( .A(y[2780]), .B(x[2780]), .Z(n10003) );
  XNOR U9976 ( .A(y[2781]), .B(x[2781]), .Z(n10002) );
  AND U9977 ( .A(n10004), .B(n10005), .Z(n9996) );
  AND U9978 ( .A(n10006), .B(n10007), .Z(n10005) );
  XNOR U9979 ( .A(y[2782]), .B(x[2782]), .Z(n10007) );
  XNOR U9980 ( .A(y[2783]), .B(x[2783]), .Z(n10006) );
  AND U9981 ( .A(n10008), .B(n10009), .Z(n10004) );
  XNOR U9982 ( .A(y[2784]), .B(x[2784]), .Z(n10009) );
  XNOR U9983 ( .A(y[2785]), .B(x[2785]), .Z(n10008) );
  AND U9984 ( .A(n10010), .B(n10011), .Z(n9946) );
  AND U9985 ( .A(n10012), .B(n10013), .Z(n10011) );
  AND U9986 ( .A(n10014), .B(n10015), .Z(n10013) );
  AND U9987 ( .A(n10016), .B(n10017), .Z(n10015) );
  AND U9988 ( .A(n10018), .B(n10019), .Z(n10017) );
  XNOR U9989 ( .A(y[2786]), .B(x[2786]), .Z(n10019) );
  XNOR U9990 ( .A(y[2787]), .B(x[2787]), .Z(n10018) );
  AND U9991 ( .A(n10020), .B(n10021), .Z(n10016) );
  XNOR U9992 ( .A(y[2788]), .B(x[2788]), .Z(n10021) );
  XNOR U9993 ( .A(y[2789]), .B(x[2789]), .Z(n10020) );
  AND U9994 ( .A(n10022), .B(n10023), .Z(n10014) );
  AND U9995 ( .A(n10024), .B(n10025), .Z(n10023) );
  XNOR U9996 ( .A(y[2790]), .B(x[2790]), .Z(n10025) );
  XNOR U9997 ( .A(y[2791]), .B(x[2791]), .Z(n10024) );
  AND U9998 ( .A(n10026), .B(n10027), .Z(n10022) );
  XNOR U9999 ( .A(y[2792]), .B(x[2792]), .Z(n10027) );
  XNOR U10000 ( .A(y[2793]), .B(x[2793]), .Z(n10026) );
  AND U10001 ( .A(n10028), .B(n10029), .Z(n10012) );
  AND U10002 ( .A(n10030), .B(n10031), .Z(n10029) );
  AND U10003 ( .A(n10032), .B(n10033), .Z(n10031) );
  XNOR U10004 ( .A(y[2794]), .B(x[2794]), .Z(n10033) );
  XNOR U10005 ( .A(y[2795]), .B(x[2795]), .Z(n10032) );
  AND U10006 ( .A(n10034), .B(n10035), .Z(n10030) );
  XNOR U10007 ( .A(y[2796]), .B(x[2796]), .Z(n10035) );
  XNOR U10008 ( .A(y[2797]), .B(x[2797]), .Z(n10034) );
  AND U10009 ( .A(n10036), .B(n10037), .Z(n10028) );
  AND U10010 ( .A(n10038), .B(n10039), .Z(n10037) );
  XNOR U10011 ( .A(y[2798]), .B(x[2798]), .Z(n10039) );
  XNOR U10012 ( .A(y[2799]), .B(x[2799]), .Z(n10038) );
  AND U10013 ( .A(n10040), .B(n10041), .Z(n10036) );
  XNOR U10014 ( .A(y[2800]), .B(x[2800]), .Z(n10041) );
  XNOR U10015 ( .A(y[2801]), .B(x[2801]), .Z(n10040) );
  AND U10016 ( .A(n10042), .B(n10043), .Z(n10010) );
  AND U10017 ( .A(n10044), .B(n10045), .Z(n10043) );
  AND U10018 ( .A(n10046), .B(n10047), .Z(n10045) );
  AND U10019 ( .A(n10048), .B(n10049), .Z(n10047) );
  XNOR U10020 ( .A(y[2802]), .B(x[2802]), .Z(n10049) );
  XNOR U10021 ( .A(y[2803]), .B(x[2803]), .Z(n10048) );
  AND U10022 ( .A(n10050), .B(n10051), .Z(n10046) );
  XNOR U10023 ( .A(y[2804]), .B(x[2804]), .Z(n10051) );
  XNOR U10024 ( .A(y[2805]), .B(x[2805]), .Z(n10050) );
  AND U10025 ( .A(n10052), .B(n10053), .Z(n10044) );
  AND U10026 ( .A(n10054), .B(n10055), .Z(n10053) );
  XNOR U10027 ( .A(y[2806]), .B(x[2806]), .Z(n10055) );
  XNOR U10028 ( .A(y[2807]), .B(x[2807]), .Z(n10054) );
  AND U10029 ( .A(n10056), .B(n10057), .Z(n10052) );
  XNOR U10030 ( .A(y[2808]), .B(x[2808]), .Z(n10057) );
  XNOR U10031 ( .A(y[2809]), .B(x[2809]), .Z(n10056) );
  AND U10032 ( .A(n10058), .B(n10059), .Z(n10042) );
  AND U10033 ( .A(n10060), .B(n10061), .Z(n10059) );
  AND U10034 ( .A(n10062), .B(n10063), .Z(n10061) );
  XNOR U10035 ( .A(y[2810]), .B(x[2810]), .Z(n10063) );
  XNOR U10036 ( .A(y[2811]), .B(x[2811]), .Z(n10062) );
  AND U10037 ( .A(n10064), .B(n10065), .Z(n10060) );
  XNOR U10038 ( .A(y[2812]), .B(x[2812]), .Z(n10065) );
  XNOR U10039 ( .A(y[2813]), .B(x[2813]), .Z(n10064) );
  AND U10040 ( .A(n10066), .B(n10067), .Z(n10058) );
  AND U10041 ( .A(n10068), .B(n10069), .Z(n10067) );
  XNOR U10042 ( .A(y[2814]), .B(x[2814]), .Z(n10069) );
  XNOR U10043 ( .A(y[2815]), .B(x[2815]), .Z(n10068) );
  AND U10044 ( .A(n10070), .B(n10071), .Z(n10066) );
  XNOR U10045 ( .A(y[2816]), .B(x[2816]), .Z(n10071) );
  XNOR U10046 ( .A(y[2817]), .B(x[2817]), .Z(n10070) );
  AND U10047 ( .A(n10072), .B(n10073), .Z(n8664) );
  AND U10048 ( .A(n10074), .B(n10075), .Z(n10073) );
  AND U10049 ( .A(n10076), .B(n10077), .Z(n10075) );
  AND U10050 ( .A(n10078), .B(n10079), .Z(n10077) );
  AND U10051 ( .A(n10080), .B(n10081), .Z(n10079) );
  AND U10052 ( .A(n10082), .B(n10083), .Z(n10081) );
  AND U10053 ( .A(n10084), .B(n10085), .Z(n10083) );
  AND U10054 ( .A(n10086), .B(n10087), .Z(n10085) );
  AND U10055 ( .A(n10088), .B(n10089), .Z(n10087) );
  XNOR U10056 ( .A(y[3330]), .B(x[3330]), .Z(n10089) );
  XNOR U10057 ( .A(y[3331]), .B(x[3331]), .Z(n10088) );
  AND U10058 ( .A(n10090), .B(n10091), .Z(n10086) );
  XNOR U10059 ( .A(y[3332]), .B(x[3332]), .Z(n10091) );
  XNOR U10060 ( .A(y[3333]), .B(x[3333]), .Z(n10090) );
  AND U10061 ( .A(n10092), .B(n10093), .Z(n10084) );
  AND U10062 ( .A(n10094), .B(n10095), .Z(n10093) );
  XNOR U10063 ( .A(y[3334]), .B(x[3334]), .Z(n10095) );
  XNOR U10064 ( .A(y[3335]), .B(x[3335]), .Z(n10094) );
  AND U10065 ( .A(n10096), .B(n10097), .Z(n10092) );
  XNOR U10066 ( .A(y[3336]), .B(x[3336]), .Z(n10097) );
  XNOR U10067 ( .A(y[3337]), .B(x[3337]), .Z(n10096) );
  AND U10068 ( .A(n10098), .B(n10099), .Z(n10082) );
  AND U10069 ( .A(n10100), .B(n10101), .Z(n10099) );
  AND U10070 ( .A(n10102), .B(n10103), .Z(n10101) );
  XNOR U10071 ( .A(y[3338]), .B(x[3338]), .Z(n10103) );
  XNOR U10072 ( .A(y[3339]), .B(x[3339]), .Z(n10102) );
  AND U10073 ( .A(n10104), .B(n10105), .Z(n10100) );
  XNOR U10074 ( .A(y[3340]), .B(x[3340]), .Z(n10105) );
  XNOR U10075 ( .A(y[3341]), .B(x[3341]), .Z(n10104) );
  AND U10076 ( .A(n10106), .B(n10107), .Z(n10098) );
  AND U10077 ( .A(n10108), .B(n10109), .Z(n10107) );
  XNOR U10078 ( .A(y[3342]), .B(x[3342]), .Z(n10109) );
  XNOR U10079 ( .A(y[3343]), .B(x[3343]), .Z(n10108) );
  AND U10080 ( .A(n10110), .B(n10111), .Z(n10106) );
  XNOR U10081 ( .A(y[3344]), .B(x[3344]), .Z(n10111) );
  XNOR U10082 ( .A(y[3345]), .B(x[3345]), .Z(n10110) );
  AND U10083 ( .A(n10112), .B(n10113), .Z(n10080) );
  AND U10084 ( .A(n10114), .B(n10115), .Z(n10113) );
  AND U10085 ( .A(n10116), .B(n10117), .Z(n10115) );
  AND U10086 ( .A(n10118), .B(n10119), .Z(n10117) );
  XNOR U10087 ( .A(y[3346]), .B(x[3346]), .Z(n10119) );
  XNOR U10088 ( .A(y[3347]), .B(x[3347]), .Z(n10118) );
  AND U10089 ( .A(n10120), .B(n10121), .Z(n10116) );
  XNOR U10090 ( .A(y[3348]), .B(x[3348]), .Z(n10121) );
  XNOR U10091 ( .A(y[3349]), .B(x[3349]), .Z(n10120) );
  AND U10092 ( .A(n10122), .B(n10123), .Z(n10114) );
  AND U10093 ( .A(n10124), .B(n10125), .Z(n10123) );
  XNOR U10094 ( .A(y[3350]), .B(x[3350]), .Z(n10125) );
  XNOR U10095 ( .A(y[3351]), .B(x[3351]), .Z(n10124) );
  AND U10096 ( .A(n10126), .B(n10127), .Z(n10122) );
  XNOR U10097 ( .A(y[3352]), .B(x[3352]), .Z(n10127) );
  XNOR U10098 ( .A(y[3353]), .B(x[3353]), .Z(n10126) );
  AND U10099 ( .A(n10128), .B(n10129), .Z(n10112) );
  AND U10100 ( .A(n10130), .B(n10131), .Z(n10129) );
  AND U10101 ( .A(n10132), .B(n10133), .Z(n10131) );
  XNOR U10102 ( .A(y[3354]), .B(x[3354]), .Z(n10133) );
  XNOR U10103 ( .A(y[3355]), .B(x[3355]), .Z(n10132) );
  AND U10104 ( .A(n10134), .B(n10135), .Z(n10130) );
  XNOR U10105 ( .A(y[3356]), .B(x[3356]), .Z(n10135) );
  XNOR U10106 ( .A(y[3357]), .B(x[3357]), .Z(n10134) );
  AND U10107 ( .A(n10136), .B(n10137), .Z(n10128) );
  AND U10108 ( .A(n10138), .B(n10139), .Z(n10137) );
  XNOR U10109 ( .A(y[3358]), .B(x[3358]), .Z(n10139) );
  XNOR U10110 ( .A(y[3359]), .B(x[3359]), .Z(n10138) );
  AND U10111 ( .A(n10140), .B(n10141), .Z(n10136) );
  XNOR U10112 ( .A(y[3360]), .B(x[3360]), .Z(n10141) );
  XNOR U10113 ( .A(y[3361]), .B(x[3361]), .Z(n10140) );
  AND U10114 ( .A(n10142), .B(n10143), .Z(n10078) );
  AND U10115 ( .A(n10144), .B(n10145), .Z(n10143) );
  AND U10116 ( .A(n10146), .B(n10147), .Z(n10145) );
  AND U10117 ( .A(n10148), .B(n10149), .Z(n10147) );
  AND U10118 ( .A(n10150), .B(n10151), .Z(n10149) );
  XNOR U10119 ( .A(y[3362]), .B(x[3362]), .Z(n10151) );
  XNOR U10120 ( .A(y[3363]), .B(x[3363]), .Z(n10150) );
  AND U10121 ( .A(n10152), .B(n10153), .Z(n10148) );
  XNOR U10122 ( .A(y[3364]), .B(x[3364]), .Z(n10153) );
  XNOR U10123 ( .A(y[3365]), .B(x[3365]), .Z(n10152) );
  AND U10124 ( .A(n10154), .B(n10155), .Z(n10146) );
  AND U10125 ( .A(n10156), .B(n10157), .Z(n10155) );
  XNOR U10126 ( .A(y[3366]), .B(x[3366]), .Z(n10157) );
  XNOR U10127 ( .A(y[3367]), .B(x[3367]), .Z(n10156) );
  AND U10128 ( .A(n10158), .B(n10159), .Z(n10154) );
  XNOR U10129 ( .A(y[3368]), .B(x[3368]), .Z(n10159) );
  XNOR U10130 ( .A(y[3369]), .B(x[3369]), .Z(n10158) );
  AND U10131 ( .A(n10160), .B(n10161), .Z(n10144) );
  AND U10132 ( .A(n10162), .B(n10163), .Z(n10161) );
  AND U10133 ( .A(n10164), .B(n10165), .Z(n10163) );
  XNOR U10134 ( .A(y[3370]), .B(x[3370]), .Z(n10165) );
  XNOR U10135 ( .A(y[3371]), .B(x[3371]), .Z(n10164) );
  AND U10136 ( .A(n10166), .B(n10167), .Z(n10162) );
  XNOR U10137 ( .A(y[3372]), .B(x[3372]), .Z(n10167) );
  XNOR U10138 ( .A(y[3373]), .B(x[3373]), .Z(n10166) );
  AND U10139 ( .A(n10168), .B(n10169), .Z(n10160) );
  AND U10140 ( .A(n10170), .B(n10171), .Z(n10169) );
  XNOR U10141 ( .A(y[3374]), .B(x[3374]), .Z(n10171) );
  XNOR U10142 ( .A(y[3375]), .B(x[3375]), .Z(n10170) );
  AND U10143 ( .A(n10172), .B(n10173), .Z(n10168) );
  XNOR U10144 ( .A(y[3376]), .B(x[3376]), .Z(n10173) );
  XNOR U10145 ( .A(y[3377]), .B(x[3377]), .Z(n10172) );
  AND U10146 ( .A(n10174), .B(n10175), .Z(n10142) );
  AND U10147 ( .A(n10176), .B(n10177), .Z(n10175) );
  AND U10148 ( .A(n10178), .B(n10179), .Z(n10177) );
  AND U10149 ( .A(n10180), .B(n10181), .Z(n10179) );
  XNOR U10150 ( .A(y[3378]), .B(x[3378]), .Z(n10181) );
  XNOR U10151 ( .A(y[3379]), .B(x[3379]), .Z(n10180) );
  AND U10152 ( .A(n10182), .B(n10183), .Z(n10178) );
  XNOR U10153 ( .A(y[3380]), .B(x[3380]), .Z(n10183) );
  XNOR U10154 ( .A(y[3381]), .B(x[3381]), .Z(n10182) );
  AND U10155 ( .A(n10184), .B(n10185), .Z(n10176) );
  AND U10156 ( .A(n10186), .B(n10187), .Z(n10185) );
  XNOR U10157 ( .A(y[3382]), .B(x[3382]), .Z(n10187) );
  XNOR U10158 ( .A(y[3383]), .B(x[3383]), .Z(n10186) );
  AND U10159 ( .A(n10188), .B(n10189), .Z(n10184) );
  XNOR U10160 ( .A(y[3384]), .B(x[3384]), .Z(n10189) );
  XNOR U10161 ( .A(y[3385]), .B(x[3385]), .Z(n10188) );
  AND U10162 ( .A(n10190), .B(n10191), .Z(n10174) );
  AND U10163 ( .A(n10192), .B(n10193), .Z(n10191) );
  AND U10164 ( .A(n10194), .B(n10195), .Z(n10193) );
  XNOR U10165 ( .A(y[3386]), .B(x[3386]), .Z(n10195) );
  XNOR U10166 ( .A(y[3387]), .B(x[3387]), .Z(n10194) );
  AND U10167 ( .A(n10196), .B(n10197), .Z(n10192) );
  XNOR U10168 ( .A(y[3388]), .B(x[3388]), .Z(n10197) );
  XNOR U10169 ( .A(y[3389]), .B(x[3389]), .Z(n10196) );
  AND U10170 ( .A(n10198), .B(n10199), .Z(n10190) );
  AND U10171 ( .A(n10200), .B(n10201), .Z(n10199) );
  XNOR U10172 ( .A(y[3390]), .B(x[3390]), .Z(n10201) );
  XNOR U10173 ( .A(y[3391]), .B(x[3391]), .Z(n10200) );
  AND U10174 ( .A(n10202), .B(n10203), .Z(n10198) );
  XNOR U10175 ( .A(y[3392]), .B(x[3392]), .Z(n10203) );
  XNOR U10176 ( .A(y[3393]), .B(x[3393]), .Z(n10202) );
  AND U10177 ( .A(n10204), .B(n10205), .Z(n10076) );
  AND U10178 ( .A(n10206), .B(n10207), .Z(n10205) );
  AND U10179 ( .A(n10208), .B(n10209), .Z(n10207) );
  AND U10180 ( .A(n10210), .B(n10211), .Z(n10209) );
  AND U10181 ( .A(n10212), .B(n10213), .Z(n10211) );
  AND U10182 ( .A(n10214), .B(n10215), .Z(n10213) );
  XNOR U10183 ( .A(y[3394]), .B(x[3394]), .Z(n10215) );
  XNOR U10184 ( .A(y[3395]), .B(x[3395]), .Z(n10214) );
  AND U10185 ( .A(n10216), .B(n10217), .Z(n10212) );
  XNOR U10186 ( .A(y[3396]), .B(x[3396]), .Z(n10217) );
  XNOR U10187 ( .A(y[3397]), .B(x[3397]), .Z(n10216) );
  AND U10188 ( .A(n10218), .B(n10219), .Z(n10210) );
  AND U10189 ( .A(n10220), .B(n10221), .Z(n10219) );
  XNOR U10190 ( .A(y[3398]), .B(x[3398]), .Z(n10221) );
  XNOR U10191 ( .A(y[3399]), .B(x[3399]), .Z(n10220) );
  AND U10192 ( .A(n10222), .B(n10223), .Z(n10218) );
  XNOR U10193 ( .A(y[3400]), .B(x[3400]), .Z(n10223) );
  XNOR U10194 ( .A(y[3401]), .B(x[3401]), .Z(n10222) );
  AND U10195 ( .A(n10224), .B(n10225), .Z(n10208) );
  AND U10196 ( .A(n10226), .B(n10227), .Z(n10225) );
  AND U10197 ( .A(n10228), .B(n10229), .Z(n10227) );
  XNOR U10198 ( .A(y[3402]), .B(x[3402]), .Z(n10229) );
  XNOR U10199 ( .A(y[3403]), .B(x[3403]), .Z(n10228) );
  AND U10200 ( .A(n10230), .B(n10231), .Z(n10226) );
  XNOR U10201 ( .A(y[3404]), .B(x[3404]), .Z(n10231) );
  XNOR U10202 ( .A(y[3405]), .B(x[3405]), .Z(n10230) );
  AND U10203 ( .A(n10232), .B(n10233), .Z(n10224) );
  AND U10204 ( .A(n10234), .B(n10235), .Z(n10233) );
  XNOR U10205 ( .A(y[3406]), .B(x[3406]), .Z(n10235) );
  XNOR U10206 ( .A(y[3407]), .B(x[3407]), .Z(n10234) );
  AND U10207 ( .A(n10236), .B(n10237), .Z(n10232) );
  XNOR U10208 ( .A(y[3408]), .B(x[3408]), .Z(n10237) );
  XNOR U10209 ( .A(y[3409]), .B(x[3409]), .Z(n10236) );
  AND U10210 ( .A(n10238), .B(n10239), .Z(n10206) );
  AND U10211 ( .A(n10240), .B(n10241), .Z(n10239) );
  AND U10212 ( .A(n10242), .B(n10243), .Z(n10241) );
  AND U10213 ( .A(n10244), .B(n10245), .Z(n10243) );
  XNOR U10214 ( .A(y[3410]), .B(x[3410]), .Z(n10245) );
  XNOR U10215 ( .A(y[3411]), .B(x[3411]), .Z(n10244) );
  AND U10216 ( .A(n10246), .B(n10247), .Z(n10242) );
  XNOR U10217 ( .A(y[3412]), .B(x[3412]), .Z(n10247) );
  XNOR U10218 ( .A(y[3413]), .B(x[3413]), .Z(n10246) );
  AND U10219 ( .A(n10248), .B(n10249), .Z(n10240) );
  AND U10220 ( .A(n10250), .B(n10251), .Z(n10249) );
  XNOR U10221 ( .A(y[3414]), .B(x[3414]), .Z(n10251) );
  XNOR U10222 ( .A(y[3415]), .B(x[3415]), .Z(n10250) );
  AND U10223 ( .A(n10252), .B(n10253), .Z(n10248) );
  XNOR U10224 ( .A(y[3416]), .B(x[3416]), .Z(n10253) );
  XNOR U10225 ( .A(y[3417]), .B(x[3417]), .Z(n10252) );
  AND U10226 ( .A(n10254), .B(n10255), .Z(n10238) );
  AND U10227 ( .A(n10256), .B(n10257), .Z(n10255) );
  AND U10228 ( .A(n10258), .B(n10259), .Z(n10257) );
  XNOR U10229 ( .A(y[3418]), .B(x[3418]), .Z(n10259) );
  XNOR U10230 ( .A(y[3419]), .B(x[3419]), .Z(n10258) );
  AND U10231 ( .A(n10260), .B(n10261), .Z(n10256) );
  XNOR U10232 ( .A(y[3420]), .B(x[3420]), .Z(n10261) );
  XNOR U10233 ( .A(y[3421]), .B(x[3421]), .Z(n10260) );
  AND U10234 ( .A(n10262), .B(n10263), .Z(n10254) );
  AND U10235 ( .A(n10264), .B(n10265), .Z(n10263) );
  XNOR U10236 ( .A(y[3422]), .B(x[3422]), .Z(n10265) );
  XNOR U10237 ( .A(y[3423]), .B(x[3423]), .Z(n10264) );
  AND U10238 ( .A(n10266), .B(n10267), .Z(n10262) );
  XNOR U10239 ( .A(y[3424]), .B(x[3424]), .Z(n10267) );
  XNOR U10240 ( .A(y[3425]), .B(x[3425]), .Z(n10266) );
  AND U10241 ( .A(n10268), .B(n10269), .Z(n10204) );
  AND U10242 ( .A(n10270), .B(n10271), .Z(n10269) );
  AND U10243 ( .A(n10272), .B(n10273), .Z(n10271) );
  AND U10244 ( .A(n10274), .B(n10275), .Z(n10273) );
  AND U10245 ( .A(n10276), .B(n10277), .Z(n10275) );
  XNOR U10246 ( .A(y[3426]), .B(x[3426]), .Z(n10277) );
  XNOR U10247 ( .A(y[3427]), .B(x[3427]), .Z(n10276) );
  AND U10248 ( .A(n10278), .B(n10279), .Z(n10274) );
  XNOR U10249 ( .A(y[3428]), .B(x[3428]), .Z(n10279) );
  XNOR U10250 ( .A(y[3429]), .B(x[3429]), .Z(n10278) );
  AND U10251 ( .A(n10280), .B(n10281), .Z(n10272) );
  AND U10252 ( .A(n10282), .B(n10283), .Z(n10281) );
  XNOR U10253 ( .A(y[3430]), .B(x[3430]), .Z(n10283) );
  XNOR U10254 ( .A(y[3431]), .B(x[3431]), .Z(n10282) );
  AND U10255 ( .A(n10284), .B(n10285), .Z(n10280) );
  XNOR U10256 ( .A(y[3432]), .B(x[3432]), .Z(n10285) );
  XNOR U10257 ( .A(y[3433]), .B(x[3433]), .Z(n10284) );
  AND U10258 ( .A(n10286), .B(n10287), .Z(n10270) );
  AND U10259 ( .A(n10288), .B(n10289), .Z(n10287) );
  AND U10260 ( .A(n10290), .B(n10291), .Z(n10289) );
  XNOR U10261 ( .A(y[3434]), .B(x[3434]), .Z(n10291) );
  XNOR U10262 ( .A(y[3435]), .B(x[3435]), .Z(n10290) );
  AND U10263 ( .A(n10292), .B(n10293), .Z(n10288) );
  XNOR U10264 ( .A(y[3436]), .B(x[3436]), .Z(n10293) );
  XNOR U10265 ( .A(y[3437]), .B(x[3437]), .Z(n10292) );
  AND U10266 ( .A(n10294), .B(n10295), .Z(n10286) );
  AND U10267 ( .A(n10296), .B(n10297), .Z(n10295) );
  XNOR U10268 ( .A(y[3438]), .B(x[3438]), .Z(n10297) );
  XNOR U10269 ( .A(y[3439]), .B(x[3439]), .Z(n10296) );
  AND U10270 ( .A(n10298), .B(n10299), .Z(n10294) );
  XNOR U10271 ( .A(y[3440]), .B(x[3440]), .Z(n10299) );
  XNOR U10272 ( .A(y[3441]), .B(x[3441]), .Z(n10298) );
  AND U10273 ( .A(n10300), .B(n10301), .Z(n10268) );
  AND U10274 ( .A(n10302), .B(n10303), .Z(n10301) );
  AND U10275 ( .A(n10304), .B(n10305), .Z(n10303) );
  AND U10276 ( .A(n10306), .B(n10307), .Z(n10305) );
  XNOR U10277 ( .A(y[3442]), .B(x[3442]), .Z(n10307) );
  XNOR U10278 ( .A(y[3443]), .B(x[3443]), .Z(n10306) );
  AND U10279 ( .A(n10308), .B(n10309), .Z(n10304) );
  XNOR U10280 ( .A(y[3444]), .B(x[3444]), .Z(n10309) );
  XNOR U10281 ( .A(y[3445]), .B(x[3445]), .Z(n10308) );
  AND U10282 ( .A(n10310), .B(n10311), .Z(n10302) );
  AND U10283 ( .A(n10312), .B(n10313), .Z(n10311) );
  XNOR U10284 ( .A(y[3446]), .B(x[3446]), .Z(n10313) );
  XNOR U10285 ( .A(y[3447]), .B(x[3447]), .Z(n10312) );
  AND U10286 ( .A(n10314), .B(n10315), .Z(n10310) );
  XNOR U10287 ( .A(y[3448]), .B(x[3448]), .Z(n10315) );
  XNOR U10288 ( .A(y[3449]), .B(x[3449]), .Z(n10314) );
  AND U10289 ( .A(n10316), .B(n10317), .Z(n10300) );
  AND U10290 ( .A(n10318), .B(n10319), .Z(n10317) );
  AND U10291 ( .A(n10320), .B(n10321), .Z(n10319) );
  XNOR U10292 ( .A(y[3450]), .B(x[3450]), .Z(n10321) );
  XNOR U10293 ( .A(y[3451]), .B(x[3451]), .Z(n10320) );
  AND U10294 ( .A(n10322), .B(n10323), .Z(n10318) );
  XNOR U10295 ( .A(y[3452]), .B(x[3452]), .Z(n10323) );
  XNOR U10296 ( .A(y[3453]), .B(x[3453]), .Z(n10322) );
  AND U10297 ( .A(n10324), .B(n10325), .Z(n10316) );
  AND U10298 ( .A(n10326), .B(n10327), .Z(n10325) );
  XNOR U10299 ( .A(y[3454]), .B(x[3454]), .Z(n10327) );
  XNOR U10300 ( .A(y[3455]), .B(x[3455]), .Z(n10326) );
  AND U10301 ( .A(n10328), .B(n10329), .Z(n10324) );
  XNOR U10302 ( .A(y[3456]), .B(x[3456]), .Z(n10329) );
  XNOR U10303 ( .A(y[3457]), .B(x[3457]), .Z(n10328) );
  AND U10304 ( .A(n10330), .B(n10331), .Z(n10074) );
  AND U10305 ( .A(n10332), .B(n10333), .Z(n10331) );
  AND U10306 ( .A(n10334), .B(n10335), .Z(n10333) );
  AND U10307 ( .A(n10336), .B(n10337), .Z(n10335) );
  AND U10308 ( .A(n10338), .B(n10339), .Z(n10337) );
  AND U10309 ( .A(n10340), .B(n10341), .Z(n10339) );
  AND U10310 ( .A(n10342), .B(n10343), .Z(n10341) );
  AND U10311 ( .A(n10344), .B(n10345), .Z(n10343) );
  XNOR U10312 ( .A(y[3074]), .B(x[3074]), .Z(n10345) );
  XNOR U10313 ( .A(y[3077]), .B(x[3077]), .Z(n10344) );
  AND U10314 ( .A(n10346), .B(n10347), .Z(n10342) );
  XNOR U10315 ( .A(y[3075]), .B(x[3075]), .Z(n10347) );
  XNOR U10316 ( .A(y[3076]), .B(x[3076]), .Z(n10346) );
  AND U10317 ( .A(n10348), .B(n10349), .Z(n10340) );
  AND U10318 ( .A(n10350), .B(n10351), .Z(n10349) );
  XNOR U10319 ( .A(y[3078]), .B(x[3078]), .Z(n10351) );
  XNOR U10320 ( .A(y[3079]), .B(x[3079]), .Z(n10350) );
  AND U10321 ( .A(n10352), .B(n10353), .Z(n10348) );
  XNOR U10322 ( .A(y[3080]), .B(x[3080]), .Z(n10353) );
  XNOR U10323 ( .A(y[3081]), .B(x[3081]), .Z(n10352) );
  AND U10324 ( .A(n10354), .B(n10355), .Z(n10338) );
  AND U10325 ( .A(n10356), .B(n10357), .Z(n10355) );
  AND U10326 ( .A(n10358), .B(n10359), .Z(n10357) );
  XNOR U10327 ( .A(y[3082]), .B(x[3082]), .Z(n10359) );
  XNOR U10328 ( .A(y[3083]), .B(x[3083]), .Z(n10358) );
  AND U10329 ( .A(n10360), .B(n10361), .Z(n10356) );
  XNOR U10330 ( .A(y[3084]), .B(x[3084]), .Z(n10361) );
  XNOR U10331 ( .A(y[3085]), .B(x[3085]), .Z(n10360) );
  AND U10332 ( .A(n10362), .B(n10363), .Z(n10354) );
  AND U10333 ( .A(n10364), .B(n10365), .Z(n10363) );
  XNOR U10334 ( .A(y[3086]), .B(x[3086]), .Z(n10365) );
  XNOR U10335 ( .A(y[3087]), .B(x[3087]), .Z(n10364) );
  AND U10336 ( .A(n10366), .B(n10367), .Z(n10362) );
  XNOR U10337 ( .A(y[3088]), .B(x[3088]), .Z(n10367) );
  XNOR U10338 ( .A(y[3089]), .B(x[3089]), .Z(n10366) );
  AND U10339 ( .A(n10368), .B(n10369), .Z(n10336) );
  AND U10340 ( .A(n10370), .B(n10371), .Z(n10369) );
  AND U10341 ( .A(n10372), .B(n10373), .Z(n10371) );
  AND U10342 ( .A(n10374), .B(n10375), .Z(n10373) );
  XNOR U10343 ( .A(y[3090]), .B(x[3090]), .Z(n10375) );
  XNOR U10344 ( .A(y[3091]), .B(x[3091]), .Z(n10374) );
  AND U10345 ( .A(n10376), .B(n10377), .Z(n10372) );
  XNOR U10346 ( .A(y[3092]), .B(x[3092]), .Z(n10377) );
  XNOR U10347 ( .A(y[3093]), .B(x[3093]), .Z(n10376) );
  AND U10348 ( .A(n10378), .B(n10379), .Z(n10370) );
  AND U10349 ( .A(n10380), .B(n10381), .Z(n10379) );
  XNOR U10350 ( .A(y[3094]), .B(x[3094]), .Z(n10381) );
  XNOR U10351 ( .A(y[3095]), .B(x[3095]), .Z(n10380) );
  AND U10352 ( .A(n10382), .B(n10383), .Z(n10378) );
  XNOR U10353 ( .A(y[3096]), .B(x[3096]), .Z(n10383) );
  XNOR U10354 ( .A(y[3097]), .B(x[3097]), .Z(n10382) );
  AND U10355 ( .A(n10384), .B(n10385), .Z(n10368) );
  AND U10356 ( .A(n10386), .B(n10387), .Z(n10385) );
  AND U10357 ( .A(n10388), .B(n10389), .Z(n10387) );
  XNOR U10358 ( .A(y[3098]), .B(x[3098]), .Z(n10389) );
  XNOR U10359 ( .A(y[3099]), .B(x[3099]), .Z(n10388) );
  AND U10360 ( .A(n10390), .B(n10391), .Z(n10386) );
  XNOR U10361 ( .A(y[3100]), .B(x[3100]), .Z(n10391) );
  XNOR U10362 ( .A(y[3101]), .B(x[3101]), .Z(n10390) );
  AND U10363 ( .A(n10392), .B(n10393), .Z(n10384) );
  AND U10364 ( .A(n10394), .B(n10395), .Z(n10393) );
  XNOR U10365 ( .A(y[3102]), .B(x[3102]), .Z(n10395) );
  XNOR U10366 ( .A(y[3103]), .B(x[3103]), .Z(n10394) );
  AND U10367 ( .A(n10396), .B(n10397), .Z(n10392) );
  XNOR U10368 ( .A(y[3104]), .B(x[3104]), .Z(n10397) );
  XNOR U10369 ( .A(y[3105]), .B(x[3105]), .Z(n10396) );
  AND U10370 ( .A(n10398), .B(n10399), .Z(n10334) );
  AND U10371 ( .A(n10400), .B(n10401), .Z(n10399) );
  AND U10372 ( .A(n10402), .B(n10403), .Z(n10401) );
  AND U10373 ( .A(n10404), .B(n10405), .Z(n10403) );
  AND U10374 ( .A(n10406), .B(n10407), .Z(n10405) );
  XNOR U10375 ( .A(y[3106]), .B(x[3106]), .Z(n10407) );
  XNOR U10376 ( .A(y[3107]), .B(x[3107]), .Z(n10406) );
  AND U10377 ( .A(n10408), .B(n10409), .Z(n10404) );
  XNOR U10378 ( .A(y[3108]), .B(x[3108]), .Z(n10409) );
  XNOR U10379 ( .A(y[3109]), .B(x[3109]), .Z(n10408) );
  AND U10380 ( .A(n10410), .B(n10411), .Z(n10402) );
  AND U10381 ( .A(n10412), .B(n10413), .Z(n10411) );
  XNOR U10382 ( .A(y[3110]), .B(x[3110]), .Z(n10413) );
  XNOR U10383 ( .A(y[3111]), .B(x[3111]), .Z(n10412) );
  AND U10384 ( .A(n10414), .B(n10415), .Z(n10410) );
  XNOR U10385 ( .A(y[3112]), .B(x[3112]), .Z(n10415) );
  XNOR U10386 ( .A(y[3113]), .B(x[3113]), .Z(n10414) );
  AND U10387 ( .A(n10416), .B(n10417), .Z(n10400) );
  AND U10388 ( .A(n10418), .B(n10419), .Z(n10417) );
  AND U10389 ( .A(n10420), .B(n10421), .Z(n10419) );
  XNOR U10390 ( .A(y[3114]), .B(x[3114]), .Z(n10421) );
  XNOR U10391 ( .A(y[3115]), .B(x[3115]), .Z(n10420) );
  AND U10392 ( .A(n10422), .B(n10423), .Z(n10418) );
  XNOR U10393 ( .A(y[3116]), .B(x[3116]), .Z(n10423) );
  XNOR U10394 ( .A(y[3117]), .B(x[3117]), .Z(n10422) );
  AND U10395 ( .A(n10424), .B(n10425), .Z(n10416) );
  AND U10396 ( .A(n10426), .B(n10427), .Z(n10425) );
  XNOR U10397 ( .A(y[3118]), .B(x[3118]), .Z(n10427) );
  XNOR U10398 ( .A(y[3119]), .B(x[3119]), .Z(n10426) );
  AND U10399 ( .A(n10428), .B(n10429), .Z(n10424) );
  XNOR U10400 ( .A(y[3120]), .B(x[3120]), .Z(n10429) );
  XNOR U10401 ( .A(y[3121]), .B(x[3121]), .Z(n10428) );
  AND U10402 ( .A(n10430), .B(n10431), .Z(n10398) );
  AND U10403 ( .A(n10432), .B(n10433), .Z(n10431) );
  AND U10404 ( .A(n10434), .B(n10435), .Z(n10433) );
  AND U10405 ( .A(n10436), .B(n10437), .Z(n10435) );
  XNOR U10406 ( .A(y[3122]), .B(x[3122]), .Z(n10437) );
  XNOR U10407 ( .A(y[3123]), .B(x[3123]), .Z(n10436) );
  AND U10408 ( .A(n10438), .B(n10439), .Z(n10434) );
  XNOR U10409 ( .A(y[3124]), .B(x[3124]), .Z(n10439) );
  XNOR U10410 ( .A(y[3125]), .B(x[3125]), .Z(n10438) );
  AND U10411 ( .A(n10440), .B(n10441), .Z(n10432) );
  AND U10412 ( .A(n10442), .B(n10443), .Z(n10441) );
  XNOR U10413 ( .A(y[3126]), .B(x[3126]), .Z(n10443) );
  XNOR U10414 ( .A(y[3127]), .B(x[3127]), .Z(n10442) );
  AND U10415 ( .A(n10444), .B(n10445), .Z(n10440) );
  XNOR U10416 ( .A(y[3128]), .B(x[3128]), .Z(n10445) );
  XNOR U10417 ( .A(y[3129]), .B(x[3129]), .Z(n10444) );
  AND U10418 ( .A(n10446), .B(n10447), .Z(n10430) );
  AND U10419 ( .A(n10448), .B(n10449), .Z(n10447) );
  AND U10420 ( .A(n10450), .B(n10451), .Z(n10449) );
  XNOR U10421 ( .A(y[3130]), .B(x[3130]), .Z(n10451) );
  XNOR U10422 ( .A(y[3131]), .B(x[3131]), .Z(n10450) );
  AND U10423 ( .A(n10452), .B(n10453), .Z(n10448) );
  XNOR U10424 ( .A(y[3132]), .B(x[3132]), .Z(n10453) );
  XNOR U10425 ( .A(y[3133]), .B(x[3133]), .Z(n10452) );
  AND U10426 ( .A(n10454), .B(n10455), .Z(n10446) );
  AND U10427 ( .A(n10456), .B(n10457), .Z(n10455) );
  XNOR U10428 ( .A(y[3134]), .B(x[3134]), .Z(n10457) );
  XNOR U10429 ( .A(y[3135]), .B(x[3135]), .Z(n10456) );
  AND U10430 ( .A(n10458), .B(n10459), .Z(n10454) );
  XNOR U10431 ( .A(y[3136]), .B(x[3136]), .Z(n10459) );
  XNOR U10432 ( .A(y[3137]), .B(x[3137]), .Z(n10458) );
  AND U10433 ( .A(n10460), .B(n10461), .Z(n10332) );
  AND U10434 ( .A(n10462), .B(n10463), .Z(n10461) );
  AND U10435 ( .A(n10464), .B(n10465), .Z(n10463) );
  AND U10436 ( .A(n10466), .B(n10467), .Z(n10465) );
  AND U10437 ( .A(n10468), .B(n10469), .Z(n10467) );
  AND U10438 ( .A(n10470), .B(n10471), .Z(n10469) );
  XNOR U10439 ( .A(y[3138]), .B(x[3138]), .Z(n10471) );
  XNOR U10440 ( .A(y[3139]), .B(x[3139]), .Z(n10470) );
  AND U10441 ( .A(n10472), .B(n10473), .Z(n10468) );
  XNOR U10442 ( .A(y[3140]), .B(x[3140]), .Z(n10473) );
  XNOR U10443 ( .A(y[3141]), .B(x[3141]), .Z(n10472) );
  AND U10444 ( .A(n10474), .B(n10475), .Z(n10466) );
  AND U10445 ( .A(n10476), .B(n10477), .Z(n10475) );
  XNOR U10446 ( .A(y[3142]), .B(x[3142]), .Z(n10477) );
  XNOR U10447 ( .A(y[3143]), .B(x[3143]), .Z(n10476) );
  AND U10448 ( .A(n10478), .B(n10479), .Z(n10474) );
  XNOR U10449 ( .A(y[3144]), .B(x[3144]), .Z(n10479) );
  XNOR U10450 ( .A(y[3145]), .B(x[3145]), .Z(n10478) );
  AND U10451 ( .A(n10480), .B(n10481), .Z(n10464) );
  AND U10452 ( .A(n10482), .B(n10483), .Z(n10481) );
  AND U10453 ( .A(n10484), .B(n10485), .Z(n10483) );
  XNOR U10454 ( .A(y[3146]), .B(x[3146]), .Z(n10485) );
  XNOR U10455 ( .A(y[3147]), .B(x[3147]), .Z(n10484) );
  AND U10456 ( .A(n10486), .B(n10487), .Z(n10482) );
  XNOR U10457 ( .A(y[3148]), .B(x[3148]), .Z(n10487) );
  XNOR U10458 ( .A(y[3149]), .B(x[3149]), .Z(n10486) );
  AND U10459 ( .A(n10488), .B(n10489), .Z(n10480) );
  AND U10460 ( .A(n10490), .B(n10491), .Z(n10489) );
  XNOR U10461 ( .A(y[3150]), .B(x[3150]), .Z(n10491) );
  XNOR U10462 ( .A(y[3151]), .B(x[3151]), .Z(n10490) );
  AND U10463 ( .A(n10492), .B(n10493), .Z(n10488) );
  XNOR U10464 ( .A(y[3152]), .B(x[3152]), .Z(n10493) );
  XNOR U10465 ( .A(y[3153]), .B(x[3153]), .Z(n10492) );
  AND U10466 ( .A(n10494), .B(n10495), .Z(n10462) );
  AND U10467 ( .A(n10496), .B(n10497), .Z(n10495) );
  AND U10468 ( .A(n10498), .B(n10499), .Z(n10497) );
  AND U10469 ( .A(n10500), .B(n10501), .Z(n10499) );
  XNOR U10470 ( .A(y[3154]), .B(x[3154]), .Z(n10501) );
  XNOR U10471 ( .A(y[3155]), .B(x[3155]), .Z(n10500) );
  AND U10472 ( .A(n10502), .B(n10503), .Z(n10498) );
  XNOR U10473 ( .A(y[3156]), .B(x[3156]), .Z(n10503) );
  XNOR U10474 ( .A(y[3157]), .B(x[3157]), .Z(n10502) );
  AND U10475 ( .A(n10504), .B(n10505), .Z(n10496) );
  AND U10476 ( .A(n10506), .B(n10507), .Z(n10505) );
  XNOR U10477 ( .A(y[3158]), .B(x[3158]), .Z(n10507) );
  XNOR U10478 ( .A(y[3159]), .B(x[3159]), .Z(n10506) );
  AND U10479 ( .A(n10508), .B(n10509), .Z(n10504) );
  XNOR U10480 ( .A(y[3160]), .B(x[3160]), .Z(n10509) );
  XNOR U10481 ( .A(y[3161]), .B(x[3161]), .Z(n10508) );
  AND U10482 ( .A(n10510), .B(n10511), .Z(n10494) );
  AND U10483 ( .A(n10512), .B(n10513), .Z(n10511) );
  AND U10484 ( .A(n10514), .B(n10515), .Z(n10513) );
  XNOR U10485 ( .A(y[3162]), .B(x[3162]), .Z(n10515) );
  XNOR U10486 ( .A(y[3163]), .B(x[3163]), .Z(n10514) );
  AND U10487 ( .A(n10516), .B(n10517), .Z(n10512) );
  XNOR U10488 ( .A(y[3164]), .B(x[3164]), .Z(n10517) );
  XNOR U10489 ( .A(y[3165]), .B(x[3165]), .Z(n10516) );
  AND U10490 ( .A(n10518), .B(n10519), .Z(n10510) );
  AND U10491 ( .A(n10520), .B(n10521), .Z(n10519) );
  XNOR U10492 ( .A(y[3166]), .B(x[3166]), .Z(n10521) );
  XNOR U10493 ( .A(y[3167]), .B(x[3167]), .Z(n10520) );
  AND U10494 ( .A(n10522), .B(n10523), .Z(n10518) );
  XNOR U10495 ( .A(y[3168]), .B(x[3168]), .Z(n10523) );
  XNOR U10496 ( .A(y[3169]), .B(x[3169]), .Z(n10522) );
  AND U10497 ( .A(n10524), .B(n10525), .Z(n10460) );
  AND U10498 ( .A(n10526), .B(n10527), .Z(n10525) );
  AND U10499 ( .A(n10528), .B(n10529), .Z(n10527) );
  AND U10500 ( .A(n10530), .B(n10531), .Z(n10529) );
  AND U10501 ( .A(n10532), .B(n10533), .Z(n10531) );
  XNOR U10502 ( .A(y[3170]), .B(x[3170]), .Z(n10533) );
  XNOR U10503 ( .A(y[3171]), .B(x[3171]), .Z(n10532) );
  AND U10504 ( .A(n10534), .B(n10535), .Z(n10530) );
  XNOR U10505 ( .A(y[3172]), .B(x[3172]), .Z(n10535) );
  XNOR U10506 ( .A(y[3173]), .B(x[3173]), .Z(n10534) );
  AND U10507 ( .A(n10536), .B(n10537), .Z(n10528) );
  AND U10508 ( .A(n10538), .B(n10539), .Z(n10537) );
  XNOR U10509 ( .A(y[3174]), .B(x[3174]), .Z(n10539) );
  XNOR U10510 ( .A(y[3175]), .B(x[3175]), .Z(n10538) );
  AND U10511 ( .A(n10540), .B(n10541), .Z(n10536) );
  XNOR U10512 ( .A(y[3176]), .B(x[3176]), .Z(n10541) );
  XNOR U10513 ( .A(y[3177]), .B(x[3177]), .Z(n10540) );
  AND U10514 ( .A(n10542), .B(n10543), .Z(n10526) );
  AND U10515 ( .A(n10544), .B(n10545), .Z(n10543) );
  AND U10516 ( .A(n10546), .B(n10547), .Z(n10545) );
  XNOR U10517 ( .A(y[3178]), .B(x[3178]), .Z(n10547) );
  XNOR U10518 ( .A(y[3179]), .B(x[3179]), .Z(n10546) );
  AND U10519 ( .A(n10548), .B(n10549), .Z(n10544) );
  XNOR U10520 ( .A(y[3180]), .B(x[3180]), .Z(n10549) );
  XNOR U10521 ( .A(y[3181]), .B(x[3181]), .Z(n10548) );
  AND U10522 ( .A(n10550), .B(n10551), .Z(n10542) );
  AND U10523 ( .A(n10552), .B(n10553), .Z(n10551) );
  XNOR U10524 ( .A(y[3182]), .B(x[3182]), .Z(n10553) );
  XNOR U10525 ( .A(y[3183]), .B(x[3183]), .Z(n10552) );
  AND U10526 ( .A(n10554), .B(n10555), .Z(n10550) );
  XNOR U10527 ( .A(y[3184]), .B(x[3184]), .Z(n10555) );
  XNOR U10528 ( .A(y[3185]), .B(x[3185]), .Z(n10554) );
  AND U10529 ( .A(n10556), .B(n10557), .Z(n10524) );
  AND U10530 ( .A(n10558), .B(n10559), .Z(n10557) );
  AND U10531 ( .A(n10560), .B(n10561), .Z(n10559) );
  AND U10532 ( .A(n10562), .B(n10563), .Z(n10561) );
  XNOR U10533 ( .A(y[3186]), .B(x[3186]), .Z(n10563) );
  XNOR U10534 ( .A(y[3187]), .B(x[3187]), .Z(n10562) );
  AND U10535 ( .A(n10564), .B(n10565), .Z(n10560) );
  XNOR U10536 ( .A(y[3188]), .B(x[3188]), .Z(n10565) );
  XNOR U10537 ( .A(y[3189]), .B(x[3189]), .Z(n10564) );
  AND U10538 ( .A(n10566), .B(n10567), .Z(n10558) );
  AND U10539 ( .A(n10568), .B(n10569), .Z(n10567) );
  XNOR U10540 ( .A(y[3190]), .B(x[3190]), .Z(n10569) );
  XNOR U10541 ( .A(y[3191]), .B(x[3191]), .Z(n10568) );
  AND U10542 ( .A(n10570), .B(n10571), .Z(n10566) );
  XNOR U10543 ( .A(y[3192]), .B(x[3192]), .Z(n10571) );
  XNOR U10544 ( .A(y[3193]), .B(x[3193]), .Z(n10570) );
  AND U10545 ( .A(n10572), .B(n10573), .Z(n10556) );
  AND U10546 ( .A(n10574), .B(n10575), .Z(n10573) );
  AND U10547 ( .A(n10576), .B(n10577), .Z(n10575) );
  XNOR U10548 ( .A(y[3194]), .B(x[3194]), .Z(n10577) );
  XNOR U10549 ( .A(y[3195]), .B(x[3195]), .Z(n10576) );
  AND U10550 ( .A(n10578), .B(n10579), .Z(n10574) );
  XNOR U10551 ( .A(y[3196]), .B(x[3196]), .Z(n10579) );
  XNOR U10552 ( .A(y[3197]), .B(x[3197]), .Z(n10578) );
  AND U10553 ( .A(n10580), .B(n10581), .Z(n10572) );
  AND U10554 ( .A(n10582), .B(n10583), .Z(n10581) );
  XNOR U10555 ( .A(y[3198]), .B(x[3198]), .Z(n10583) );
  XNOR U10556 ( .A(y[3199]), .B(x[3199]), .Z(n10582) );
  AND U10557 ( .A(n10584), .B(n10585), .Z(n10580) );
  XNOR U10558 ( .A(y[3200]), .B(x[3200]), .Z(n10585) );
  XNOR U10559 ( .A(y[3201]), .B(x[3201]), .Z(n10584) );
  AND U10560 ( .A(n10586), .B(n10587), .Z(n10330) );
  AND U10561 ( .A(n10588), .B(n10589), .Z(n10587) );
  AND U10562 ( .A(n10590), .B(n10591), .Z(n10589) );
  AND U10563 ( .A(n10592), .B(n10593), .Z(n10591) );
  AND U10564 ( .A(n10594), .B(n10595), .Z(n10593) );
  AND U10565 ( .A(n10596), .B(n10597), .Z(n10595) );
  AND U10566 ( .A(n10598), .B(n10599), .Z(n10597) );
  XNOR U10567 ( .A(y[3202]), .B(x[3202]), .Z(n10599) );
  XNOR U10568 ( .A(y[3203]), .B(x[3203]), .Z(n10598) );
  AND U10569 ( .A(n10600), .B(n10601), .Z(n10596) );
  XNOR U10570 ( .A(y[3204]), .B(x[3204]), .Z(n10601) );
  XNOR U10571 ( .A(y[3205]), .B(x[3205]), .Z(n10600) );
  AND U10572 ( .A(n10602), .B(n10603), .Z(n10594) );
  AND U10573 ( .A(n10604), .B(n10605), .Z(n10603) );
  XNOR U10574 ( .A(y[3206]), .B(x[3206]), .Z(n10605) );
  XNOR U10575 ( .A(y[3207]), .B(x[3207]), .Z(n10604) );
  AND U10576 ( .A(n10606), .B(n10607), .Z(n10602) );
  XNOR U10577 ( .A(y[3208]), .B(x[3208]), .Z(n10607) );
  XNOR U10578 ( .A(y[3209]), .B(x[3209]), .Z(n10606) );
  AND U10579 ( .A(n10608), .B(n10609), .Z(n10592) );
  AND U10580 ( .A(n10610), .B(n10611), .Z(n10609) );
  AND U10581 ( .A(n10612), .B(n10613), .Z(n10611) );
  XNOR U10582 ( .A(y[3210]), .B(x[3210]), .Z(n10613) );
  XNOR U10583 ( .A(y[3211]), .B(x[3211]), .Z(n10612) );
  AND U10584 ( .A(n10614), .B(n10615), .Z(n10610) );
  XNOR U10585 ( .A(y[3212]), .B(x[3212]), .Z(n10615) );
  XNOR U10586 ( .A(y[3213]), .B(x[3213]), .Z(n10614) );
  AND U10587 ( .A(n10616), .B(n10617), .Z(n10608) );
  AND U10588 ( .A(n10618), .B(n10619), .Z(n10617) );
  XNOR U10589 ( .A(y[3214]), .B(x[3214]), .Z(n10619) );
  XNOR U10590 ( .A(y[3215]), .B(x[3215]), .Z(n10618) );
  AND U10591 ( .A(n10620), .B(n10621), .Z(n10616) );
  XNOR U10592 ( .A(y[3216]), .B(x[3216]), .Z(n10621) );
  XNOR U10593 ( .A(y[3217]), .B(x[3217]), .Z(n10620) );
  AND U10594 ( .A(n10622), .B(n10623), .Z(n10590) );
  AND U10595 ( .A(n10624), .B(n10625), .Z(n10623) );
  AND U10596 ( .A(n10626), .B(n10627), .Z(n10625) );
  AND U10597 ( .A(n10628), .B(n10629), .Z(n10627) );
  XNOR U10598 ( .A(y[3218]), .B(x[3218]), .Z(n10629) );
  XNOR U10599 ( .A(y[3219]), .B(x[3219]), .Z(n10628) );
  AND U10600 ( .A(n10630), .B(n10631), .Z(n10626) );
  XNOR U10601 ( .A(y[3220]), .B(x[3220]), .Z(n10631) );
  XNOR U10602 ( .A(y[3221]), .B(x[3221]), .Z(n10630) );
  AND U10603 ( .A(n10632), .B(n10633), .Z(n10624) );
  AND U10604 ( .A(n10634), .B(n10635), .Z(n10633) );
  XNOR U10605 ( .A(y[3222]), .B(x[3222]), .Z(n10635) );
  XNOR U10606 ( .A(y[3223]), .B(x[3223]), .Z(n10634) );
  AND U10607 ( .A(n10636), .B(n10637), .Z(n10632) );
  XNOR U10608 ( .A(y[3224]), .B(x[3224]), .Z(n10637) );
  XNOR U10609 ( .A(y[3225]), .B(x[3225]), .Z(n10636) );
  AND U10610 ( .A(n10638), .B(n10639), .Z(n10622) );
  AND U10611 ( .A(n10640), .B(n10641), .Z(n10639) );
  AND U10612 ( .A(n10642), .B(n10643), .Z(n10641) );
  XNOR U10613 ( .A(y[3226]), .B(x[3226]), .Z(n10643) );
  XNOR U10614 ( .A(y[3227]), .B(x[3227]), .Z(n10642) );
  AND U10615 ( .A(n10644), .B(n10645), .Z(n10640) );
  XNOR U10616 ( .A(y[3228]), .B(x[3228]), .Z(n10645) );
  XNOR U10617 ( .A(y[3229]), .B(x[3229]), .Z(n10644) );
  AND U10618 ( .A(n10646), .B(n10647), .Z(n10638) );
  AND U10619 ( .A(n10648), .B(n10649), .Z(n10647) );
  XNOR U10620 ( .A(y[3230]), .B(x[3230]), .Z(n10649) );
  XNOR U10621 ( .A(y[3231]), .B(x[3231]), .Z(n10648) );
  AND U10622 ( .A(n10650), .B(n10651), .Z(n10646) );
  XNOR U10623 ( .A(y[3232]), .B(x[3232]), .Z(n10651) );
  XNOR U10624 ( .A(y[3233]), .B(x[3233]), .Z(n10650) );
  AND U10625 ( .A(n10652), .B(n10653), .Z(n10588) );
  AND U10626 ( .A(n10654), .B(n10655), .Z(n10653) );
  AND U10627 ( .A(n10656), .B(n10657), .Z(n10655) );
  AND U10628 ( .A(n10658), .B(n10659), .Z(n10657) );
  AND U10629 ( .A(n10660), .B(n10661), .Z(n10659) );
  XNOR U10630 ( .A(y[3234]), .B(x[3234]), .Z(n10661) );
  XNOR U10631 ( .A(y[3235]), .B(x[3235]), .Z(n10660) );
  AND U10632 ( .A(n10662), .B(n10663), .Z(n10658) );
  XNOR U10633 ( .A(y[3236]), .B(x[3236]), .Z(n10663) );
  XNOR U10634 ( .A(y[3237]), .B(x[3237]), .Z(n10662) );
  AND U10635 ( .A(n10664), .B(n10665), .Z(n10656) );
  AND U10636 ( .A(n10666), .B(n10667), .Z(n10665) );
  XNOR U10637 ( .A(y[3238]), .B(x[3238]), .Z(n10667) );
  XNOR U10638 ( .A(y[3239]), .B(x[3239]), .Z(n10666) );
  AND U10639 ( .A(n10668), .B(n10669), .Z(n10664) );
  XNOR U10640 ( .A(y[3240]), .B(x[3240]), .Z(n10669) );
  XNOR U10641 ( .A(y[3241]), .B(x[3241]), .Z(n10668) );
  AND U10642 ( .A(n10670), .B(n10671), .Z(n10654) );
  AND U10643 ( .A(n10672), .B(n10673), .Z(n10671) );
  AND U10644 ( .A(n10674), .B(n10675), .Z(n10673) );
  XNOR U10645 ( .A(y[3242]), .B(x[3242]), .Z(n10675) );
  XNOR U10646 ( .A(y[3243]), .B(x[3243]), .Z(n10674) );
  AND U10647 ( .A(n10676), .B(n10677), .Z(n10672) );
  XNOR U10648 ( .A(y[3244]), .B(x[3244]), .Z(n10677) );
  XNOR U10649 ( .A(y[3245]), .B(x[3245]), .Z(n10676) );
  AND U10650 ( .A(n10678), .B(n10679), .Z(n10670) );
  AND U10651 ( .A(n10680), .B(n10681), .Z(n10679) );
  XNOR U10652 ( .A(y[3246]), .B(x[3246]), .Z(n10681) );
  XNOR U10653 ( .A(y[3247]), .B(x[3247]), .Z(n10680) );
  AND U10654 ( .A(n10682), .B(n10683), .Z(n10678) );
  XNOR U10655 ( .A(y[3248]), .B(x[3248]), .Z(n10683) );
  XNOR U10656 ( .A(y[3249]), .B(x[3249]), .Z(n10682) );
  AND U10657 ( .A(n10684), .B(n10685), .Z(n10652) );
  AND U10658 ( .A(n10686), .B(n10687), .Z(n10685) );
  AND U10659 ( .A(n10688), .B(n10689), .Z(n10687) );
  AND U10660 ( .A(n10690), .B(n10691), .Z(n10689) );
  XNOR U10661 ( .A(y[3250]), .B(x[3250]), .Z(n10691) );
  XNOR U10662 ( .A(y[3251]), .B(x[3251]), .Z(n10690) );
  AND U10663 ( .A(n10692), .B(n10693), .Z(n10688) );
  XNOR U10664 ( .A(y[3252]), .B(x[3252]), .Z(n10693) );
  XNOR U10665 ( .A(y[3253]), .B(x[3253]), .Z(n10692) );
  AND U10666 ( .A(n10694), .B(n10695), .Z(n10686) );
  AND U10667 ( .A(n10696), .B(n10697), .Z(n10695) );
  XNOR U10668 ( .A(y[3254]), .B(x[3254]), .Z(n10697) );
  XNOR U10669 ( .A(y[3255]), .B(x[3255]), .Z(n10696) );
  AND U10670 ( .A(n10698), .B(n10699), .Z(n10694) );
  XNOR U10671 ( .A(y[3256]), .B(x[3256]), .Z(n10699) );
  XNOR U10672 ( .A(y[3257]), .B(x[3257]), .Z(n10698) );
  AND U10673 ( .A(n10700), .B(n10701), .Z(n10684) );
  AND U10674 ( .A(n10702), .B(n10703), .Z(n10701) );
  AND U10675 ( .A(n10704), .B(n10705), .Z(n10703) );
  XNOR U10676 ( .A(y[3258]), .B(x[3258]), .Z(n10705) );
  XNOR U10677 ( .A(y[3259]), .B(x[3259]), .Z(n10704) );
  AND U10678 ( .A(n10706), .B(n10707), .Z(n10702) );
  XNOR U10679 ( .A(y[3260]), .B(x[3260]), .Z(n10707) );
  XNOR U10680 ( .A(y[3261]), .B(x[3261]), .Z(n10706) );
  AND U10681 ( .A(n10708), .B(n10709), .Z(n10700) );
  AND U10682 ( .A(n10710), .B(n10711), .Z(n10709) );
  XNOR U10683 ( .A(y[3262]), .B(x[3262]), .Z(n10711) );
  XNOR U10684 ( .A(y[3263]), .B(x[3263]), .Z(n10710) );
  AND U10685 ( .A(n10712), .B(n10713), .Z(n10708) );
  XNOR U10686 ( .A(y[3264]), .B(x[3264]), .Z(n10713) );
  XNOR U10687 ( .A(y[3265]), .B(x[3265]), .Z(n10712) );
  AND U10688 ( .A(n10714), .B(n10715), .Z(n10586) );
  AND U10689 ( .A(n10716), .B(n10717), .Z(n10715) );
  AND U10690 ( .A(n10718), .B(n10719), .Z(n10717) );
  AND U10691 ( .A(n10720), .B(n10721), .Z(n10719) );
  AND U10692 ( .A(n10722), .B(n10723), .Z(n10721) );
  AND U10693 ( .A(n10724), .B(n10725), .Z(n10723) );
  XNOR U10694 ( .A(y[3266]), .B(x[3266]), .Z(n10725) );
  XNOR U10695 ( .A(y[3267]), .B(x[3267]), .Z(n10724) );
  AND U10696 ( .A(n10726), .B(n10727), .Z(n10722) );
  XNOR U10697 ( .A(y[3268]), .B(x[3268]), .Z(n10727) );
  XNOR U10698 ( .A(y[3269]), .B(x[3269]), .Z(n10726) );
  AND U10699 ( .A(n10728), .B(n10729), .Z(n10720) );
  AND U10700 ( .A(n10730), .B(n10731), .Z(n10729) );
  XNOR U10701 ( .A(y[3270]), .B(x[3270]), .Z(n10731) );
  XNOR U10702 ( .A(y[3271]), .B(x[3271]), .Z(n10730) );
  AND U10703 ( .A(n10732), .B(n10733), .Z(n10728) );
  XNOR U10704 ( .A(y[3272]), .B(x[3272]), .Z(n10733) );
  XNOR U10705 ( .A(y[3273]), .B(x[3273]), .Z(n10732) );
  AND U10706 ( .A(n10734), .B(n10735), .Z(n10718) );
  AND U10707 ( .A(n10736), .B(n10737), .Z(n10735) );
  AND U10708 ( .A(n10738), .B(n10739), .Z(n10737) );
  XNOR U10709 ( .A(y[3274]), .B(x[3274]), .Z(n10739) );
  XNOR U10710 ( .A(y[3275]), .B(x[3275]), .Z(n10738) );
  AND U10711 ( .A(n10740), .B(n10741), .Z(n10736) );
  XNOR U10712 ( .A(y[3276]), .B(x[3276]), .Z(n10741) );
  XNOR U10713 ( .A(y[3277]), .B(x[3277]), .Z(n10740) );
  AND U10714 ( .A(n10742), .B(n10743), .Z(n10734) );
  AND U10715 ( .A(n10744), .B(n10745), .Z(n10743) );
  XNOR U10716 ( .A(y[3278]), .B(x[3278]), .Z(n10745) );
  XNOR U10717 ( .A(y[3279]), .B(x[3279]), .Z(n10744) );
  AND U10718 ( .A(n10746), .B(n10747), .Z(n10742) );
  XNOR U10719 ( .A(y[3280]), .B(x[3280]), .Z(n10747) );
  XNOR U10720 ( .A(y[3281]), .B(x[3281]), .Z(n10746) );
  AND U10721 ( .A(n10748), .B(n10749), .Z(n10716) );
  AND U10722 ( .A(n10750), .B(n10751), .Z(n10749) );
  AND U10723 ( .A(n10752), .B(n10753), .Z(n10751) );
  AND U10724 ( .A(n10754), .B(n10755), .Z(n10753) );
  XNOR U10725 ( .A(y[3282]), .B(x[3282]), .Z(n10755) );
  XNOR U10726 ( .A(y[3283]), .B(x[3283]), .Z(n10754) );
  AND U10727 ( .A(n10756), .B(n10757), .Z(n10752) );
  XNOR U10728 ( .A(y[3284]), .B(x[3284]), .Z(n10757) );
  XNOR U10729 ( .A(y[3285]), .B(x[3285]), .Z(n10756) );
  AND U10730 ( .A(n10758), .B(n10759), .Z(n10750) );
  AND U10731 ( .A(n10760), .B(n10761), .Z(n10759) );
  XNOR U10732 ( .A(y[3286]), .B(x[3286]), .Z(n10761) );
  XNOR U10733 ( .A(y[3287]), .B(x[3287]), .Z(n10760) );
  AND U10734 ( .A(n10762), .B(n10763), .Z(n10758) );
  XNOR U10735 ( .A(y[3288]), .B(x[3288]), .Z(n10763) );
  XNOR U10736 ( .A(y[3289]), .B(x[3289]), .Z(n10762) );
  AND U10737 ( .A(n10764), .B(n10765), .Z(n10748) );
  AND U10738 ( .A(n10766), .B(n10767), .Z(n10765) );
  AND U10739 ( .A(n10768), .B(n10769), .Z(n10767) );
  XNOR U10740 ( .A(y[3290]), .B(x[3290]), .Z(n10769) );
  XNOR U10741 ( .A(y[3291]), .B(x[3291]), .Z(n10768) );
  AND U10742 ( .A(n10770), .B(n10771), .Z(n10766) );
  XNOR U10743 ( .A(y[3292]), .B(x[3292]), .Z(n10771) );
  XNOR U10744 ( .A(y[3293]), .B(x[3293]), .Z(n10770) );
  AND U10745 ( .A(n10772), .B(n10773), .Z(n10764) );
  AND U10746 ( .A(n10774), .B(n10775), .Z(n10773) );
  XNOR U10747 ( .A(y[3294]), .B(x[3294]), .Z(n10775) );
  XNOR U10748 ( .A(y[3295]), .B(x[3295]), .Z(n10774) );
  AND U10749 ( .A(n10776), .B(n10777), .Z(n10772) );
  XNOR U10750 ( .A(y[3296]), .B(x[3296]), .Z(n10777) );
  XNOR U10751 ( .A(y[3297]), .B(x[3297]), .Z(n10776) );
  AND U10752 ( .A(n10778), .B(n10779), .Z(n10714) );
  AND U10753 ( .A(n10780), .B(n10781), .Z(n10779) );
  AND U10754 ( .A(n10782), .B(n10783), .Z(n10781) );
  AND U10755 ( .A(n10784), .B(n10785), .Z(n10783) );
  AND U10756 ( .A(n10786), .B(n10787), .Z(n10785) );
  XNOR U10757 ( .A(y[3298]), .B(x[3298]), .Z(n10787) );
  XNOR U10758 ( .A(y[3299]), .B(x[3299]), .Z(n10786) );
  AND U10759 ( .A(n10788), .B(n10789), .Z(n10784) );
  XNOR U10760 ( .A(y[3300]), .B(x[3300]), .Z(n10789) );
  XNOR U10761 ( .A(y[3301]), .B(x[3301]), .Z(n10788) );
  AND U10762 ( .A(n10790), .B(n10791), .Z(n10782) );
  AND U10763 ( .A(n10792), .B(n10793), .Z(n10791) );
  XNOR U10764 ( .A(y[3302]), .B(x[3302]), .Z(n10793) );
  XNOR U10765 ( .A(y[3303]), .B(x[3303]), .Z(n10792) );
  AND U10766 ( .A(n10794), .B(n10795), .Z(n10790) );
  XNOR U10767 ( .A(y[3304]), .B(x[3304]), .Z(n10795) );
  XNOR U10768 ( .A(y[3305]), .B(x[3305]), .Z(n10794) );
  AND U10769 ( .A(n10796), .B(n10797), .Z(n10780) );
  AND U10770 ( .A(n10798), .B(n10799), .Z(n10797) );
  AND U10771 ( .A(n10800), .B(n10801), .Z(n10799) );
  XNOR U10772 ( .A(y[3306]), .B(x[3306]), .Z(n10801) );
  XNOR U10773 ( .A(y[3307]), .B(x[3307]), .Z(n10800) );
  AND U10774 ( .A(n10802), .B(n10803), .Z(n10798) );
  XNOR U10775 ( .A(y[3308]), .B(x[3308]), .Z(n10803) );
  XNOR U10776 ( .A(y[3309]), .B(x[3309]), .Z(n10802) );
  AND U10777 ( .A(n10804), .B(n10805), .Z(n10796) );
  AND U10778 ( .A(n10806), .B(n10807), .Z(n10805) );
  XNOR U10779 ( .A(y[3310]), .B(x[3310]), .Z(n10807) );
  XNOR U10780 ( .A(y[3311]), .B(x[3311]), .Z(n10806) );
  AND U10781 ( .A(n10808), .B(n10809), .Z(n10804) );
  XNOR U10782 ( .A(y[3312]), .B(x[3312]), .Z(n10809) );
  XNOR U10783 ( .A(y[3313]), .B(x[3313]), .Z(n10808) );
  AND U10784 ( .A(n10810), .B(n10811), .Z(n10778) );
  AND U10785 ( .A(n10812), .B(n10813), .Z(n10811) );
  AND U10786 ( .A(n10814), .B(n10815), .Z(n10813) );
  AND U10787 ( .A(n10816), .B(n10817), .Z(n10815) );
  XNOR U10788 ( .A(y[3314]), .B(x[3314]), .Z(n10817) );
  XNOR U10789 ( .A(y[3315]), .B(x[3315]), .Z(n10816) );
  AND U10790 ( .A(n10818), .B(n10819), .Z(n10814) );
  XNOR U10791 ( .A(y[3316]), .B(x[3316]), .Z(n10819) );
  XNOR U10792 ( .A(y[3317]), .B(x[3317]), .Z(n10818) );
  AND U10793 ( .A(n10820), .B(n10821), .Z(n10812) );
  AND U10794 ( .A(n10822), .B(n10823), .Z(n10821) );
  XNOR U10795 ( .A(y[3318]), .B(x[3318]), .Z(n10823) );
  XNOR U10796 ( .A(y[3319]), .B(x[3319]), .Z(n10822) );
  AND U10797 ( .A(n10824), .B(n10825), .Z(n10820) );
  XNOR U10798 ( .A(y[3320]), .B(x[3320]), .Z(n10825) );
  XNOR U10799 ( .A(y[3321]), .B(x[3321]), .Z(n10824) );
  AND U10800 ( .A(n10826), .B(n10827), .Z(n10810) );
  AND U10801 ( .A(n10828), .B(n10829), .Z(n10827) );
  AND U10802 ( .A(n10830), .B(n10831), .Z(n10829) );
  XNOR U10803 ( .A(y[3322]), .B(x[3322]), .Z(n10831) );
  XNOR U10804 ( .A(y[3323]), .B(x[3323]), .Z(n10830) );
  AND U10805 ( .A(n10832), .B(n10833), .Z(n10828) );
  XNOR U10806 ( .A(y[3324]), .B(x[3324]), .Z(n10833) );
  XNOR U10807 ( .A(y[3325]), .B(x[3325]), .Z(n10832) );
  AND U10808 ( .A(n10834), .B(n10835), .Z(n10826) );
  AND U10809 ( .A(n10836), .B(n10837), .Z(n10835) );
  XNOR U10810 ( .A(y[3326]), .B(x[3326]), .Z(n10837) );
  XNOR U10811 ( .A(y[3327]), .B(x[3327]), .Z(n10836) );
  AND U10812 ( .A(n10838), .B(n10839), .Z(n10834) );
  XNOR U10813 ( .A(y[3328]), .B(x[3328]), .Z(n10839) );
  XNOR U10814 ( .A(y[3329]), .B(x[3329]), .Z(n10838) );
  AND U10815 ( .A(n10840), .B(n10841), .Z(n10072) );
  AND U10816 ( .A(n10842), .B(n10843), .Z(n10841) );
  AND U10817 ( .A(n10844), .B(n10845), .Z(n10843) );
  AND U10818 ( .A(n10846), .B(n10847), .Z(n10845) );
  AND U10819 ( .A(n10848), .B(n10849), .Z(n10847) );
  AND U10820 ( .A(n10850), .B(n10851), .Z(n10849) );
  AND U10821 ( .A(n10852), .B(n10853), .Z(n10851) );
  AND U10822 ( .A(n10854), .B(n10855), .Z(n10853) );
  AND U10823 ( .A(n10856), .B(n10857), .Z(n10855) );
  XNOR U10824 ( .A(y[3840]), .B(x[3840]), .Z(n10857) );
  XNOR U10825 ( .A(y[3841]), .B(x[3841]), .Z(n10856) );
  AND U10826 ( .A(n10858), .B(n10859), .Z(n10854) );
  XNOR U10827 ( .A(y[3842]), .B(x[3842]), .Z(n10859) );
  XNOR U10828 ( .A(y[3843]), .B(x[3843]), .Z(n10858) );
  AND U10829 ( .A(n10860), .B(n10861), .Z(n10852) );
  AND U10830 ( .A(n10862), .B(n10863), .Z(n10861) );
  XNOR U10831 ( .A(y[3844]), .B(x[3844]), .Z(n10863) );
  XNOR U10832 ( .A(y[3845]), .B(x[3845]), .Z(n10862) );
  AND U10833 ( .A(n10864), .B(n10865), .Z(n10860) );
  XNOR U10834 ( .A(y[3846]), .B(x[3846]), .Z(n10865) );
  XNOR U10835 ( .A(y[3847]), .B(x[3847]), .Z(n10864) );
  AND U10836 ( .A(n10866), .B(n10867), .Z(n10850) );
  AND U10837 ( .A(n10868), .B(n10869), .Z(n10867) );
  AND U10838 ( .A(n10870), .B(n10871), .Z(n10869) );
  XNOR U10839 ( .A(y[3848]), .B(x[3848]), .Z(n10871) );
  XNOR U10840 ( .A(y[3849]), .B(x[3849]), .Z(n10870) );
  AND U10841 ( .A(n10872), .B(n10873), .Z(n10868) );
  XNOR U10842 ( .A(y[3850]), .B(x[3850]), .Z(n10873) );
  XNOR U10843 ( .A(y[3851]), .B(x[3851]), .Z(n10872) );
  AND U10844 ( .A(n10874), .B(n10875), .Z(n10866) );
  AND U10845 ( .A(n10876), .B(n10877), .Z(n10875) );
  XNOR U10846 ( .A(y[3852]), .B(x[3852]), .Z(n10877) );
  XNOR U10847 ( .A(y[3853]), .B(x[3853]), .Z(n10876) );
  AND U10848 ( .A(n10878), .B(n10879), .Z(n10874) );
  XNOR U10849 ( .A(y[3854]), .B(x[3854]), .Z(n10879) );
  XNOR U10850 ( .A(y[3855]), .B(x[3855]), .Z(n10878) );
  AND U10851 ( .A(n10880), .B(n10881), .Z(n10848) );
  AND U10852 ( .A(n10882), .B(n10883), .Z(n10881) );
  AND U10853 ( .A(n10884), .B(n10885), .Z(n10883) );
  AND U10854 ( .A(n10886), .B(n10887), .Z(n10885) );
  XNOR U10855 ( .A(y[3856]), .B(x[3856]), .Z(n10887) );
  XNOR U10856 ( .A(y[3857]), .B(x[3857]), .Z(n10886) );
  AND U10857 ( .A(n10888), .B(n10889), .Z(n10884) );
  XNOR U10858 ( .A(y[3858]), .B(x[3858]), .Z(n10889) );
  XNOR U10859 ( .A(y[3859]), .B(x[3859]), .Z(n10888) );
  AND U10860 ( .A(n10890), .B(n10891), .Z(n10882) );
  AND U10861 ( .A(n10892), .B(n10893), .Z(n10891) );
  XNOR U10862 ( .A(y[3860]), .B(x[3860]), .Z(n10893) );
  XNOR U10863 ( .A(y[3861]), .B(x[3861]), .Z(n10892) );
  AND U10864 ( .A(n10894), .B(n10895), .Z(n10890) );
  XNOR U10865 ( .A(y[3862]), .B(x[3862]), .Z(n10895) );
  XNOR U10866 ( .A(y[3863]), .B(x[3863]), .Z(n10894) );
  AND U10867 ( .A(n10896), .B(n10897), .Z(n10880) );
  AND U10868 ( .A(n10898), .B(n10899), .Z(n10897) );
  AND U10869 ( .A(n10900), .B(n10901), .Z(n10899) );
  XNOR U10870 ( .A(y[3864]), .B(x[3864]), .Z(n10901) );
  XNOR U10871 ( .A(y[3865]), .B(x[3865]), .Z(n10900) );
  AND U10872 ( .A(n10902), .B(n10903), .Z(n10898) );
  XNOR U10873 ( .A(y[3866]), .B(x[3866]), .Z(n10903) );
  XNOR U10874 ( .A(y[3867]), .B(x[3867]), .Z(n10902) );
  AND U10875 ( .A(n10904), .B(n10905), .Z(n10896) );
  AND U10876 ( .A(n10906), .B(n10907), .Z(n10905) );
  XNOR U10877 ( .A(y[3868]), .B(x[3868]), .Z(n10907) );
  XNOR U10878 ( .A(y[3869]), .B(x[3869]), .Z(n10906) );
  AND U10879 ( .A(n10908), .B(n10909), .Z(n10904) );
  XNOR U10880 ( .A(y[3870]), .B(x[3870]), .Z(n10909) );
  XNOR U10881 ( .A(y[3871]), .B(x[3871]), .Z(n10908) );
  AND U10882 ( .A(n10910), .B(n10911), .Z(n10846) );
  AND U10883 ( .A(n10912), .B(n10913), .Z(n10911) );
  AND U10884 ( .A(n10914), .B(n10915), .Z(n10913) );
  AND U10885 ( .A(n10916), .B(n10917), .Z(n10915) );
  AND U10886 ( .A(n10918), .B(n10919), .Z(n10917) );
  XNOR U10887 ( .A(y[3872]), .B(x[3872]), .Z(n10919) );
  XNOR U10888 ( .A(y[3873]), .B(x[3873]), .Z(n10918) );
  AND U10889 ( .A(n10920), .B(n10921), .Z(n10916) );
  XNOR U10890 ( .A(y[3874]), .B(x[3874]), .Z(n10921) );
  XNOR U10891 ( .A(y[3875]), .B(x[3875]), .Z(n10920) );
  AND U10892 ( .A(n10922), .B(n10923), .Z(n10914) );
  AND U10893 ( .A(n10924), .B(n10925), .Z(n10923) );
  XNOR U10894 ( .A(y[3876]), .B(x[3876]), .Z(n10925) );
  XNOR U10895 ( .A(y[3877]), .B(x[3877]), .Z(n10924) );
  AND U10896 ( .A(n10926), .B(n10927), .Z(n10922) );
  XNOR U10897 ( .A(y[3878]), .B(x[3878]), .Z(n10927) );
  XNOR U10898 ( .A(y[3879]), .B(x[3879]), .Z(n10926) );
  AND U10899 ( .A(n10928), .B(n10929), .Z(n10912) );
  AND U10900 ( .A(n10930), .B(n10931), .Z(n10929) );
  AND U10901 ( .A(n10932), .B(n10933), .Z(n10931) );
  XNOR U10902 ( .A(y[3880]), .B(x[3880]), .Z(n10933) );
  XNOR U10903 ( .A(y[3881]), .B(x[3881]), .Z(n10932) );
  AND U10904 ( .A(n10934), .B(n10935), .Z(n10930) );
  XNOR U10905 ( .A(y[3882]), .B(x[3882]), .Z(n10935) );
  XNOR U10906 ( .A(y[3883]), .B(x[3883]), .Z(n10934) );
  AND U10907 ( .A(n10936), .B(n10937), .Z(n10928) );
  AND U10908 ( .A(n10938), .B(n10939), .Z(n10937) );
  XNOR U10909 ( .A(y[3884]), .B(x[3884]), .Z(n10939) );
  XNOR U10910 ( .A(y[3885]), .B(x[3885]), .Z(n10938) );
  AND U10911 ( .A(n10940), .B(n10941), .Z(n10936) );
  XNOR U10912 ( .A(y[3886]), .B(x[3886]), .Z(n10941) );
  XNOR U10913 ( .A(y[3887]), .B(x[3887]), .Z(n10940) );
  AND U10914 ( .A(n10942), .B(n10943), .Z(n10910) );
  AND U10915 ( .A(n10944), .B(n10945), .Z(n10943) );
  AND U10916 ( .A(n10946), .B(n10947), .Z(n10945) );
  AND U10917 ( .A(n10948), .B(n10949), .Z(n10947) );
  XNOR U10918 ( .A(y[3888]), .B(x[3888]), .Z(n10949) );
  XNOR U10919 ( .A(y[3889]), .B(x[3889]), .Z(n10948) );
  AND U10920 ( .A(n10950), .B(n10951), .Z(n10946) );
  XNOR U10921 ( .A(y[3890]), .B(x[3890]), .Z(n10951) );
  XNOR U10922 ( .A(y[3891]), .B(x[3891]), .Z(n10950) );
  AND U10923 ( .A(n10952), .B(n10953), .Z(n10944) );
  AND U10924 ( .A(n10954), .B(n10955), .Z(n10953) );
  XNOR U10925 ( .A(y[3892]), .B(x[3892]), .Z(n10955) );
  XNOR U10926 ( .A(y[3893]), .B(x[3893]), .Z(n10954) );
  AND U10927 ( .A(n10956), .B(n10957), .Z(n10952) );
  XNOR U10928 ( .A(y[3894]), .B(x[3894]), .Z(n10957) );
  XNOR U10929 ( .A(y[3895]), .B(x[3895]), .Z(n10956) );
  AND U10930 ( .A(n10958), .B(n10959), .Z(n10942) );
  AND U10931 ( .A(n10960), .B(n10961), .Z(n10959) );
  AND U10932 ( .A(n10962), .B(n10963), .Z(n10961) );
  XNOR U10933 ( .A(y[3896]), .B(x[3896]), .Z(n10963) );
  XNOR U10934 ( .A(y[3897]), .B(x[3897]), .Z(n10962) );
  AND U10935 ( .A(n10964), .B(n10965), .Z(n10960) );
  XNOR U10936 ( .A(y[3898]), .B(x[3898]), .Z(n10965) );
  XNOR U10937 ( .A(y[3899]), .B(x[3899]), .Z(n10964) );
  AND U10938 ( .A(n10966), .B(n10967), .Z(n10958) );
  AND U10939 ( .A(n10968), .B(n10969), .Z(n10967) );
  XNOR U10940 ( .A(y[3900]), .B(x[3900]), .Z(n10969) );
  XNOR U10941 ( .A(y[3901]), .B(x[3901]), .Z(n10968) );
  AND U10942 ( .A(n10970), .B(n10971), .Z(n10966) );
  XNOR U10943 ( .A(y[3902]), .B(x[3902]), .Z(n10971) );
  XNOR U10944 ( .A(y[3903]), .B(x[3903]), .Z(n10970) );
  AND U10945 ( .A(n10972), .B(n10973), .Z(n10844) );
  AND U10946 ( .A(n10974), .B(n10975), .Z(n10973) );
  AND U10947 ( .A(n10976), .B(n10977), .Z(n10975) );
  AND U10948 ( .A(n10978), .B(n10979), .Z(n10977) );
  AND U10949 ( .A(n10980), .B(n10981), .Z(n10979) );
  AND U10950 ( .A(n10982), .B(n10983), .Z(n10981) );
  XNOR U10951 ( .A(y[3904]), .B(x[3904]), .Z(n10983) );
  XNOR U10952 ( .A(y[3905]), .B(x[3905]), .Z(n10982) );
  AND U10953 ( .A(n10984), .B(n10985), .Z(n10980) );
  XNOR U10954 ( .A(y[3906]), .B(x[3906]), .Z(n10985) );
  XNOR U10955 ( .A(y[3907]), .B(x[3907]), .Z(n10984) );
  AND U10956 ( .A(n10986), .B(n10987), .Z(n10978) );
  AND U10957 ( .A(n10988), .B(n10989), .Z(n10987) );
  XNOR U10958 ( .A(y[3908]), .B(x[3908]), .Z(n10989) );
  XNOR U10959 ( .A(y[3909]), .B(x[3909]), .Z(n10988) );
  AND U10960 ( .A(n10990), .B(n10991), .Z(n10986) );
  XNOR U10961 ( .A(y[3910]), .B(x[3910]), .Z(n10991) );
  XNOR U10962 ( .A(y[3911]), .B(x[3911]), .Z(n10990) );
  AND U10963 ( .A(n10992), .B(n10993), .Z(n10976) );
  AND U10964 ( .A(n10994), .B(n10995), .Z(n10993) );
  AND U10965 ( .A(n10996), .B(n10997), .Z(n10995) );
  XNOR U10966 ( .A(y[3912]), .B(x[3912]), .Z(n10997) );
  XNOR U10967 ( .A(y[3913]), .B(x[3913]), .Z(n10996) );
  AND U10968 ( .A(n10998), .B(n10999), .Z(n10994) );
  XNOR U10969 ( .A(y[3914]), .B(x[3914]), .Z(n10999) );
  XNOR U10970 ( .A(y[3915]), .B(x[3915]), .Z(n10998) );
  AND U10971 ( .A(n11000), .B(n11001), .Z(n10992) );
  AND U10972 ( .A(n11002), .B(n11003), .Z(n11001) );
  XNOR U10973 ( .A(y[3916]), .B(x[3916]), .Z(n11003) );
  XNOR U10974 ( .A(y[3917]), .B(x[3917]), .Z(n11002) );
  AND U10975 ( .A(n11004), .B(n11005), .Z(n11000) );
  XNOR U10976 ( .A(y[3918]), .B(x[3918]), .Z(n11005) );
  XNOR U10977 ( .A(y[3919]), .B(x[3919]), .Z(n11004) );
  AND U10978 ( .A(n11006), .B(n11007), .Z(n10974) );
  AND U10979 ( .A(n11008), .B(n11009), .Z(n11007) );
  AND U10980 ( .A(n11010), .B(n11011), .Z(n11009) );
  AND U10981 ( .A(n11012), .B(n11013), .Z(n11011) );
  XNOR U10982 ( .A(y[3920]), .B(x[3920]), .Z(n11013) );
  XNOR U10983 ( .A(y[3921]), .B(x[3921]), .Z(n11012) );
  AND U10984 ( .A(n11014), .B(n11015), .Z(n11010) );
  XNOR U10985 ( .A(y[3922]), .B(x[3922]), .Z(n11015) );
  XNOR U10986 ( .A(y[3923]), .B(x[3923]), .Z(n11014) );
  AND U10987 ( .A(n11016), .B(n11017), .Z(n11008) );
  AND U10988 ( .A(n11018), .B(n11019), .Z(n11017) );
  XNOR U10989 ( .A(y[3924]), .B(x[3924]), .Z(n11019) );
  XNOR U10990 ( .A(y[3925]), .B(x[3925]), .Z(n11018) );
  AND U10991 ( .A(n11020), .B(n11021), .Z(n11016) );
  XNOR U10992 ( .A(y[3926]), .B(x[3926]), .Z(n11021) );
  XNOR U10993 ( .A(y[3927]), .B(x[3927]), .Z(n11020) );
  AND U10994 ( .A(n11022), .B(n11023), .Z(n11006) );
  AND U10995 ( .A(n11024), .B(n11025), .Z(n11023) );
  AND U10996 ( .A(n11026), .B(n11027), .Z(n11025) );
  XNOR U10997 ( .A(y[3928]), .B(x[3928]), .Z(n11027) );
  XNOR U10998 ( .A(y[3929]), .B(x[3929]), .Z(n11026) );
  AND U10999 ( .A(n11028), .B(n11029), .Z(n11024) );
  XNOR U11000 ( .A(y[3930]), .B(x[3930]), .Z(n11029) );
  XNOR U11001 ( .A(y[3931]), .B(x[3931]), .Z(n11028) );
  AND U11002 ( .A(n11030), .B(n11031), .Z(n11022) );
  AND U11003 ( .A(n11032), .B(n11033), .Z(n11031) );
  XNOR U11004 ( .A(y[3932]), .B(x[3932]), .Z(n11033) );
  XNOR U11005 ( .A(y[3933]), .B(x[3933]), .Z(n11032) );
  AND U11006 ( .A(n11034), .B(n11035), .Z(n11030) );
  XNOR U11007 ( .A(y[3934]), .B(x[3934]), .Z(n11035) );
  XNOR U11008 ( .A(y[3935]), .B(x[3935]), .Z(n11034) );
  AND U11009 ( .A(n11036), .B(n11037), .Z(n10972) );
  AND U11010 ( .A(n11038), .B(n11039), .Z(n11037) );
  AND U11011 ( .A(n11040), .B(n11041), .Z(n11039) );
  AND U11012 ( .A(n11042), .B(n11043), .Z(n11041) );
  AND U11013 ( .A(n11044), .B(n11045), .Z(n11043) );
  XNOR U11014 ( .A(y[3936]), .B(x[3936]), .Z(n11045) );
  XNOR U11015 ( .A(y[3937]), .B(x[3937]), .Z(n11044) );
  AND U11016 ( .A(n11046), .B(n11047), .Z(n11042) );
  XNOR U11017 ( .A(y[3938]), .B(x[3938]), .Z(n11047) );
  XNOR U11018 ( .A(y[3939]), .B(x[3939]), .Z(n11046) );
  AND U11019 ( .A(n11048), .B(n11049), .Z(n11040) );
  AND U11020 ( .A(n11050), .B(n11051), .Z(n11049) );
  XNOR U11021 ( .A(y[3940]), .B(x[3940]), .Z(n11051) );
  XNOR U11022 ( .A(y[3941]), .B(x[3941]), .Z(n11050) );
  AND U11023 ( .A(n11052), .B(n11053), .Z(n11048) );
  XNOR U11024 ( .A(y[3942]), .B(x[3942]), .Z(n11053) );
  XNOR U11025 ( .A(y[3943]), .B(x[3943]), .Z(n11052) );
  AND U11026 ( .A(n11054), .B(n11055), .Z(n11038) );
  AND U11027 ( .A(n11056), .B(n11057), .Z(n11055) );
  AND U11028 ( .A(n11058), .B(n11059), .Z(n11057) );
  XNOR U11029 ( .A(y[3944]), .B(x[3944]), .Z(n11059) );
  XNOR U11030 ( .A(y[3945]), .B(x[3945]), .Z(n11058) );
  AND U11031 ( .A(n11060), .B(n11061), .Z(n11056) );
  XNOR U11032 ( .A(y[3946]), .B(x[3946]), .Z(n11061) );
  XNOR U11033 ( .A(y[3947]), .B(x[3947]), .Z(n11060) );
  AND U11034 ( .A(n11062), .B(n11063), .Z(n11054) );
  AND U11035 ( .A(n11064), .B(n11065), .Z(n11063) );
  XNOR U11036 ( .A(y[3948]), .B(x[3948]), .Z(n11065) );
  XNOR U11037 ( .A(y[3949]), .B(x[3949]), .Z(n11064) );
  AND U11038 ( .A(n11066), .B(n11067), .Z(n11062) );
  XNOR U11039 ( .A(y[3950]), .B(x[3950]), .Z(n11067) );
  XNOR U11040 ( .A(y[3951]), .B(x[3951]), .Z(n11066) );
  AND U11041 ( .A(n11068), .B(n11069), .Z(n11036) );
  AND U11042 ( .A(n11070), .B(n11071), .Z(n11069) );
  AND U11043 ( .A(n11072), .B(n11073), .Z(n11071) );
  AND U11044 ( .A(n11074), .B(n11075), .Z(n11073) );
  XNOR U11045 ( .A(y[3952]), .B(x[3952]), .Z(n11075) );
  XNOR U11046 ( .A(y[3953]), .B(x[3953]), .Z(n11074) );
  AND U11047 ( .A(n11076), .B(n11077), .Z(n11072) );
  XNOR U11048 ( .A(y[3954]), .B(x[3954]), .Z(n11077) );
  XNOR U11049 ( .A(y[3955]), .B(x[3955]), .Z(n11076) );
  AND U11050 ( .A(n11078), .B(n11079), .Z(n11070) );
  AND U11051 ( .A(n11080), .B(n11081), .Z(n11079) );
  XNOR U11052 ( .A(y[3956]), .B(x[3956]), .Z(n11081) );
  XNOR U11053 ( .A(y[3957]), .B(x[3957]), .Z(n11080) );
  AND U11054 ( .A(n11082), .B(n11083), .Z(n11078) );
  XNOR U11055 ( .A(y[3958]), .B(x[3958]), .Z(n11083) );
  XNOR U11056 ( .A(y[3959]), .B(x[3959]), .Z(n11082) );
  AND U11057 ( .A(n11084), .B(n11085), .Z(n11068) );
  AND U11058 ( .A(n11086), .B(n11087), .Z(n11085) );
  AND U11059 ( .A(n11088), .B(n11089), .Z(n11087) );
  XNOR U11060 ( .A(y[3960]), .B(x[3960]), .Z(n11089) );
  XNOR U11061 ( .A(y[3961]), .B(x[3961]), .Z(n11088) );
  AND U11062 ( .A(n11090), .B(n11091), .Z(n11086) );
  XNOR U11063 ( .A(y[3962]), .B(x[3962]), .Z(n11091) );
  XNOR U11064 ( .A(y[3963]), .B(x[3963]), .Z(n11090) );
  AND U11065 ( .A(n11092), .B(n11093), .Z(n11084) );
  AND U11066 ( .A(n11094), .B(n11095), .Z(n11093) );
  XNOR U11067 ( .A(y[3964]), .B(x[3964]), .Z(n11095) );
  XNOR U11068 ( .A(y[3965]), .B(x[3965]), .Z(n11094) );
  AND U11069 ( .A(n11096), .B(n11097), .Z(n11092) );
  XNOR U11070 ( .A(y[3966]), .B(x[3966]), .Z(n11097) );
  XNOR U11071 ( .A(y[3967]), .B(x[3967]), .Z(n11096) );
  AND U11072 ( .A(n11098), .B(n11099), .Z(n10842) );
  AND U11073 ( .A(n11100), .B(n11101), .Z(n11099) );
  AND U11074 ( .A(n11102), .B(n11103), .Z(n11101) );
  AND U11075 ( .A(n11104), .B(n11105), .Z(n11103) );
  AND U11076 ( .A(n11106), .B(n11107), .Z(n11105) );
  AND U11077 ( .A(n11108), .B(n11109), .Z(n11107) );
  AND U11078 ( .A(n11110), .B(n11111), .Z(n11109) );
  XNOR U11079 ( .A(y[3968]), .B(x[3968]), .Z(n11111) );
  XNOR U11080 ( .A(y[3969]), .B(x[3969]), .Z(n11110) );
  AND U11081 ( .A(n11112), .B(n11113), .Z(n11108) );
  XNOR U11082 ( .A(y[3970]), .B(x[3970]), .Z(n11113) );
  XNOR U11083 ( .A(y[3971]), .B(x[3971]), .Z(n11112) );
  AND U11084 ( .A(n11114), .B(n11115), .Z(n11106) );
  AND U11085 ( .A(n11116), .B(n11117), .Z(n11115) );
  XNOR U11086 ( .A(y[3972]), .B(x[3972]), .Z(n11117) );
  XNOR U11087 ( .A(y[3973]), .B(x[3973]), .Z(n11116) );
  AND U11088 ( .A(n11118), .B(n11119), .Z(n11114) );
  XNOR U11089 ( .A(y[3974]), .B(x[3974]), .Z(n11119) );
  XNOR U11090 ( .A(y[3975]), .B(x[3975]), .Z(n11118) );
  AND U11091 ( .A(n11120), .B(n11121), .Z(n11104) );
  AND U11092 ( .A(n11122), .B(n11123), .Z(n11121) );
  AND U11093 ( .A(n11124), .B(n11125), .Z(n11123) );
  XNOR U11094 ( .A(y[3976]), .B(x[3976]), .Z(n11125) );
  XNOR U11095 ( .A(y[3977]), .B(x[3977]), .Z(n11124) );
  AND U11096 ( .A(n11126), .B(n11127), .Z(n11122) );
  XNOR U11097 ( .A(y[3978]), .B(x[3978]), .Z(n11127) );
  XNOR U11098 ( .A(y[3979]), .B(x[3979]), .Z(n11126) );
  AND U11099 ( .A(n11128), .B(n11129), .Z(n11120) );
  AND U11100 ( .A(n11130), .B(n11131), .Z(n11129) );
  XNOR U11101 ( .A(y[3980]), .B(x[3980]), .Z(n11131) );
  XNOR U11102 ( .A(y[3981]), .B(x[3981]), .Z(n11130) );
  AND U11103 ( .A(n11132), .B(n11133), .Z(n11128) );
  XNOR U11104 ( .A(y[3982]), .B(x[3982]), .Z(n11133) );
  XNOR U11105 ( .A(y[3983]), .B(x[3983]), .Z(n11132) );
  AND U11106 ( .A(n11134), .B(n11135), .Z(n11102) );
  AND U11107 ( .A(n11136), .B(n11137), .Z(n11135) );
  AND U11108 ( .A(n11138), .B(n11139), .Z(n11137) );
  AND U11109 ( .A(n11140), .B(n11141), .Z(n11139) );
  XNOR U11110 ( .A(y[3984]), .B(x[3984]), .Z(n11141) );
  XNOR U11111 ( .A(y[3985]), .B(x[3985]), .Z(n11140) );
  AND U11112 ( .A(n11142), .B(n11143), .Z(n11138) );
  XNOR U11113 ( .A(y[3986]), .B(x[3986]), .Z(n11143) );
  XNOR U11114 ( .A(y[3987]), .B(x[3987]), .Z(n11142) );
  AND U11115 ( .A(n11144), .B(n11145), .Z(n11136) );
  AND U11116 ( .A(n11146), .B(n11147), .Z(n11145) );
  XNOR U11117 ( .A(y[3988]), .B(x[3988]), .Z(n11147) );
  XNOR U11118 ( .A(y[3989]), .B(x[3989]), .Z(n11146) );
  AND U11119 ( .A(n11148), .B(n11149), .Z(n11144) );
  XNOR U11120 ( .A(y[3990]), .B(x[3990]), .Z(n11149) );
  XNOR U11121 ( .A(y[3991]), .B(x[3991]), .Z(n11148) );
  AND U11122 ( .A(n11150), .B(n11151), .Z(n11134) );
  AND U11123 ( .A(n11152), .B(n11153), .Z(n11151) );
  AND U11124 ( .A(n11154), .B(n11155), .Z(n11153) );
  XNOR U11125 ( .A(y[3992]), .B(x[3992]), .Z(n11155) );
  XNOR U11126 ( .A(y[3993]), .B(x[3993]), .Z(n11154) );
  AND U11127 ( .A(n11156), .B(n11157), .Z(n11152) );
  XNOR U11128 ( .A(y[3994]), .B(x[3994]), .Z(n11157) );
  XNOR U11129 ( .A(y[3995]), .B(x[3995]), .Z(n11156) );
  AND U11130 ( .A(n11158), .B(n11159), .Z(n11150) );
  AND U11131 ( .A(n11160), .B(n11161), .Z(n11159) );
  XNOR U11132 ( .A(y[3996]), .B(x[3996]), .Z(n11161) );
  XNOR U11133 ( .A(y[3997]), .B(x[3997]), .Z(n11160) );
  AND U11134 ( .A(n11162), .B(n11163), .Z(n11158) );
  XNOR U11135 ( .A(y[3998]), .B(x[3998]), .Z(n11163) );
  XNOR U11136 ( .A(y[3999]), .B(x[3999]), .Z(n11162) );
  AND U11137 ( .A(n11164), .B(n11165), .Z(n11100) );
  AND U11138 ( .A(n11166), .B(n11167), .Z(n11165) );
  AND U11139 ( .A(n11168), .B(n11169), .Z(n11167) );
  AND U11140 ( .A(n11170), .B(n11171), .Z(n11169) );
  AND U11141 ( .A(n11172), .B(n11173), .Z(n11171) );
  XNOR U11142 ( .A(y[4000]), .B(x[4000]), .Z(n11173) );
  XNOR U11143 ( .A(y[4001]), .B(x[4001]), .Z(n11172) );
  AND U11144 ( .A(n11174), .B(n11175), .Z(n11170) );
  XNOR U11145 ( .A(y[4002]), .B(x[4002]), .Z(n11175) );
  XNOR U11146 ( .A(y[4003]), .B(x[4003]), .Z(n11174) );
  AND U11147 ( .A(n11176), .B(n11177), .Z(n11168) );
  AND U11148 ( .A(n11178), .B(n11179), .Z(n11177) );
  XNOR U11149 ( .A(y[4004]), .B(x[4004]), .Z(n11179) );
  XNOR U11150 ( .A(y[4005]), .B(x[4005]), .Z(n11178) );
  AND U11151 ( .A(n11180), .B(n11181), .Z(n11176) );
  XNOR U11152 ( .A(y[4006]), .B(x[4006]), .Z(n11181) );
  XNOR U11153 ( .A(y[4007]), .B(x[4007]), .Z(n11180) );
  AND U11154 ( .A(n11182), .B(n11183), .Z(n11166) );
  AND U11155 ( .A(n11184), .B(n11185), .Z(n11183) );
  AND U11156 ( .A(n11186), .B(n11187), .Z(n11185) );
  XNOR U11157 ( .A(y[4008]), .B(x[4008]), .Z(n11187) );
  XNOR U11158 ( .A(y[4009]), .B(x[4009]), .Z(n11186) );
  AND U11159 ( .A(n11188), .B(n11189), .Z(n11184) );
  XNOR U11160 ( .A(y[4010]), .B(x[4010]), .Z(n11189) );
  XNOR U11161 ( .A(y[4011]), .B(x[4011]), .Z(n11188) );
  AND U11162 ( .A(n11190), .B(n11191), .Z(n11182) );
  AND U11163 ( .A(n11192), .B(n11193), .Z(n11191) );
  XNOR U11164 ( .A(y[4012]), .B(x[4012]), .Z(n11193) );
  XNOR U11165 ( .A(y[4013]), .B(x[4013]), .Z(n11192) );
  AND U11166 ( .A(n11194), .B(n11195), .Z(n11190) );
  XNOR U11167 ( .A(y[4014]), .B(x[4014]), .Z(n11195) );
  XNOR U11168 ( .A(y[4015]), .B(x[4015]), .Z(n11194) );
  AND U11169 ( .A(n11196), .B(n11197), .Z(n11164) );
  AND U11170 ( .A(n11198), .B(n11199), .Z(n11197) );
  AND U11171 ( .A(n11200), .B(n11201), .Z(n11199) );
  AND U11172 ( .A(n11202), .B(n11203), .Z(n11201) );
  XNOR U11173 ( .A(y[4016]), .B(x[4016]), .Z(n11203) );
  XNOR U11174 ( .A(y[4017]), .B(x[4017]), .Z(n11202) );
  AND U11175 ( .A(n11204), .B(n11205), .Z(n11200) );
  XNOR U11176 ( .A(y[4018]), .B(x[4018]), .Z(n11205) );
  XNOR U11177 ( .A(y[4019]), .B(x[4019]), .Z(n11204) );
  AND U11178 ( .A(n11206), .B(n11207), .Z(n11198) );
  AND U11179 ( .A(n11208), .B(n11209), .Z(n11207) );
  XNOR U11180 ( .A(y[4020]), .B(x[4020]), .Z(n11209) );
  XNOR U11181 ( .A(y[4021]), .B(x[4021]), .Z(n11208) );
  AND U11182 ( .A(n11210), .B(n11211), .Z(n11206) );
  XNOR U11183 ( .A(y[4022]), .B(x[4022]), .Z(n11211) );
  XNOR U11184 ( .A(y[4023]), .B(x[4023]), .Z(n11210) );
  AND U11185 ( .A(n11212), .B(n11213), .Z(n11196) );
  AND U11186 ( .A(n11214), .B(n11215), .Z(n11213) );
  AND U11187 ( .A(n11216), .B(n11217), .Z(n11215) );
  XNOR U11188 ( .A(y[4024]), .B(x[4024]), .Z(n11217) );
  XNOR U11189 ( .A(y[4025]), .B(x[4025]), .Z(n11216) );
  AND U11190 ( .A(n11218), .B(n11219), .Z(n11214) );
  XNOR U11191 ( .A(y[4026]), .B(x[4026]), .Z(n11219) );
  XNOR U11192 ( .A(y[4027]), .B(x[4027]), .Z(n11218) );
  AND U11193 ( .A(n11220), .B(n11221), .Z(n11212) );
  AND U11194 ( .A(n11222), .B(n11223), .Z(n11221) );
  XNOR U11195 ( .A(y[4028]), .B(x[4028]), .Z(n11223) );
  XNOR U11196 ( .A(y[4029]), .B(x[4029]), .Z(n11222) );
  AND U11197 ( .A(n11224), .B(n11225), .Z(n11220) );
  XNOR U11198 ( .A(y[4030]), .B(x[4030]), .Z(n11225) );
  XNOR U11199 ( .A(y[4031]), .B(x[4031]), .Z(n11224) );
  AND U11200 ( .A(n11226), .B(n11227), .Z(n11098) );
  AND U11201 ( .A(n11228), .B(n11229), .Z(n11227) );
  AND U11202 ( .A(n11230), .B(n11231), .Z(n11229) );
  AND U11203 ( .A(n11232), .B(n11233), .Z(n11231) );
  AND U11204 ( .A(n11234), .B(n11235), .Z(n11233) );
  AND U11205 ( .A(n11236), .B(n11237), .Z(n11235) );
  XNOR U11206 ( .A(y[4032]), .B(x[4032]), .Z(n11237) );
  XNOR U11207 ( .A(y[4033]), .B(x[4033]), .Z(n11236) );
  AND U11208 ( .A(n11238), .B(n11239), .Z(n11234) );
  XNOR U11209 ( .A(y[4034]), .B(x[4034]), .Z(n11239) );
  XNOR U11210 ( .A(y[4035]), .B(x[4035]), .Z(n11238) );
  AND U11211 ( .A(n11240), .B(n11241), .Z(n11232) );
  AND U11212 ( .A(n11242), .B(n11243), .Z(n11241) );
  XNOR U11213 ( .A(y[4036]), .B(x[4036]), .Z(n11243) );
  XNOR U11214 ( .A(y[4037]), .B(x[4037]), .Z(n11242) );
  AND U11215 ( .A(n11244), .B(n11245), .Z(n11240) );
  XNOR U11216 ( .A(y[4038]), .B(x[4038]), .Z(n11245) );
  XNOR U11217 ( .A(y[4039]), .B(x[4039]), .Z(n11244) );
  AND U11218 ( .A(n11246), .B(n11247), .Z(n11230) );
  AND U11219 ( .A(n11248), .B(n11249), .Z(n11247) );
  AND U11220 ( .A(n11250), .B(n11251), .Z(n11249) );
  XNOR U11221 ( .A(y[4040]), .B(x[4040]), .Z(n11251) );
  XNOR U11222 ( .A(y[4041]), .B(x[4041]), .Z(n11250) );
  AND U11223 ( .A(n11252), .B(n11253), .Z(n11248) );
  XNOR U11224 ( .A(y[4042]), .B(x[4042]), .Z(n11253) );
  XNOR U11225 ( .A(y[4043]), .B(x[4043]), .Z(n11252) );
  AND U11226 ( .A(n11254), .B(n11255), .Z(n11246) );
  AND U11227 ( .A(n11256), .B(n11257), .Z(n11255) );
  XNOR U11228 ( .A(y[4044]), .B(x[4044]), .Z(n11257) );
  XNOR U11229 ( .A(y[4045]), .B(x[4045]), .Z(n11256) );
  AND U11230 ( .A(n11258), .B(n11259), .Z(n11254) );
  XNOR U11231 ( .A(y[4046]), .B(x[4046]), .Z(n11259) );
  XNOR U11232 ( .A(y[4047]), .B(x[4047]), .Z(n11258) );
  AND U11233 ( .A(n11260), .B(n11261), .Z(n11228) );
  AND U11234 ( .A(n11262), .B(n11263), .Z(n11261) );
  AND U11235 ( .A(n11264), .B(n11265), .Z(n11263) );
  AND U11236 ( .A(n11266), .B(n11267), .Z(n11265) );
  XNOR U11237 ( .A(y[4048]), .B(x[4048]), .Z(n11267) );
  XNOR U11238 ( .A(y[4049]), .B(x[4049]), .Z(n11266) );
  AND U11239 ( .A(n11268), .B(n11269), .Z(n11264) );
  XNOR U11240 ( .A(y[4050]), .B(x[4050]), .Z(n11269) );
  XNOR U11241 ( .A(y[4051]), .B(x[4051]), .Z(n11268) );
  AND U11242 ( .A(n11270), .B(n11271), .Z(n11262) );
  AND U11243 ( .A(n11272), .B(n11273), .Z(n11271) );
  XNOR U11244 ( .A(y[4052]), .B(x[4052]), .Z(n11273) );
  XNOR U11245 ( .A(y[4053]), .B(x[4053]), .Z(n11272) );
  AND U11246 ( .A(n11274), .B(n11275), .Z(n11270) );
  XNOR U11247 ( .A(y[4054]), .B(x[4054]), .Z(n11275) );
  XNOR U11248 ( .A(y[4055]), .B(x[4055]), .Z(n11274) );
  AND U11249 ( .A(n11276), .B(n11277), .Z(n11260) );
  AND U11250 ( .A(n11278), .B(n11279), .Z(n11277) );
  AND U11251 ( .A(n11280), .B(n11281), .Z(n11279) );
  XNOR U11252 ( .A(y[4056]), .B(x[4056]), .Z(n11281) );
  XNOR U11253 ( .A(y[4057]), .B(x[4057]), .Z(n11280) );
  AND U11254 ( .A(n11282), .B(n11283), .Z(n11278) );
  XNOR U11255 ( .A(y[4058]), .B(x[4058]), .Z(n11283) );
  XNOR U11256 ( .A(y[4059]), .B(x[4059]), .Z(n11282) );
  AND U11257 ( .A(n11284), .B(n11285), .Z(n11276) );
  AND U11258 ( .A(n11286), .B(n11287), .Z(n11285) );
  XNOR U11259 ( .A(y[4060]), .B(x[4060]), .Z(n11287) );
  XNOR U11260 ( .A(y[4061]), .B(x[4061]), .Z(n11286) );
  AND U11261 ( .A(n11288), .B(n11289), .Z(n11284) );
  XNOR U11262 ( .A(y[4062]), .B(x[4062]), .Z(n11289) );
  XNOR U11263 ( .A(y[4063]), .B(x[4063]), .Z(n11288) );
  AND U11264 ( .A(n11290), .B(n11291), .Z(n11226) );
  AND U11265 ( .A(n11292), .B(n11293), .Z(n11291) );
  AND U11266 ( .A(n11294), .B(n11295), .Z(n11293) );
  AND U11267 ( .A(n11296), .B(n11297), .Z(n11295) );
  AND U11268 ( .A(n11298), .B(n11299), .Z(n11297) );
  XNOR U11269 ( .A(y[4064]), .B(x[4064]), .Z(n11299) );
  XNOR U11270 ( .A(y[4065]), .B(x[4065]), .Z(n11298) );
  AND U11271 ( .A(n11300), .B(n11301), .Z(n11296) );
  XNOR U11272 ( .A(y[4066]), .B(x[4066]), .Z(n11301) );
  XNOR U11273 ( .A(y[4067]), .B(x[4067]), .Z(n11300) );
  AND U11274 ( .A(n11302), .B(n11303), .Z(n11294) );
  AND U11275 ( .A(n11304), .B(n11305), .Z(n11303) );
  XNOR U11276 ( .A(y[4068]), .B(x[4068]), .Z(n11305) );
  XNOR U11277 ( .A(y[4069]), .B(x[4069]), .Z(n11304) );
  AND U11278 ( .A(n11306), .B(n11307), .Z(n11302) );
  XNOR U11279 ( .A(y[4070]), .B(x[4070]), .Z(n11307) );
  XNOR U11280 ( .A(y[4071]), .B(x[4071]), .Z(n11306) );
  AND U11281 ( .A(n11308), .B(n11309), .Z(n11292) );
  AND U11282 ( .A(n11310), .B(n11311), .Z(n11309) );
  AND U11283 ( .A(n11312), .B(n11313), .Z(n11311) );
  XNOR U11284 ( .A(y[4072]), .B(x[4072]), .Z(n11313) );
  XNOR U11285 ( .A(y[4073]), .B(x[4073]), .Z(n11312) );
  AND U11286 ( .A(n11314), .B(n11315), .Z(n11310) );
  XNOR U11287 ( .A(y[4074]), .B(x[4074]), .Z(n11315) );
  XNOR U11288 ( .A(y[4075]), .B(x[4075]), .Z(n11314) );
  AND U11289 ( .A(n11316), .B(n11317), .Z(n11308) );
  AND U11290 ( .A(n11318), .B(n11319), .Z(n11317) );
  XNOR U11291 ( .A(y[4076]), .B(x[4076]), .Z(n11319) );
  XNOR U11292 ( .A(y[4077]), .B(x[4077]), .Z(n11318) );
  AND U11293 ( .A(n11320), .B(n11321), .Z(n11316) );
  XNOR U11294 ( .A(y[4078]), .B(x[4078]), .Z(n11321) );
  XNOR U11295 ( .A(y[4079]), .B(x[4079]), .Z(n11320) );
  AND U11296 ( .A(n11322), .B(n11323), .Z(n11290) );
  AND U11297 ( .A(n11324), .B(n11325), .Z(n11323) );
  AND U11298 ( .A(n11326), .B(n11327), .Z(n11325) );
  AND U11299 ( .A(n11328), .B(n11329), .Z(n11327) );
  XNOR U11300 ( .A(y[4080]), .B(x[4080]), .Z(n11329) );
  XNOR U11301 ( .A(y[4081]), .B(x[4081]), .Z(n11328) );
  AND U11302 ( .A(n11330), .B(n11331), .Z(n11326) );
  XNOR U11303 ( .A(y[4082]), .B(x[4082]), .Z(n11331) );
  XNOR U11304 ( .A(y[4083]), .B(x[4083]), .Z(n11330) );
  AND U11305 ( .A(n11332), .B(n11333), .Z(n11324) );
  AND U11306 ( .A(n11334), .B(n11335), .Z(n11333) );
  XNOR U11307 ( .A(y[4084]), .B(x[4084]), .Z(n11335) );
  XNOR U11308 ( .A(y[4085]), .B(x[4085]), .Z(n11334) );
  AND U11309 ( .A(n11336), .B(n11337), .Z(n11332) );
  XNOR U11310 ( .A(y[4086]), .B(x[4086]), .Z(n11337) );
  XNOR U11311 ( .A(y[4087]), .B(x[4087]), .Z(n11336) );
  AND U11312 ( .A(n11338), .B(n11339), .Z(n11322) );
  AND U11313 ( .A(n11340), .B(n11341), .Z(n11339) );
  AND U11314 ( .A(n11342), .B(n11343), .Z(n11341) );
  XNOR U11315 ( .A(y[4088]), .B(x[4088]), .Z(n11343) );
  XNOR U11316 ( .A(y[4089]), .B(x[4089]), .Z(n11342) );
  AND U11317 ( .A(n11344), .B(n11345), .Z(n11340) );
  XNOR U11318 ( .A(y[4090]), .B(x[4090]), .Z(n11345) );
  XNOR U11319 ( .A(y[4091]), .B(x[4091]), .Z(n11344) );
  AND U11320 ( .A(n11346), .B(n11347), .Z(n11338) );
  AND U11321 ( .A(n11348), .B(n11349), .Z(n11347) );
  XNOR U11322 ( .A(y[4092]), .B(x[4092]), .Z(n11349) );
  XNOR U11323 ( .A(y[4093]), .B(x[4093]), .Z(n11348) );
  AND U11324 ( .A(n11350), .B(n11351), .Z(n11346) );
  XNOR U11325 ( .A(y[4094]), .B(x[4094]), .Z(n11351) );
  XNOR U11326 ( .A(y[4095]), .B(x[4095]), .Z(n11350) );
  AND U11327 ( .A(n11352), .B(n11353), .Z(n10840) );
  AND U11328 ( .A(n11354), .B(n11355), .Z(n11353) );
  AND U11329 ( .A(n11356), .B(n11357), .Z(n11355) );
  AND U11330 ( .A(n11358), .B(n11359), .Z(n11357) );
  AND U11331 ( .A(n11360), .B(n11361), .Z(n11359) );
  AND U11332 ( .A(n11362), .B(n11363), .Z(n11361) );
  AND U11333 ( .A(n11364), .B(n11365), .Z(n11363) );
  AND U11334 ( .A(n11366), .B(n11367), .Z(n11365) );
  XNOR U11335 ( .A(y[3584]), .B(x[3584]), .Z(n11367) );
  XNOR U11336 ( .A(y[3587]), .B(x[3587]), .Z(n11366) );
  AND U11337 ( .A(n11368), .B(n11369), .Z(n11364) );
  XNOR U11338 ( .A(y[3585]), .B(x[3585]), .Z(n11369) );
  XNOR U11339 ( .A(y[3586]), .B(x[3586]), .Z(n11368) );
  AND U11340 ( .A(n11370), .B(n11371), .Z(n11362) );
  AND U11341 ( .A(n11372), .B(n11373), .Z(n11371) );
  XNOR U11342 ( .A(y[3588]), .B(x[3588]), .Z(n11373) );
  XNOR U11343 ( .A(y[3589]), .B(x[3589]), .Z(n11372) );
  AND U11344 ( .A(n11374), .B(n11375), .Z(n11370) );
  XNOR U11345 ( .A(y[3590]), .B(x[3590]), .Z(n11375) );
  XNOR U11346 ( .A(y[3591]), .B(x[3591]), .Z(n11374) );
  AND U11347 ( .A(n11376), .B(n11377), .Z(n11360) );
  AND U11348 ( .A(n11378), .B(n11379), .Z(n11377) );
  AND U11349 ( .A(n11380), .B(n11381), .Z(n11379) );
  XNOR U11350 ( .A(y[3592]), .B(x[3592]), .Z(n11381) );
  XNOR U11351 ( .A(y[3593]), .B(x[3593]), .Z(n11380) );
  AND U11352 ( .A(n11382), .B(n11383), .Z(n11378) );
  XNOR U11353 ( .A(y[3594]), .B(x[3594]), .Z(n11383) );
  XNOR U11354 ( .A(y[3595]), .B(x[3595]), .Z(n11382) );
  AND U11355 ( .A(n11384), .B(n11385), .Z(n11376) );
  AND U11356 ( .A(n11386), .B(n11387), .Z(n11385) );
  XNOR U11357 ( .A(y[3596]), .B(x[3596]), .Z(n11387) );
  XNOR U11358 ( .A(y[3597]), .B(x[3597]), .Z(n11386) );
  AND U11359 ( .A(n11388), .B(n11389), .Z(n11384) );
  XNOR U11360 ( .A(y[3598]), .B(x[3598]), .Z(n11389) );
  XNOR U11361 ( .A(y[3599]), .B(x[3599]), .Z(n11388) );
  AND U11362 ( .A(n11390), .B(n11391), .Z(n11358) );
  AND U11363 ( .A(n11392), .B(n11393), .Z(n11391) );
  AND U11364 ( .A(n11394), .B(n11395), .Z(n11393) );
  AND U11365 ( .A(n11396), .B(n11397), .Z(n11395) );
  XNOR U11366 ( .A(y[3600]), .B(x[3600]), .Z(n11397) );
  XNOR U11367 ( .A(y[3601]), .B(x[3601]), .Z(n11396) );
  AND U11368 ( .A(n11398), .B(n11399), .Z(n11394) );
  XNOR U11369 ( .A(y[3602]), .B(x[3602]), .Z(n11399) );
  XNOR U11370 ( .A(y[3603]), .B(x[3603]), .Z(n11398) );
  AND U11371 ( .A(n11400), .B(n11401), .Z(n11392) );
  AND U11372 ( .A(n11402), .B(n11403), .Z(n11401) );
  XNOR U11373 ( .A(y[3604]), .B(x[3604]), .Z(n11403) );
  XNOR U11374 ( .A(y[3605]), .B(x[3605]), .Z(n11402) );
  AND U11375 ( .A(n11404), .B(n11405), .Z(n11400) );
  XNOR U11376 ( .A(y[3606]), .B(x[3606]), .Z(n11405) );
  XNOR U11377 ( .A(y[3607]), .B(x[3607]), .Z(n11404) );
  AND U11378 ( .A(n11406), .B(n11407), .Z(n11390) );
  AND U11379 ( .A(n11408), .B(n11409), .Z(n11407) );
  AND U11380 ( .A(n11410), .B(n11411), .Z(n11409) );
  XNOR U11381 ( .A(y[3608]), .B(x[3608]), .Z(n11411) );
  XNOR U11382 ( .A(y[3609]), .B(x[3609]), .Z(n11410) );
  AND U11383 ( .A(n11412), .B(n11413), .Z(n11408) );
  XNOR U11384 ( .A(y[3610]), .B(x[3610]), .Z(n11413) );
  XNOR U11385 ( .A(y[3611]), .B(x[3611]), .Z(n11412) );
  AND U11386 ( .A(n11414), .B(n11415), .Z(n11406) );
  AND U11387 ( .A(n11416), .B(n11417), .Z(n11415) );
  XNOR U11388 ( .A(y[3612]), .B(x[3612]), .Z(n11417) );
  XNOR U11389 ( .A(y[3613]), .B(x[3613]), .Z(n11416) );
  AND U11390 ( .A(n11418), .B(n11419), .Z(n11414) );
  XNOR U11391 ( .A(y[3614]), .B(x[3614]), .Z(n11419) );
  XNOR U11392 ( .A(y[3615]), .B(x[3615]), .Z(n11418) );
  AND U11393 ( .A(n11420), .B(n11421), .Z(n11356) );
  AND U11394 ( .A(n11422), .B(n11423), .Z(n11421) );
  AND U11395 ( .A(n11424), .B(n11425), .Z(n11423) );
  AND U11396 ( .A(n11426), .B(n11427), .Z(n11425) );
  AND U11397 ( .A(n11428), .B(n11429), .Z(n11427) );
  XNOR U11398 ( .A(y[3616]), .B(x[3616]), .Z(n11429) );
  XNOR U11399 ( .A(y[3617]), .B(x[3617]), .Z(n11428) );
  AND U11400 ( .A(n11430), .B(n11431), .Z(n11426) );
  XNOR U11401 ( .A(y[3618]), .B(x[3618]), .Z(n11431) );
  XNOR U11402 ( .A(y[3619]), .B(x[3619]), .Z(n11430) );
  AND U11403 ( .A(n11432), .B(n11433), .Z(n11424) );
  AND U11404 ( .A(n11434), .B(n11435), .Z(n11433) );
  XNOR U11405 ( .A(y[3620]), .B(x[3620]), .Z(n11435) );
  XNOR U11406 ( .A(y[3621]), .B(x[3621]), .Z(n11434) );
  AND U11407 ( .A(n11436), .B(n11437), .Z(n11432) );
  XNOR U11408 ( .A(y[3622]), .B(x[3622]), .Z(n11437) );
  XNOR U11409 ( .A(y[3623]), .B(x[3623]), .Z(n11436) );
  AND U11410 ( .A(n11438), .B(n11439), .Z(n11422) );
  AND U11411 ( .A(n11440), .B(n11441), .Z(n11439) );
  AND U11412 ( .A(n11442), .B(n11443), .Z(n11441) );
  XNOR U11413 ( .A(y[3624]), .B(x[3624]), .Z(n11443) );
  XNOR U11414 ( .A(y[3625]), .B(x[3625]), .Z(n11442) );
  AND U11415 ( .A(n11444), .B(n11445), .Z(n11440) );
  XNOR U11416 ( .A(y[3626]), .B(x[3626]), .Z(n11445) );
  XNOR U11417 ( .A(y[3627]), .B(x[3627]), .Z(n11444) );
  AND U11418 ( .A(n11446), .B(n11447), .Z(n11438) );
  AND U11419 ( .A(n11448), .B(n11449), .Z(n11447) );
  XNOR U11420 ( .A(y[3628]), .B(x[3628]), .Z(n11449) );
  XNOR U11421 ( .A(y[3629]), .B(x[3629]), .Z(n11448) );
  AND U11422 ( .A(n11450), .B(n11451), .Z(n11446) );
  XNOR U11423 ( .A(y[3630]), .B(x[3630]), .Z(n11451) );
  XNOR U11424 ( .A(y[3631]), .B(x[3631]), .Z(n11450) );
  AND U11425 ( .A(n11452), .B(n11453), .Z(n11420) );
  AND U11426 ( .A(n11454), .B(n11455), .Z(n11453) );
  AND U11427 ( .A(n11456), .B(n11457), .Z(n11455) );
  AND U11428 ( .A(n11458), .B(n11459), .Z(n11457) );
  XNOR U11429 ( .A(y[3632]), .B(x[3632]), .Z(n11459) );
  XNOR U11430 ( .A(y[3633]), .B(x[3633]), .Z(n11458) );
  AND U11431 ( .A(n11460), .B(n11461), .Z(n11456) );
  XNOR U11432 ( .A(y[3634]), .B(x[3634]), .Z(n11461) );
  XNOR U11433 ( .A(y[3635]), .B(x[3635]), .Z(n11460) );
  AND U11434 ( .A(n11462), .B(n11463), .Z(n11454) );
  AND U11435 ( .A(n11464), .B(n11465), .Z(n11463) );
  XNOR U11436 ( .A(y[3636]), .B(x[3636]), .Z(n11465) );
  XNOR U11437 ( .A(y[3637]), .B(x[3637]), .Z(n11464) );
  AND U11438 ( .A(n11466), .B(n11467), .Z(n11462) );
  XNOR U11439 ( .A(y[3638]), .B(x[3638]), .Z(n11467) );
  XNOR U11440 ( .A(y[3639]), .B(x[3639]), .Z(n11466) );
  AND U11441 ( .A(n11468), .B(n11469), .Z(n11452) );
  AND U11442 ( .A(n11470), .B(n11471), .Z(n11469) );
  AND U11443 ( .A(n11472), .B(n11473), .Z(n11471) );
  XNOR U11444 ( .A(y[3640]), .B(x[3640]), .Z(n11473) );
  XNOR U11445 ( .A(y[3641]), .B(x[3641]), .Z(n11472) );
  AND U11446 ( .A(n11474), .B(n11475), .Z(n11470) );
  XNOR U11447 ( .A(y[3642]), .B(x[3642]), .Z(n11475) );
  XNOR U11448 ( .A(y[3643]), .B(x[3643]), .Z(n11474) );
  AND U11449 ( .A(n11476), .B(n11477), .Z(n11468) );
  AND U11450 ( .A(n11478), .B(n11479), .Z(n11477) );
  XNOR U11451 ( .A(y[3644]), .B(x[3644]), .Z(n11479) );
  XNOR U11452 ( .A(y[3645]), .B(x[3645]), .Z(n11478) );
  AND U11453 ( .A(n11480), .B(n11481), .Z(n11476) );
  XNOR U11454 ( .A(y[3646]), .B(x[3646]), .Z(n11481) );
  XNOR U11455 ( .A(y[3647]), .B(x[3647]), .Z(n11480) );
  AND U11456 ( .A(n11482), .B(n11483), .Z(n11354) );
  AND U11457 ( .A(n11484), .B(n11485), .Z(n11483) );
  AND U11458 ( .A(n11486), .B(n11487), .Z(n11485) );
  AND U11459 ( .A(n11488), .B(n11489), .Z(n11487) );
  AND U11460 ( .A(n11490), .B(n11491), .Z(n11489) );
  AND U11461 ( .A(n11492), .B(n11493), .Z(n11491) );
  XNOR U11462 ( .A(y[3648]), .B(x[3648]), .Z(n11493) );
  XNOR U11463 ( .A(y[3649]), .B(x[3649]), .Z(n11492) );
  AND U11464 ( .A(n11494), .B(n11495), .Z(n11490) );
  XNOR U11465 ( .A(y[3650]), .B(x[3650]), .Z(n11495) );
  XNOR U11466 ( .A(y[3651]), .B(x[3651]), .Z(n11494) );
  AND U11467 ( .A(n11496), .B(n11497), .Z(n11488) );
  AND U11468 ( .A(n11498), .B(n11499), .Z(n11497) );
  XNOR U11469 ( .A(y[3652]), .B(x[3652]), .Z(n11499) );
  XNOR U11470 ( .A(y[3653]), .B(x[3653]), .Z(n11498) );
  AND U11471 ( .A(n11500), .B(n11501), .Z(n11496) );
  XNOR U11472 ( .A(y[3654]), .B(x[3654]), .Z(n11501) );
  XNOR U11473 ( .A(y[3655]), .B(x[3655]), .Z(n11500) );
  AND U11474 ( .A(n11502), .B(n11503), .Z(n11486) );
  AND U11475 ( .A(n11504), .B(n11505), .Z(n11503) );
  AND U11476 ( .A(n11506), .B(n11507), .Z(n11505) );
  XNOR U11477 ( .A(y[3656]), .B(x[3656]), .Z(n11507) );
  XNOR U11478 ( .A(y[3657]), .B(x[3657]), .Z(n11506) );
  AND U11479 ( .A(n11508), .B(n11509), .Z(n11504) );
  XNOR U11480 ( .A(y[3658]), .B(x[3658]), .Z(n11509) );
  XNOR U11481 ( .A(y[3659]), .B(x[3659]), .Z(n11508) );
  AND U11482 ( .A(n11510), .B(n11511), .Z(n11502) );
  AND U11483 ( .A(n11512), .B(n11513), .Z(n11511) );
  XNOR U11484 ( .A(y[3660]), .B(x[3660]), .Z(n11513) );
  XNOR U11485 ( .A(y[3661]), .B(x[3661]), .Z(n11512) );
  AND U11486 ( .A(n11514), .B(n11515), .Z(n11510) );
  XNOR U11487 ( .A(y[3662]), .B(x[3662]), .Z(n11515) );
  XNOR U11488 ( .A(y[3663]), .B(x[3663]), .Z(n11514) );
  AND U11489 ( .A(n11516), .B(n11517), .Z(n11484) );
  AND U11490 ( .A(n11518), .B(n11519), .Z(n11517) );
  AND U11491 ( .A(n11520), .B(n11521), .Z(n11519) );
  AND U11492 ( .A(n11522), .B(n11523), .Z(n11521) );
  XNOR U11493 ( .A(y[3664]), .B(x[3664]), .Z(n11523) );
  XNOR U11494 ( .A(y[3665]), .B(x[3665]), .Z(n11522) );
  AND U11495 ( .A(n11524), .B(n11525), .Z(n11520) );
  XNOR U11496 ( .A(y[3666]), .B(x[3666]), .Z(n11525) );
  XNOR U11497 ( .A(y[3667]), .B(x[3667]), .Z(n11524) );
  AND U11498 ( .A(n11526), .B(n11527), .Z(n11518) );
  AND U11499 ( .A(n11528), .B(n11529), .Z(n11527) );
  XNOR U11500 ( .A(y[3668]), .B(x[3668]), .Z(n11529) );
  XNOR U11501 ( .A(y[3669]), .B(x[3669]), .Z(n11528) );
  AND U11502 ( .A(n11530), .B(n11531), .Z(n11526) );
  XNOR U11503 ( .A(y[3670]), .B(x[3670]), .Z(n11531) );
  XNOR U11504 ( .A(y[3671]), .B(x[3671]), .Z(n11530) );
  AND U11505 ( .A(n11532), .B(n11533), .Z(n11516) );
  AND U11506 ( .A(n11534), .B(n11535), .Z(n11533) );
  AND U11507 ( .A(n11536), .B(n11537), .Z(n11535) );
  XNOR U11508 ( .A(y[3672]), .B(x[3672]), .Z(n11537) );
  XNOR U11509 ( .A(y[3673]), .B(x[3673]), .Z(n11536) );
  AND U11510 ( .A(n11538), .B(n11539), .Z(n11534) );
  XNOR U11511 ( .A(y[3674]), .B(x[3674]), .Z(n11539) );
  XNOR U11512 ( .A(y[3675]), .B(x[3675]), .Z(n11538) );
  AND U11513 ( .A(n11540), .B(n11541), .Z(n11532) );
  AND U11514 ( .A(n11542), .B(n11543), .Z(n11541) );
  XNOR U11515 ( .A(y[3676]), .B(x[3676]), .Z(n11543) );
  XNOR U11516 ( .A(y[3677]), .B(x[3677]), .Z(n11542) );
  AND U11517 ( .A(n11544), .B(n11545), .Z(n11540) );
  XNOR U11518 ( .A(y[3678]), .B(x[3678]), .Z(n11545) );
  XNOR U11519 ( .A(y[3679]), .B(x[3679]), .Z(n11544) );
  AND U11520 ( .A(n11546), .B(n11547), .Z(n11482) );
  AND U11521 ( .A(n11548), .B(n11549), .Z(n11547) );
  AND U11522 ( .A(n11550), .B(n11551), .Z(n11549) );
  AND U11523 ( .A(n11552), .B(n11553), .Z(n11551) );
  AND U11524 ( .A(n11554), .B(n11555), .Z(n11553) );
  XNOR U11525 ( .A(y[3680]), .B(x[3680]), .Z(n11555) );
  XNOR U11526 ( .A(y[3681]), .B(x[3681]), .Z(n11554) );
  AND U11527 ( .A(n11556), .B(n11557), .Z(n11552) );
  XNOR U11528 ( .A(y[3682]), .B(x[3682]), .Z(n11557) );
  XNOR U11529 ( .A(y[3683]), .B(x[3683]), .Z(n11556) );
  AND U11530 ( .A(n11558), .B(n11559), .Z(n11550) );
  AND U11531 ( .A(n11560), .B(n11561), .Z(n11559) );
  XNOR U11532 ( .A(y[3684]), .B(x[3684]), .Z(n11561) );
  XNOR U11533 ( .A(y[3685]), .B(x[3685]), .Z(n11560) );
  AND U11534 ( .A(n11562), .B(n11563), .Z(n11558) );
  XNOR U11535 ( .A(y[3686]), .B(x[3686]), .Z(n11563) );
  XNOR U11536 ( .A(y[3687]), .B(x[3687]), .Z(n11562) );
  AND U11537 ( .A(n11564), .B(n11565), .Z(n11548) );
  AND U11538 ( .A(n11566), .B(n11567), .Z(n11565) );
  AND U11539 ( .A(n11568), .B(n11569), .Z(n11567) );
  XNOR U11540 ( .A(y[3688]), .B(x[3688]), .Z(n11569) );
  XNOR U11541 ( .A(y[3689]), .B(x[3689]), .Z(n11568) );
  AND U11542 ( .A(n11570), .B(n11571), .Z(n11566) );
  XNOR U11543 ( .A(y[3690]), .B(x[3690]), .Z(n11571) );
  XNOR U11544 ( .A(y[3691]), .B(x[3691]), .Z(n11570) );
  AND U11545 ( .A(n11572), .B(n11573), .Z(n11564) );
  AND U11546 ( .A(n11574), .B(n11575), .Z(n11573) );
  XNOR U11547 ( .A(y[3692]), .B(x[3692]), .Z(n11575) );
  XNOR U11548 ( .A(y[3693]), .B(x[3693]), .Z(n11574) );
  AND U11549 ( .A(n11576), .B(n11577), .Z(n11572) );
  XNOR U11550 ( .A(y[3694]), .B(x[3694]), .Z(n11577) );
  XNOR U11551 ( .A(y[3695]), .B(x[3695]), .Z(n11576) );
  AND U11552 ( .A(n11578), .B(n11579), .Z(n11546) );
  AND U11553 ( .A(n11580), .B(n11581), .Z(n11579) );
  AND U11554 ( .A(n11582), .B(n11583), .Z(n11581) );
  AND U11555 ( .A(n11584), .B(n11585), .Z(n11583) );
  XNOR U11556 ( .A(y[3696]), .B(x[3696]), .Z(n11585) );
  XNOR U11557 ( .A(y[3697]), .B(x[3697]), .Z(n11584) );
  AND U11558 ( .A(n11586), .B(n11587), .Z(n11582) );
  XNOR U11559 ( .A(y[3698]), .B(x[3698]), .Z(n11587) );
  XNOR U11560 ( .A(y[3699]), .B(x[3699]), .Z(n11586) );
  AND U11561 ( .A(n11588), .B(n11589), .Z(n11580) );
  AND U11562 ( .A(n11590), .B(n11591), .Z(n11589) );
  XNOR U11563 ( .A(y[3700]), .B(x[3700]), .Z(n11591) );
  XNOR U11564 ( .A(y[3701]), .B(x[3701]), .Z(n11590) );
  AND U11565 ( .A(n11592), .B(n11593), .Z(n11588) );
  XNOR U11566 ( .A(y[3702]), .B(x[3702]), .Z(n11593) );
  XNOR U11567 ( .A(y[3703]), .B(x[3703]), .Z(n11592) );
  AND U11568 ( .A(n11594), .B(n11595), .Z(n11578) );
  AND U11569 ( .A(n11596), .B(n11597), .Z(n11595) );
  AND U11570 ( .A(n11598), .B(n11599), .Z(n11597) );
  XNOR U11571 ( .A(y[3704]), .B(x[3704]), .Z(n11599) );
  XNOR U11572 ( .A(y[3705]), .B(x[3705]), .Z(n11598) );
  AND U11573 ( .A(n11600), .B(n11601), .Z(n11596) );
  XNOR U11574 ( .A(y[3706]), .B(x[3706]), .Z(n11601) );
  XNOR U11575 ( .A(y[3707]), .B(x[3707]), .Z(n11600) );
  AND U11576 ( .A(n11602), .B(n11603), .Z(n11594) );
  AND U11577 ( .A(n11604), .B(n11605), .Z(n11603) );
  XNOR U11578 ( .A(y[3708]), .B(x[3708]), .Z(n11605) );
  XNOR U11579 ( .A(y[3709]), .B(x[3709]), .Z(n11604) );
  AND U11580 ( .A(n11606), .B(n11607), .Z(n11602) );
  XNOR U11581 ( .A(y[3710]), .B(x[3710]), .Z(n11607) );
  XNOR U11582 ( .A(y[3711]), .B(x[3711]), .Z(n11606) );
  AND U11583 ( .A(n11608), .B(n11609), .Z(n11352) );
  AND U11584 ( .A(n11610), .B(n11611), .Z(n11609) );
  AND U11585 ( .A(n11612), .B(n11613), .Z(n11611) );
  AND U11586 ( .A(n11614), .B(n11615), .Z(n11613) );
  AND U11587 ( .A(n11616), .B(n11617), .Z(n11615) );
  AND U11588 ( .A(n11618), .B(n11619), .Z(n11617) );
  AND U11589 ( .A(n11620), .B(n11621), .Z(n11619) );
  XNOR U11590 ( .A(y[3712]), .B(x[3712]), .Z(n11621) );
  XNOR U11591 ( .A(y[3713]), .B(x[3713]), .Z(n11620) );
  AND U11592 ( .A(n11622), .B(n11623), .Z(n11618) );
  XNOR U11593 ( .A(y[3714]), .B(x[3714]), .Z(n11623) );
  XNOR U11594 ( .A(y[3715]), .B(x[3715]), .Z(n11622) );
  AND U11595 ( .A(n11624), .B(n11625), .Z(n11616) );
  AND U11596 ( .A(n11626), .B(n11627), .Z(n11625) );
  XNOR U11597 ( .A(y[3716]), .B(x[3716]), .Z(n11627) );
  XNOR U11598 ( .A(y[3717]), .B(x[3717]), .Z(n11626) );
  AND U11599 ( .A(n11628), .B(n11629), .Z(n11624) );
  XNOR U11600 ( .A(y[3718]), .B(x[3718]), .Z(n11629) );
  XNOR U11601 ( .A(y[3719]), .B(x[3719]), .Z(n11628) );
  AND U11602 ( .A(n11630), .B(n11631), .Z(n11614) );
  AND U11603 ( .A(n11632), .B(n11633), .Z(n11631) );
  AND U11604 ( .A(n11634), .B(n11635), .Z(n11633) );
  XNOR U11605 ( .A(y[3720]), .B(x[3720]), .Z(n11635) );
  XNOR U11606 ( .A(y[3721]), .B(x[3721]), .Z(n11634) );
  AND U11607 ( .A(n11636), .B(n11637), .Z(n11632) );
  XNOR U11608 ( .A(y[3722]), .B(x[3722]), .Z(n11637) );
  XNOR U11609 ( .A(y[3723]), .B(x[3723]), .Z(n11636) );
  AND U11610 ( .A(n11638), .B(n11639), .Z(n11630) );
  AND U11611 ( .A(n11640), .B(n11641), .Z(n11639) );
  XNOR U11612 ( .A(y[3724]), .B(x[3724]), .Z(n11641) );
  XNOR U11613 ( .A(y[3725]), .B(x[3725]), .Z(n11640) );
  AND U11614 ( .A(n11642), .B(n11643), .Z(n11638) );
  XNOR U11615 ( .A(y[3726]), .B(x[3726]), .Z(n11643) );
  XNOR U11616 ( .A(y[3727]), .B(x[3727]), .Z(n11642) );
  AND U11617 ( .A(n11644), .B(n11645), .Z(n11612) );
  AND U11618 ( .A(n11646), .B(n11647), .Z(n11645) );
  AND U11619 ( .A(n11648), .B(n11649), .Z(n11647) );
  AND U11620 ( .A(n11650), .B(n11651), .Z(n11649) );
  XNOR U11621 ( .A(y[3728]), .B(x[3728]), .Z(n11651) );
  XNOR U11622 ( .A(y[3729]), .B(x[3729]), .Z(n11650) );
  AND U11623 ( .A(n11652), .B(n11653), .Z(n11648) );
  XNOR U11624 ( .A(y[3730]), .B(x[3730]), .Z(n11653) );
  XNOR U11625 ( .A(y[3731]), .B(x[3731]), .Z(n11652) );
  AND U11626 ( .A(n11654), .B(n11655), .Z(n11646) );
  AND U11627 ( .A(n11656), .B(n11657), .Z(n11655) );
  XNOR U11628 ( .A(y[3732]), .B(x[3732]), .Z(n11657) );
  XNOR U11629 ( .A(y[3733]), .B(x[3733]), .Z(n11656) );
  AND U11630 ( .A(n11658), .B(n11659), .Z(n11654) );
  XNOR U11631 ( .A(y[3734]), .B(x[3734]), .Z(n11659) );
  XNOR U11632 ( .A(y[3735]), .B(x[3735]), .Z(n11658) );
  AND U11633 ( .A(n11660), .B(n11661), .Z(n11644) );
  AND U11634 ( .A(n11662), .B(n11663), .Z(n11661) );
  AND U11635 ( .A(n11664), .B(n11665), .Z(n11663) );
  XNOR U11636 ( .A(y[3736]), .B(x[3736]), .Z(n11665) );
  XNOR U11637 ( .A(y[3737]), .B(x[3737]), .Z(n11664) );
  AND U11638 ( .A(n11666), .B(n11667), .Z(n11662) );
  XNOR U11639 ( .A(y[3738]), .B(x[3738]), .Z(n11667) );
  XNOR U11640 ( .A(y[3739]), .B(x[3739]), .Z(n11666) );
  AND U11641 ( .A(n11668), .B(n11669), .Z(n11660) );
  AND U11642 ( .A(n11670), .B(n11671), .Z(n11669) );
  XNOR U11643 ( .A(y[3740]), .B(x[3740]), .Z(n11671) );
  XNOR U11644 ( .A(y[3741]), .B(x[3741]), .Z(n11670) );
  AND U11645 ( .A(n11672), .B(n11673), .Z(n11668) );
  XNOR U11646 ( .A(y[3742]), .B(x[3742]), .Z(n11673) );
  XNOR U11647 ( .A(y[3743]), .B(x[3743]), .Z(n11672) );
  AND U11648 ( .A(n11674), .B(n11675), .Z(n11610) );
  AND U11649 ( .A(n11676), .B(n11677), .Z(n11675) );
  AND U11650 ( .A(n11678), .B(n11679), .Z(n11677) );
  AND U11651 ( .A(n11680), .B(n11681), .Z(n11679) );
  AND U11652 ( .A(n11682), .B(n11683), .Z(n11681) );
  XNOR U11653 ( .A(y[3744]), .B(x[3744]), .Z(n11683) );
  XNOR U11654 ( .A(y[3745]), .B(x[3745]), .Z(n11682) );
  AND U11655 ( .A(n11684), .B(n11685), .Z(n11680) );
  XNOR U11656 ( .A(y[3746]), .B(x[3746]), .Z(n11685) );
  XNOR U11657 ( .A(y[3747]), .B(x[3747]), .Z(n11684) );
  AND U11658 ( .A(n11686), .B(n11687), .Z(n11678) );
  AND U11659 ( .A(n11688), .B(n11689), .Z(n11687) );
  XNOR U11660 ( .A(y[3748]), .B(x[3748]), .Z(n11689) );
  XNOR U11661 ( .A(y[3749]), .B(x[3749]), .Z(n11688) );
  AND U11662 ( .A(n11690), .B(n11691), .Z(n11686) );
  XNOR U11663 ( .A(y[3750]), .B(x[3750]), .Z(n11691) );
  XNOR U11664 ( .A(y[3751]), .B(x[3751]), .Z(n11690) );
  AND U11665 ( .A(n11692), .B(n11693), .Z(n11676) );
  AND U11666 ( .A(n11694), .B(n11695), .Z(n11693) );
  AND U11667 ( .A(n11696), .B(n11697), .Z(n11695) );
  XNOR U11668 ( .A(y[3752]), .B(x[3752]), .Z(n11697) );
  XNOR U11669 ( .A(y[3753]), .B(x[3753]), .Z(n11696) );
  AND U11670 ( .A(n11698), .B(n11699), .Z(n11694) );
  XNOR U11671 ( .A(y[3754]), .B(x[3754]), .Z(n11699) );
  XNOR U11672 ( .A(y[3755]), .B(x[3755]), .Z(n11698) );
  AND U11673 ( .A(n11700), .B(n11701), .Z(n11692) );
  AND U11674 ( .A(n11702), .B(n11703), .Z(n11701) );
  XNOR U11675 ( .A(y[3756]), .B(x[3756]), .Z(n11703) );
  XNOR U11676 ( .A(y[3757]), .B(x[3757]), .Z(n11702) );
  AND U11677 ( .A(n11704), .B(n11705), .Z(n11700) );
  XNOR U11678 ( .A(y[3758]), .B(x[3758]), .Z(n11705) );
  XNOR U11679 ( .A(y[3759]), .B(x[3759]), .Z(n11704) );
  AND U11680 ( .A(n11706), .B(n11707), .Z(n11674) );
  AND U11681 ( .A(n11708), .B(n11709), .Z(n11707) );
  AND U11682 ( .A(n11710), .B(n11711), .Z(n11709) );
  AND U11683 ( .A(n11712), .B(n11713), .Z(n11711) );
  XNOR U11684 ( .A(y[3760]), .B(x[3760]), .Z(n11713) );
  XNOR U11685 ( .A(y[3761]), .B(x[3761]), .Z(n11712) );
  AND U11686 ( .A(n11714), .B(n11715), .Z(n11710) );
  XNOR U11687 ( .A(y[3762]), .B(x[3762]), .Z(n11715) );
  XNOR U11688 ( .A(y[3763]), .B(x[3763]), .Z(n11714) );
  AND U11689 ( .A(n11716), .B(n11717), .Z(n11708) );
  AND U11690 ( .A(n11718), .B(n11719), .Z(n11717) );
  XNOR U11691 ( .A(y[3764]), .B(x[3764]), .Z(n11719) );
  XNOR U11692 ( .A(y[3765]), .B(x[3765]), .Z(n11718) );
  AND U11693 ( .A(n11720), .B(n11721), .Z(n11716) );
  XNOR U11694 ( .A(y[3766]), .B(x[3766]), .Z(n11721) );
  XNOR U11695 ( .A(y[3767]), .B(x[3767]), .Z(n11720) );
  AND U11696 ( .A(n11722), .B(n11723), .Z(n11706) );
  AND U11697 ( .A(n11724), .B(n11725), .Z(n11723) );
  AND U11698 ( .A(n11726), .B(n11727), .Z(n11725) );
  XNOR U11699 ( .A(y[3768]), .B(x[3768]), .Z(n11727) );
  XNOR U11700 ( .A(y[3769]), .B(x[3769]), .Z(n11726) );
  AND U11701 ( .A(n11728), .B(n11729), .Z(n11724) );
  XNOR U11702 ( .A(y[3770]), .B(x[3770]), .Z(n11729) );
  XNOR U11703 ( .A(y[3771]), .B(x[3771]), .Z(n11728) );
  AND U11704 ( .A(n11730), .B(n11731), .Z(n11722) );
  AND U11705 ( .A(n11732), .B(n11733), .Z(n11731) );
  XNOR U11706 ( .A(y[3772]), .B(x[3772]), .Z(n11733) );
  XNOR U11707 ( .A(y[3773]), .B(x[3773]), .Z(n11732) );
  AND U11708 ( .A(n11734), .B(n11735), .Z(n11730) );
  XNOR U11709 ( .A(y[3774]), .B(x[3774]), .Z(n11735) );
  XNOR U11710 ( .A(y[3775]), .B(x[3775]), .Z(n11734) );
  AND U11711 ( .A(n11736), .B(n11737), .Z(n11608) );
  AND U11712 ( .A(n11738), .B(n11739), .Z(n11737) );
  AND U11713 ( .A(n11740), .B(n11741), .Z(n11739) );
  AND U11714 ( .A(n11742), .B(n11743), .Z(n11741) );
  AND U11715 ( .A(n11744), .B(n11745), .Z(n11743) );
  AND U11716 ( .A(n11746), .B(n11747), .Z(n11745) );
  XNOR U11717 ( .A(y[3776]), .B(x[3776]), .Z(n11747) );
  XNOR U11718 ( .A(y[3777]), .B(x[3777]), .Z(n11746) );
  AND U11719 ( .A(n11748), .B(n11749), .Z(n11744) );
  XNOR U11720 ( .A(y[3778]), .B(x[3778]), .Z(n11749) );
  XNOR U11721 ( .A(y[3779]), .B(x[3779]), .Z(n11748) );
  AND U11722 ( .A(n11750), .B(n11751), .Z(n11742) );
  AND U11723 ( .A(n11752), .B(n11753), .Z(n11751) );
  XNOR U11724 ( .A(y[3780]), .B(x[3780]), .Z(n11753) );
  XNOR U11725 ( .A(y[3781]), .B(x[3781]), .Z(n11752) );
  AND U11726 ( .A(n11754), .B(n11755), .Z(n11750) );
  XNOR U11727 ( .A(y[3782]), .B(x[3782]), .Z(n11755) );
  XNOR U11728 ( .A(y[3783]), .B(x[3783]), .Z(n11754) );
  AND U11729 ( .A(n11756), .B(n11757), .Z(n11740) );
  AND U11730 ( .A(n11758), .B(n11759), .Z(n11757) );
  AND U11731 ( .A(n11760), .B(n11761), .Z(n11759) );
  XNOR U11732 ( .A(y[3784]), .B(x[3784]), .Z(n11761) );
  XNOR U11733 ( .A(y[3785]), .B(x[3785]), .Z(n11760) );
  AND U11734 ( .A(n11762), .B(n11763), .Z(n11758) );
  XNOR U11735 ( .A(y[3786]), .B(x[3786]), .Z(n11763) );
  XNOR U11736 ( .A(y[3787]), .B(x[3787]), .Z(n11762) );
  AND U11737 ( .A(n11764), .B(n11765), .Z(n11756) );
  AND U11738 ( .A(n11766), .B(n11767), .Z(n11765) );
  XNOR U11739 ( .A(y[3788]), .B(x[3788]), .Z(n11767) );
  XNOR U11740 ( .A(y[3789]), .B(x[3789]), .Z(n11766) );
  AND U11741 ( .A(n11768), .B(n11769), .Z(n11764) );
  XNOR U11742 ( .A(y[3790]), .B(x[3790]), .Z(n11769) );
  XNOR U11743 ( .A(y[3791]), .B(x[3791]), .Z(n11768) );
  AND U11744 ( .A(n11770), .B(n11771), .Z(n11738) );
  AND U11745 ( .A(n11772), .B(n11773), .Z(n11771) );
  AND U11746 ( .A(n11774), .B(n11775), .Z(n11773) );
  AND U11747 ( .A(n11776), .B(n11777), .Z(n11775) );
  XNOR U11748 ( .A(y[3792]), .B(x[3792]), .Z(n11777) );
  XNOR U11749 ( .A(y[3793]), .B(x[3793]), .Z(n11776) );
  AND U11750 ( .A(n11778), .B(n11779), .Z(n11774) );
  XNOR U11751 ( .A(y[3794]), .B(x[3794]), .Z(n11779) );
  XNOR U11752 ( .A(y[3795]), .B(x[3795]), .Z(n11778) );
  AND U11753 ( .A(n11780), .B(n11781), .Z(n11772) );
  AND U11754 ( .A(n11782), .B(n11783), .Z(n11781) );
  XNOR U11755 ( .A(y[3796]), .B(x[3796]), .Z(n11783) );
  XNOR U11756 ( .A(y[3797]), .B(x[3797]), .Z(n11782) );
  AND U11757 ( .A(n11784), .B(n11785), .Z(n11780) );
  XNOR U11758 ( .A(y[3798]), .B(x[3798]), .Z(n11785) );
  XNOR U11759 ( .A(y[3799]), .B(x[3799]), .Z(n11784) );
  AND U11760 ( .A(n11786), .B(n11787), .Z(n11770) );
  AND U11761 ( .A(n11788), .B(n11789), .Z(n11787) );
  AND U11762 ( .A(n11790), .B(n11791), .Z(n11789) );
  XNOR U11763 ( .A(y[3800]), .B(x[3800]), .Z(n11791) );
  XNOR U11764 ( .A(y[3801]), .B(x[3801]), .Z(n11790) );
  AND U11765 ( .A(n11792), .B(n11793), .Z(n11788) );
  XNOR U11766 ( .A(y[3802]), .B(x[3802]), .Z(n11793) );
  XNOR U11767 ( .A(y[3803]), .B(x[3803]), .Z(n11792) );
  AND U11768 ( .A(n11794), .B(n11795), .Z(n11786) );
  AND U11769 ( .A(n11796), .B(n11797), .Z(n11795) );
  XNOR U11770 ( .A(y[3804]), .B(x[3804]), .Z(n11797) );
  XNOR U11771 ( .A(y[3805]), .B(x[3805]), .Z(n11796) );
  AND U11772 ( .A(n11798), .B(n11799), .Z(n11794) );
  XNOR U11773 ( .A(y[3806]), .B(x[3806]), .Z(n11799) );
  XNOR U11774 ( .A(y[3807]), .B(x[3807]), .Z(n11798) );
  AND U11775 ( .A(n11800), .B(n11801), .Z(n11736) );
  AND U11776 ( .A(n11802), .B(n11803), .Z(n11801) );
  AND U11777 ( .A(n11804), .B(n11805), .Z(n11803) );
  AND U11778 ( .A(n11806), .B(n11807), .Z(n11805) );
  AND U11779 ( .A(n11808), .B(n11809), .Z(n11807) );
  XNOR U11780 ( .A(y[3808]), .B(x[3808]), .Z(n11809) );
  XNOR U11781 ( .A(y[3809]), .B(x[3809]), .Z(n11808) );
  AND U11782 ( .A(n11810), .B(n11811), .Z(n11806) );
  XNOR U11783 ( .A(y[3810]), .B(x[3810]), .Z(n11811) );
  XNOR U11784 ( .A(y[3811]), .B(x[3811]), .Z(n11810) );
  AND U11785 ( .A(n11812), .B(n11813), .Z(n11804) );
  AND U11786 ( .A(n11814), .B(n11815), .Z(n11813) );
  XNOR U11787 ( .A(y[3812]), .B(x[3812]), .Z(n11815) );
  XNOR U11788 ( .A(y[3813]), .B(x[3813]), .Z(n11814) );
  AND U11789 ( .A(n11816), .B(n11817), .Z(n11812) );
  XNOR U11790 ( .A(y[3814]), .B(x[3814]), .Z(n11817) );
  XNOR U11791 ( .A(y[3815]), .B(x[3815]), .Z(n11816) );
  AND U11792 ( .A(n11818), .B(n11819), .Z(n11802) );
  AND U11793 ( .A(n11820), .B(n11821), .Z(n11819) );
  AND U11794 ( .A(n11822), .B(n11823), .Z(n11821) );
  XNOR U11795 ( .A(y[3816]), .B(x[3816]), .Z(n11823) );
  XNOR U11796 ( .A(y[3817]), .B(x[3817]), .Z(n11822) );
  AND U11797 ( .A(n11824), .B(n11825), .Z(n11820) );
  XNOR U11798 ( .A(y[3818]), .B(x[3818]), .Z(n11825) );
  XNOR U11799 ( .A(y[3819]), .B(x[3819]), .Z(n11824) );
  AND U11800 ( .A(n11826), .B(n11827), .Z(n11818) );
  AND U11801 ( .A(n11828), .B(n11829), .Z(n11827) );
  XNOR U11802 ( .A(y[3820]), .B(x[3820]), .Z(n11829) );
  XNOR U11803 ( .A(y[3821]), .B(x[3821]), .Z(n11828) );
  AND U11804 ( .A(n11830), .B(n11831), .Z(n11826) );
  XNOR U11805 ( .A(y[3822]), .B(x[3822]), .Z(n11831) );
  XNOR U11806 ( .A(y[3823]), .B(x[3823]), .Z(n11830) );
  AND U11807 ( .A(n11832), .B(n11833), .Z(n11800) );
  AND U11808 ( .A(n11834), .B(n11835), .Z(n11833) );
  AND U11809 ( .A(n11836), .B(n11837), .Z(n11835) );
  AND U11810 ( .A(n11838), .B(n11839), .Z(n11837) );
  XNOR U11811 ( .A(y[3824]), .B(x[3824]), .Z(n11839) );
  XNOR U11812 ( .A(y[3825]), .B(x[3825]), .Z(n11838) );
  AND U11813 ( .A(n11840), .B(n11841), .Z(n11836) );
  XNOR U11814 ( .A(y[3826]), .B(x[3826]), .Z(n11841) );
  XNOR U11815 ( .A(y[3827]), .B(x[3827]), .Z(n11840) );
  AND U11816 ( .A(n11842), .B(n11843), .Z(n11834) );
  AND U11817 ( .A(n11844), .B(n11845), .Z(n11843) );
  XNOR U11818 ( .A(y[3828]), .B(x[3828]), .Z(n11845) );
  XNOR U11819 ( .A(y[3829]), .B(x[3829]), .Z(n11844) );
  AND U11820 ( .A(n11846), .B(n11847), .Z(n11842) );
  XNOR U11821 ( .A(y[3830]), .B(x[3830]), .Z(n11847) );
  XNOR U11822 ( .A(y[3831]), .B(x[3831]), .Z(n11846) );
  AND U11823 ( .A(n11848), .B(n11849), .Z(n11832) );
  AND U11824 ( .A(n11850), .B(n11851), .Z(n11849) );
  AND U11825 ( .A(n11852), .B(n11853), .Z(n11851) );
  XNOR U11826 ( .A(y[3832]), .B(x[3832]), .Z(n11853) );
  XNOR U11827 ( .A(y[3833]), .B(x[3833]), .Z(n11852) );
  AND U11828 ( .A(n11854), .B(n11855), .Z(n11850) );
  XNOR U11829 ( .A(y[3834]), .B(x[3834]), .Z(n11855) );
  XNOR U11830 ( .A(y[3835]), .B(x[3835]), .Z(n11854) );
  AND U11831 ( .A(n11856), .B(n11857), .Z(n11848) );
  AND U11832 ( .A(n11858), .B(n11859), .Z(n11857) );
  XNOR U11833 ( .A(y[3836]), .B(x[3836]), .Z(n11859) );
  XNOR U11834 ( .A(y[3837]), .B(x[3837]), .Z(n11858) );
  AND U11835 ( .A(n11860), .B(n11861), .Z(n11856) );
  XNOR U11836 ( .A(y[3838]), .B(x[3838]), .Z(n11861) );
  XNOR U11837 ( .A(y[3839]), .B(x[3839]), .Z(n11860) );
  AND U11838 ( .A(n11862), .B(n11863), .Z(n8662) );
  AND U11839 ( .A(n11864), .B(n11865), .Z(n11863) );
  AND U11840 ( .A(n11866), .B(n11867), .Z(n11865) );
  XNOR U11841 ( .A(y[2034]), .B(x[2034]), .Z(n11867) );
  XNOR U11842 ( .A(y[2035]), .B(x[2035]), .Z(n11866) );
  AND U11843 ( .A(n11868), .B(n11869), .Z(n11864) );
  XNOR U11844 ( .A(y[2036]), .B(x[2036]), .Z(n11869) );
  XNOR U11845 ( .A(y[2037]), .B(x[2037]), .Z(n11868) );
  AND U11846 ( .A(n11870), .B(n11871), .Z(n11862) );
  AND U11847 ( .A(n11872), .B(n11873), .Z(n11871) );
  XNOR U11848 ( .A(y[2496]), .B(x[2496]), .Z(n11873) );
  XNOR U11849 ( .A(y[2497]), .B(x[2497]), .Z(n11872) );
  AND U11850 ( .A(n11874), .B(n11875), .Z(n11870) );
  XNOR U11851 ( .A(y[2498]), .B(x[2498]), .Z(n11875) );
  XNOR U11852 ( .A(y[2499]), .B(x[2499]), .Z(n11874) );
  AND U11853 ( .A(n11876), .B(n11877), .Z(n8660) );
  AND U11854 ( .A(n11878), .B(n11879), .Z(n11877) );
  AND U11855 ( .A(n11880), .B(n11881), .Z(n11879) );
  AND U11856 ( .A(n11882), .B(n11883), .Z(n11881) );
  XNOR U11857 ( .A(y[2500]), .B(x[2500]), .Z(n11883) );
  XNOR U11858 ( .A(y[2501]), .B(x[2501]), .Z(n11882) );
  AND U11859 ( .A(n11884), .B(n11885), .Z(n11880) );
  XNOR U11860 ( .A(y[2502]), .B(x[2502]), .Z(n11885) );
  XNOR U11861 ( .A(y[2503]), .B(x[2503]), .Z(n11884) );
  AND U11862 ( .A(n11886), .B(n11887), .Z(n11878) );
  AND U11863 ( .A(n11888), .B(n11889), .Z(n11887) );
  XNOR U11864 ( .A(y[2504]), .B(x[2504]), .Z(n11889) );
  XNOR U11865 ( .A(y[2505]), .B(x[2505]), .Z(n11888) );
  AND U11866 ( .A(n11890), .B(n11891), .Z(n11886) );
  XNOR U11867 ( .A(y[2506]), .B(x[2506]), .Z(n11891) );
  XNOR U11868 ( .A(y[2507]), .B(x[2507]), .Z(n11890) );
  AND U11869 ( .A(n11892), .B(n11893), .Z(n11876) );
  AND U11870 ( .A(n11894), .B(n11895), .Z(n11893) );
  AND U11871 ( .A(n11896), .B(n11897), .Z(n11895) );
  XNOR U11872 ( .A(y[2508]), .B(x[2508]), .Z(n11897) );
  XNOR U11873 ( .A(y[2509]), .B(x[2509]), .Z(n11896) );
  AND U11874 ( .A(n11898), .B(n11899), .Z(n11894) );
  XNOR U11875 ( .A(y[2510]), .B(x[2510]), .Z(n11899) );
  XNOR U11876 ( .A(y[2511]), .B(x[2511]), .Z(n11898) );
  AND U11877 ( .A(n11900), .B(n11901), .Z(n11892) );
  XNOR U11878 ( .A(y[2514]), .B(x[2514]), .Z(n11901) );
  AND U11879 ( .A(n11902), .B(n11903), .Z(n11900) );
  XNOR U11880 ( .A(y[2512]), .B(x[2512]), .Z(n11903) );
  XNOR U11881 ( .A(y[2513]), .B(x[2513]), .Z(n11902) );
  AND U11882 ( .A(n11904), .B(n11905), .Z(n8658) );
  AND U11883 ( .A(n11906), .B(n11907), .Z(n11905) );
  AND U11884 ( .A(n11908), .B(n11909), .Z(n11907) );
  AND U11885 ( .A(n11910), .B(n11911), .Z(n11909) );
  AND U11886 ( .A(n11912), .B(n11913), .Z(n11911) );
  XNOR U11887 ( .A(y[2515]), .B(x[2515]), .Z(n11913) );
  XNOR U11888 ( .A(y[2516]), .B(x[2516]), .Z(n11912) );
  AND U11889 ( .A(n11914), .B(n11915), .Z(n11910) );
  XNOR U11890 ( .A(y[2517]), .B(x[2517]), .Z(n11915) );
  XNOR U11891 ( .A(y[2518]), .B(x[2518]), .Z(n11914) );
  AND U11892 ( .A(n11916), .B(n11917), .Z(n11908) );
  AND U11893 ( .A(n11918), .B(n11919), .Z(n11917) );
  XNOR U11894 ( .A(y[2519]), .B(x[2519]), .Z(n11919) );
  XNOR U11895 ( .A(y[2520]), .B(x[2520]), .Z(n11918) );
  AND U11896 ( .A(n11920), .B(n11921), .Z(n11916) );
  XNOR U11897 ( .A(y[2521]), .B(x[2521]), .Z(n11921) );
  XNOR U11898 ( .A(y[2522]), .B(x[2522]), .Z(n11920) );
  AND U11899 ( .A(n11922), .B(n11923), .Z(n11906) );
  AND U11900 ( .A(n11924), .B(n11925), .Z(n11923) );
  AND U11901 ( .A(n11926), .B(n11927), .Z(n11925) );
  XNOR U11902 ( .A(y[2523]), .B(x[2523]), .Z(n11927) );
  XNOR U11903 ( .A(y[2524]), .B(x[2524]), .Z(n11926) );
  AND U11904 ( .A(n11928), .B(n11929), .Z(n11924) );
  XNOR U11905 ( .A(y[2525]), .B(x[2525]), .Z(n11929) );
  XNOR U11906 ( .A(y[2526]), .B(x[2526]), .Z(n11928) );
  AND U11907 ( .A(n11930), .B(n11931), .Z(n11922) );
  XNOR U11908 ( .A(y[2433]), .B(x[2433]), .Z(n11931) );
  AND U11909 ( .A(n11932), .B(n11933), .Z(n11930) );
  XNOR U11910 ( .A(y[2527]), .B(x[2527]), .Z(n11933) );
  XNOR U11911 ( .A(y[2432]), .B(x[2432]), .Z(n11932) );
  AND U11912 ( .A(n11934), .B(n11935), .Z(n11904) );
  AND U11913 ( .A(n11936), .B(n11937), .Z(n11935) );
  AND U11914 ( .A(n11938), .B(n11939), .Z(n11937) );
  AND U11915 ( .A(n11940), .B(n11941), .Z(n11939) );
  XNOR U11916 ( .A(y[2434]), .B(x[2434]), .Z(n11941) );
  XNOR U11917 ( .A(y[2435]), .B(x[2435]), .Z(n11940) );
  AND U11918 ( .A(n11942), .B(n11943), .Z(n11938) );
  XNOR U11919 ( .A(y[2436]), .B(x[2436]), .Z(n11943) );
  XNOR U11920 ( .A(y[2437]), .B(x[2437]), .Z(n11942) );
  AND U11921 ( .A(n11944), .B(n11945), .Z(n11936) );
  AND U11922 ( .A(n11946), .B(n11947), .Z(n11945) );
  XNOR U11923 ( .A(y[2438]), .B(x[2438]), .Z(n11947) );
  XNOR U11924 ( .A(y[2439]), .B(x[2439]), .Z(n11946) );
  AND U11925 ( .A(n11948), .B(n11949), .Z(n11944) );
  XNOR U11926 ( .A(y[2440]), .B(x[2440]), .Z(n11949) );
  XNOR U11927 ( .A(y[2441]), .B(x[2441]), .Z(n11948) );
  AND U11928 ( .A(n11950), .B(n11951), .Z(n11934) );
  AND U11929 ( .A(n11952), .B(n11953), .Z(n11951) );
  AND U11930 ( .A(n11954), .B(n11955), .Z(n11953) );
  XNOR U11931 ( .A(y[2442]), .B(x[2442]), .Z(n11955) );
  XNOR U11932 ( .A(y[2443]), .B(x[2443]), .Z(n11954) );
  AND U11933 ( .A(n11956), .B(n11957), .Z(n11952) );
  XNOR U11934 ( .A(y[2444]), .B(x[2444]), .Z(n11957) );
  XNOR U11935 ( .A(y[2445]), .B(x[2445]), .Z(n11956) );
  AND U11936 ( .A(n11958), .B(n11959), .Z(n11950) );
  XNOR U11937 ( .A(y[2448]), .B(x[2448]), .Z(n11959) );
  AND U11938 ( .A(n11960), .B(n11961), .Z(n11958) );
  XNOR U11939 ( .A(y[2446]), .B(x[2446]), .Z(n11961) );
  XNOR U11940 ( .A(y[2447]), .B(x[2447]), .Z(n11960) );
  AND U11941 ( .A(n11962), .B(n11963), .Z(n8656) );
  AND U11942 ( .A(n11964), .B(n11965), .Z(n11963) );
  AND U11943 ( .A(n11966), .B(n11967), .Z(n11965) );
  AND U11944 ( .A(n11968), .B(n11969), .Z(n11967) );
  AND U11945 ( .A(n11970), .B(n11971), .Z(n11969) );
  AND U11946 ( .A(n11972), .B(n11973), .Z(n11971) );
  XNOR U11947 ( .A(y[2449]), .B(x[2449]), .Z(n11973) );
  XNOR U11948 ( .A(y[2450]), .B(x[2450]), .Z(n11972) );
  AND U11949 ( .A(n11974), .B(n11975), .Z(n11970) );
  XNOR U11950 ( .A(y[2451]), .B(x[2451]), .Z(n11975) );
  XNOR U11951 ( .A(y[2452]), .B(x[2452]), .Z(n11974) );
  AND U11952 ( .A(n11976), .B(n11977), .Z(n11968) );
  AND U11953 ( .A(n11978), .B(n11979), .Z(n11977) );
  XNOR U11954 ( .A(y[2453]), .B(x[2453]), .Z(n11979) );
  XNOR U11955 ( .A(y[2454]), .B(x[2454]), .Z(n11978) );
  AND U11956 ( .A(n11980), .B(n11981), .Z(n11976) );
  XNOR U11957 ( .A(y[2455]), .B(x[2455]), .Z(n11981) );
  XNOR U11958 ( .A(y[2456]), .B(x[2456]), .Z(n11980) );
  AND U11959 ( .A(n11982), .B(n11983), .Z(n11966) );
  AND U11960 ( .A(n11984), .B(n11985), .Z(n11983) );
  AND U11961 ( .A(n11986), .B(n11987), .Z(n11985) );
  XNOR U11962 ( .A(y[2457]), .B(x[2457]), .Z(n11987) );
  XNOR U11963 ( .A(y[2458]), .B(x[2458]), .Z(n11986) );
  AND U11964 ( .A(n11988), .B(n11989), .Z(n11984) );
  XNOR U11965 ( .A(y[2459]), .B(x[2459]), .Z(n11989) );
  XNOR U11966 ( .A(y[2460]), .B(x[2460]), .Z(n11988) );
  AND U11967 ( .A(n11990), .B(n11991), .Z(n11982) );
  AND U11968 ( .A(n11992), .B(n11993), .Z(n11991) );
  XNOR U11969 ( .A(y[2461]), .B(x[2461]), .Z(n11993) );
  XNOR U11970 ( .A(y[2462]), .B(x[2462]), .Z(n11992) );
  AND U11971 ( .A(n11994), .B(n11995), .Z(n11990) );
  XNOR U11972 ( .A(y[2463]), .B(x[2463]), .Z(n11995) );
  XNOR U11973 ( .A(y[2464]), .B(x[2464]), .Z(n11994) );
  AND U11974 ( .A(n11996), .B(n11997), .Z(n11964) );
  AND U11975 ( .A(n11998), .B(n11999), .Z(n11997) );
  AND U11976 ( .A(n12000), .B(n12001), .Z(n11999) );
  AND U11977 ( .A(n12002), .B(n12003), .Z(n12001) );
  XNOR U11978 ( .A(y[2465]), .B(x[2465]), .Z(n12003) );
  XNOR U11979 ( .A(y[2466]), .B(x[2466]), .Z(n12002) );
  AND U11980 ( .A(n12004), .B(n12005), .Z(n12000) );
  XNOR U11981 ( .A(y[2467]), .B(x[2467]), .Z(n12005) );
  XNOR U11982 ( .A(y[2468]), .B(x[2468]), .Z(n12004) );
  AND U11983 ( .A(n12006), .B(n12007), .Z(n11998) );
  AND U11984 ( .A(n12008), .B(n12009), .Z(n12007) );
  XNOR U11985 ( .A(y[2469]), .B(x[2469]), .Z(n12009) );
  XNOR U11986 ( .A(y[2470]), .B(x[2470]), .Z(n12008) );
  AND U11987 ( .A(n12010), .B(n12011), .Z(n12006) );
  XNOR U11988 ( .A(y[2471]), .B(x[2471]), .Z(n12011) );
  XNOR U11989 ( .A(y[2472]), .B(x[2472]), .Z(n12010) );
  AND U11990 ( .A(n12012), .B(n12013), .Z(n11996) );
  AND U11991 ( .A(n12014), .B(n12015), .Z(n12013) );
  AND U11992 ( .A(n12016), .B(n12017), .Z(n12015) );
  XNOR U11993 ( .A(y[2473]), .B(x[2473]), .Z(n12017) );
  XNOR U11994 ( .A(y[2474]), .B(x[2474]), .Z(n12016) );
  AND U11995 ( .A(n12018), .B(n12019), .Z(n12014) );
  XNOR U11996 ( .A(y[2475]), .B(x[2475]), .Z(n12019) );
  XNOR U11997 ( .A(y[2476]), .B(x[2476]), .Z(n12018) );
  AND U11998 ( .A(n12020), .B(n12021), .Z(n12012) );
  XNOR U11999 ( .A(y[2479]), .B(x[2479]), .Z(n12021) );
  AND U12000 ( .A(n12022), .B(n12023), .Z(n12020) );
  XNOR U12001 ( .A(y[2477]), .B(x[2477]), .Z(n12023) );
  XNOR U12002 ( .A(y[2478]), .B(x[2478]), .Z(n12022) );
  AND U12003 ( .A(n12024), .B(n12025), .Z(n11962) );
  AND U12004 ( .A(n12026), .B(n12027), .Z(n12025) );
  AND U12005 ( .A(n12028), .B(n12029), .Z(n12027) );
  AND U12006 ( .A(n12030), .B(n12031), .Z(n12029) );
  AND U12007 ( .A(n12032), .B(n12033), .Z(n12031) );
  XNOR U12008 ( .A(y[2480]), .B(x[2480]), .Z(n12033) );
  XNOR U12009 ( .A(y[2481]), .B(x[2481]), .Z(n12032) );
  AND U12010 ( .A(n12034), .B(n12035), .Z(n12030) );
  XNOR U12011 ( .A(y[2482]), .B(x[2482]), .Z(n12035) );
  XNOR U12012 ( .A(y[2483]), .B(x[2483]), .Z(n12034) );
  AND U12013 ( .A(n12036), .B(n12037), .Z(n12028) );
  AND U12014 ( .A(n12038), .B(n12039), .Z(n12037) );
  XNOR U12015 ( .A(y[2484]), .B(x[2484]), .Z(n12039) );
  XNOR U12016 ( .A(y[2485]), .B(x[2485]), .Z(n12038) );
  AND U12017 ( .A(n12040), .B(n12041), .Z(n12036) );
  XNOR U12018 ( .A(y[2486]), .B(x[2486]), .Z(n12041) );
  XNOR U12019 ( .A(y[2487]), .B(x[2487]), .Z(n12040) );
  AND U12020 ( .A(n12042), .B(n12043), .Z(n12026) );
  AND U12021 ( .A(n12044), .B(n12045), .Z(n12043) );
  AND U12022 ( .A(n12046), .B(n12047), .Z(n12045) );
  XNOR U12023 ( .A(y[2488]), .B(x[2488]), .Z(n12047) );
  XNOR U12024 ( .A(y[2489]), .B(x[2489]), .Z(n12046) );
  AND U12025 ( .A(n12048), .B(n12049), .Z(n12044) );
  XNOR U12026 ( .A(y[2490]), .B(x[2490]), .Z(n12049) );
  XNOR U12027 ( .A(y[2491]), .B(x[2491]), .Z(n12048) );
  AND U12028 ( .A(n12050), .B(n12051), .Z(n12042) );
  XNOR U12029 ( .A(y[2494]), .B(x[2494]), .Z(n12051) );
  AND U12030 ( .A(n12052), .B(n12053), .Z(n12050) );
  XNOR U12031 ( .A(y[2492]), .B(x[2492]), .Z(n12053) );
  XNOR U12032 ( .A(y[2493]), .B(x[2493]), .Z(n12052) );
  AND U12033 ( .A(n12054), .B(n12055), .Z(n12024) );
  AND U12034 ( .A(n12056), .B(n12057), .Z(n12055) );
  AND U12035 ( .A(n12058), .B(n12059), .Z(n12057) );
  AND U12036 ( .A(n12060), .B(n12061), .Z(n12059) );
  XNOR U12037 ( .A(y[2495]), .B(x[2495]), .Z(n12061) );
  XNOR U12038 ( .A(y[2304]), .B(x[2304]), .Z(n12060) );
  AND U12039 ( .A(n12062), .B(n12063), .Z(n12058) );
  XNOR U12040 ( .A(y[2305]), .B(x[2305]), .Z(n12063) );
  XNOR U12041 ( .A(y[2306]), .B(x[2306]), .Z(n12062) );
  AND U12042 ( .A(n12064), .B(n12065), .Z(n12056) );
  AND U12043 ( .A(n12066), .B(n12067), .Z(n12065) );
  XNOR U12044 ( .A(y[2307]), .B(x[2307]), .Z(n12067) );
  XNOR U12045 ( .A(y[2308]), .B(x[2308]), .Z(n12066) );
  AND U12046 ( .A(n12068), .B(n12069), .Z(n12064) );
  XNOR U12047 ( .A(y[2309]), .B(x[2309]), .Z(n12069) );
  XNOR U12048 ( .A(y[2310]), .B(x[2310]), .Z(n12068) );
  AND U12049 ( .A(n12070), .B(n12071), .Z(n12054) );
  AND U12050 ( .A(n12072), .B(n12073), .Z(n12071) );
  AND U12051 ( .A(n12074), .B(n12075), .Z(n12073) );
  XNOR U12052 ( .A(y[2311]), .B(x[2311]), .Z(n12075) );
  XNOR U12053 ( .A(y[2312]), .B(x[2312]), .Z(n12074) );
  AND U12054 ( .A(n12076), .B(n12077), .Z(n12072) );
  XNOR U12055 ( .A(y[2313]), .B(x[2313]), .Z(n12077) );
  XNOR U12056 ( .A(y[2314]), .B(x[2314]), .Z(n12076) );
  AND U12057 ( .A(n12078), .B(n12079), .Z(n12070) );
  XNOR U12058 ( .A(y[2317]), .B(x[2317]), .Z(n12079) );
  AND U12059 ( .A(n12080), .B(n12081), .Z(n12078) );
  XNOR U12060 ( .A(y[2315]), .B(x[2315]), .Z(n12081) );
  XNOR U12061 ( .A(y[2316]), .B(x[2316]), .Z(n12080) );
  AND U12062 ( .A(n12082), .B(n12083), .Z(n8654) );
  AND U12063 ( .A(n12084), .B(n12085), .Z(n12083) );
  AND U12064 ( .A(n12086), .B(n12087), .Z(n12085) );
  AND U12065 ( .A(n12088), .B(n12089), .Z(n12087) );
  AND U12066 ( .A(n12090), .B(n12091), .Z(n12089) );
  AND U12067 ( .A(n12092), .B(n12093), .Z(n12091) );
  AND U12068 ( .A(n12094), .B(n12095), .Z(n12093) );
  XNOR U12069 ( .A(y[2318]), .B(x[2318]), .Z(n12095) );
  XNOR U12070 ( .A(y[2319]), .B(x[2319]), .Z(n12094) );
  AND U12071 ( .A(n12096), .B(n12097), .Z(n12092) );
  XNOR U12072 ( .A(y[2320]), .B(x[2320]), .Z(n12097) );
  XNOR U12073 ( .A(y[2321]), .B(x[2321]), .Z(n12096) );
  AND U12074 ( .A(n12098), .B(n12099), .Z(n12090) );
  AND U12075 ( .A(n12100), .B(n12101), .Z(n12099) );
  XNOR U12076 ( .A(y[2322]), .B(x[2322]), .Z(n12101) );
  XNOR U12077 ( .A(y[2323]), .B(x[2323]), .Z(n12100) );
  AND U12078 ( .A(n12102), .B(n12103), .Z(n12098) );
  XNOR U12079 ( .A(y[2324]), .B(x[2324]), .Z(n12103) );
  XNOR U12080 ( .A(y[2325]), .B(x[2325]), .Z(n12102) );
  AND U12081 ( .A(n12104), .B(n12105), .Z(n12088) );
  AND U12082 ( .A(n12106), .B(n12107), .Z(n12105) );
  AND U12083 ( .A(n12108), .B(n12109), .Z(n12107) );
  XNOR U12084 ( .A(y[2326]), .B(x[2326]), .Z(n12109) );
  XNOR U12085 ( .A(y[2327]), .B(x[2327]), .Z(n12108) );
  AND U12086 ( .A(n12110), .B(n12111), .Z(n12106) );
  XNOR U12087 ( .A(y[2328]), .B(x[2328]), .Z(n12111) );
  XNOR U12088 ( .A(y[2329]), .B(x[2329]), .Z(n12110) );
  AND U12089 ( .A(n12112), .B(n12113), .Z(n12104) );
  AND U12090 ( .A(n12114), .B(n12115), .Z(n12113) );
  XNOR U12091 ( .A(y[2330]), .B(x[2330]), .Z(n12115) );
  XNOR U12092 ( .A(y[2331]), .B(x[2331]), .Z(n12114) );
  AND U12093 ( .A(n12116), .B(n12117), .Z(n12112) );
  XNOR U12094 ( .A(y[2332]), .B(x[2332]), .Z(n12117) );
  XNOR U12095 ( .A(y[2333]), .B(x[2333]), .Z(n12116) );
  AND U12096 ( .A(n12118), .B(n12119), .Z(n12086) );
  AND U12097 ( .A(n12120), .B(n12121), .Z(n12119) );
  AND U12098 ( .A(n12122), .B(n12123), .Z(n12121) );
  AND U12099 ( .A(n12124), .B(n12125), .Z(n12123) );
  XNOR U12100 ( .A(y[2334]), .B(x[2334]), .Z(n12125) );
  XNOR U12101 ( .A(y[2335]), .B(x[2335]), .Z(n12124) );
  AND U12102 ( .A(n12126), .B(n12127), .Z(n12122) );
  XNOR U12103 ( .A(y[2336]), .B(x[2336]), .Z(n12127) );
  XNOR U12104 ( .A(y[2337]), .B(x[2337]), .Z(n12126) );
  AND U12105 ( .A(n12128), .B(n12129), .Z(n12120) );
  AND U12106 ( .A(n12130), .B(n12131), .Z(n12129) );
  XNOR U12107 ( .A(y[2338]), .B(x[2338]), .Z(n12131) );
  XNOR U12108 ( .A(y[2339]), .B(x[2339]), .Z(n12130) );
  AND U12109 ( .A(n12132), .B(n12133), .Z(n12128) );
  XNOR U12110 ( .A(y[2340]), .B(x[2340]), .Z(n12133) );
  XNOR U12111 ( .A(y[2341]), .B(x[2341]), .Z(n12132) );
  AND U12112 ( .A(n12134), .B(n12135), .Z(n12118) );
  AND U12113 ( .A(n12136), .B(n12137), .Z(n12135) );
  AND U12114 ( .A(n12138), .B(n12139), .Z(n12137) );
  XNOR U12115 ( .A(y[2342]), .B(x[2342]), .Z(n12139) );
  XNOR U12116 ( .A(y[2343]), .B(x[2343]), .Z(n12138) );
  AND U12117 ( .A(n12140), .B(n12141), .Z(n12136) );
  XNOR U12118 ( .A(y[2344]), .B(x[2344]), .Z(n12141) );
  XNOR U12119 ( .A(y[2345]), .B(x[2345]), .Z(n12140) );
  AND U12120 ( .A(n12142), .B(n12143), .Z(n12134) );
  XNOR U12121 ( .A(y[2348]), .B(x[2348]), .Z(n12143) );
  AND U12122 ( .A(n12144), .B(n12145), .Z(n12142) );
  XNOR U12123 ( .A(y[2346]), .B(x[2346]), .Z(n12145) );
  XNOR U12124 ( .A(y[2347]), .B(x[2347]), .Z(n12144) );
  AND U12125 ( .A(n12146), .B(n12147), .Z(n12084) );
  AND U12126 ( .A(n12148), .B(n12149), .Z(n12147) );
  AND U12127 ( .A(n12150), .B(n12151), .Z(n12149) );
  AND U12128 ( .A(n12152), .B(n12153), .Z(n12151) );
  AND U12129 ( .A(n12154), .B(n12155), .Z(n12153) );
  XNOR U12130 ( .A(y[2349]), .B(x[2349]), .Z(n12155) );
  XNOR U12131 ( .A(y[2350]), .B(x[2350]), .Z(n12154) );
  AND U12132 ( .A(n12156), .B(n12157), .Z(n12152) );
  XNOR U12133 ( .A(y[2351]), .B(x[2351]), .Z(n12157) );
  XNOR U12134 ( .A(y[2352]), .B(x[2352]), .Z(n12156) );
  AND U12135 ( .A(n12158), .B(n12159), .Z(n12150) );
  AND U12136 ( .A(n12160), .B(n12161), .Z(n12159) );
  XNOR U12137 ( .A(y[2353]), .B(x[2353]), .Z(n12161) );
  XNOR U12138 ( .A(y[2354]), .B(x[2354]), .Z(n12160) );
  AND U12139 ( .A(n12162), .B(n12163), .Z(n12158) );
  XNOR U12140 ( .A(y[2355]), .B(x[2355]), .Z(n12163) );
  XNOR U12141 ( .A(y[2356]), .B(x[2356]), .Z(n12162) );
  AND U12142 ( .A(n12164), .B(n12165), .Z(n12148) );
  AND U12143 ( .A(n12166), .B(n12167), .Z(n12165) );
  AND U12144 ( .A(n12168), .B(n12169), .Z(n12167) );
  XNOR U12145 ( .A(y[2357]), .B(x[2357]), .Z(n12169) );
  XNOR U12146 ( .A(y[2358]), .B(x[2358]), .Z(n12168) );
  AND U12147 ( .A(n12170), .B(n12171), .Z(n12166) );
  XNOR U12148 ( .A(y[2359]), .B(x[2359]), .Z(n12171) );
  XNOR U12149 ( .A(y[2360]), .B(x[2360]), .Z(n12170) );
  AND U12150 ( .A(n12172), .B(n12173), .Z(n12164) );
  XNOR U12151 ( .A(y[2363]), .B(x[2363]), .Z(n12173) );
  AND U12152 ( .A(n12174), .B(n12175), .Z(n12172) );
  XNOR U12153 ( .A(y[2361]), .B(x[2361]), .Z(n12175) );
  XNOR U12154 ( .A(y[2362]), .B(x[2362]), .Z(n12174) );
  AND U12155 ( .A(n12176), .B(n12177), .Z(n12146) );
  AND U12156 ( .A(n12178), .B(n12179), .Z(n12177) );
  AND U12157 ( .A(n12180), .B(n12181), .Z(n12179) );
  AND U12158 ( .A(n12182), .B(n12183), .Z(n12181) );
  XNOR U12159 ( .A(y[2364]), .B(x[2364]), .Z(n12183) );
  XNOR U12160 ( .A(y[2365]), .B(x[2365]), .Z(n12182) );
  AND U12161 ( .A(n12184), .B(n12185), .Z(n12180) );
  XNOR U12162 ( .A(y[2366]), .B(x[2366]), .Z(n12185) );
  XNOR U12163 ( .A(y[2367]), .B(x[2367]), .Z(n12184) );
  AND U12164 ( .A(n12186), .B(n12187), .Z(n12178) );
  AND U12165 ( .A(n12188), .B(n12189), .Z(n12187) );
  XNOR U12166 ( .A(y[2368]), .B(x[2368]), .Z(n12189) );
  XNOR U12167 ( .A(y[2369]), .B(x[2369]), .Z(n12188) );
  AND U12168 ( .A(n12190), .B(n12191), .Z(n12186) );
  XNOR U12169 ( .A(y[2370]), .B(x[2370]), .Z(n12191) );
  XNOR U12170 ( .A(y[2371]), .B(x[2371]), .Z(n12190) );
  AND U12171 ( .A(n12192), .B(n12193), .Z(n12176) );
  AND U12172 ( .A(n12194), .B(n12195), .Z(n12193) );
  AND U12173 ( .A(n12196), .B(n12197), .Z(n12195) );
  XNOR U12174 ( .A(y[2372]), .B(x[2372]), .Z(n12197) );
  XNOR U12175 ( .A(y[2373]), .B(x[2373]), .Z(n12196) );
  AND U12176 ( .A(n12198), .B(n12199), .Z(n12194) );
  XNOR U12177 ( .A(y[2374]), .B(x[2374]), .Z(n12199) );
  XNOR U12178 ( .A(y[2375]), .B(x[2375]), .Z(n12198) );
  AND U12179 ( .A(n12200), .B(n12201), .Z(n12192) );
  XNOR U12180 ( .A(y[2378]), .B(x[2378]), .Z(n12201) );
  AND U12181 ( .A(n12202), .B(n12203), .Z(n12200) );
  XNOR U12182 ( .A(y[2376]), .B(x[2376]), .Z(n12203) );
  XNOR U12183 ( .A(y[2377]), .B(x[2377]), .Z(n12202) );
  AND U12184 ( .A(n12204), .B(n12205), .Z(n12082) );
  AND U12185 ( .A(n12206), .B(n12207), .Z(n12205) );
  AND U12186 ( .A(n12208), .B(n12209), .Z(n12207) );
  AND U12187 ( .A(n12210), .B(n12211), .Z(n12209) );
  AND U12188 ( .A(n12212), .B(n12213), .Z(n12211) );
  AND U12189 ( .A(n12214), .B(n12215), .Z(n12213) );
  XNOR U12190 ( .A(y[2379]), .B(x[2379]), .Z(n12215) );
  XNOR U12191 ( .A(y[2380]), .B(x[2380]), .Z(n12214) );
  AND U12192 ( .A(n12216), .B(n12217), .Z(n12212) );
  XNOR U12193 ( .A(y[2381]), .B(x[2381]), .Z(n12217) );
  XNOR U12194 ( .A(y[2382]), .B(x[2382]), .Z(n12216) );
  AND U12195 ( .A(n12218), .B(n12219), .Z(n12210) );
  AND U12196 ( .A(n12220), .B(n12221), .Z(n12219) );
  XNOR U12197 ( .A(y[2383]), .B(x[2383]), .Z(n12221) );
  XNOR U12198 ( .A(y[2384]), .B(x[2384]), .Z(n12220) );
  AND U12199 ( .A(n12222), .B(n12223), .Z(n12218) );
  XNOR U12200 ( .A(y[2385]), .B(x[2385]), .Z(n12223) );
  XNOR U12201 ( .A(y[2386]), .B(x[2386]), .Z(n12222) );
  AND U12202 ( .A(n12224), .B(n12225), .Z(n12208) );
  AND U12203 ( .A(n12226), .B(n12227), .Z(n12225) );
  AND U12204 ( .A(n12228), .B(n12229), .Z(n12227) );
  XNOR U12205 ( .A(y[2387]), .B(x[2387]), .Z(n12229) );
  XNOR U12206 ( .A(y[2388]), .B(x[2388]), .Z(n12228) );
  AND U12207 ( .A(n12230), .B(n12231), .Z(n12226) );
  XNOR U12208 ( .A(y[2389]), .B(x[2389]), .Z(n12231) );
  XNOR U12209 ( .A(y[2390]), .B(x[2390]), .Z(n12230) );
  AND U12210 ( .A(n12232), .B(n12233), .Z(n12224) );
  XNOR U12211 ( .A(y[2393]), .B(x[2393]), .Z(n12233) );
  AND U12212 ( .A(n12234), .B(n12235), .Z(n12232) );
  XNOR U12213 ( .A(y[2391]), .B(x[2391]), .Z(n12235) );
  XNOR U12214 ( .A(y[2392]), .B(x[2392]), .Z(n12234) );
  AND U12215 ( .A(n12236), .B(n12237), .Z(n12206) );
  AND U12216 ( .A(n12238), .B(n12239), .Z(n12237) );
  AND U12217 ( .A(n12240), .B(n12241), .Z(n12239) );
  AND U12218 ( .A(n12242), .B(n12243), .Z(n12241) );
  XNOR U12219 ( .A(y[2394]), .B(x[2394]), .Z(n12243) );
  XNOR U12220 ( .A(y[2395]), .B(x[2395]), .Z(n12242) );
  AND U12221 ( .A(n12244), .B(n12245), .Z(n12240) );
  XNOR U12222 ( .A(y[2396]), .B(x[2396]), .Z(n12245) );
  XNOR U12223 ( .A(y[2397]), .B(x[2397]), .Z(n12244) );
  AND U12224 ( .A(n12246), .B(n12247), .Z(n12238) );
  AND U12225 ( .A(n12248), .B(n12249), .Z(n12247) );
  XNOR U12226 ( .A(y[2398]), .B(x[2398]), .Z(n12249) );
  XNOR U12227 ( .A(y[2399]), .B(x[2399]), .Z(n12248) );
  AND U12228 ( .A(n12250), .B(n12251), .Z(n12246) );
  XNOR U12229 ( .A(y[2400]), .B(x[2400]), .Z(n12251) );
  XNOR U12230 ( .A(y[2401]), .B(x[2401]), .Z(n12250) );
  AND U12231 ( .A(n12252), .B(n12253), .Z(n12236) );
  AND U12232 ( .A(n12254), .B(n12255), .Z(n12253) );
  AND U12233 ( .A(n12256), .B(n12257), .Z(n12255) );
  XNOR U12234 ( .A(y[2402]), .B(x[2402]), .Z(n12257) );
  XNOR U12235 ( .A(y[2403]), .B(x[2403]), .Z(n12256) );
  AND U12236 ( .A(n12258), .B(n12259), .Z(n12254) );
  XNOR U12237 ( .A(y[2404]), .B(x[2404]), .Z(n12259) );
  XNOR U12238 ( .A(y[2405]), .B(x[2405]), .Z(n12258) );
  AND U12239 ( .A(n12260), .B(n12261), .Z(n12252) );
  XNOR U12240 ( .A(y[2408]), .B(x[2408]), .Z(n12261) );
  AND U12241 ( .A(n12262), .B(n12263), .Z(n12260) );
  XNOR U12242 ( .A(y[2406]), .B(x[2406]), .Z(n12263) );
  XNOR U12243 ( .A(y[2407]), .B(x[2407]), .Z(n12262) );
  AND U12244 ( .A(n12264), .B(n12265), .Z(n12204) );
  AND U12245 ( .A(n12266), .B(n12267), .Z(n12265) );
  AND U12246 ( .A(n12268), .B(n12269), .Z(n12267) );
  AND U12247 ( .A(n12270), .B(n12271), .Z(n12269) );
  AND U12248 ( .A(n12272), .B(n12273), .Z(n12271) );
  XNOR U12249 ( .A(y[2409]), .B(x[2409]), .Z(n12273) );
  XNOR U12250 ( .A(y[2410]), .B(x[2410]), .Z(n12272) );
  AND U12251 ( .A(n12274), .B(n12275), .Z(n12270) );
  XNOR U12252 ( .A(y[2411]), .B(x[2411]), .Z(n12275) );
  XNOR U12253 ( .A(y[2412]), .B(x[2412]), .Z(n12274) );
  AND U12254 ( .A(n12276), .B(n12277), .Z(n12268) );
  AND U12255 ( .A(n12278), .B(n12279), .Z(n12277) );
  XNOR U12256 ( .A(y[2413]), .B(x[2413]), .Z(n12279) );
  XNOR U12257 ( .A(y[2414]), .B(x[2414]), .Z(n12278) );
  AND U12258 ( .A(n12280), .B(n12281), .Z(n12276) );
  XNOR U12259 ( .A(y[2415]), .B(x[2415]), .Z(n12281) );
  XNOR U12260 ( .A(y[2416]), .B(x[2416]), .Z(n12280) );
  AND U12261 ( .A(n12282), .B(n12283), .Z(n12266) );
  AND U12262 ( .A(n12284), .B(n12285), .Z(n12283) );
  AND U12263 ( .A(n12286), .B(n12287), .Z(n12285) );
  XNOR U12264 ( .A(y[2417]), .B(x[2417]), .Z(n12287) );
  XNOR U12265 ( .A(y[2418]), .B(x[2418]), .Z(n12286) );
  AND U12266 ( .A(n12288), .B(n12289), .Z(n12284) );
  XNOR U12267 ( .A(y[2419]), .B(x[2419]), .Z(n12289) );
  XNOR U12268 ( .A(y[2420]), .B(x[2420]), .Z(n12288) );
  AND U12269 ( .A(n12290), .B(n12291), .Z(n12282) );
  XNOR U12270 ( .A(y[2423]), .B(x[2423]), .Z(n12291) );
  AND U12271 ( .A(n12292), .B(n12293), .Z(n12290) );
  XNOR U12272 ( .A(y[2421]), .B(x[2421]), .Z(n12293) );
  XNOR U12273 ( .A(y[2422]), .B(x[2422]), .Z(n12292) );
  AND U12274 ( .A(n12294), .B(n12295), .Z(n12264) );
  AND U12275 ( .A(n12296), .B(n12297), .Z(n12295) );
  AND U12276 ( .A(n12298), .B(n12299), .Z(n12297) );
  AND U12277 ( .A(n12300), .B(n12301), .Z(n12299) );
  XNOR U12278 ( .A(y[2424]), .B(x[2424]), .Z(n12301) );
  XNOR U12279 ( .A(y[2425]), .B(x[2425]), .Z(n12300) );
  AND U12280 ( .A(n12302), .B(n12303), .Z(n12298) );
  XNOR U12281 ( .A(y[2426]), .B(x[2426]), .Z(n12303) );
  XNOR U12282 ( .A(y[2427]), .B(x[2427]), .Z(n12302) );
  AND U12283 ( .A(n12304), .B(n12305), .Z(n12296) );
  AND U12284 ( .A(n12306), .B(n12307), .Z(n12305) );
  XNOR U12285 ( .A(y[2428]), .B(x[2428]), .Z(n12307) );
  XNOR U12286 ( .A(y[2429]), .B(x[2429]), .Z(n12306) );
  AND U12287 ( .A(n12308), .B(n12309), .Z(n12304) );
  XNOR U12288 ( .A(y[2430]), .B(x[2430]), .Z(n12309) );
  XNOR U12289 ( .A(y[2431]), .B(x[2431]), .Z(n12308) );
  AND U12290 ( .A(n12310), .B(n12311), .Z(n12294) );
  AND U12291 ( .A(n12312), .B(n12313), .Z(n12311) );
  AND U12292 ( .A(n12314), .B(n12315), .Z(n12313) );
  XNOR U12293 ( .A(y[2038]), .B(x[2038]), .Z(n12315) );
  XNOR U12294 ( .A(y[2039]), .B(x[2039]), .Z(n12314) );
  AND U12295 ( .A(n12316), .B(n12317), .Z(n12312) );
  XNOR U12296 ( .A(y[1514]), .B(x[1514]), .Z(n12317) );
  XNOR U12297 ( .A(y[1515]), .B(x[1515]), .Z(n12316) );
  AND U12298 ( .A(n12318), .B(n12319), .Z(n12310) );
  XNOR U12299 ( .A(y[1518]), .B(x[1518]), .Z(n12319) );
  AND U12300 ( .A(n12320), .B(n12321), .Z(n12318) );
  XNOR U12301 ( .A(y[1516]), .B(x[1516]), .Z(n12321) );
  XNOR U12302 ( .A(y[1517]), .B(x[1517]), .Z(n12320) );
  AND U12303 ( .A(n12322), .B(n12323), .Z(n8652) );
  AND U12304 ( .A(n12324), .B(n12325), .Z(n12323) );
  AND U12305 ( .A(n12326), .B(n12327), .Z(n12325) );
  AND U12306 ( .A(n12328), .B(n12329), .Z(n12327) );
  AND U12307 ( .A(n12330), .B(n12331), .Z(n12329) );
  AND U12308 ( .A(n12332), .B(n12333), .Z(n12331) );
  AND U12309 ( .A(n12334), .B(n12335), .Z(n12333) );
  AND U12310 ( .A(n12336), .B(n12337), .Z(n12335) );
  XNOR U12311 ( .A(y[1519]), .B(x[1519]), .Z(n12337) );
  XNOR U12312 ( .A(y[1520]), .B(x[1520]), .Z(n12336) );
  AND U12313 ( .A(n12338), .B(n12339), .Z(n12334) );
  XNOR U12314 ( .A(y[1521]), .B(x[1521]), .Z(n12339) );
  XNOR U12315 ( .A(y[1522]), .B(x[1522]), .Z(n12338) );
  AND U12316 ( .A(n12340), .B(n12341), .Z(n12332) );
  AND U12317 ( .A(n12342), .B(n12343), .Z(n12341) );
  XNOR U12318 ( .A(y[1523]), .B(x[1523]), .Z(n12343) );
  XNOR U12319 ( .A(y[1524]), .B(x[1524]), .Z(n12342) );
  AND U12320 ( .A(n12344), .B(n12345), .Z(n12340) );
  XNOR U12321 ( .A(y[1525]), .B(x[1525]), .Z(n12345) );
  XNOR U12322 ( .A(y[1526]), .B(x[1526]), .Z(n12344) );
  AND U12323 ( .A(n12346), .B(n12347), .Z(n12330) );
  AND U12324 ( .A(n12348), .B(n12349), .Z(n12347) );
  AND U12325 ( .A(n12350), .B(n12351), .Z(n12349) );
  XNOR U12326 ( .A(y[1527]), .B(x[1527]), .Z(n12351) );
  XNOR U12327 ( .A(y[1528]), .B(x[1528]), .Z(n12350) );
  AND U12328 ( .A(n12352), .B(n12353), .Z(n12348) );
  XNOR U12329 ( .A(y[1529]), .B(x[1529]), .Z(n12353) );
  XNOR U12330 ( .A(y[2528]), .B(x[2528]), .Z(n12352) );
  AND U12331 ( .A(n12354), .B(n12355), .Z(n12346) );
  AND U12332 ( .A(n12356), .B(n12357), .Z(n12355) );
  XNOR U12333 ( .A(y[2529]), .B(x[2529]), .Z(n12357) );
  XNOR U12334 ( .A(y[2530]), .B(x[2530]), .Z(n12356) );
  AND U12335 ( .A(n12358), .B(n12359), .Z(n12354) );
  XNOR U12336 ( .A(y[2531]), .B(x[2531]), .Z(n12359) );
  XNOR U12337 ( .A(y[2532]), .B(x[2532]), .Z(n12358) );
  AND U12338 ( .A(n12360), .B(n12361), .Z(n12328) );
  AND U12339 ( .A(n12362), .B(n12363), .Z(n12361) );
  AND U12340 ( .A(n12364), .B(n12365), .Z(n12363) );
  AND U12341 ( .A(n12366), .B(n12367), .Z(n12365) );
  XNOR U12342 ( .A(y[2533]), .B(x[2533]), .Z(n12367) );
  XNOR U12343 ( .A(y[2534]), .B(x[2534]), .Z(n12366) );
  AND U12344 ( .A(n12368), .B(n12369), .Z(n12364) );
  XNOR U12345 ( .A(y[2535]), .B(x[2535]), .Z(n12369) );
  XNOR U12346 ( .A(y[2536]), .B(x[2536]), .Z(n12368) );
  AND U12347 ( .A(n12370), .B(n12371), .Z(n12362) );
  AND U12348 ( .A(n12372), .B(n12373), .Z(n12371) );
  XNOR U12349 ( .A(y[2537]), .B(x[2537]), .Z(n12373) );
  XNOR U12350 ( .A(y[2538]), .B(x[2538]), .Z(n12372) );
  AND U12351 ( .A(n12374), .B(n12375), .Z(n12370) );
  XNOR U12352 ( .A(y[2539]), .B(x[2539]), .Z(n12375) );
  XNOR U12353 ( .A(y[2540]), .B(x[2540]), .Z(n12374) );
  AND U12354 ( .A(n12376), .B(n12377), .Z(n12360) );
  AND U12355 ( .A(n12378), .B(n12379), .Z(n12377) );
  AND U12356 ( .A(n12380), .B(n12381), .Z(n12379) );
  XNOR U12357 ( .A(y[2541]), .B(x[2541]), .Z(n12381) );
  XNOR U12358 ( .A(y[2542]), .B(x[2542]), .Z(n12380) );
  AND U12359 ( .A(n12382), .B(n12383), .Z(n12378) );
  XNOR U12360 ( .A(y[2543]), .B(x[2543]), .Z(n12383) );
  XNOR U12361 ( .A(y[2544]), .B(x[2544]), .Z(n12382) );
  AND U12362 ( .A(n12384), .B(n12385), .Z(n12376) );
  XNOR U12363 ( .A(y[2547]), .B(x[2547]), .Z(n12385) );
  AND U12364 ( .A(n12386), .B(n12387), .Z(n12384) );
  XNOR U12365 ( .A(y[2545]), .B(x[2545]), .Z(n12387) );
  XNOR U12366 ( .A(y[2546]), .B(x[2546]), .Z(n12386) );
  AND U12367 ( .A(n12388), .B(n12389), .Z(n12326) );
  AND U12368 ( .A(n12390), .B(n12391), .Z(n12389) );
  AND U12369 ( .A(n12392), .B(n12393), .Z(n12391) );
  AND U12370 ( .A(n12394), .B(n12395), .Z(n12393) );
  AND U12371 ( .A(n12396), .B(n12397), .Z(n12395) );
  XNOR U12372 ( .A(y[2548]), .B(x[2548]), .Z(n12397) );
  XNOR U12373 ( .A(y[2549]), .B(x[2549]), .Z(n12396) );
  AND U12374 ( .A(n12398), .B(n12399), .Z(n12394) );
  XNOR U12375 ( .A(y[2550]), .B(x[2550]), .Z(n12399) );
  XNOR U12376 ( .A(y[2551]), .B(x[2551]), .Z(n12398) );
  AND U12377 ( .A(n12400), .B(n12401), .Z(n12392) );
  AND U12378 ( .A(n12402), .B(n12403), .Z(n12401) );
  XNOR U12379 ( .A(y[2552]), .B(x[2552]), .Z(n12403) );
  XNOR U12380 ( .A(y[2553]), .B(x[2553]), .Z(n12402) );
  AND U12381 ( .A(n12404), .B(n12405), .Z(n12400) );
  XNOR U12382 ( .A(y[2554]), .B(x[2554]), .Z(n12405) );
  XNOR U12383 ( .A(y[2555]), .B(x[2555]), .Z(n12404) );
  AND U12384 ( .A(n12406), .B(n12407), .Z(n12390) );
  AND U12385 ( .A(n12408), .B(n12409), .Z(n12407) );
  AND U12386 ( .A(n12410), .B(n12411), .Z(n12409) );
  XNOR U12387 ( .A(y[2556]), .B(x[2556]), .Z(n12411) );
  XNOR U12388 ( .A(y[2557]), .B(x[2557]), .Z(n12410) );
  AND U12389 ( .A(n12412), .B(n12413), .Z(n12408) );
  XNOR U12390 ( .A(y[2040]), .B(x[2040]), .Z(n12413) );
  XNOR U12391 ( .A(y[2041]), .B(x[2041]), .Z(n12412) );
  AND U12392 ( .A(n12414), .B(n12415), .Z(n12406) );
  XNOR U12393 ( .A(y[2044]), .B(x[2044]), .Z(n12415) );
  AND U12394 ( .A(n12416), .B(n12417), .Z(n12414) );
  XNOR U12395 ( .A(y[2042]), .B(x[2042]), .Z(n12417) );
  XNOR U12396 ( .A(y[2043]), .B(x[2043]), .Z(n12416) );
  AND U12397 ( .A(n12418), .B(n12419), .Z(n12388) );
  AND U12398 ( .A(n12420), .B(n12421), .Z(n12419) );
  AND U12399 ( .A(n12422), .B(n12423), .Z(n12421) );
  AND U12400 ( .A(n12424), .B(n12425), .Z(n12423) );
  XNOR U12401 ( .A(y[2045]), .B(x[2045]), .Z(n12425) );
  XNOR U12402 ( .A(y[2046]), .B(x[2046]), .Z(n12424) );
  AND U12403 ( .A(n12426), .B(n12427), .Z(n12422) );
  XNOR U12404 ( .A(y[2047]), .B(x[2047]), .Z(n12427) );
  XNOR U12405 ( .A(y[3010]), .B(x[3010]), .Z(n12426) );
  AND U12406 ( .A(n12428), .B(n12429), .Z(n12420) );
  AND U12407 ( .A(n12430), .B(n12431), .Z(n12429) );
  XNOR U12408 ( .A(y[3011]), .B(x[3011]), .Z(n12431) );
  XNOR U12409 ( .A(y[3012]), .B(x[3012]), .Z(n12430) );
  AND U12410 ( .A(n12432), .B(n12433), .Z(n12428) );
  XNOR U12411 ( .A(y[3013]), .B(x[3013]), .Z(n12433) );
  XNOR U12412 ( .A(y[3014]), .B(x[3014]), .Z(n12432) );
  AND U12413 ( .A(n12434), .B(n12435), .Z(n12418) );
  AND U12414 ( .A(n12436), .B(n12437), .Z(n12435) );
  AND U12415 ( .A(n12438), .B(n12439), .Z(n12437) );
  XNOR U12416 ( .A(y[3015]), .B(x[3015]), .Z(n12439) );
  XNOR U12417 ( .A(y[3016]), .B(x[3016]), .Z(n12438) );
  AND U12418 ( .A(n12440), .B(n12441), .Z(n12436) );
  XNOR U12419 ( .A(y[3017]), .B(x[3017]), .Z(n12441) );
  XNOR U12420 ( .A(y[3018]), .B(x[3018]), .Z(n12440) );
  AND U12421 ( .A(n12442), .B(n12443), .Z(n12434) );
  XNOR U12422 ( .A(y[3021]), .B(x[3021]), .Z(n12443) );
  AND U12423 ( .A(n12444), .B(n12445), .Z(n12442) );
  XNOR U12424 ( .A(y[3019]), .B(x[3019]), .Z(n12445) );
  XNOR U12425 ( .A(y[3020]), .B(x[3020]), .Z(n12444) );
  AND U12426 ( .A(n12446), .B(n12447), .Z(n12324) );
  AND U12427 ( .A(n12448), .B(n12449), .Z(n12447) );
  AND U12428 ( .A(n12450), .B(n12451), .Z(n12449) );
  AND U12429 ( .A(n12452), .B(n12453), .Z(n12451) );
  AND U12430 ( .A(n12454), .B(n12455), .Z(n12453) );
  AND U12431 ( .A(n12456), .B(n12457), .Z(n12455) );
  XNOR U12432 ( .A(y[3022]), .B(x[3022]), .Z(n12457) );
  XNOR U12433 ( .A(y[3023]), .B(x[3023]), .Z(n12456) );
  AND U12434 ( .A(n12458), .B(n12459), .Z(n12454) );
  XNOR U12435 ( .A(y[3024]), .B(x[3024]), .Z(n12459) );
  XNOR U12436 ( .A(y[3025]), .B(x[3025]), .Z(n12458) );
  AND U12437 ( .A(n12460), .B(n12461), .Z(n12452) );
  AND U12438 ( .A(n12462), .B(n12463), .Z(n12461) );
  XNOR U12439 ( .A(y[3026]), .B(x[3026]), .Z(n12463) );
  XNOR U12440 ( .A(y[3027]), .B(x[3027]), .Z(n12462) );
  AND U12441 ( .A(n12464), .B(n12465), .Z(n12460) );
  XNOR U12442 ( .A(y[3028]), .B(x[3028]), .Z(n12465) );
  XNOR U12443 ( .A(y[3029]), .B(x[3029]), .Z(n12464) );
  AND U12444 ( .A(n12466), .B(n12467), .Z(n12450) );
  AND U12445 ( .A(n12468), .B(n12469), .Z(n12467) );
  AND U12446 ( .A(n12470), .B(n12471), .Z(n12469) );
  XNOR U12447 ( .A(y[3030]), .B(x[3030]), .Z(n12471) );
  XNOR U12448 ( .A(y[3031]), .B(x[3031]), .Z(n12470) );
  AND U12449 ( .A(n12472), .B(n12473), .Z(n12468) );
  XNOR U12450 ( .A(y[3032]), .B(x[3032]), .Z(n12473) );
  XNOR U12451 ( .A(y[3033]), .B(x[3033]), .Z(n12472) );
  AND U12452 ( .A(n12474), .B(n12475), .Z(n12466) );
  AND U12453 ( .A(n12476), .B(n12477), .Z(n12475) );
  XNOR U12454 ( .A(y[3034]), .B(x[3034]), .Z(n12477) );
  XNOR U12455 ( .A(y[3035]), .B(x[3035]), .Z(n12476) );
  AND U12456 ( .A(n12478), .B(n12479), .Z(n12474) );
  XNOR U12457 ( .A(y[3036]), .B(x[3036]), .Z(n12479) );
  XNOR U12458 ( .A(y[3037]), .B(x[3037]), .Z(n12478) );
  AND U12459 ( .A(n12480), .B(n12481), .Z(n12448) );
  AND U12460 ( .A(n12482), .B(n12483), .Z(n12481) );
  AND U12461 ( .A(n12484), .B(n12485), .Z(n12483) );
  AND U12462 ( .A(n12486), .B(n12487), .Z(n12485) );
  XNOR U12463 ( .A(y[3038]), .B(x[3038]), .Z(n12487) );
  XNOR U12464 ( .A(y[3039]), .B(x[3039]), .Z(n12486) );
  AND U12465 ( .A(n12488), .B(n12489), .Z(n12484) );
  XNOR U12466 ( .A(y[3040]), .B(x[3040]), .Z(n12489) );
  XNOR U12467 ( .A(y[3041]), .B(x[3041]), .Z(n12488) );
  AND U12468 ( .A(n12490), .B(n12491), .Z(n12482) );
  AND U12469 ( .A(n12492), .B(n12493), .Z(n12491) );
  XNOR U12470 ( .A(y[3042]), .B(x[3042]), .Z(n12493) );
  XNOR U12471 ( .A(y[3043]), .B(x[3043]), .Z(n12492) );
  AND U12472 ( .A(n12494), .B(n12495), .Z(n12490) );
  XNOR U12473 ( .A(y[3044]), .B(x[3044]), .Z(n12495) );
  XNOR U12474 ( .A(y[3045]), .B(x[3045]), .Z(n12494) );
  AND U12475 ( .A(n12496), .B(n12497), .Z(n12480) );
  AND U12476 ( .A(n12498), .B(n12499), .Z(n12497) );
  AND U12477 ( .A(n12500), .B(n12501), .Z(n12499) );
  XNOR U12478 ( .A(y[3046]), .B(x[3046]), .Z(n12501) );
  XNOR U12479 ( .A(y[3047]), .B(x[3047]), .Z(n12500) );
  AND U12480 ( .A(n12502), .B(n12503), .Z(n12498) );
  XNOR U12481 ( .A(y[3048]), .B(x[3048]), .Z(n12503) );
  XNOR U12482 ( .A(y[3049]), .B(x[3049]), .Z(n12502) );
  AND U12483 ( .A(n12504), .B(n12505), .Z(n12496) );
  XNOR U12484 ( .A(y[3052]), .B(x[3052]), .Z(n12505) );
  AND U12485 ( .A(n12506), .B(n12507), .Z(n12504) );
  XNOR U12486 ( .A(y[3050]), .B(x[3050]), .Z(n12507) );
  XNOR U12487 ( .A(y[3051]), .B(x[3051]), .Z(n12506) );
  AND U12488 ( .A(n12508), .B(n12509), .Z(n12446) );
  AND U12489 ( .A(n12510), .B(n12511), .Z(n12509) );
  AND U12490 ( .A(n12512), .B(n12513), .Z(n12511) );
  AND U12491 ( .A(n12514), .B(n12515), .Z(n12513) );
  AND U12492 ( .A(n12516), .B(n12517), .Z(n12515) );
  XNOR U12493 ( .A(y[3053]), .B(x[3053]), .Z(n12517) );
  XNOR U12494 ( .A(y[3054]), .B(x[3054]), .Z(n12516) );
  AND U12495 ( .A(n12518), .B(n12519), .Z(n12514) );
  XNOR U12496 ( .A(y[3055]), .B(x[3055]), .Z(n12519) );
  XNOR U12497 ( .A(y[3056]), .B(x[3056]), .Z(n12518) );
  AND U12498 ( .A(n12520), .B(n12521), .Z(n12512) );
  AND U12499 ( .A(n12522), .B(n12523), .Z(n12521) );
  XNOR U12500 ( .A(y[3057]), .B(x[3057]), .Z(n12523) );
  XNOR U12501 ( .A(y[3058]), .B(x[3058]), .Z(n12522) );
  AND U12502 ( .A(n12524), .B(n12525), .Z(n12520) );
  XNOR U12503 ( .A(y[3059]), .B(x[3059]), .Z(n12525) );
  XNOR U12504 ( .A(y[3060]), .B(x[3060]), .Z(n12524) );
  AND U12505 ( .A(n12526), .B(n12527), .Z(n12510) );
  AND U12506 ( .A(n12528), .B(n12529), .Z(n12527) );
  AND U12507 ( .A(n12530), .B(n12531), .Z(n12529) );
  XNOR U12508 ( .A(y[3061]), .B(x[3061]), .Z(n12531) );
  XNOR U12509 ( .A(y[3062]), .B(x[3062]), .Z(n12530) );
  AND U12510 ( .A(n12532), .B(n12533), .Z(n12528) );
  XNOR U12511 ( .A(y[3063]), .B(x[3063]), .Z(n12533) );
  XNOR U12512 ( .A(y[3064]), .B(x[3064]), .Z(n12532) );
  AND U12513 ( .A(n12534), .B(n12535), .Z(n12526) );
  XNOR U12514 ( .A(y[3067]), .B(x[3067]), .Z(n12535) );
  AND U12515 ( .A(n12536), .B(n12537), .Z(n12534) );
  XNOR U12516 ( .A(y[3065]), .B(x[3065]), .Z(n12537) );
  XNOR U12517 ( .A(y[3066]), .B(x[3066]), .Z(n12536) );
  AND U12518 ( .A(n12538), .B(n12539), .Z(n12508) );
  AND U12519 ( .A(n12540), .B(n12541), .Z(n12539) );
  AND U12520 ( .A(n12542), .B(n12543), .Z(n12541) );
  AND U12521 ( .A(n12544), .B(n12545), .Z(n12543) );
  XNOR U12522 ( .A(y[3068]), .B(x[3068]), .Z(n12545) );
  XNOR U12523 ( .A(y[3069]), .B(x[3069]), .Z(n12544) );
  AND U12524 ( .A(n12546), .B(n12547), .Z(n12542) );
  XNOR U12525 ( .A(y[3070]), .B(x[3070]), .Z(n12547) );
  XNOR U12526 ( .A(y[3071]), .B(x[3071]), .Z(n12546) );
  AND U12527 ( .A(n12548), .B(n12549), .Z(n12540) );
  AND U12528 ( .A(n12550), .B(n12551), .Z(n12549) );
  XNOR U12529 ( .A(y[2558]), .B(x[2558]), .Z(n12551) );
  XNOR U12530 ( .A(y[2559]), .B(x[2559]), .Z(n12550) );
  AND U12531 ( .A(n12552), .B(n12553), .Z(n12548) );
  XNOR U12532 ( .A(y[2560]), .B(x[2560]), .Z(n12553) );
  XNOR U12533 ( .A(y[2561]), .B(x[2561]), .Z(n12552) );
  AND U12534 ( .A(n12554), .B(n12555), .Z(n12538) );
  AND U12535 ( .A(n12556), .B(n12557), .Z(n12555) );
  AND U12536 ( .A(n12558), .B(n12559), .Z(n12557) );
  XNOR U12537 ( .A(y[3458]), .B(x[3458]), .Z(n12559) );
  XNOR U12538 ( .A(y[3459]), .B(x[3459]), .Z(n12558) );
  AND U12539 ( .A(n12560), .B(n12561), .Z(n12556) );
  XNOR U12540 ( .A(y[3460]), .B(x[3460]), .Z(n12561) );
  XNOR U12541 ( .A(y[3461]), .B(x[3461]), .Z(n12560) );
  AND U12542 ( .A(n12562), .B(n12563), .Z(n12554) );
  XNOR U12543 ( .A(y[3464]), .B(x[3464]), .Z(n12563) );
  AND U12544 ( .A(n12564), .B(n12565), .Z(n12562) );
  XNOR U12545 ( .A(y[3462]), .B(x[3462]), .Z(n12565) );
  XNOR U12546 ( .A(y[3463]), .B(x[3463]), .Z(n12564) );
  AND U12547 ( .A(n12566), .B(n12567), .Z(n12322) );
  AND U12548 ( .A(n12568), .B(n12569), .Z(n12567) );
  AND U12549 ( .A(n12570), .B(n12571), .Z(n12569) );
  AND U12550 ( .A(n12572), .B(n12573), .Z(n12571) );
  AND U12551 ( .A(n12574), .B(n12575), .Z(n12573) );
  AND U12552 ( .A(n12576), .B(n12577), .Z(n12575) );
  AND U12553 ( .A(n12578), .B(n12579), .Z(n12577) );
  XNOR U12554 ( .A(y[3465]), .B(x[3465]), .Z(n12579) );
  XNOR U12555 ( .A(y[3466]), .B(x[3466]), .Z(n12578) );
  AND U12556 ( .A(n12580), .B(n12581), .Z(n12576) );
  XNOR U12557 ( .A(y[3467]), .B(x[3467]), .Z(n12581) );
  XNOR U12558 ( .A(y[3468]), .B(x[3468]), .Z(n12580) );
  AND U12559 ( .A(n12582), .B(n12583), .Z(n12574) );
  AND U12560 ( .A(n12584), .B(n12585), .Z(n12583) );
  XNOR U12561 ( .A(y[3469]), .B(x[3469]), .Z(n12585) );
  XNOR U12562 ( .A(y[3470]), .B(x[3470]), .Z(n12584) );
  AND U12563 ( .A(n12586), .B(n12587), .Z(n12582) );
  XNOR U12564 ( .A(y[3471]), .B(x[3471]), .Z(n12587) );
  XNOR U12565 ( .A(y[3472]), .B(x[3472]), .Z(n12586) );
  AND U12566 ( .A(n12588), .B(n12589), .Z(n12572) );
  AND U12567 ( .A(n12590), .B(n12591), .Z(n12589) );
  AND U12568 ( .A(n12592), .B(n12593), .Z(n12591) );
  XNOR U12569 ( .A(y[3473]), .B(x[3473]), .Z(n12593) );
  XNOR U12570 ( .A(y[3474]), .B(x[3474]), .Z(n12592) );
  AND U12571 ( .A(n12594), .B(n12595), .Z(n12590) );
  XNOR U12572 ( .A(y[3475]), .B(x[3475]), .Z(n12595) );
  XNOR U12573 ( .A(y[3476]), .B(x[3476]), .Z(n12594) );
  AND U12574 ( .A(n12596), .B(n12597), .Z(n12588) );
  AND U12575 ( .A(n12598), .B(n12599), .Z(n12597) );
  XNOR U12576 ( .A(y[3477]), .B(x[3477]), .Z(n12599) );
  XNOR U12577 ( .A(y[3478]), .B(x[3478]), .Z(n12598) );
  AND U12578 ( .A(n12600), .B(n12601), .Z(n12596) );
  XNOR U12579 ( .A(y[3479]), .B(x[3479]), .Z(n12601) );
  XNOR U12580 ( .A(y[3480]), .B(x[3480]), .Z(n12600) );
  AND U12581 ( .A(n12602), .B(n12603), .Z(n12570) );
  AND U12582 ( .A(n12604), .B(n12605), .Z(n12603) );
  AND U12583 ( .A(n12606), .B(n12607), .Z(n12605) );
  AND U12584 ( .A(n12608), .B(n12609), .Z(n12607) );
  XNOR U12585 ( .A(y[3481]), .B(x[3481]), .Z(n12609) );
  XNOR U12586 ( .A(y[3482]), .B(x[3482]), .Z(n12608) );
  AND U12587 ( .A(n12610), .B(n12611), .Z(n12606) );
  XNOR U12588 ( .A(y[3483]), .B(x[3483]), .Z(n12611) );
  XNOR U12589 ( .A(y[3484]), .B(x[3484]), .Z(n12610) );
  AND U12590 ( .A(n12612), .B(n12613), .Z(n12604) );
  AND U12591 ( .A(n12614), .B(n12615), .Z(n12613) );
  XNOR U12592 ( .A(y[3485]), .B(x[3485]), .Z(n12615) );
  XNOR U12593 ( .A(y[3486]), .B(x[3486]), .Z(n12614) );
  AND U12594 ( .A(n12616), .B(n12617), .Z(n12612) );
  XNOR U12595 ( .A(y[3487]), .B(x[3487]), .Z(n12617) );
  XNOR U12596 ( .A(y[3488]), .B(x[3488]), .Z(n12616) );
  AND U12597 ( .A(n12618), .B(n12619), .Z(n12602) );
  AND U12598 ( .A(n12620), .B(n12621), .Z(n12619) );
  AND U12599 ( .A(n12622), .B(n12623), .Z(n12621) );
  XNOR U12600 ( .A(y[3489]), .B(x[3489]), .Z(n12623) );
  XNOR U12601 ( .A(y[3490]), .B(x[3490]), .Z(n12622) );
  AND U12602 ( .A(n12624), .B(n12625), .Z(n12620) );
  XNOR U12603 ( .A(y[3491]), .B(x[3491]), .Z(n12625) );
  XNOR U12604 ( .A(y[3492]), .B(x[3492]), .Z(n12624) );
  AND U12605 ( .A(n12626), .B(n12627), .Z(n12618) );
  XNOR U12606 ( .A(y[3495]), .B(x[3495]), .Z(n12627) );
  AND U12607 ( .A(n12628), .B(n12629), .Z(n12626) );
  XNOR U12608 ( .A(y[3493]), .B(x[3493]), .Z(n12629) );
  XNOR U12609 ( .A(y[3494]), .B(x[3494]), .Z(n12628) );
  AND U12610 ( .A(n12630), .B(n12631), .Z(n12568) );
  AND U12611 ( .A(n12632), .B(n12633), .Z(n12631) );
  AND U12612 ( .A(n12634), .B(n12635), .Z(n12633) );
  AND U12613 ( .A(n12636), .B(n12637), .Z(n12635) );
  AND U12614 ( .A(n12638), .B(n12639), .Z(n12637) );
  XNOR U12615 ( .A(y[3496]), .B(x[3496]), .Z(n12639) );
  XNOR U12616 ( .A(y[3497]), .B(x[3497]), .Z(n12638) );
  AND U12617 ( .A(n12640), .B(n12641), .Z(n12636) );
  XNOR U12618 ( .A(y[3498]), .B(x[3498]), .Z(n12641) );
  XNOR U12619 ( .A(y[3499]), .B(x[3499]), .Z(n12640) );
  AND U12620 ( .A(n12642), .B(n12643), .Z(n12634) );
  AND U12621 ( .A(n12644), .B(n12645), .Z(n12643) );
  XNOR U12622 ( .A(y[3500]), .B(x[3500]), .Z(n12645) );
  XNOR U12623 ( .A(y[3501]), .B(x[3501]), .Z(n12644) );
  AND U12624 ( .A(n12646), .B(n12647), .Z(n12642) );
  XNOR U12625 ( .A(y[3502]), .B(x[3502]), .Z(n12647) );
  XNOR U12626 ( .A(y[3503]), .B(x[3503]), .Z(n12646) );
  AND U12627 ( .A(n12648), .B(n12649), .Z(n12632) );
  AND U12628 ( .A(n12650), .B(n12651), .Z(n12649) );
  AND U12629 ( .A(n12652), .B(n12653), .Z(n12651) );
  XNOR U12630 ( .A(y[3504]), .B(x[3504]), .Z(n12653) );
  XNOR U12631 ( .A(y[3505]), .B(x[3505]), .Z(n12652) );
  AND U12632 ( .A(n12654), .B(n12655), .Z(n12650) );
  XNOR U12633 ( .A(y[3506]), .B(x[3506]), .Z(n12655) );
  XNOR U12634 ( .A(y[3507]), .B(x[3507]), .Z(n12654) );
  AND U12635 ( .A(n12656), .B(n12657), .Z(n12648) );
  XNOR U12636 ( .A(y[3510]), .B(x[3510]), .Z(n12657) );
  AND U12637 ( .A(n12658), .B(n12659), .Z(n12656) );
  XNOR U12638 ( .A(y[3508]), .B(x[3508]), .Z(n12659) );
  XNOR U12639 ( .A(y[3509]), .B(x[3509]), .Z(n12658) );
  AND U12640 ( .A(n12660), .B(n12661), .Z(n12630) );
  AND U12641 ( .A(n12662), .B(n12663), .Z(n12661) );
  AND U12642 ( .A(n12664), .B(n12665), .Z(n12663) );
  AND U12643 ( .A(n12666), .B(n12667), .Z(n12665) );
  XNOR U12644 ( .A(y[3511]), .B(x[3511]), .Z(n12667) );
  XNOR U12645 ( .A(y[3512]), .B(x[3512]), .Z(n12666) );
  AND U12646 ( .A(n12668), .B(n12669), .Z(n12664) );
  XNOR U12647 ( .A(y[3513]), .B(x[3513]), .Z(n12669) );
  XNOR U12648 ( .A(y[3514]), .B(x[3514]), .Z(n12668) );
  AND U12649 ( .A(n12670), .B(n12671), .Z(n12662) );
  AND U12650 ( .A(n12672), .B(n12673), .Z(n12671) );
  XNOR U12651 ( .A(y[3515]), .B(x[3515]), .Z(n12673) );
  XNOR U12652 ( .A(y[3516]), .B(x[3516]), .Z(n12672) );
  AND U12653 ( .A(n12674), .B(n12675), .Z(n12670) );
  XNOR U12654 ( .A(y[3517]), .B(x[3517]), .Z(n12675) );
  XNOR U12655 ( .A(y[3518]), .B(x[3518]), .Z(n12674) );
  AND U12656 ( .A(n12676), .B(n12677), .Z(n12660) );
  AND U12657 ( .A(n12678), .B(n12679), .Z(n12677) );
  AND U12658 ( .A(n12680), .B(n12681), .Z(n12679) );
  XNOR U12659 ( .A(y[3519]), .B(x[3519]), .Z(n12681) );
  XNOR U12660 ( .A(y[3520]), .B(x[3520]), .Z(n12680) );
  AND U12661 ( .A(n12682), .B(n12683), .Z(n12678) );
  XNOR U12662 ( .A(y[3521]), .B(x[3521]), .Z(n12683) );
  XNOR U12663 ( .A(y[3522]), .B(x[3522]), .Z(n12682) );
  AND U12664 ( .A(n12684), .B(n12685), .Z(n12676) );
  XNOR U12665 ( .A(y[3525]), .B(x[3525]), .Z(n12685) );
  AND U12666 ( .A(n12686), .B(n12687), .Z(n12684) );
  XNOR U12667 ( .A(y[3523]), .B(x[3523]), .Z(n12687) );
  XNOR U12668 ( .A(y[3524]), .B(x[3524]), .Z(n12686) );
  AND U12669 ( .A(n12688), .B(n12689), .Z(n12566) );
  AND U12670 ( .A(n12690), .B(n12691), .Z(n12689) );
  AND U12671 ( .A(n12692), .B(n12693), .Z(n12691) );
  AND U12672 ( .A(n12694), .B(n12695), .Z(n12693) );
  AND U12673 ( .A(n12696), .B(n12697), .Z(n12695) );
  AND U12674 ( .A(n12698), .B(n12699), .Z(n12697) );
  XNOR U12675 ( .A(y[3526]), .B(x[3526]), .Z(n12699) );
  XNOR U12676 ( .A(y[3527]), .B(x[3527]), .Z(n12698) );
  AND U12677 ( .A(n12700), .B(n12701), .Z(n12696) );
  XNOR U12678 ( .A(y[3528]), .B(x[3528]), .Z(n12701) );
  XNOR U12679 ( .A(y[3529]), .B(x[3529]), .Z(n12700) );
  AND U12680 ( .A(n12702), .B(n12703), .Z(n12694) );
  AND U12681 ( .A(n12704), .B(n12705), .Z(n12703) );
  XNOR U12682 ( .A(y[3530]), .B(x[3530]), .Z(n12705) );
  XNOR U12683 ( .A(y[3531]), .B(x[3531]), .Z(n12704) );
  AND U12684 ( .A(n12706), .B(n12707), .Z(n12702) );
  XNOR U12685 ( .A(y[3532]), .B(x[3532]), .Z(n12707) );
  XNOR U12686 ( .A(y[3533]), .B(x[3533]), .Z(n12706) );
  AND U12687 ( .A(n12708), .B(n12709), .Z(n12692) );
  AND U12688 ( .A(n12710), .B(n12711), .Z(n12709) );
  AND U12689 ( .A(n12712), .B(n12713), .Z(n12711) );
  XNOR U12690 ( .A(y[3534]), .B(x[3534]), .Z(n12713) );
  XNOR U12691 ( .A(y[3535]), .B(x[3535]), .Z(n12712) );
  AND U12692 ( .A(n12714), .B(n12715), .Z(n12710) );
  XNOR U12693 ( .A(y[3536]), .B(x[3536]), .Z(n12715) );
  XNOR U12694 ( .A(y[3537]), .B(x[3537]), .Z(n12714) );
  AND U12695 ( .A(n12716), .B(n12717), .Z(n12708) );
  XNOR U12696 ( .A(y[3540]), .B(x[3540]), .Z(n12717) );
  AND U12697 ( .A(n12718), .B(n12719), .Z(n12716) );
  XNOR U12698 ( .A(y[3538]), .B(x[3538]), .Z(n12719) );
  XNOR U12699 ( .A(y[3539]), .B(x[3539]), .Z(n12718) );
  AND U12700 ( .A(n12720), .B(n12721), .Z(n12690) );
  AND U12701 ( .A(n12722), .B(n12723), .Z(n12721) );
  AND U12702 ( .A(n12724), .B(n12725), .Z(n12723) );
  AND U12703 ( .A(n12726), .B(n12727), .Z(n12725) );
  XNOR U12704 ( .A(y[3541]), .B(x[3541]), .Z(n12727) );
  XNOR U12705 ( .A(y[3542]), .B(x[3542]), .Z(n12726) );
  AND U12706 ( .A(n12728), .B(n12729), .Z(n12724) );
  XNOR U12707 ( .A(y[3543]), .B(x[3543]), .Z(n12729) );
  XNOR U12708 ( .A(y[3544]), .B(x[3544]), .Z(n12728) );
  AND U12709 ( .A(n12730), .B(n12731), .Z(n12722) );
  AND U12710 ( .A(n12732), .B(n12733), .Z(n12731) );
  XNOR U12711 ( .A(y[3545]), .B(x[3545]), .Z(n12733) );
  XNOR U12712 ( .A(y[3546]), .B(x[3546]), .Z(n12732) );
  AND U12713 ( .A(n12734), .B(n12735), .Z(n12730) );
  XNOR U12714 ( .A(y[3547]), .B(x[3547]), .Z(n12735) );
  XNOR U12715 ( .A(y[3548]), .B(x[3548]), .Z(n12734) );
  AND U12716 ( .A(n12736), .B(n12737), .Z(n12720) );
  AND U12717 ( .A(n12738), .B(n12739), .Z(n12737) );
  AND U12718 ( .A(n12740), .B(n12741), .Z(n12739) );
  XNOR U12719 ( .A(y[3549]), .B(x[3549]), .Z(n12741) );
  XNOR U12720 ( .A(y[3550]), .B(x[3550]), .Z(n12740) );
  AND U12721 ( .A(n12742), .B(n12743), .Z(n12738) );
  XNOR U12722 ( .A(y[3551]), .B(x[3551]), .Z(n12743) );
  XNOR U12723 ( .A(y[3552]), .B(x[3552]), .Z(n12742) );
  AND U12724 ( .A(n12744), .B(n12745), .Z(n12736) );
  XNOR U12725 ( .A(y[3555]), .B(x[3555]), .Z(n12745) );
  AND U12726 ( .A(n12746), .B(n12747), .Z(n12744) );
  XNOR U12727 ( .A(y[3553]), .B(x[3553]), .Z(n12747) );
  XNOR U12728 ( .A(y[3554]), .B(x[3554]), .Z(n12746) );
  AND U12729 ( .A(n12748), .B(n12749), .Z(n12688) );
  AND U12730 ( .A(n12750), .B(n12751), .Z(n12749) );
  AND U12731 ( .A(n12752), .B(n12753), .Z(n12751) );
  AND U12732 ( .A(n12754), .B(n12755), .Z(n12753) );
  AND U12733 ( .A(n12756), .B(n12757), .Z(n12755) );
  XNOR U12734 ( .A(y[3556]), .B(x[3556]), .Z(n12757) );
  XNOR U12735 ( .A(y[3557]), .B(x[3557]), .Z(n12756) );
  AND U12736 ( .A(n12758), .B(n12759), .Z(n12754) );
  XNOR U12737 ( .A(y[3558]), .B(x[3558]), .Z(n12759) );
  XNOR U12738 ( .A(y[3559]), .B(x[3559]), .Z(n12758) );
  AND U12739 ( .A(n12760), .B(n12761), .Z(n12752) );
  AND U12740 ( .A(n12762), .B(n12763), .Z(n12761) );
  XNOR U12741 ( .A(y[3560]), .B(x[3560]), .Z(n12763) );
  XNOR U12742 ( .A(y[3561]), .B(x[3561]), .Z(n12762) );
  AND U12743 ( .A(n12764), .B(n12765), .Z(n12760) );
  XNOR U12744 ( .A(y[3562]), .B(x[3562]), .Z(n12765) );
  XNOR U12745 ( .A(y[3563]), .B(x[3563]), .Z(n12764) );
  AND U12746 ( .A(n12766), .B(n12767), .Z(n12750) );
  AND U12747 ( .A(n12768), .B(n12769), .Z(n12767) );
  AND U12748 ( .A(n12770), .B(n12771), .Z(n12769) );
  XNOR U12749 ( .A(y[3564]), .B(x[3564]), .Z(n12771) );
  XNOR U12750 ( .A(y[3565]), .B(x[3565]), .Z(n12770) );
  AND U12751 ( .A(n12772), .B(n12773), .Z(n12768) );
  XNOR U12752 ( .A(y[3566]), .B(x[3566]), .Z(n12773) );
  XNOR U12753 ( .A(y[3567]), .B(x[3567]), .Z(n12772) );
  AND U12754 ( .A(n12774), .B(n12775), .Z(n12766) );
  XNOR U12755 ( .A(y[3570]), .B(x[3570]), .Z(n12775) );
  AND U12756 ( .A(n12776), .B(n12777), .Z(n12774) );
  XNOR U12757 ( .A(y[3568]), .B(x[3568]), .Z(n12777) );
  XNOR U12758 ( .A(y[3569]), .B(x[3569]), .Z(n12776) );
  AND U12759 ( .A(n12778), .B(n12779), .Z(n12748) );
  AND U12760 ( .A(n12780), .B(n12781), .Z(n12779) );
  AND U12761 ( .A(n12782), .B(n12783), .Z(n12781) );
  AND U12762 ( .A(n12784), .B(n12785), .Z(n12783) );
  XNOR U12763 ( .A(y[3571]), .B(x[3571]), .Z(n12785) );
  XNOR U12764 ( .A(y[3572]), .B(x[3572]), .Z(n12784) );
  AND U12765 ( .A(n12786), .B(n12787), .Z(n12782) );
  XNOR U12766 ( .A(y[3573]), .B(x[3573]), .Z(n12787) );
  XNOR U12767 ( .A(y[3574]), .B(x[3574]), .Z(n12786) );
  AND U12768 ( .A(n12788), .B(n12789), .Z(n12780) );
  AND U12769 ( .A(n12790), .B(n12791), .Z(n12789) );
  XNOR U12770 ( .A(y[3575]), .B(x[3575]), .Z(n12791) );
  XNOR U12771 ( .A(y[3576]), .B(x[3576]), .Z(n12790) );
  AND U12772 ( .A(n12792), .B(n12793), .Z(n12788) );
  XNOR U12773 ( .A(y[3577]), .B(x[3577]), .Z(n12793) );
  XNOR U12774 ( .A(y[3578]), .B(x[3578]), .Z(n12792) );
  AND U12775 ( .A(n12794), .B(n12795), .Z(n12778) );
  AND U12776 ( .A(n12796), .B(n12797), .Z(n12795) );
  AND U12777 ( .A(n12798), .B(n12799), .Z(n12797) );
  XNOR U12778 ( .A(y[3579]), .B(x[3579]), .Z(n12799) );
  XNOR U12779 ( .A(y[3580]), .B(x[3580]), .Z(n12798) );
  AND U12780 ( .A(n12800), .B(n12801), .Z(n12796) );
  XNOR U12781 ( .A(y[3581]), .B(x[3581]), .Z(n12801) );
  XNOR U12782 ( .A(y[3582]), .B(x[3582]), .Z(n12800) );
  AND U12783 ( .A(n12802), .B(n12803), .Z(n12794) );
  XNOR U12784 ( .A(y[3073]), .B(x[3073]), .Z(n12803) );
  AND U12785 ( .A(n12804), .B(n12805), .Z(n12802) );
  XNOR U12786 ( .A(y[3583]), .B(x[3583]), .Z(n12805) );
  XNOR U12787 ( .A(y[3072]), .B(x[3072]), .Z(n12804) );
  AND U12788 ( .A(n12806), .B(n12807), .Z(n8650) );
  AND U12789 ( .A(n12808), .B(n12809), .Z(n12807) );
  AND U12790 ( .A(n12810), .B(n12811), .Z(n12809) );
  AND U12791 ( .A(n12812), .B(n12813), .Z(n12811) );
  AND U12792 ( .A(n12814), .B(n12815), .Z(n12813) );
  AND U12793 ( .A(n12816), .B(n12817), .Z(n12815) );
  AND U12794 ( .A(n12818), .B(n12819), .Z(n12817) );
  AND U12795 ( .A(n12820), .B(n12821), .Z(n12819) );
  XNOR U12796 ( .A(y[1530]), .B(x[1530]), .Z(n12821) );
  XNOR U12797 ( .A(y[1531]), .B(x[1531]), .Z(n12820) );
  AND U12798 ( .A(n12822), .B(n12823), .Z(n12818) );
  XNOR U12799 ( .A(y[1532]), .B(x[1532]), .Z(n12823) );
  XNOR U12800 ( .A(y[1533]), .B(x[1533]), .Z(n12822) );
  AND U12801 ( .A(n12824), .B(n12825), .Z(n12816) );
  AND U12802 ( .A(n12826), .B(n12827), .Z(n12825) );
  XNOR U12803 ( .A(y[1534]), .B(x[1534]), .Z(n12827) );
  XNOR U12804 ( .A(y[1535]), .B(x[1535]), .Z(n12826) );
  AND U12805 ( .A(n12828), .B(n12829), .Z(n12824) );
  XNOR U12806 ( .A(y[1536]), .B(x[1536]), .Z(n12829) );
  XNOR U12807 ( .A(y[1537]), .B(x[1537]), .Z(n12828) );
  AND U12808 ( .A(n12830), .B(n12831), .Z(n12814) );
  AND U12809 ( .A(n12832), .B(n12833), .Z(n12831) );
  AND U12810 ( .A(n12834), .B(n12835), .Z(n12833) );
  XNOR U12811 ( .A(y[1538]), .B(x[1538]), .Z(n12835) );
  XNOR U12812 ( .A(y[1539]), .B(x[1539]), .Z(n12834) );
  AND U12813 ( .A(n12836), .B(n12837), .Z(n12832) );
  XNOR U12814 ( .A(y[1540]), .B(x[1540]), .Z(n12837) );
  XNOR U12815 ( .A(y[1541]), .B(x[1541]), .Z(n12836) );
  AND U12816 ( .A(n12838), .B(n12839), .Z(n12830) );
  AND U12817 ( .A(n12840), .B(n12841), .Z(n12839) );
  XNOR U12818 ( .A(y[1542]), .B(x[1542]), .Z(n12841) );
  XNOR U12819 ( .A(y[1543]), .B(x[1543]), .Z(n12840) );
  AND U12820 ( .A(n12842), .B(n12843), .Z(n12838) );
  XNOR U12821 ( .A(y[1544]), .B(x[1544]), .Z(n12843) );
  XNOR U12822 ( .A(y[1547]), .B(x[1547]), .Z(n12842) );
  AND U12823 ( .A(n12844), .B(n12845), .Z(n12812) );
  AND U12824 ( .A(n12846), .B(n12847), .Z(n12845) );
  AND U12825 ( .A(n12848), .B(n12849), .Z(n12847) );
  AND U12826 ( .A(n12850), .B(n12851), .Z(n12849) );
  XNOR U12827 ( .A(y[1545]), .B(x[1545]), .Z(n12851) );
  XNOR U12828 ( .A(y[1546]), .B(x[1546]), .Z(n12850) );
  AND U12829 ( .A(n12852), .B(n12853), .Z(n12848) );
  XNOR U12830 ( .A(y[1548]), .B(x[1548]), .Z(n12853) );
  XNOR U12831 ( .A(y[1549]), .B(x[1549]), .Z(n12852) );
  AND U12832 ( .A(n12854), .B(n12855), .Z(n12846) );
  AND U12833 ( .A(n12856), .B(n12857), .Z(n12855) );
  XNOR U12834 ( .A(y[1550]), .B(x[1550]), .Z(n12857) );
  XNOR U12835 ( .A(y[1551]), .B(x[1551]), .Z(n12856) );
  AND U12836 ( .A(n12858), .B(n12859), .Z(n12854) );
  XNOR U12837 ( .A(y[1552]), .B(x[1552]), .Z(n12859) );
  XNOR U12838 ( .A(y[1553]), .B(x[1553]), .Z(n12858) );
  AND U12839 ( .A(n12860), .B(n12861), .Z(n12844) );
  AND U12840 ( .A(n12862), .B(n12863), .Z(n12861) );
  AND U12841 ( .A(n12864), .B(n12865), .Z(n12863) );
  XNOR U12842 ( .A(y[1554]), .B(x[1554]), .Z(n12865) );
  XNOR U12843 ( .A(y[1555]), .B(x[1555]), .Z(n12864) );
  AND U12844 ( .A(n12866), .B(n12867), .Z(n12862) );
  XNOR U12845 ( .A(y[1556]), .B(x[1556]), .Z(n12867) );
  XNOR U12846 ( .A(y[1557]), .B(x[1557]), .Z(n12866) );
  AND U12847 ( .A(n12868), .B(n12869), .Z(n12860) );
  AND U12848 ( .A(n12870), .B(n12871), .Z(n12869) );
  XNOR U12849 ( .A(y[1558]), .B(x[1558]), .Z(n12871) );
  XNOR U12850 ( .A(y[1559]), .B(x[1559]), .Z(n12870) );
  AND U12851 ( .A(n12872), .B(n12873), .Z(n12868) );
  XNOR U12852 ( .A(y[1560]), .B(x[1560]), .Z(n12873) );
  XNOR U12853 ( .A(y[1561]), .B(x[1561]), .Z(n12872) );
  AND U12854 ( .A(n12874), .B(n12875), .Z(n12810) );
  AND U12855 ( .A(n12876), .B(n12877), .Z(n12875) );
  AND U12856 ( .A(n12878), .B(n12879), .Z(n12877) );
  AND U12857 ( .A(n12880), .B(n12881), .Z(n12879) );
  AND U12858 ( .A(n12882), .B(n12883), .Z(n12881) );
  XNOR U12859 ( .A(y[1562]), .B(x[1562]), .Z(n12883) );
  XNOR U12860 ( .A(y[1563]), .B(x[1563]), .Z(n12882) );
  AND U12861 ( .A(n12884), .B(n12885), .Z(n12880) );
  XNOR U12862 ( .A(y[1564]), .B(x[1564]), .Z(n12885) );
  XNOR U12863 ( .A(y[1565]), .B(x[1565]), .Z(n12884) );
  AND U12864 ( .A(n12886), .B(n12887), .Z(n12878) );
  AND U12865 ( .A(n12888), .B(n12889), .Z(n12887) );
  XNOR U12866 ( .A(y[1566]), .B(x[1566]), .Z(n12889) );
  XNOR U12867 ( .A(y[1567]), .B(x[1567]), .Z(n12888) );
  AND U12868 ( .A(n12890), .B(n12891), .Z(n12886) );
  XNOR U12869 ( .A(y[1568]), .B(x[1568]), .Z(n12891) );
  XNOR U12870 ( .A(y[1569]), .B(x[1569]), .Z(n12890) );
  AND U12871 ( .A(n12892), .B(n12893), .Z(n12876) );
  AND U12872 ( .A(n12894), .B(n12895), .Z(n12893) );
  AND U12873 ( .A(n12896), .B(n12897), .Z(n12895) );
  XNOR U12874 ( .A(y[1570]), .B(x[1570]), .Z(n12897) );
  XNOR U12875 ( .A(y[1571]), .B(x[1571]), .Z(n12896) );
  AND U12876 ( .A(n12898), .B(n12899), .Z(n12894) );
  XNOR U12877 ( .A(y[1572]), .B(x[1572]), .Z(n12899) );
  XNOR U12878 ( .A(y[1573]), .B(x[1573]), .Z(n12898) );
  AND U12879 ( .A(n12900), .B(n12901), .Z(n12892) );
  AND U12880 ( .A(n12902), .B(n12903), .Z(n12901) );
  XNOR U12881 ( .A(y[1574]), .B(x[1574]), .Z(n12903) );
  XNOR U12882 ( .A(y[1575]), .B(x[1575]), .Z(n12902) );
  AND U12883 ( .A(n12904), .B(n12905), .Z(n12900) );
  XNOR U12884 ( .A(y[1576]), .B(x[1576]), .Z(n12905) );
  XNOR U12885 ( .A(y[1577]), .B(x[1577]), .Z(n12904) );
  AND U12886 ( .A(n12906), .B(n12907), .Z(n12874) );
  AND U12887 ( .A(n12908), .B(n12909), .Z(n12907) );
  AND U12888 ( .A(n12910), .B(n12911), .Z(n12909) );
  AND U12889 ( .A(n12912), .B(n12913), .Z(n12911) );
  XNOR U12890 ( .A(y[1578]), .B(x[1578]), .Z(n12913) );
  XNOR U12891 ( .A(y[1579]), .B(x[1579]), .Z(n12912) );
  AND U12892 ( .A(n12914), .B(n12915), .Z(n12910) );
  XNOR U12893 ( .A(y[1580]), .B(x[1580]), .Z(n12915) );
  XNOR U12894 ( .A(y[1581]), .B(x[1581]), .Z(n12914) );
  AND U12895 ( .A(n12916), .B(n12917), .Z(n12908) );
  AND U12896 ( .A(n12918), .B(n12919), .Z(n12917) );
  XNOR U12897 ( .A(y[1582]), .B(x[1582]), .Z(n12919) );
  XNOR U12898 ( .A(y[1583]), .B(x[1583]), .Z(n12918) );
  AND U12899 ( .A(n12920), .B(n12921), .Z(n12916) );
  XNOR U12900 ( .A(y[1584]), .B(x[1584]), .Z(n12921) );
  XNOR U12901 ( .A(y[1585]), .B(x[1585]), .Z(n12920) );
  AND U12902 ( .A(n12922), .B(n12923), .Z(n12906) );
  AND U12903 ( .A(n12924), .B(n12925), .Z(n12923) );
  AND U12904 ( .A(n12926), .B(n12927), .Z(n12925) );
  XNOR U12905 ( .A(y[1586]), .B(x[1586]), .Z(n12927) );
  XNOR U12906 ( .A(y[1587]), .B(x[1587]), .Z(n12926) );
  AND U12907 ( .A(n12928), .B(n12929), .Z(n12924) );
  XNOR U12908 ( .A(y[1588]), .B(x[1588]), .Z(n12929) );
  XNOR U12909 ( .A(y[1589]), .B(x[1589]), .Z(n12928) );
  AND U12910 ( .A(n12930), .B(n12931), .Z(n12922) );
  AND U12911 ( .A(n12932), .B(n12933), .Z(n12931) );
  XNOR U12912 ( .A(y[1590]), .B(x[1590]), .Z(n12933) );
  XNOR U12913 ( .A(y[1591]), .B(x[1591]), .Z(n12932) );
  AND U12914 ( .A(n12934), .B(n12935), .Z(n12930) );
  XNOR U12915 ( .A(y[1592]), .B(x[1592]), .Z(n12935) );
  XNOR U12916 ( .A(y[1593]), .B(x[1593]), .Z(n12934) );
  AND U12917 ( .A(n12936), .B(n12937), .Z(n12808) );
  AND U12918 ( .A(n12938), .B(n12939), .Z(n12937) );
  AND U12919 ( .A(n12940), .B(n12941), .Z(n12939) );
  AND U12920 ( .A(n12942), .B(n12943), .Z(n12941) );
  AND U12921 ( .A(n12944), .B(n12945), .Z(n12943) );
  AND U12922 ( .A(n12946), .B(n12947), .Z(n12945) );
  XNOR U12923 ( .A(y[1594]), .B(x[1594]), .Z(n12947) );
  XNOR U12924 ( .A(y[1595]), .B(x[1595]), .Z(n12946) );
  AND U12925 ( .A(n12948), .B(n12949), .Z(n12944) );
  XNOR U12926 ( .A(y[1596]), .B(x[1596]), .Z(n12949) );
  XNOR U12927 ( .A(y[1597]), .B(x[1597]), .Z(n12948) );
  AND U12928 ( .A(n12950), .B(n12951), .Z(n12942) );
  AND U12929 ( .A(n12952), .B(n12953), .Z(n12951) );
  XNOR U12930 ( .A(y[1598]), .B(x[1598]), .Z(n12953) );
  XNOR U12931 ( .A(y[1599]), .B(x[1599]), .Z(n12952) );
  AND U12932 ( .A(n12954), .B(n12955), .Z(n12950) );
  XNOR U12933 ( .A(y[1600]), .B(x[1600]), .Z(n12955) );
  XNOR U12934 ( .A(y[1601]), .B(x[1601]), .Z(n12954) );
  AND U12935 ( .A(n12956), .B(n12957), .Z(n12940) );
  AND U12936 ( .A(n12958), .B(n12959), .Z(n12957) );
  AND U12937 ( .A(n12960), .B(n12961), .Z(n12959) );
  XNOR U12938 ( .A(y[1602]), .B(x[1602]), .Z(n12961) );
  XNOR U12939 ( .A(y[1603]), .B(x[1603]), .Z(n12960) );
  AND U12940 ( .A(n12962), .B(n12963), .Z(n12958) );
  XNOR U12941 ( .A(y[1604]), .B(x[1604]), .Z(n12963) );
  XNOR U12942 ( .A(y[1605]), .B(x[1605]), .Z(n12962) );
  AND U12943 ( .A(n12964), .B(n12965), .Z(n12956) );
  AND U12944 ( .A(n12966), .B(n12967), .Z(n12965) );
  XNOR U12945 ( .A(y[1606]), .B(x[1606]), .Z(n12967) );
  XNOR U12946 ( .A(y[1607]), .B(x[1607]), .Z(n12966) );
  AND U12947 ( .A(n12968), .B(n12969), .Z(n12964) );
  XNOR U12948 ( .A(y[1608]), .B(x[1608]), .Z(n12969) );
  XNOR U12949 ( .A(y[1609]), .B(x[1609]), .Z(n12968) );
  AND U12950 ( .A(n12970), .B(n12971), .Z(n12938) );
  AND U12951 ( .A(n12972), .B(n12973), .Z(n12971) );
  AND U12952 ( .A(n12974), .B(n12975), .Z(n12973) );
  AND U12953 ( .A(n12976), .B(n12977), .Z(n12975) );
  XNOR U12954 ( .A(y[1610]), .B(x[1610]), .Z(n12977) );
  XNOR U12955 ( .A(y[1611]), .B(x[1611]), .Z(n12976) );
  AND U12956 ( .A(n12978), .B(n12979), .Z(n12974) );
  XNOR U12957 ( .A(y[1612]), .B(x[1612]), .Z(n12979) );
  XNOR U12958 ( .A(y[1613]), .B(x[1613]), .Z(n12978) );
  AND U12959 ( .A(n12980), .B(n12981), .Z(n12972) );
  AND U12960 ( .A(n12982), .B(n12983), .Z(n12981) );
  XNOR U12961 ( .A(y[1614]), .B(x[1614]), .Z(n12983) );
  XNOR U12962 ( .A(y[1615]), .B(x[1615]), .Z(n12982) );
  AND U12963 ( .A(n12984), .B(n12985), .Z(n12980) );
  XNOR U12964 ( .A(y[1616]), .B(x[1616]), .Z(n12985) );
  XNOR U12965 ( .A(y[1617]), .B(x[1617]), .Z(n12984) );
  AND U12966 ( .A(n12986), .B(n12987), .Z(n12970) );
  AND U12967 ( .A(n12988), .B(n12989), .Z(n12987) );
  AND U12968 ( .A(n12990), .B(n12991), .Z(n12989) );
  XNOR U12969 ( .A(y[1618]), .B(x[1618]), .Z(n12991) );
  XNOR U12970 ( .A(y[1619]), .B(x[1619]), .Z(n12990) );
  AND U12971 ( .A(n12992), .B(n12993), .Z(n12988) );
  XNOR U12972 ( .A(y[1620]), .B(x[1620]), .Z(n12993) );
  XNOR U12973 ( .A(y[1621]), .B(x[1621]), .Z(n12992) );
  AND U12974 ( .A(n12994), .B(n12995), .Z(n12986) );
  AND U12975 ( .A(n12996), .B(n12997), .Z(n12995) );
  XNOR U12976 ( .A(y[1622]), .B(x[1622]), .Z(n12997) );
  XNOR U12977 ( .A(y[1623]), .B(x[1623]), .Z(n12996) );
  AND U12978 ( .A(n12998), .B(n12999), .Z(n12994) );
  XNOR U12979 ( .A(y[1624]), .B(x[1624]), .Z(n12999) );
  XNOR U12980 ( .A(y[1625]), .B(x[1625]), .Z(n12998) );
  AND U12981 ( .A(n13000), .B(n13001), .Z(n12936) );
  AND U12982 ( .A(n13002), .B(n13003), .Z(n13001) );
  AND U12983 ( .A(n13004), .B(n13005), .Z(n13003) );
  AND U12984 ( .A(n13006), .B(n13007), .Z(n13005) );
  AND U12985 ( .A(n13008), .B(n13009), .Z(n13007) );
  XNOR U12986 ( .A(y[1626]), .B(x[1626]), .Z(n13009) );
  XNOR U12987 ( .A(y[1627]), .B(x[1627]), .Z(n13008) );
  AND U12988 ( .A(n13010), .B(n13011), .Z(n13006) );
  XNOR U12989 ( .A(y[1628]), .B(x[1628]), .Z(n13011) );
  XNOR U12990 ( .A(y[1629]), .B(x[1629]), .Z(n13010) );
  AND U12991 ( .A(n13012), .B(n13013), .Z(n13004) );
  AND U12992 ( .A(n13014), .B(n13015), .Z(n13013) );
  XNOR U12993 ( .A(y[1630]), .B(x[1630]), .Z(n13015) );
  XNOR U12994 ( .A(y[1631]), .B(x[1631]), .Z(n13014) );
  AND U12995 ( .A(n13016), .B(n13017), .Z(n13012) );
  XNOR U12996 ( .A(y[1632]), .B(x[1632]), .Z(n13017) );
  XNOR U12997 ( .A(y[1633]), .B(x[1633]), .Z(n13016) );
  AND U12998 ( .A(n13018), .B(n13019), .Z(n13002) );
  AND U12999 ( .A(n13020), .B(n13021), .Z(n13019) );
  AND U13000 ( .A(n13022), .B(n13023), .Z(n13021) );
  XNOR U13001 ( .A(y[1634]), .B(x[1634]), .Z(n13023) );
  XNOR U13002 ( .A(y[1635]), .B(x[1635]), .Z(n13022) );
  AND U13003 ( .A(n13024), .B(n13025), .Z(n13020) );
  XNOR U13004 ( .A(y[1636]), .B(x[1636]), .Z(n13025) );
  XNOR U13005 ( .A(y[1637]), .B(x[1637]), .Z(n13024) );
  AND U13006 ( .A(n13026), .B(n13027), .Z(n13018) );
  AND U13007 ( .A(n13028), .B(n13029), .Z(n13027) );
  XNOR U13008 ( .A(y[1638]), .B(x[1638]), .Z(n13029) );
  XNOR U13009 ( .A(y[1639]), .B(x[1639]), .Z(n13028) );
  AND U13010 ( .A(n13030), .B(n13031), .Z(n13026) );
  XNOR U13011 ( .A(y[1640]), .B(x[1640]), .Z(n13031) );
  XNOR U13012 ( .A(y[1641]), .B(x[1641]), .Z(n13030) );
  AND U13013 ( .A(n13032), .B(n13033), .Z(n13000) );
  AND U13014 ( .A(n13034), .B(n13035), .Z(n13033) );
  AND U13015 ( .A(n13036), .B(n13037), .Z(n13035) );
  AND U13016 ( .A(n13038), .B(n13039), .Z(n13037) );
  XNOR U13017 ( .A(y[1642]), .B(x[1642]), .Z(n13039) );
  XNOR U13018 ( .A(y[1643]), .B(x[1643]), .Z(n13038) );
  AND U13019 ( .A(n13040), .B(n13041), .Z(n13036) );
  XNOR U13020 ( .A(y[1644]), .B(x[1644]), .Z(n13041) );
  XNOR U13021 ( .A(y[1645]), .B(x[1645]), .Z(n13040) );
  AND U13022 ( .A(n13042), .B(n13043), .Z(n13034) );
  AND U13023 ( .A(n13044), .B(n13045), .Z(n13043) );
  XNOR U13024 ( .A(y[1646]), .B(x[1646]), .Z(n13045) );
  XNOR U13025 ( .A(y[1647]), .B(x[1647]), .Z(n13044) );
  AND U13026 ( .A(n13046), .B(n13047), .Z(n13042) );
  XNOR U13027 ( .A(y[1648]), .B(x[1648]), .Z(n13047) );
  XNOR U13028 ( .A(y[1649]), .B(x[1649]), .Z(n13046) );
  AND U13029 ( .A(n13048), .B(n13049), .Z(n13032) );
  AND U13030 ( .A(n13050), .B(n13051), .Z(n13049) );
  AND U13031 ( .A(n13052), .B(n13053), .Z(n13051) );
  XNOR U13032 ( .A(y[1650]), .B(x[1650]), .Z(n13053) );
  XNOR U13033 ( .A(y[1651]), .B(x[1651]), .Z(n13052) );
  AND U13034 ( .A(n13054), .B(n13055), .Z(n13050) );
  XNOR U13035 ( .A(y[1652]), .B(x[1652]), .Z(n13055) );
  XNOR U13036 ( .A(y[1653]), .B(x[1653]), .Z(n13054) );
  AND U13037 ( .A(n13056), .B(n13057), .Z(n13048) );
  AND U13038 ( .A(n13058), .B(n13059), .Z(n13057) );
  XNOR U13039 ( .A(y[1654]), .B(x[1654]), .Z(n13059) );
  XNOR U13040 ( .A(y[1655]), .B(x[1655]), .Z(n13058) );
  AND U13041 ( .A(n13060), .B(n13061), .Z(n13056) );
  XNOR U13042 ( .A(y[1656]), .B(x[1656]), .Z(n13061) );
  XNOR U13043 ( .A(y[1657]), .B(x[1657]), .Z(n13060) );
  AND U13044 ( .A(n13062), .B(n13063), .Z(n12806) );
  AND U13045 ( .A(n13064), .B(n13065), .Z(n13063) );
  AND U13046 ( .A(n13066), .B(n13067), .Z(n13065) );
  AND U13047 ( .A(n13068), .B(n13069), .Z(n13067) );
  AND U13048 ( .A(n13070), .B(n13071), .Z(n13069) );
  AND U13049 ( .A(n13072), .B(n13073), .Z(n13071) );
  AND U13050 ( .A(n13074), .B(n13075), .Z(n13073) );
  XNOR U13051 ( .A(y[1658]), .B(x[1658]), .Z(n13075) );
  XNOR U13052 ( .A(y[1659]), .B(x[1659]), .Z(n13074) );
  AND U13053 ( .A(n13076), .B(n13077), .Z(n13072) );
  XNOR U13054 ( .A(y[1660]), .B(x[1660]), .Z(n13077) );
  XNOR U13055 ( .A(y[1661]), .B(x[1661]), .Z(n13076) );
  AND U13056 ( .A(n13078), .B(n13079), .Z(n13070) );
  AND U13057 ( .A(n13080), .B(n13081), .Z(n13079) );
  XNOR U13058 ( .A(y[1662]), .B(x[1662]), .Z(n13081) );
  XNOR U13059 ( .A(y[1663]), .B(x[1663]), .Z(n13080) );
  AND U13060 ( .A(n13082), .B(n13083), .Z(n13078) );
  XNOR U13061 ( .A(y[1664]), .B(x[1664]), .Z(n13083) );
  XNOR U13062 ( .A(y[1665]), .B(x[1665]), .Z(n13082) );
  AND U13063 ( .A(n13084), .B(n13085), .Z(n13068) );
  AND U13064 ( .A(n13086), .B(n13087), .Z(n13085) );
  AND U13065 ( .A(n13088), .B(n13089), .Z(n13087) );
  XNOR U13066 ( .A(y[1666]), .B(x[1666]), .Z(n13089) );
  XNOR U13067 ( .A(y[1667]), .B(x[1667]), .Z(n13088) );
  AND U13068 ( .A(n13090), .B(n13091), .Z(n13086) );
  XNOR U13069 ( .A(y[1668]), .B(x[1668]), .Z(n13091) );
  XNOR U13070 ( .A(y[1669]), .B(x[1669]), .Z(n13090) );
  AND U13071 ( .A(n13092), .B(n13093), .Z(n13084) );
  AND U13072 ( .A(n13094), .B(n13095), .Z(n13093) );
  XNOR U13073 ( .A(y[1670]), .B(x[1670]), .Z(n13095) );
  XNOR U13074 ( .A(y[1671]), .B(x[1671]), .Z(n13094) );
  AND U13075 ( .A(n13096), .B(n13097), .Z(n13092) );
  XNOR U13076 ( .A(y[1672]), .B(x[1672]), .Z(n13097) );
  XNOR U13077 ( .A(y[1673]), .B(x[1673]), .Z(n13096) );
  AND U13078 ( .A(n13098), .B(n13099), .Z(n13066) );
  AND U13079 ( .A(n13100), .B(n13101), .Z(n13099) );
  AND U13080 ( .A(n13102), .B(n13103), .Z(n13101) );
  AND U13081 ( .A(n13104), .B(n13105), .Z(n13103) );
  XNOR U13082 ( .A(y[1674]), .B(x[1674]), .Z(n13105) );
  XNOR U13083 ( .A(y[1675]), .B(x[1675]), .Z(n13104) );
  AND U13084 ( .A(n13106), .B(n13107), .Z(n13102) );
  XNOR U13085 ( .A(y[1676]), .B(x[1676]), .Z(n13107) );
  XNOR U13086 ( .A(y[1677]), .B(x[1677]), .Z(n13106) );
  AND U13087 ( .A(n13108), .B(n13109), .Z(n13100) );
  AND U13088 ( .A(n13110), .B(n13111), .Z(n13109) );
  XNOR U13089 ( .A(y[1678]), .B(x[1678]), .Z(n13111) );
  XNOR U13090 ( .A(y[1679]), .B(x[1679]), .Z(n13110) );
  AND U13091 ( .A(n13112), .B(n13113), .Z(n13108) );
  XNOR U13092 ( .A(y[1680]), .B(x[1680]), .Z(n13113) );
  XNOR U13093 ( .A(y[1681]), .B(x[1681]), .Z(n13112) );
  AND U13094 ( .A(n13114), .B(n13115), .Z(n13098) );
  AND U13095 ( .A(n13116), .B(n13117), .Z(n13115) );
  AND U13096 ( .A(n13118), .B(n13119), .Z(n13117) );
  XNOR U13097 ( .A(y[1682]), .B(x[1682]), .Z(n13119) );
  XNOR U13098 ( .A(y[1683]), .B(x[1683]), .Z(n13118) );
  AND U13099 ( .A(n13120), .B(n13121), .Z(n13116) );
  XNOR U13100 ( .A(y[1684]), .B(x[1684]), .Z(n13121) );
  XNOR U13101 ( .A(y[1685]), .B(x[1685]), .Z(n13120) );
  AND U13102 ( .A(n13122), .B(n13123), .Z(n13114) );
  AND U13103 ( .A(n13124), .B(n13125), .Z(n13123) );
  XNOR U13104 ( .A(y[1686]), .B(x[1686]), .Z(n13125) );
  XNOR U13105 ( .A(y[1687]), .B(x[1687]), .Z(n13124) );
  AND U13106 ( .A(n13126), .B(n13127), .Z(n13122) );
  XNOR U13107 ( .A(y[1688]), .B(x[1688]), .Z(n13127) );
  XNOR U13108 ( .A(y[1689]), .B(x[1689]), .Z(n13126) );
  AND U13109 ( .A(n13128), .B(n13129), .Z(n13064) );
  AND U13110 ( .A(n13130), .B(n13131), .Z(n13129) );
  AND U13111 ( .A(n13132), .B(n13133), .Z(n13131) );
  AND U13112 ( .A(n13134), .B(n13135), .Z(n13133) );
  AND U13113 ( .A(n13136), .B(n13137), .Z(n13135) );
  XNOR U13114 ( .A(y[1690]), .B(x[1690]), .Z(n13137) );
  XNOR U13115 ( .A(y[1691]), .B(x[1691]), .Z(n13136) );
  AND U13116 ( .A(n13138), .B(n13139), .Z(n13134) );
  XNOR U13117 ( .A(y[1692]), .B(x[1692]), .Z(n13139) );
  XNOR U13118 ( .A(y[1693]), .B(x[1693]), .Z(n13138) );
  AND U13119 ( .A(n13140), .B(n13141), .Z(n13132) );
  AND U13120 ( .A(n13142), .B(n13143), .Z(n13141) );
  XNOR U13121 ( .A(y[1694]), .B(x[1694]), .Z(n13143) );
  XNOR U13122 ( .A(y[1695]), .B(x[1695]), .Z(n13142) );
  AND U13123 ( .A(n13144), .B(n13145), .Z(n13140) );
  XNOR U13124 ( .A(y[1696]), .B(x[1696]), .Z(n13145) );
  XNOR U13125 ( .A(y[1697]), .B(x[1697]), .Z(n13144) );
  AND U13126 ( .A(n13146), .B(n13147), .Z(n13130) );
  AND U13127 ( .A(n13148), .B(n13149), .Z(n13147) );
  AND U13128 ( .A(n13150), .B(n13151), .Z(n13149) );
  XNOR U13129 ( .A(y[1698]), .B(x[1698]), .Z(n13151) );
  XNOR U13130 ( .A(y[1699]), .B(x[1699]), .Z(n13150) );
  AND U13131 ( .A(n13152), .B(n13153), .Z(n13148) );
  XNOR U13132 ( .A(y[1700]), .B(x[1700]), .Z(n13153) );
  XNOR U13133 ( .A(y[1701]), .B(x[1701]), .Z(n13152) );
  AND U13134 ( .A(n13154), .B(n13155), .Z(n13146) );
  AND U13135 ( .A(n13156), .B(n13157), .Z(n13155) );
  XNOR U13136 ( .A(y[1702]), .B(x[1702]), .Z(n13157) );
  XNOR U13137 ( .A(y[1703]), .B(x[1703]), .Z(n13156) );
  AND U13138 ( .A(n13158), .B(n13159), .Z(n13154) );
  XNOR U13139 ( .A(y[1704]), .B(x[1704]), .Z(n13159) );
  XNOR U13140 ( .A(y[1705]), .B(x[1705]), .Z(n13158) );
  AND U13141 ( .A(n13160), .B(n13161), .Z(n13128) );
  AND U13142 ( .A(n13162), .B(n13163), .Z(n13161) );
  AND U13143 ( .A(n13164), .B(n13165), .Z(n13163) );
  AND U13144 ( .A(n13166), .B(n13167), .Z(n13165) );
  XNOR U13145 ( .A(y[1706]), .B(x[1706]), .Z(n13167) );
  XNOR U13146 ( .A(y[1707]), .B(x[1707]), .Z(n13166) );
  AND U13147 ( .A(n13168), .B(n13169), .Z(n13164) );
  XNOR U13148 ( .A(y[1708]), .B(x[1708]), .Z(n13169) );
  XNOR U13149 ( .A(y[1709]), .B(x[1709]), .Z(n13168) );
  AND U13150 ( .A(n13170), .B(n13171), .Z(n13162) );
  AND U13151 ( .A(n13172), .B(n13173), .Z(n13171) );
  XNOR U13152 ( .A(y[1710]), .B(x[1710]), .Z(n13173) );
  XNOR U13153 ( .A(y[1711]), .B(x[1711]), .Z(n13172) );
  AND U13154 ( .A(n13174), .B(n13175), .Z(n13170) );
  XNOR U13155 ( .A(y[1712]), .B(x[1712]), .Z(n13175) );
  XNOR U13156 ( .A(y[1713]), .B(x[1713]), .Z(n13174) );
  AND U13157 ( .A(n13176), .B(n13177), .Z(n13160) );
  AND U13158 ( .A(n13178), .B(n13179), .Z(n13177) );
  AND U13159 ( .A(n13180), .B(n13181), .Z(n13179) );
  XNOR U13160 ( .A(y[1714]), .B(x[1714]), .Z(n13181) );
  XNOR U13161 ( .A(y[1715]), .B(x[1715]), .Z(n13180) );
  AND U13162 ( .A(n13182), .B(n13183), .Z(n13178) );
  XNOR U13163 ( .A(y[1716]), .B(x[1716]), .Z(n13183) );
  XNOR U13164 ( .A(y[1717]), .B(x[1717]), .Z(n13182) );
  AND U13165 ( .A(n13184), .B(n13185), .Z(n13176) );
  AND U13166 ( .A(n13186), .B(n13187), .Z(n13185) );
  XNOR U13167 ( .A(y[1718]), .B(x[1718]), .Z(n13187) );
  XNOR U13168 ( .A(y[1719]), .B(x[1719]), .Z(n13186) );
  AND U13169 ( .A(n13188), .B(n13189), .Z(n13184) );
  XNOR U13170 ( .A(y[1720]), .B(x[1720]), .Z(n13189) );
  XNOR U13171 ( .A(y[1721]), .B(x[1721]), .Z(n13188) );
  AND U13172 ( .A(n13190), .B(n13191), .Z(n13062) );
  AND U13173 ( .A(n13192), .B(n13193), .Z(n13191) );
  AND U13174 ( .A(n13194), .B(n13195), .Z(n13193) );
  AND U13175 ( .A(n13196), .B(n13197), .Z(n13195) );
  AND U13176 ( .A(n13198), .B(n13199), .Z(n13197) );
  AND U13177 ( .A(n13200), .B(n13201), .Z(n13199) );
  XNOR U13178 ( .A(y[1722]), .B(x[1722]), .Z(n13201) );
  XNOR U13179 ( .A(y[1723]), .B(x[1723]), .Z(n13200) );
  AND U13180 ( .A(n13202), .B(n13203), .Z(n13198) );
  XNOR U13181 ( .A(y[1724]), .B(x[1724]), .Z(n13203) );
  XNOR U13182 ( .A(y[1725]), .B(x[1725]), .Z(n13202) );
  AND U13183 ( .A(n13204), .B(n13205), .Z(n13196) );
  AND U13184 ( .A(n13206), .B(n13207), .Z(n13205) );
  XNOR U13185 ( .A(y[1726]), .B(x[1726]), .Z(n13207) );
  XNOR U13186 ( .A(y[1727]), .B(x[1727]), .Z(n13206) );
  AND U13187 ( .A(n13208), .B(n13209), .Z(n13204) );
  XNOR U13188 ( .A(y[1728]), .B(x[1728]), .Z(n13209) );
  XNOR U13189 ( .A(y[1729]), .B(x[1729]), .Z(n13208) );
  AND U13190 ( .A(n13210), .B(n13211), .Z(n13194) );
  AND U13191 ( .A(n13212), .B(n13213), .Z(n13211) );
  AND U13192 ( .A(n13214), .B(n13215), .Z(n13213) );
  XNOR U13193 ( .A(y[1730]), .B(x[1730]), .Z(n13215) );
  XNOR U13194 ( .A(y[1731]), .B(x[1731]), .Z(n13214) );
  AND U13195 ( .A(n13216), .B(n13217), .Z(n13212) );
  XNOR U13196 ( .A(y[1732]), .B(x[1732]), .Z(n13217) );
  XNOR U13197 ( .A(y[1733]), .B(x[1733]), .Z(n13216) );
  AND U13198 ( .A(n13218), .B(n13219), .Z(n13210) );
  AND U13199 ( .A(n13220), .B(n13221), .Z(n13219) );
  XNOR U13200 ( .A(y[1734]), .B(x[1734]), .Z(n13221) );
  XNOR U13201 ( .A(y[1735]), .B(x[1735]), .Z(n13220) );
  AND U13202 ( .A(n13222), .B(n13223), .Z(n13218) );
  XNOR U13203 ( .A(y[1736]), .B(x[1736]), .Z(n13223) );
  XNOR U13204 ( .A(y[1737]), .B(x[1737]), .Z(n13222) );
  AND U13205 ( .A(n13224), .B(n13225), .Z(n13192) );
  AND U13206 ( .A(n13226), .B(n13227), .Z(n13225) );
  AND U13207 ( .A(n13228), .B(n13229), .Z(n13227) );
  AND U13208 ( .A(n13230), .B(n13231), .Z(n13229) );
  XNOR U13209 ( .A(y[1738]), .B(x[1738]), .Z(n13231) );
  XNOR U13210 ( .A(y[1739]), .B(x[1739]), .Z(n13230) );
  AND U13211 ( .A(n13232), .B(n13233), .Z(n13228) );
  XNOR U13212 ( .A(y[1740]), .B(x[1740]), .Z(n13233) );
  XNOR U13213 ( .A(y[1741]), .B(x[1741]), .Z(n13232) );
  AND U13214 ( .A(n13234), .B(n13235), .Z(n13226) );
  AND U13215 ( .A(n13236), .B(n13237), .Z(n13235) );
  XNOR U13216 ( .A(y[1742]), .B(x[1742]), .Z(n13237) );
  XNOR U13217 ( .A(y[1743]), .B(x[1743]), .Z(n13236) );
  AND U13218 ( .A(n13238), .B(n13239), .Z(n13234) );
  XNOR U13219 ( .A(y[1744]), .B(x[1744]), .Z(n13239) );
  XNOR U13220 ( .A(y[1745]), .B(x[1745]), .Z(n13238) );
  AND U13221 ( .A(n13240), .B(n13241), .Z(n13224) );
  AND U13222 ( .A(n13242), .B(n13243), .Z(n13241) );
  AND U13223 ( .A(n13244), .B(n13245), .Z(n13243) );
  XNOR U13224 ( .A(y[1746]), .B(x[1746]), .Z(n13245) );
  XNOR U13225 ( .A(y[1747]), .B(x[1747]), .Z(n13244) );
  AND U13226 ( .A(n13246), .B(n13247), .Z(n13242) );
  XNOR U13227 ( .A(y[1748]), .B(x[1748]), .Z(n13247) );
  XNOR U13228 ( .A(y[1749]), .B(x[1749]), .Z(n13246) );
  AND U13229 ( .A(n13248), .B(n13249), .Z(n13240) );
  AND U13230 ( .A(n13250), .B(n13251), .Z(n13249) );
  XNOR U13231 ( .A(y[1750]), .B(x[1750]), .Z(n13251) );
  XNOR U13232 ( .A(y[1751]), .B(x[1751]), .Z(n13250) );
  AND U13233 ( .A(n13252), .B(n13253), .Z(n13248) );
  XNOR U13234 ( .A(y[1752]), .B(x[1752]), .Z(n13253) );
  XNOR U13235 ( .A(y[1753]), .B(x[1753]), .Z(n13252) );
  AND U13236 ( .A(n13254), .B(n13255), .Z(n13190) );
  AND U13237 ( .A(n13256), .B(n13257), .Z(n13255) );
  AND U13238 ( .A(n13258), .B(n13259), .Z(n13257) );
  AND U13239 ( .A(n13260), .B(n13261), .Z(n13259) );
  AND U13240 ( .A(n13262), .B(n13263), .Z(n13261) );
  XNOR U13241 ( .A(y[1754]), .B(x[1754]), .Z(n13263) );
  XNOR U13242 ( .A(y[1755]), .B(x[1755]), .Z(n13262) );
  AND U13243 ( .A(n13264), .B(n13265), .Z(n13260) );
  XNOR U13244 ( .A(y[1756]), .B(x[1756]), .Z(n13265) );
  XNOR U13245 ( .A(y[1757]), .B(x[1757]), .Z(n13264) );
  AND U13246 ( .A(n13266), .B(n13267), .Z(n13258) );
  AND U13247 ( .A(n13268), .B(n13269), .Z(n13267) );
  XNOR U13248 ( .A(y[1758]), .B(x[1758]), .Z(n13269) );
  XNOR U13249 ( .A(y[1759]), .B(x[1759]), .Z(n13268) );
  AND U13250 ( .A(n13270), .B(n13271), .Z(n13266) );
  XNOR U13251 ( .A(y[1760]), .B(x[1760]), .Z(n13271) );
  XNOR U13252 ( .A(y[1761]), .B(x[1761]), .Z(n13270) );
  AND U13253 ( .A(n13272), .B(n13273), .Z(n13256) );
  AND U13254 ( .A(n13274), .B(n13275), .Z(n13273) );
  AND U13255 ( .A(n13276), .B(n13277), .Z(n13275) );
  XNOR U13256 ( .A(y[1762]), .B(x[1762]), .Z(n13277) );
  XNOR U13257 ( .A(y[1763]), .B(x[1763]), .Z(n13276) );
  AND U13258 ( .A(n13278), .B(n13279), .Z(n13274) );
  XNOR U13259 ( .A(y[1764]), .B(x[1764]), .Z(n13279) );
  XNOR U13260 ( .A(y[1765]), .B(x[1765]), .Z(n13278) );
  AND U13261 ( .A(n13280), .B(n13281), .Z(n13272) );
  AND U13262 ( .A(n13282), .B(n13283), .Z(n13281) );
  XNOR U13263 ( .A(y[1766]), .B(x[1766]), .Z(n13283) );
  XNOR U13264 ( .A(y[1767]), .B(x[1767]), .Z(n13282) );
  AND U13265 ( .A(n13284), .B(n13285), .Z(n13280) );
  XNOR U13266 ( .A(y[1768]), .B(x[1768]), .Z(n13285) );
  XNOR U13267 ( .A(y[1769]), .B(x[1769]), .Z(n13284) );
  AND U13268 ( .A(n13286), .B(n13287), .Z(n13254) );
  AND U13269 ( .A(n13288), .B(n13289), .Z(n13287) );
  AND U13270 ( .A(n13290), .B(n13291), .Z(n13289) );
  AND U13271 ( .A(n13292), .B(n13293), .Z(n13291) );
  XNOR U13272 ( .A(y[1770]), .B(x[1770]), .Z(n13293) );
  XNOR U13273 ( .A(y[1771]), .B(x[1771]), .Z(n13292) );
  AND U13274 ( .A(n13294), .B(n13295), .Z(n13290) );
  XNOR U13275 ( .A(y[1772]), .B(x[1772]), .Z(n13295) );
  XNOR U13276 ( .A(y[1773]), .B(x[1773]), .Z(n13294) );
  AND U13277 ( .A(n13296), .B(n13297), .Z(n13288) );
  AND U13278 ( .A(n13298), .B(n13299), .Z(n13297) );
  XNOR U13279 ( .A(y[1774]), .B(x[1774]), .Z(n13299) );
  XNOR U13280 ( .A(y[1775]), .B(x[1775]), .Z(n13298) );
  AND U13281 ( .A(n13300), .B(n13301), .Z(n13296) );
  XNOR U13282 ( .A(y[1776]), .B(x[1776]), .Z(n13301) );
  XNOR U13283 ( .A(y[1777]), .B(x[1777]), .Z(n13300) );
  AND U13284 ( .A(n13302), .B(n13303), .Z(n13286) );
  AND U13285 ( .A(n13304), .B(n13305), .Z(n13303) );
  AND U13286 ( .A(n13306), .B(n13307), .Z(n13305) );
  XNOR U13287 ( .A(y[1778]), .B(x[1778]), .Z(n13307) );
  XNOR U13288 ( .A(y[1779]), .B(x[1779]), .Z(n13306) );
  AND U13289 ( .A(n13308), .B(n13309), .Z(n13304) );
  XNOR U13290 ( .A(y[1780]), .B(x[1780]), .Z(n13309) );
  XNOR U13291 ( .A(y[1781]), .B(x[1781]), .Z(n13308) );
  AND U13292 ( .A(n13310), .B(n13311), .Z(n13302) );
  AND U13293 ( .A(n13312), .B(n13313), .Z(n13311) );
  XNOR U13294 ( .A(y[1782]), .B(x[1782]), .Z(n13313) );
  XNOR U13295 ( .A(y[1783]), .B(x[1783]), .Z(n13312) );
  AND U13296 ( .A(n13314), .B(n13315), .Z(n13310) );
  XNOR U13297 ( .A(y[1784]), .B(x[1784]), .Z(n13315) );
  XNOR U13298 ( .A(y[1785]), .B(x[1785]), .Z(n13314) );
  AND U13299 ( .A(n13316), .B(n13317), .Z(n8646) );
  XNOR U13300 ( .A(y[1501]), .B(x[1501]), .Z(n13317) );
  XNOR U13301 ( .A(y[1502]), .B(x[1502]), .Z(n13316) );
  AND U13302 ( .A(n13318), .B(n13319), .Z(n8644) );
  AND U13303 ( .A(n13320), .B(n13321), .Z(n13319) );
  XNOR U13304 ( .A(y[1505]), .B(x[1505]), .Z(n13321) );
  AND U13305 ( .A(n13322), .B(n13323), .Z(n13320) );
  XNOR U13306 ( .A(y[1503]), .B(x[1503]), .Z(n13323) );
  XNOR U13307 ( .A(y[1504]), .B(x[1504]), .Z(n13322) );
  AND U13308 ( .A(n13324), .B(n13325), .Z(n13318) );
  XNOR U13309 ( .A(y[1506]), .B(x[1506]), .Z(n13325) );
  XNOR U13310 ( .A(y[1507]), .B(x[1507]), .Z(n13324) );
  AND U13311 ( .A(n13326), .B(n13327), .Z(n8642) );
  AND U13312 ( .A(n13328), .B(n13329), .Z(n13327) );
  AND U13313 ( .A(n13330), .B(n13331), .Z(n13329) );
  XNOR U13314 ( .A(y[974]), .B(x[974]), .Z(n13331) );
  AND U13315 ( .A(n13332), .B(n13333), .Z(n13330) );
  XNOR U13316 ( .A(y[972]), .B(x[972]), .Z(n13333) );
  XNOR U13317 ( .A(y[973]), .B(x[973]), .Z(n13332) );
  AND U13318 ( .A(n13334), .B(n13335), .Z(n13328) );
  XNOR U13319 ( .A(y[975]), .B(x[975]), .Z(n13335) );
  XNOR U13320 ( .A(y[976]), .B(x[976]), .Z(n13334) );
  AND U13321 ( .A(n13336), .B(n13337), .Z(n13326) );
  AND U13322 ( .A(n13338), .B(n13339), .Z(n13337) );
  XNOR U13323 ( .A(y[977]), .B(x[977]), .Z(n13339) );
  XNOR U13324 ( .A(y[978]), .B(x[978]), .Z(n13338) );
  AND U13325 ( .A(n13340), .B(n13341), .Z(n13336) );
  XNOR U13326 ( .A(y[979]), .B(x[979]), .Z(n13341) );
  XNOR U13327 ( .A(y[980]), .B(x[980]), .Z(n13340) );
  AND U13328 ( .A(n13342), .B(n13343), .Z(n8640) );
  AND U13329 ( .A(n13344), .B(n13345), .Z(n13343) );
  AND U13330 ( .A(n13346), .B(n13347), .Z(n13345) );
  AND U13331 ( .A(n13348), .B(n13349), .Z(n13347) );
  XNOR U13332 ( .A(y[983]), .B(x[983]), .Z(n13349) );
  AND U13333 ( .A(n13350), .B(n13351), .Z(n13348) );
  XNOR U13334 ( .A(y[981]), .B(x[981]), .Z(n13351) );
  XNOR U13335 ( .A(y[982]), .B(x[982]), .Z(n13350) );
  AND U13336 ( .A(n13352), .B(n13353), .Z(n13346) );
  XNOR U13337 ( .A(y[984]), .B(x[984]), .Z(n13353) );
  XNOR U13338 ( .A(y[985]), .B(x[985]), .Z(n13352) );
  AND U13339 ( .A(n13354), .B(n13355), .Z(n13344) );
  AND U13340 ( .A(n13356), .B(n13357), .Z(n13355) );
  XNOR U13341 ( .A(y[986]), .B(x[986]), .Z(n13357) );
  XNOR U13342 ( .A(y[987]), .B(x[987]), .Z(n13356) );
  AND U13343 ( .A(n13358), .B(n13359), .Z(n13354) );
  XNOR U13344 ( .A(y[988]), .B(x[988]), .Z(n13359) );
  XNOR U13345 ( .A(y[989]), .B(x[989]), .Z(n13358) );
  AND U13346 ( .A(n13360), .B(n13361), .Z(n13342) );
  AND U13347 ( .A(n13362), .B(n13363), .Z(n13361) );
  AND U13348 ( .A(n13364), .B(n13365), .Z(n13363) );
  XNOR U13349 ( .A(y[992]), .B(x[992]), .Z(n13365) );
  AND U13350 ( .A(n13366), .B(n13367), .Z(n13364) );
  XNOR U13351 ( .A(y[990]), .B(x[990]), .Z(n13367) );
  XNOR U13352 ( .A(y[991]), .B(x[991]), .Z(n13366) );
  AND U13353 ( .A(n13368), .B(n13369), .Z(n13362) );
  XNOR U13354 ( .A(y[993]), .B(x[993]), .Z(n13369) );
  XNOR U13355 ( .A(y[994]), .B(x[994]), .Z(n13368) );
  AND U13356 ( .A(n13370), .B(n13371), .Z(n13360) );
  AND U13357 ( .A(n13372), .B(n13373), .Z(n13371) );
  XNOR U13358 ( .A(y[995]), .B(x[995]), .Z(n13373) );
  XNOR U13359 ( .A(y[996]), .B(x[996]), .Z(n13372) );
  AND U13360 ( .A(n13374), .B(n13375), .Z(n13370) );
  XNOR U13361 ( .A(y[997]), .B(x[997]), .Z(n13375) );
  XNOR U13362 ( .A(y[998]), .B(x[998]), .Z(n13374) );
  AND U13363 ( .A(n13376), .B(n13377), .Z(n8638) );
  AND U13364 ( .A(n13378), .B(n13379), .Z(n13377) );
  AND U13365 ( .A(n13380), .B(n13381), .Z(n13379) );
  AND U13366 ( .A(n13382), .B(n13383), .Z(n13381) );
  AND U13367 ( .A(n13384), .B(n13385), .Z(n13383) );
  XNOR U13368 ( .A(y[1001]), .B(x[1001]), .Z(n13385) );
  AND U13369 ( .A(n13386), .B(n13387), .Z(n13384) );
  XNOR U13370 ( .A(y[999]), .B(x[999]), .Z(n13387) );
  XNOR U13371 ( .A(y[1000]), .B(x[1000]), .Z(n13386) );
  AND U13372 ( .A(n13388), .B(n13389), .Z(n13382) );
  XNOR U13373 ( .A(y[1002]), .B(x[1002]), .Z(n13389) );
  XNOR U13374 ( .A(y[1003]), .B(x[1003]), .Z(n13388) );
  AND U13375 ( .A(n13390), .B(n13391), .Z(n13380) );
  AND U13376 ( .A(n13392), .B(n13393), .Z(n13391) );
  XNOR U13377 ( .A(y[1510]), .B(x[1510]), .Z(n13393) );
  AND U13378 ( .A(n13394), .B(n13395), .Z(n13392) );
  XNOR U13379 ( .A(y[1508]), .B(x[1508]), .Z(n13395) );
  XNOR U13380 ( .A(y[1509]), .B(x[1509]), .Z(n13394) );
  AND U13381 ( .A(n13396), .B(n13397), .Z(n13390) );
  XNOR U13382 ( .A(y[1511]), .B(x[1511]), .Z(n13397) );
  XNOR U13383 ( .A(y[1512]), .B(x[1512]), .Z(n13396) );
  AND U13384 ( .A(n13398), .B(n13399), .Z(n13378) );
  AND U13385 ( .A(n13400), .B(n13401), .Z(n13399) );
  AND U13386 ( .A(n13402), .B(n13403), .Z(n13401) );
  XNOR U13387 ( .A(y[1787]), .B(x[1787]), .Z(n13403) );
  AND U13388 ( .A(n13404), .B(n13405), .Z(n13402) );
  XNOR U13389 ( .A(y[1513]), .B(x[1513]), .Z(n13405) );
  XNOR U13390 ( .A(y[1786]), .B(x[1786]), .Z(n13404) );
  AND U13391 ( .A(n13406), .B(n13407), .Z(n13400) );
  XNOR U13392 ( .A(y[1788]), .B(x[1788]), .Z(n13407) );
  XNOR U13393 ( .A(y[1789]), .B(x[1789]), .Z(n13406) );
  AND U13394 ( .A(n13408), .B(n13409), .Z(n13398) );
  AND U13395 ( .A(n13410), .B(n13411), .Z(n13409) );
  XNOR U13396 ( .A(y[1790]), .B(x[1790]), .Z(n13411) );
  XNOR U13397 ( .A(y[1791]), .B(x[1791]), .Z(n13410) );
  AND U13398 ( .A(n13412), .B(n13413), .Z(n13408) );
  XNOR U13399 ( .A(y[1792]), .B(x[1792]), .Z(n13413) );
  XNOR U13400 ( .A(y[1793]), .B(x[1793]), .Z(n13412) );
  AND U13401 ( .A(n13414), .B(n13415), .Z(n13376) );
  AND U13402 ( .A(n13416), .B(n13417), .Z(n13415) );
  AND U13403 ( .A(n13418), .B(n13419), .Z(n13417) );
  AND U13404 ( .A(n13420), .B(n13421), .Z(n13419) );
  XNOR U13405 ( .A(y[1796]), .B(x[1796]), .Z(n13421) );
  AND U13406 ( .A(n13422), .B(n13423), .Z(n13420) );
  XNOR U13407 ( .A(y[1794]), .B(x[1794]), .Z(n13423) );
  XNOR U13408 ( .A(y[1795]), .B(x[1795]), .Z(n13422) );
  AND U13409 ( .A(n13424), .B(n13425), .Z(n13418) );
  XNOR U13410 ( .A(y[1797]), .B(x[1797]), .Z(n13425) );
  XNOR U13411 ( .A(y[1798]), .B(x[1798]), .Z(n13424) );
  AND U13412 ( .A(n13426), .B(n13427), .Z(n13416) );
  AND U13413 ( .A(n13428), .B(n13429), .Z(n13427) );
  XNOR U13414 ( .A(y[1799]), .B(x[1799]), .Z(n13429) );
  XNOR U13415 ( .A(y[1800]), .B(x[1800]), .Z(n13428) );
  AND U13416 ( .A(n13430), .B(n13431), .Z(n13426) );
  XNOR U13417 ( .A(y[1801]), .B(x[1801]), .Z(n13431) );
  XNOR U13418 ( .A(y[1802]), .B(x[1802]), .Z(n13430) );
  AND U13419 ( .A(n13432), .B(n13433), .Z(n13414) );
  AND U13420 ( .A(n13434), .B(n13435), .Z(n13433) );
  AND U13421 ( .A(n13436), .B(n13437), .Z(n13435) );
  XNOR U13422 ( .A(y[1805]), .B(x[1805]), .Z(n13437) );
  AND U13423 ( .A(n13438), .B(n13439), .Z(n13436) );
  XNOR U13424 ( .A(y[1803]), .B(x[1803]), .Z(n13439) );
  XNOR U13425 ( .A(y[1804]), .B(x[1804]), .Z(n13438) );
  AND U13426 ( .A(n13440), .B(n13441), .Z(n13434) );
  XNOR U13427 ( .A(y[1806]), .B(x[1806]), .Z(n13441) );
  XNOR U13428 ( .A(y[1807]), .B(x[1807]), .Z(n13440) );
  AND U13429 ( .A(n13442), .B(n13443), .Z(n13432) );
  AND U13430 ( .A(n13444), .B(n13445), .Z(n13443) );
  XNOR U13431 ( .A(y[1808]), .B(x[1808]), .Z(n13445) );
  XNOR U13432 ( .A(y[1809]), .B(x[1809]), .Z(n13444) );
  AND U13433 ( .A(n13446), .B(n13447), .Z(n13442) );
  XNOR U13434 ( .A(y[1810]), .B(x[1810]), .Z(n13447) );
  XNOR U13435 ( .A(y[1811]), .B(x[1811]), .Z(n13446) );
  AND U13436 ( .A(n13448), .B(n13449), .Z(n8636) );
  AND U13437 ( .A(n13450), .B(n13451), .Z(n13449) );
  AND U13438 ( .A(n13452), .B(n13453), .Z(n13451) );
  AND U13439 ( .A(n13454), .B(n13455), .Z(n13453) );
  AND U13440 ( .A(n13456), .B(n13457), .Z(n13455) );
  AND U13441 ( .A(n13458), .B(n13459), .Z(n13457) );
  XNOR U13442 ( .A(y[1814]), .B(x[1814]), .Z(n13459) );
  AND U13443 ( .A(n13460), .B(n13461), .Z(n13458) );
  XNOR U13444 ( .A(y[1812]), .B(x[1812]), .Z(n13461) );
  XNOR U13445 ( .A(y[1813]), .B(x[1813]), .Z(n13460) );
  AND U13446 ( .A(n13462), .B(n13463), .Z(n13456) );
  XNOR U13447 ( .A(y[1815]), .B(x[1815]), .Z(n13463) );
  XNOR U13448 ( .A(y[1816]), .B(x[1816]), .Z(n13462) );
  AND U13449 ( .A(n13464), .B(n13465), .Z(n13454) );
  AND U13450 ( .A(n13466), .B(n13467), .Z(n13465) );
  XNOR U13451 ( .A(y[1819]), .B(x[1819]), .Z(n13467) );
  AND U13452 ( .A(n13468), .B(n13469), .Z(n13466) );
  XNOR U13453 ( .A(y[1817]), .B(x[1817]), .Z(n13469) );
  XNOR U13454 ( .A(y[1818]), .B(x[1818]), .Z(n13468) );
  AND U13455 ( .A(n13470), .B(n13471), .Z(n13464) );
  XNOR U13456 ( .A(y[1820]), .B(x[1820]), .Z(n13471) );
  XNOR U13457 ( .A(y[1821]), .B(x[1821]), .Z(n13470) );
  AND U13458 ( .A(n13472), .B(n13473), .Z(n13452) );
  AND U13459 ( .A(n13474), .B(n13475), .Z(n13473) );
  AND U13460 ( .A(n13476), .B(n13477), .Z(n13475) );
  XNOR U13461 ( .A(y[1824]), .B(x[1824]), .Z(n13477) );
  AND U13462 ( .A(n13478), .B(n13479), .Z(n13476) );
  XNOR U13463 ( .A(y[1822]), .B(x[1822]), .Z(n13479) );
  XNOR U13464 ( .A(y[1823]), .B(x[1823]), .Z(n13478) );
  AND U13465 ( .A(n13480), .B(n13481), .Z(n13474) );
  XNOR U13466 ( .A(y[1825]), .B(x[1825]), .Z(n13481) );
  XNOR U13467 ( .A(y[1826]), .B(x[1826]), .Z(n13480) );
  AND U13468 ( .A(n13482), .B(n13483), .Z(n13472) );
  AND U13469 ( .A(n13484), .B(n13485), .Z(n13483) );
  XNOR U13470 ( .A(y[1827]), .B(x[1827]), .Z(n13485) );
  XNOR U13471 ( .A(y[1828]), .B(x[1828]), .Z(n13484) );
  AND U13472 ( .A(n13486), .B(n13487), .Z(n13482) );
  XNOR U13473 ( .A(y[1829]), .B(x[1829]), .Z(n13487) );
  XNOR U13474 ( .A(y[1830]), .B(x[1830]), .Z(n13486) );
  AND U13475 ( .A(n13488), .B(n13489), .Z(n13450) );
  AND U13476 ( .A(n13490), .B(n13491), .Z(n13489) );
  AND U13477 ( .A(n13492), .B(n13493), .Z(n13491) );
  AND U13478 ( .A(n13494), .B(n13495), .Z(n13493) );
  XNOR U13479 ( .A(y[1833]), .B(x[1833]), .Z(n13495) );
  AND U13480 ( .A(n13496), .B(n13497), .Z(n13494) );
  XNOR U13481 ( .A(y[1831]), .B(x[1831]), .Z(n13497) );
  XNOR U13482 ( .A(y[1832]), .B(x[1832]), .Z(n13496) );
  AND U13483 ( .A(n13498), .B(n13499), .Z(n13492) );
  XNOR U13484 ( .A(y[1834]), .B(x[1834]), .Z(n13499) );
  XNOR U13485 ( .A(y[1835]), .B(x[1835]), .Z(n13498) );
  AND U13486 ( .A(n13500), .B(n13501), .Z(n13490) );
  AND U13487 ( .A(n13502), .B(n13503), .Z(n13501) );
  XNOR U13488 ( .A(y[1836]), .B(x[1836]), .Z(n13503) );
  XNOR U13489 ( .A(y[1837]), .B(x[1837]), .Z(n13502) );
  AND U13490 ( .A(n13504), .B(n13505), .Z(n13500) );
  XNOR U13491 ( .A(y[1838]), .B(x[1838]), .Z(n13505) );
  XNOR U13492 ( .A(y[1839]), .B(x[1839]), .Z(n13504) );
  AND U13493 ( .A(n13506), .B(n13507), .Z(n13488) );
  AND U13494 ( .A(n13508), .B(n13509), .Z(n13507) );
  AND U13495 ( .A(n13510), .B(n13511), .Z(n13509) );
  XNOR U13496 ( .A(y[1842]), .B(x[1842]), .Z(n13511) );
  AND U13497 ( .A(n13512), .B(n13513), .Z(n13510) );
  XNOR U13498 ( .A(y[1840]), .B(x[1840]), .Z(n13513) );
  XNOR U13499 ( .A(y[1841]), .B(x[1841]), .Z(n13512) );
  AND U13500 ( .A(n13514), .B(n13515), .Z(n13508) );
  XNOR U13501 ( .A(y[1843]), .B(x[1843]), .Z(n13515) );
  XNOR U13502 ( .A(y[1844]), .B(x[1844]), .Z(n13514) );
  AND U13503 ( .A(n13516), .B(n13517), .Z(n13506) );
  AND U13504 ( .A(n13518), .B(n13519), .Z(n13517) );
  XNOR U13505 ( .A(y[1845]), .B(x[1845]), .Z(n13519) );
  XNOR U13506 ( .A(y[1846]), .B(x[1846]), .Z(n13518) );
  AND U13507 ( .A(n13520), .B(n13521), .Z(n13516) );
  XNOR U13508 ( .A(y[1847]), .B(x[1847]), .Z(n13521) );
  XNOR U13509 ( .A(y[1848]), .B(x[1848]), .Z(n13520) );
  AND U13510 ( .A(n13522), .B(n13523), .Z(n13448) );
  AND U13511 ( .A(n13524), .B(n13525), .Z(n13523) );
  AND U13512 ( .A(n13526), .B(n13527), .Z(n13525) );
  AND U13513 ( .A(n13528), .B(n13529), .Z(n13527) );
  AND U13514 ( .A(n13530), .B(n13531), .Z(n13529) );
  XNOR U13515 ( .A(y[1851]), .B(x[1851]), .Z(n13531) );
  AND U13516 ( .A(n13532), .B(n13533), .Z(n13530) );
  XNOR U13517 ( .A(y[1849]), .B(x[1849]), .Z(n13533) );
  XNOR U13518 ( .A(y[1850]), .B(x[1850]), .Z(n13532) );
  AND U13519 ( .A(n13534), .B(n13535), .Z(n13528) );
  XNOR U13520 ( .A(y[1852]), .B(x[1852]), .Z(n13535) );
  XNOR U13521 ( .A(y[1853]), .B(x[1853]), .Z(n13534) );
  AND U13522 ( .A(n13536), .B(n13537), .Z(n13526) );
  AND U13523 ( .A(n13538), .B(n13539), .Z(n13537) );
  XNOR U13524 ( .A(y[1856]), .B(x[1856]), .Z(n13539) );
  AND U13525 ( .A(n13540), .B(n13541), .Z(n13538) );
  XNOR U13526 ( .A(y[1854]), .B(x[1854]), .Z(n13541) );
  XNOR U13527 ( .A(y[1855]), .B(x[1855]), .Z(n13540) );
  AND U13528 ( .A(n13542), .B(n13543), .Z(n13536) );
  XNOR U13529 ( .A(y[1857]), .B(x[1857]), .Z(n13543) );
  XNOR U13530 ( .A(y[1858]), .B(x[1858]), .Z(n13542) );
  AND U13531 ( .A(n13544), .B(n13545), .Z(n13524) );
  AND U13532 ( .A(n13546), .B(n13547), .Z(n13545) );
  AND U13533 ( .A(n13548), .B(n13549), .Z(n13547) );
  XNOR U13534 ( .A(y[1861]), .B(x[1861]), .Z(n13549) );
  AND U13535 ( .A(n13550), .B(n13551), .Z(n13548) );
  XNOR U13536 ( .A(y[1859]), .B(x[1859]), .Z(n13551) );
  XNOR U13537 ( .A(y[1860]), .B(x[1860]), .Z(n13550) );
  AND U13538 ( .A(n13552), .B(n13553), .Z(n13546) );
  XNOR U13539 ( .A(y[1862]), .B(x[1862]), .Z(n13553) );
  XNOR U13540 ( .A(y[1863]), .B(x[1863]), .Z(n13552) );
  AND U13541 ( .A(n13554), .B(n13555), .Z(n13544) );
  AND U13542 ( .A(n13556), .B(n13557), .Z(n13555) );
  XNOR U13543 ( .A(y[1864]), .B(x[1864]), .Z(n13557) );
  XNOR U13544 ( .A(y[1865]), .B(x[1865]), .Z(n13556) );
  AND U13545 ( .A(n13558), .B(n13559), .Z(n13554) );
  XNOR U13546 ( .A(y[1866]), .B(x[1866]), .Z(n13559) );
  XNOR U13547 ( .A(y[1867]), .B(x[1867]), .Z(n13558) );
  AND U13548 ( .A(n13560), .B(n13561), .Z(n13522) );
  AND U13549 ( .A(n13562), .B(n13563), .Z(n13561) );
  AND U13550 ( .A(n13564), .B(n13565), .Z(n13563) );
  AND U13551 ( .A(n13566), .B(n13567), .Z(n13565) );
  XNOR U13552 ( .A(y[1870]), .B(x[1870]), .Z(n13567) );
  AND U13553 ( .A(n13568), .B(n13569), .Z(n13566) );
  XNOR U13554 ( .A(y[1868]), .B(x[1868]), .Z(n13569) );
  XNOR U13555 ( .A(y[1869]), .B(x[1869]), .Z(n13568) );
  AND U13556 ( .A(n13570), .B(n13571), .Z(n13564) );
  XNOR U13557 ( .A(y[1871]), .B(x[1871]), .Z(n13571) );
  XNOR U13558 ( .A(y[1872]), .B(x[1872]), .Z(n13570) );
  AND U13559 ( .A(n13572), .B(n13573), .Z(n13562) );
  AND U13560 ( .A(n13574), .B(n13575), .Z(n13573) );
  XNOR U13561 ( .A(y[1873]), .B(x[1873]), .Z(n13575) );
  XNOR U13562 ( .A(y[1874]), .B(x[1874]), .Z(n13574) );
  AND U13563 ( .A(n13576), .B(n13577), .Z(n13572) );
  XNOR U13564 ( .A(y[1875]), .B(x[1875]), .Z(n13577) );
  XNOR U13565 ( .A(y[1876]), .B(x[1876]), .Z(n13576) );
  AND U13566 ( .A(n13578), .B(n13579), .Z(n13560) );
  AND U13567 ( .A(n13580), .B(n13581), .Z(n13579) );
  AND U13568 ( .A(n13582), .B(n13583), .Z(n13581) );
  XNOR U13569 ( .A(y[1879]), .B(x[1879]), .Z(n13583) );
  AND U13570 ( .A(n13584), .B(n13585), .Z(n13582) );
  XNOR U13571 ( .A(y[1877]), .B(x[1877]), .Z(n13585) );
  XNOR U13572 ( .A(y[1878]), .B(x[1878]), .Z(n13584) );
  AND U13573 ( .A(n13586), .B(n13587), .Z(n13580) );
  XNOR U13574 ( .A(y[1880]), .B(x[1880]), .Z(n13587) );
  XNOR U13575 ( .A(y[1881]), .B(x[1881]), .Z(n13586) );
  AND U13576 ( .A(n13588), .B(n13589), .Z(n13578) );
  AND U13577 ( .A(n13590), .B(n13591), .Z(n13589) );
  XNOR U13578 ( .A(y[1882]), .B(x[1882]), .Z(n13591) );
  XNOR U13579 ( .A(y[1883]), .B(x[1883]), .Z(n13590) );
  AND U13580 ( .A(n13592), .B(n13593), .Z(n13588) );
  XNOR U13581 ( .A(y[1884]), .B(x[1884]), .Z(n13593) );
  XNOR U13582 ( .A(y[1885]), .B(x[1885]), .Z(n13592) );
  AND U13583 ( .A(n13594), .B(n13595), .Z(n8634) );
  AND U13584 ( .A(n13596), .B(n13597), .Z(n13595) );
  AND U13585 ( .A(n13598), .B(n13599), .Z(n13597) );
  AND U13586 ( .A(n13600), .B(n13601), .Z(n13599) );
  AND U13587 ( .A(n13602), .B(n13603), .Z(n13601) );
  AND U13588 ( .A(n13604), .B(n13605), .Z(n13603) );
  AND U13589 ( .A(n13606), .B(n13607), .Z(n13605) );
  XNOR U13590 ( .A(y[1888]), .B(x[1888]), .Z(n13607) );
  AND U13591 ( .A(n13608), .B(n13609), .Z(n13606) );
  XNOR U13592 ( .A(y[1886]), .B(x[1886]), .Z(n13609) );
  XNOR U13593 ( .A(y[1887]), .B(x[1887]), .Z(n13608) );
  AND U13594 ( .A(n13610), .B(n13611), .Z(n13604) );
  XNOR U13595 ( .A(y[1889]), .B(x[1889]), .Z(n13611) );
  XNOR U13596 ( .A(y[1890]), .B(x[1890]), .Z(n13610) );
  AND U13597 ( .A(n13612), .B(n13613), .Z(n13602) );
  AND U13598 ( .A(n13614), .B(n13615), .Z(n13613) );
  XNOR U13599 ( .A(y[1893]), .B(x[1893]), .Z(n13615) );
  AND U13600 ( .A(n13616), .B(n13617), .Z(n13614) );
  XNOR U13601 ( .A(y[1891]), .B(x[1891]), .Z(n13617) );
  XNOR U13602 ( .A(y[1892]), .B(x[1892]), .Z(n13616) );
  AND U13603 ( .A(n13618), .B(n13619), .Z(n13612) );
  XNOR U13604 ( .A(y[1894]), .B(x[1894]), .Z(n13619) );
  XNOR U13605 ( .A(y[1895]), .B(x[1895]), .Z(n13618) );
  AND U13606 ( .A(n13620), .B(n13621), .Z(n13600) );
  AND U13607 ( .A(n13622), .B(n13623), .Z(n13621) );
  AND U13608 ( .A(n13624), .B(n13625), .Z(n13623) );
  XNOR U13609 ( .A(y[1898]), .B(x[1898]), .Z(n13625) );
  AND U13610 ( .A(n13626), .B(n13627), .Z(n13624) );
  XNOR U13611 ( .A(y[1896]), .B(x[1896]), .Z(n13627) );
  XNOR U13612 ( .A(y[1897]), .B(x[1897]), .Z(n13626) );
  AND U13613 ( .A(n13628), .B(n13629), .Z(n13622) );
  XNOR U13614 ( .A(y[1899]), .B(x[1899]), .Z(n13629) );
  XNOR U13615 ( .A(y[1900]), .B(x[1900]), .Z(n13628) );
  AND U13616 ( .A(n13630), .B(n13631), .Z(n13620) );
  AND U13617 ( .A(n13632), .B(n13633), .Z(n13631) );
  XNOR U13618 ( .A(y[1901]), .B(x[1901]), .Z(n13633) );
  XNOR U13619 ( .A(y[1902]), .B(x[1902]), .Z(n13632) );
  AND U13620 ( .A(n13634), .B(n13635), .Z(n13630) );
  XNOR U13621 ( .A(y[1903]), .B(x[1903]), .Z(n13635) );
  XNOR U13622 ( .A(y[1904]), .B(x[1904]), .Z(n13634) );
  AND U13623 ( .A(n13636), .B(n13637), .Z(n13598) );
  AND U13624 ( .A(n13638), .B(n13639), .Z(n13637) );
  AND U13625 ( .A(n13640), .B(n13641), .Z(n13639) );
  AND U13626 ( .A(n13642), .B(n13643), .Z(n13641) );
  XNOR U13627 ( .A(y[1907]), .B(x[1907]), .Z(n13643) );
  AND U13628 ( .A(n13644), .B(n13645), .Z(n13642) );
  XNOR U13629 ( .A(y[1905]), .B(x[1905]), .Z(n13645) );
  XNOR U13630 ( .A(y[1906]), .B(x[1906]), .Z(n13644) );
  AND U13631 ( .A(n13646), .B(n13647), .Z(n13640) );
  XNOR U13632 ( .A(y[1908]), .B(x[1908]), .Z(n13647) );
  XNOR U13633 ( .A(y[1909]), .B(x[1909]), .Z(n13646) );
  AND U13634 ( .A(n13648), .B(n13649), .Z(n13638) );
  AND U13635 ( .A(n13650), .B(n13651), .Z(n13649) );
  XNOR U13636 ( .A(y[1910]), .B(x[1910]), .Z(n13651) );
  XNOR U13637 ( .A(y[1911]), .B(x[1911]), .Z(n13650) );
  AND U13638 ( .A(n13652), .B(n13653), .Z(n13648) );
  XNOR U13639 ( .A(y[1912]), .B(x[1912]), .Z(n13653) );
  XNOR U13640 ( .A(y[1913]), .B(x[1913]), .Z(n13652) );
  AND U13641 ( .A(n13654), .B(n13655), .Z(n13636) );
  AND U13642 ( .A(n13656), .B(n13657), .Z(n13655) );
  AND U13643 ( .A(n13658), .B(n13659), .Z(n13657) );
  XNOR U13644 ( .A(y[1916]), .B(x[1916]), .Z(n13659) );
  AND U13645 ( .A(n13660), .B(n13661), .Z(n13658) );
  XNOR U13646 ( .A(y[1914]), .B(x[1914]), .Z(n13661) );
  XNOR U13647 ( .A(y[1915]), .B(x[1915]), .Z(n13660) );
  AND U13648 ( .A(n13662), .B(n13663), .Z(n13656) );
  XNOR U13649 ( .A(y[1917]), .B(x[1917]), .Z(n13663) );
  XNOR U13650 ( .A(y[1918]), .B(x[1918]), .Z(n13662) );
  AND U13651 ( .A(n13664), .B(n13665), .Z(n13654) );
  AND U13652 ( .A(n13666), .B(n13667), .Z(n13665) );
  XNOR U13653 ( .A(y[1919]), .B(x[1919]), .Z(n13667) );
  XNOR U13654 ( .A(y[1920]), .B(x[1920]), .Z(n13666) );
  AND U13655 ( .A(n13668), .B(n13669), .Z(n13664) );
  XNOR U13656 ( .A(y[1921]), .B(x[1921]), .Z(n13669) );
  XNOR U13657 ( .A(y[1922]), .B(x[1922]), .Z(n13668) );
  AND U13658 ( .A(n13670), .B(n13671), .Z(n13596) );
  AND U13659 ( .A(n13672), .B(n13673), .Z(n13671) );
  AND U13660 ( .A(n13674), .B(n13675), .Z(n13673) );
  AND U13661 ( .A(n13676), .B(n13677), .Z(n13675) );
  AND U13662 ( .A(n13678), .B(n13679), .Z(n13677) );
  XNOR U13663 ( .A(y[1925]), .B(x[1925]), .Z(n13679) );
  AND U13664 ( .A(n13680), .B(n13681), .Z(n13678) );
  XNOR U13665 ( .A(y[1923]), .B(x[1923]), .Z(n13681) );
  XNOR U13666 ( .A(y[1924]), .B(x[1924]), .Z(n13680) );
  AND U13667 ( .A(n13682), .B(n13683), .Z(n13676) );
  XNOR U13668 ( .A(y[1926]), .B(x[1926]), .Z(n13683) );
  XNOR U13669 ( .A(y[1927]), .B(x[1927]), .Z(n13682) );
  AND U13670 ( .A(n13684), .B(n13685), .Z(n13674) );
  AND U13671 ( .A(n13686), .B(n13687), .Z(n13685) );
  XNOR U13672 ( .A(y[1930]), .B(x[1930]), .Z(n13687) );
  AND U13673 ( .A(n13688), .B(n13689), .Z(n13686) );
  XNOR U13674 ( .A(y[1928]), .B(x[1928]), .Z(n13689) );
  XNOR U13675 ( .A(y[1929]), .B(x[1929]), .Z(n13688) );
  AND U13676 ( .A(n13690), .B(n13691), .Z(n13684) );
  XNOR U13677 ( .A(y[1931]), .B(x[1931]), .Z(n13691) );
  XNOR U13678 ( .A(y[1932]), .B(x[1932]), .Z(n13690) );
  AND U13679 ( .A(n13692), .B(n13693), .Z(n13672) );
  AND U13680 ( .A(n13694), .B(n13695), .Z(n13693) );
  AND U13681 ( .A(n13696), .B(n13697), .Z(n13695) );
  XNOR U13682 ( .A(y[1935]), .B(x[1935]), .Z(n13697) );
  AND U13683 ( .A(n13698), .B(n13699), .Z(n13696) );
  XNOR U13684 ( .A(y[1933]), .B(x[1933]), .Z(n13699) );
  XNOR U13685 ( .A(y[1934]), .B(x[1934]), .Z(n13698) );
  AND U13686 ( .A(n13700), .B(n13701), .Z(n13694) );
  XNOR U13687 ( .A(y[1936]), .B(x[1936]), .Z(n13701) );
  XNOR U13688 ( .A(y[1937]), .B(x[1937]), .Z(n13700) );
  AND U13689 ( .A(n13702), .B(n13703), .Z(n13692) );
  AND U13690 ( .A(n13704), .B(n13705), .Z(n13703) );
  XNOR U13691 ( .A(y[1938]), .B(x[1938]), .Z(n13705) );
  XNOR U13692 ( .A(y[1939]), .B(x[1939]), .Z(n13704) );
  AND U13693 ( .A(n13706), .B(n13707), .Z(n13702) );
  XNOR U13694 ( .A(y[1940]), .B(x[1940]), .Z(n13707) );
  XNOR U13695 ( .A(y[1941]), .B(x[1941]), .Z(n13706) );
  AND U13696 ( .A(n13708), .B(n13709), .Z(n13670) );
  AND U13697 ( .A(n13710), .B(n13711), .Z(n13709) );
  AND U13698 ( .A(n13712), .B(n13713), .Z(n13711) );
  AND U13699 ( .A(n13714), .B(n13715), .Z(n13713) );
  XNOR U13700 ( .A(y[1944]), .B(x[1944]), .Z(n13715) );
  AND U13701 ( .A(n13716), .B(n13717), .Z(n13714) );
  XNOR U13702 ( .A(y[1942]), .B(x[1942]), .Z(n13717) );
  XNOR U13703 ( .A(y[1943]), .B(x[1943]), .Z(n13716) );
  AND U13704 ( .A(n13718), .B(n13719), .Z(n13712) );
  XNOR U13705 ( .A(y[1945]), .B(x[1945]), .Z(n13719) );
  XNOR U13706 ( .A(y[1946]), .B(x[1946]), .Z(n13718) );
  AND U13707 ( .A(n13720), .B(n13721), .Z(n13710) );
  AND U13708 ( .A(n13722), .B(n13723), .Z(n13721) );
  XNOR U13709 ( .A(y[1947]), .B(x[1947]), .Z(n13723) );
  XNOR U13710 ( .A(y[1948]), .B(x[1948]), .Z(n13722) );
  AND U13711 ( .A(n13724), .B(n13725), .Z(n13720) );
  XNOR U13712 ( .A(y[1949]), .B(x[1949]), .Z(n13725) );
  XNOR U13713 ( .A(y[1950]), .B(x[1950]), .Z(n13724) );
  AND U13714 ( .A(n13726), .B(n13727), .Z(n13708) );
  AND U13715 ( .A(n13728), .B(n13729), .Z(n13727) );
  AND U13716 ( .A(n13730), .B(n13731), .Z(n13729) );
  XNOR U13717 ( .A(y[1953]), .B(x[1953]), .Z(n13731) );
  AND U13718 ( .A(n13732), .B(n13733), .Z(n13730) );
  XNOR U13719 ( .A(y[1951]), .B(x[1951]), .Z(n13733) );
  XNOR U13720 ( .A(y[1952]), .B(x[1952]), .Z(n13732) );
  AND U13721 ( .A(n13734), .B(n13735), .Z(n13728) );
  XNOR U13722 ( .A(y[1954]), .B(x[1954]), .Z(n13735) );
  XNOR U13723 ( .A(y[1955]), .B(x[1955]), .Z(n13734) );
  AND U13724 ( .A(n13736), .B(n13737), .Z(n13726) );
  AND U13725 ( .A(n13738), .B(n13739), .Z(n13737) );
  XNOR U13726 ( .A(y[1956]), .B(x[1956]), .Z(n13739) );
  XNOR U13727 ( .A(y[1957]), .B(x[1957]), .Z(n13738) );
  AND U13728 ( .A(n13740), .B(n13741), .Z(n13736) );
  XNOR U13729 ( .A(y[1958]), .B(x[1958]), .Z(n13741) );
  XNOR U13730 ( .A(y[1959]), .B(x[1959]), .Z(n13740) );
  AND U13731 ( .A(n13742), .B(n13743), .Z(n13594) );
  AND U13732 ( .A(n13744), .B(n13745), .Z(n13743) );
  AND U13733 ( .A(n13746), .B(n13747), .Z(n13745) );
  AND U13734 ( .A(n13748), .B(n13749), .Z(n13747) );
  AND U13735 ( .A(n13750), .B(n13751), .Z(n13749) );
  AND U13736 ( .A(n13752), .B(n13753), .Z(n13751) );
  XNOR U13737 ( .A(y[1962]), .B(x[1962]), .Z(n13753) );
  AND U13738 ( .A(n13754), .B(n13755), .Z(n13752) );
  XNOR U13739 ( .A(y[1960]), .B(x[1960]), .Z(n13755) );
  XNOR U13740 ( .A(y[1961]), .B(x[1961]), .Z(n13754) );
  AND U13741 ( .A(n13756), .B(n13757), .Z(n13750) );
  XNOR U13742 ( .A(y[1963]), .B(x[1963]), .Z(n13757) );
  XNOR U13743 ( .A(y[1964]), .B(x[1964]), .Z(n13756) );
  AND U13744 ( .A(n13758), .B(n13759), .Z(n13748) );
  AND U13745 ( .A(n13760), .B(n13761), .Z(n13759) );
  XNOR U13746 ( .A(y[1967]), .B(x[1967]), .Z(n13761) );
  AND U13747 ( .A(n13762), .B(n13763), .Z(n13760) );
  XNOR U13748 ( .A(y[1965]), .B(x[1965]), .Z(n13763) );
  XNOR U13749 ( .A(y[1966]), .B(x[1966]), .Z(n13762) );
  AND U13750 ( .A(n13764), .B(n13765), .Z(n13758) );
  XNOR U13751 ( .A(y[1968]), .B(x[1968]), .Z(n13765) );
  XNOR U13752 ( .A(y[1969]), .B(x[1969]), .Z(n13764) );
  AND U13753 ( .A(n13766), .B(n13767), .Z(n13746) );
  AND U13754 ( .A(n13768), .B(n13769), .Z(n13767) );
  AND U13755 ( .A(n13770), .B(n13771), .Z(n13769) );
  XNOR U13756 ( .A(y[1972]), .B(x[1972]), .Z(n13771) );
  AND U13757 ( .A(n13772), .B(n13773), .Z(n13770) );
  XNOR U13758 ( .A(y[1970]), .B(x[1970]), .Z(n13773) );
  XNOR U13759 ( .A(y[1971]), .B(x[1971]), .Z(n13772) );
  AND U13760 ( .A(n13774), .B(n13775), .Z(n13768) );
  XNOR U13761 ( .A(y[1973]), .B(x[1973]), .Z(n13775) );
  XNOR U13762 ( .A(y[1974]), .B(x[1974]), .Z(n13774) );
  AND U13763 ( .A(n13776), .B(n13777), .Z(n13766) );
  AND U13764 ( .A(n13778), .B(n13779), .Z(n13777) );
  XNOR U13765 ( .A(y[1975]), .B(x[1975]), .Z(n13779) );
  XNOR U13766 ( .A(y[1976]), .B(x[1976]), .Z(n13778) );
  AND U13767 ( .A(n13780), .B(n13781), .Z(n13776) );
  XNOR U13768 ( .A(y[1977]), .B(x[1977]), .Z(n13781) );
  XNOR U13769 ( .A(y[1978]), .B(x[1978]), .Z(n13780) );
  AND U13770 ( .A(n13782), .B(n13783), .Z(n13744) );
  AND U13771 ( .A(n13784), .B(n13785), .Z(n13783) );
  AND U13772 ( .A(n13786), .B(n13787), .Z(n13785) );
  AND U13773 ( .A(n13788), .B(n13789), .Z(n13787) );
  XNOR U13774 ( .A(y[1981]), .B(x[1981]), .Z(n13789) );
  AND U13775 ( .A(n13790), .B(n13791), .Z(n13788) );
  XNOR U13776 ( .A(y[1979]), .B(x[1979]), .Z(n13791) );
  XNOR U13777 ( .A(y[1980]), .B(x[1980]), .Z(n13790) );
  AND U13778 ( .A(n13792), .B(n13793), .Z(n13786) );
  XNOR U13779 ( .A(y[1982]), .B(x[1982]), .Z(n13793) );
  XNOR U13780 ( .A(y[1983]), .B(x[1983]), .Z(n13792) );
  AND U13781 ( .A(n13794), .B(n13795), .Z(n13784) );
  AND U13782 ( .A(n13796), .B(n13797), .Z(n13795) );
  XNOR U13783 ( .A(y[1984]), .B(x[1984]), .Z(n13797) );
  XNOR U13784 ( .A(y[1985]), .B(x[1985]), .Z(n13796) );
  AND U13785 ( .A(n13798), .B(n13799), .Z(n13794) );
  XNOR U13786 ( .A(y[1986]), .B(x[1986]), .Z(n13799) );
  XNOR U13787 ( .A(y[1987]), .B(x[1987]), .Z(n13798) );
  AND U13788 ( .A(n13800), .B(n13801), .Z(n13782) );
  AND U13789 ( .A(n13802), .B(n13803), .Z(n13801) );
  AND U13790 ( .A(n13804), .B(n13805), .Z(n13803) );
  XNOR U13791 ( .A(y[1990]), .B(x[1990]), .Z(n13805) );
  AND U13792 ( .A(n13806), .B(n13807), .Z(n13804) );
  XNOR U13793 ( .A(y[1988]), .B(x[1988]), .Z(n13807) );
  XNOR U13794 ( .A(y[1989]), .B(x[1989]), .Z(n13806) );
  AND U13795 ( .A(n13808), .B(n13809), .Z(n13802) );
  XNOR U13796 ( .A(y[1991]), .B(x[1991]), .Z(n13809) );
  XNOR U13797 ( .A(y[1992]), .B(x[1992]), .Z(n13808) );
  AND U13798 ( .A(n13810), .B(n13811), .Z(n13800) );
  AND U13799 ( .A(n13812), .B(n13813), .Z(n13811) );
  XNOR U13800 ( .A(y[1993]), .B(x[1993]), .Z(n13813) );
  XNOR U13801 ( .A(y[1994]), .B(x[1994]), .Z(n13812) );
  AND U13802 ( .A(n13814), .B(n13815), .Z(n13810) );
  XNOR U13803 ( .A(y[1995]), .B(x[1995]), .Z(n13815) );
  XNOR U13804 ( .A(y[1996]), .B(x[1996]), .Z(n13814) );
  AND U13805 ( .A(n13816), .B(n13817), .Z(n13742) );
  AND U13806 ( .A(n13818), .B(n13819), .Z(n13817) );
  AND U13807 ( .A(n13820), .B(n13821), .Z(n13819) );
  AND U13808 ( .A(n13822), .B(n13823), .Z(n13821) );
  AND U13809 ( .A(n13824), .B(n13825), .Z(n13823) );
  XNOR U13810 ( .A(y[1999]), .B(x[1999]), .Z(n13825) );
  AND U13811 ( .A(n13826), .B(n13827), .Z(n13824) );
  XNOR U13812 ( .A(y[1997]), .B(x[1997]), .Z(n13827) );
  XNOR U13813 ( .A(y[1998]), .B(x[1998]), .Z(n13826) );
  AND U13814 ( .A(n13828), .B(n13829), .Z(n13822) );
  XNOR U13815 ( .A(y[2000]), .B(x[2000]), .Z(n13829) );
  XNOR U13816 ( .A(y[2001]), .B(x[2001]), .Z(n13828) );
  AND U13817 ( .A(n13830), .B(n13831), .Z(n13820) );
  AND U13818 ( .A(n13832), .B(n13833), .Z(n13831) );
  XNOR U13819 ( .A(y[2004]), .B(x[2004]), .Z(n13833) );
  AND U13820 ( .A(n13834), .B(n13835), .Z(n13832) );
  XNOR U13821 ( .A(y[2002]), .B(x[2002]), .Z(n13835) );
  XNOR U13822 ( .A(y[2003]), .B(x[2003]), .Z(n13834) );
  AND U13823 ( .A(n13836), .B(n13837), .Z(n13830) );
  XNOR U13824 ( .A(y[2005]), .B(x[2005]), .Z(n13837) );
  XNOR U13825 ( .A(y[2006]), .B(x[2006]), .Z(n13836) );
  AND U13826 ( .A(n13838), .B(n13839), .Z(n13818) );
  AND U13827 ( .A(n13840), .B(n13841), .Z(n13839) );
  AND U13828 ( .A(n13842), .B(n13843), .Z(n13841) );
  XNOR U13829 ( .A(y[2009]), .B(x[2009]), .Z(n13843) );
  AND U13830 ( .A(n13844), .B(n13845), .Z(n13842) );
  XNOR U13831 ( .A(y[2007]), .B(x[2007]), .Z(n13845) );
  XNOR U13832 ( .A(y[2008]), .B(x[2008]), .Z(n13844) );
  AND U13833 ( .A(n13846), .B(n13847), .Z(n13840) );
  XNOR U13834 ( .A(y[2010]), .B(x[2010]), .Z(n13847) );
  XNOR U13835 ( .A(y[2011]), .B(x[2011]), .Z(n13846) );
  AND U13836 ( .A(n13848), .B(n13849), .Z(n13838) );
  AND U13837 ( .A(n13850), .B(n13851), .Z(n13849) );
  XNOR U13838 ( .A(y[2012]), .B(x[2012]), .Z(n13851) );
  XNOR U13839 ( .A(y[2013]), .B(x[2013]), .Z(n13850) );
  AND U13840 ( .A(n13852), .B(n13853), .Z(n13848) );
  XNOR U13841 ( .A(y[2014]), .B(x[2014]), .Z(n13853) );
  XNOR U13842 ( .A(y[2015]), .B(x[2015]), .Z(n13852) );
  AND U13843 ( .A(n13854), .B(n13855), .Z(n13816) );
  AND U13844 ( .A(n13856), .B(n13857), .Z(n13855) );
  AND U13845 ( .A(n13858), .B(n13859), .Z(n13857) );
  AND U13846 ( .A(n13860), .B(n13861), .Z(n13859) );
  XNOR U13847 ( .A(y[2018]), .B(x[2018]), .Z(n13861) );
  AND U13848 ( .A(n13862), .B(n13863), .Z(n13860) );
  XNOR U13849 ( .A(y[2016]), .B(x[2016]), .Z(n13863) );
  XNOR U13850 ( .A(y[2017]), .B(x[2017]), .Z(n13862) );
  AND U13851 ( .A(n13864), .B(n13865), .Z(n13858) );
  XNOR U13852 ( .A(y[2019]), .B(x[2019]), .Z(n13865) );
  XNOR U13853 ( .A(y[2020]), .B(x[2020]), .Z(n13864) );
  AND U13854 ( .A(n13866), .B(n13867), .Z(n13856) );
  AND U13855 ( .A(n13868), .B(n13869), .Z(n13867) );
  XNOR U13856 ( .A(y[2021]), .B(x[2021]), .Z(n13869) );
  XNOR U13857 ( .A(y[2022]), .B(x[2022]), .Z(n13868) );
  AND U13858 ( .A(n13870), .B(n13871), .Z(n13866) );
  XNOR U13859 ( .A(y[2023]), .B(x[2023]), .Z(n13871) );
  XNOR U13860 ( .A(y[2024]), .B(x[2024]), .Z(n13870) );
  AND U13861 ( .A(n13872), .B(n13873), .Z(n13854) );
  AND U13862 ( .A(n13874), .B(n13875), .Z(n13873) );
  AND U13863 ( .A(n13876), .B(n13877), .Z(n13875) );
  XNOR U13864 ( .A(y[2027]), .B(x[2027]), .Z(n13877) );
  AND U13865 ( .A(n13878), .B(n13879), .Z(n13876) );
  XNOR U13866 ( .A(y[2025]), .B(x[2025]), .Z(n13879) );
  XNOR U13867 ( .A(y[2026]), .B(x[2026]), .Z(n13878) );
  AND U13868 ( .A(n13880), .B(n13881), .Z(n13874) );
  XNOR U13869 ( .A(y[2028]), .B(x[2028]), .Z(n13881) );
  XNOR U13870 ( .A(y[2029]), .B(x[2029]), .Z(n13880) );
  AND U13871 ( .A(n13882), .B(n13883), .Z(n13872) );
  AND U13872 ( .A(n13884), .B(n13885), .Z(n13883) );
  XNOR U13873 ( .A(y[2030]), .B(x[2030]), .Z(n13885) );
  XNOR U13874 ( .A(y[2031]), .B(x[2031]), .Z(n13884) );
  AND U13875 ( .A(n13886), .B(n13887), .Z(n13882) );
  XNOR U13876 ( .A(y[2032]), .B(x[2032]), .Z(n13887) );
  XNOR U13877 ( .A(y[2033]), .B(x[2033]), .Z(n13886) );
  AND U13878 ( .A(n13888), .B(n13889), .Z(n8632) );
  AND U13879 ( .A(n13890), .B(n13891), .Z(n13889) );
  AND U13880 ( .A(n13892), .B(n13893), .Z(n13891) );
  AND U13881 ( .A(n13894), .B(n13895), .Z(n13893) );
  AND U13882 ( .A(n13896), .B(n13897), .Z(n13895) );
  AND U13883 ( .A(n13898), .B(n13899), .Z(n13897) );
  AND U13884 ( .A(n13900), .B(n13901), .Z(n13899) );
  AND U13885 ( .A(n13902), .B(n13903), .Z(n13901) );
  XNOR U13886 ( .A(y[1004]), .B(x[1004]), .Z(n13903) );
  XNOR U13887 ( .A(y[1005]), .B(x[1005]), .Z(n13902) );
  AND U13888 ( .A(n13904), .B(n13905), .Z(n13900) );
  XNOR U13889 ( .A(y[1006]), .B(x[1006]), .Z(n13905) );
  XNOR U13890 ( .A(y[1007]), .B(x[1007]), .Z(n13904) );
  AND U13891 ( .A(n13906), .B(n13907), .Z(n13898) );
  AND U13892 ( .A(n13908), .B(n13909), .Z(n13907) );
  XNOR U13893 ( .A(y[1008]), .B(x[1008]), .Z(n13909) );
  XNOR U13894 ( .A(y[1009]), .B(x[1009]), .Z(n13908) );
  AND U13895 ( .A(n13910), .B(n13911), .Z(n13906) );
  XNOR U13896 ( .A(y[1010]), .B(x[1010]), .Z(n13911) );
  XNOR U13897 ( .A(y[1011]), .B(x[1011]), .Z(n13910) );
  AND U13898 ( .A(n13912), .B(n13913), .Z(n13896) );
  AND U13899 ( .A(n13914), .B(n13915), .Z(n13913) );
  AND U13900 ( .A(n13916), .B(n13917), .Z(n13915) );
  XNOR U13901 ( .A(y[1012]), .B(x[1012]), .Z(n13917) );
  XNOR U13902 ( .A(y[1013]), .B(x[1013]), .Z(n13916) );
  AND U13903 ( .A(n13918), .B(n13919), .Z(n13914) );
  XNOR U13904 ( .A(y[1014]), .B(x[1014]), .Z(n13919) );
  XNOR U13905 ( .A(y[1015]), .B(x[1015]), .Z(n13918) );
  AND U13906 ( .A(n13920), .B(n13921), .Z(n13912) );
  AND U13907 ( .A(n13922), .B(n13923), .Z(n13921) );
  XNOR U13908 ( .A(y[1016]), .B(x[1016]), .Z(n13923) );
  XNOR U13909 ( .A(y[1017]), .B(x[1017]), .Z(n13922) );
  AND U13910 ( .A(n13924), .B(n13925), .Z(n13920) );
  XNOR U13911 ( .A(y[1018]), .B(x[1018]), .Z(n13925) );
  XNOR U13912 ( .A(y[1019]), .B(x[1019]), .Z(n13924) );
  AND U13913 ( .A(n13926), .B(n13927), .Z(n13894) );
  AND U13914 ( .A(n13928), .B(n13929), .Z(n13927) );
  AND U13915 ( .A(n13930), .B(n13931), .Z(n13929) );
  AND U13916 ( .A(n13932), .B(n13933), .Z(n13931) );
  XNOR U13917 ( .A(y[1020]), .B(x[1020]), .Z(n13933) );
  XNOR U13918 ( .A(y[1021]), .B(x[1021]), .Z(n13932) );
  AND U13919 ( .A(n13934), .B(n13935), .Z(n13930) );
  XNOR U13920 ( .A(y[1022]), .B(x[1022]), .Z(n13935) );
  XNOR U13921 ( .A(y[1023]), .B(x[1023]), .Z(n13934) );
  AND U13922 ( .A(n13936), .B(n13937), .Z(n13928) );
  AND U13923 ( .A(n13938), .B(n13939), .Z(n13937) );
  XNOR U13924 ( .A(y[1024]), .B(x[1024]), .Z(n13939) );
  XNOR U13925 ( .A(y[1025]), .B(x[1025]), .Z(n13938) );
  AND U13926 ( .A(n13940), .B(n13941), .Z(n13936) );
  XNOR U13927 ( .A(y[1026]), .B(x[1026]), .Z(n13941) );
  XNOR U13928 ( .A(y[1027]), .B(x[1027]), .Z(n13940) );
  AND U13929 ( .A(n13942), .B(n13943), .Z(n13926) );
  AND U13930 ( .A(n13944), .B(n13945), .Z(n13943) );
  AND U13931 ( .A(n13946), .B(n13947), .Z(n13945) );
  XNOR U13932 ( .A(y[1028]), .B(x[1028]), .Z(n13947) );
  XNOR U13933 ( .A(y[1029]), .B(x[1029]), .Z(n13946) );
  AND U13934 ( .A(n13948), .B(n13949), .Z(n13944) );
  XNOR U13935 ( .A(y[1030]), .B(x[1030]), .Z(n13949) );
  XNOR U13936 ( .A(y[1031]), .B(x[1031]), .Z(n13948) );
  AND U13937 ( .A(n13950), .B(n13951), .Z(n13942) );
  AND U13938 ( .A(n13952), .B(n13953), .Z(n13951) );
  XNOR U13939 ( .A(y[1032]), .B(x[1032]), .Z(n13953) );
  XNOR U13940 ( .A(y[1033]), .B(x[1033]), .Z(n13952) );
  AND U13941 ( .A(n13954), .B(n13955), .Z(n13950) );
  XNOR U13942 ( .A(y[1034]), .B(x[1034]), .Z(n13955) );
  XNOR U13943 ( .A(y[1037]), .B(x[1037]), .Z(n13954) );
  AND U13944 ( .A(n13956), .B(n13957), .Z(n13892) );
  AND U13945 ( .A(n13958), .B(n13959), .Z(n13957) );
  AND U13946 ( .A(n13960), .B(n13961), .Z(n13959) );
  AND U13947 ( .A(n13962), .B(n13963), .Z(n13961) );
  AND U13948 ( .A(n13964), .B(n13965), .Z(n13963) );
  XNOR U13949 ( .A(y[1035]), .B(x[1035]), .Z(n13965) );
  XNOR U13950 ( .A(y[1036]), .B(x[1036]), .Z(n13964) );
  AND U13951 ( .A(n13966), .B(n13967), .Z(n13962) );
  XNOR U13952 ( .A(y[1038]), .B(x[1038]), .Z(n13967) );
  XNOR U13953 ( .A(y[1039]), .B(x[1039]), .Z(n13966) );
  AND U13954 ( .A(n13968), .B(n13969), .Z(n13960) );
  AND U13955 ( .A(n13970), .B(n13971), .Z(n13969) );
  XNOR U13956 ( .A(y[1040]), .B(x[1040]), .Z(n13971) );
  XNOR U13957 ( .A(y[1041]), .B(x[1041]), .Z(n13970) );
  AND U13958 ( .A(n13972), .B(n13973), .Z(n13968) );
  XNOR U13959 ( .A(y[1042]), .B(x[1042]), .Z(n13973) );
  XNOR U13960 ( .A(y[1043]), .B(x[1043]), .Z(n13972) );
  AND U13961 ( .A(n13974), .B(n13975), .Z(n13958) );
  AND U13962 ( .A(n13976), .B(n13977), .Z(n13975) );
  AND U13963 ( .A(n13978), .B(n13979), .Z(n13977) );
  XNOR U13964 ( .A(y[1044]), .B(x[1044]), .Z(n13979) );
  XNOR U13965 ( .A(y[1045]), .B(x[1045]), .Z(n13978) );
  AND U13966 ( .A(n13980), .B(n13981), .Z(n13976) );
  XNOR U13967 ( .A(y[1046]), .B(x[1046]), .Z(n13981) );
  XNOR U13968 ( .A(y[1047]), .B(x[1047]), .Z(n13980) );
  AND U13969 ( .A(n13982), .B(n13983), .Z(n13974) );
  AND U13970 ( .A(n13984), .B(n13985), .Z(n13983) );
  XNOR U13971 ( .A(y[1048]), .B(x[1048]), .Z(n13985) );
  XNOR U13972 ( .A(y[1049]), .B(x[1049]), .Z(n13984) );
  AND U13973 ( .A(n13986), .B(n13987), .Z(n13982) );
  XNOR U13974 ( .A(y[1050]), .B(x[1050]), .Z(n13987) );
  XNOR U13975 ( .A(y[1051]), .B(x[1051]), .Z(n13986) );
  AND U13976 ( .A(n13988), .B(n13989), .Z(n13956) );
  AND U13977 ( .A(n13990), .B(n13991), .Z(n13989) );
  AND U13978 ( .A(n13992), .B(n13993), .Z(n13991) );
  AND U13979 ( .A(n13994), .B(n13995), .Z(n13993) );
  XNOR U13980 ( .A(y[1052]), .B(x[1052]), .Z(n13995) );
  XNOR U13981 ( .A(y[1053]), .B(x[1053]), .Z(n13994) );
  AND U13982 ( .A(n13996), .B(n13997), .Z(n13992) );
  XNOR U13983 ( .A(y[1054]), .B(x[1054]), .Z(n13997) );
  XNOR U13984 ( .A(y[1055]), .B(x[1055]), .Z(n13996) );
  AND U13985 ( .A(n13998), .B(n13999), .Z(n13990) );
  AND U13986 ( .A(n14000), .B(n14001), .Z(n13999) );
  XNOR U13987 ( .A(y[1056]), .B(x[1056]), .Z(n14001) );
  XNOR U13988 ( .A(y[1057]), .B(x[1057]), .Z(n14000) );
  AND U13989 ( .A(n14002), .B(n14003), .Z(n13998) );
  XNOR U13990 ( .A(y[1058]), .B(x[1058]), .Z(n14003) );
  XNOR U13991 ( .A(y[1059]), .B(x[1059]), .Z(n14002) );
  AND U13992 ( .A(n14004), .B(n14005), .Z(n13988) );
  AND U13993 ( .A(n14006), .B(n14007), .Z(n14005) );
  AND U13994 ( .A(n14008), .B(n14009), .Z(n14007) );
  XNOR U13995 ( .A(y[1060]), .B(x[1060]), .Z(n14009) );
  XNOR U13996 ( .A(y[1061]), .B(x[1061]), .Z(n14008) );
  AND U13997 ( .A(n14010), .B(n14011), .Z(n14006) );
  XNOR U13998 ( .A(y[1062]), .B(x[1062]), .Z(n14011) );
  XNOR U13999 ( .A(y[1063]), .B(x[1063]), .Z(n14010) );
  AND U14000 ( .A(n14012), .B(n14013), .Z(n14004) );
  AND U14001 ( .A(n14014), .B(n14015), .Z(n14013) );
  XNOR U14002 ( .A(y[1064]), .B(x[1064]), .Z(n14015) );
  XNOR U14003 ( .A(y[1065]), .B(x[1065]), .Z(n14014) );
  AND U14004 ( .A(n14016), .B(n14017), .Z(n14012) );
  XNOR U14005 ( .A(y[1066]), .B(x[1066]), .Z(n14017) );
  XNOR U14006 ( .A(y[1067]), .B(x[1067]), .Z(n14016) );
  AND U14007 ( .A(n14018), .B(n14019), .Z(n13890) );
  AND U14008 ( .A(n14020), .B(n14021), .Z(n14019) );
  AND U14009 ( .A(n14022), .B(n14023), .Z(n14021) );
  AND U14010 ( .A(n14024), .B(n14025), .Z(n14023) );
  AND U14011 ( .A(n14026), .B(n14027), .Z(n14025) );
  AND U14012 ( .A(n14028), .B(n14029), .Z(n14027) );
  XNOR U14013 ( .A(y[1068]), .B(x[1068]), .Z(n14029) );
  XNOR U14014 ( .A(y[1069]), .B(x[1069]), .Z(n14028) );
  AND U14015 ( .A(n14030), .B(n14031), .Z(n14026) );
  XNOR U14016 ( .A(y[1070]), .B(x[1070]), .Z(n14031) );
  XNOR U14017 ( .A(y[1071]), .B(x[1071]), .Z(n14030) );
  AND U14018 ( .A(n14032), .B(n14033), .Z(n14024) );
  AND U14019 ( .A(n14034), .B(n14035), .Z(n14033) );
  XNOR U14020 ( .A(y[1072]), .B(x[1072]), .Z(n14035) );
  XNOR U14021 ( .A(y[1073]), .B(x[1073]), .Z(n14034) );
  AND U14022 ( .A(n14036), .B(n14037), .Z(n14032) );
  XNOR U14023 ( .A(y[1074]), .B(x[1074]), .Z(n14037) );
  XNOR U14024 ( .A(y[1075]), .B(x[1075]), .Z(n14036) );
  AND U14025 ( .A(n14038), .B(n14039), .Z(n14022) );
  AND U14026 ( .A(n14040), .B(n14041), .Z(n14039) );
  AND U14027 ( .A(n14042), .B(n14043), .Z(n14041) );
  XNOR U14028 ( .A(y[1076]), .B(x[1076]), .Z(n14043) );
  XNOR U14029 ( .A(y[1077]), .B(x[1077]), .Z(n14042) );
  AND U14030 ( .A(n14044), .B(n14045), .Z(n14040) );
  XNOR U14031 ( .A(y[1078]), .B(x[1078]), .Z(n14045) );
  XNOR U14032 ( .A(y[1079]), .B(x[1079]), .Z(n14044) );
  AND U14033 ( .A(n14046), .B(n14047), .Z(n14038) );
  AND U14034 ( .A(n14048), .B(n14049), .Z(n14047) );
  XNOR U14035 ( .A(y[1080]), .B(x[1080]), .Z(n14049) );
  XNOR U14036 ( .A(y[1081]), .B(x[1081]), .Z(n14048) );
  AND U14037 ( .A(n14050), .B(n14051), .Z(n14046) );
  XNOR U14038 ( .A(y[1082]), .B(x[1082]), .Z(n14051) );
  XNOR U14039 ( .A(y[1083]), .B(x[1083]), .Z(n14050) );
  AND U14040 ( .A(n14052), .B(n14053), .Z(n14020) );
  AND U14041 ( .A(n14054), .B(n14055), .Z(n14053) );
  AND U14042 ( .A(n14056), .B(n14057), .Z(n14055) );
  AND U14043 ( .A(n14058), .B(n14059), .Z(n14057) );
  XNOR U14044 ( .A(y[1084]), .B(x[1084]), .Z(n14059) );
  XNOR U14045 ( .A(y[1085]), .B(x[1085]), .Z(n14058) );
  AND U14046 ( .A(n14060), .B(n14061), .Z(n14056) );
  XNOR U14047 ( .A(y[1086]), .B(x[1086]), .Z(n14061) );
  XNOR U14048 ( .A(y[1087]), .B(x[1087]), .Z(n14060) );
  AND U14049 ( .A(n14062), .B(n14063), .Z(n14054) );
  AND U14050 ( .A(n14064), .B(n14065), .Z(n14063) );
  XNOR U14051 ( .A(y[1088]), .B(x[1088]), .Z(n14065) );
  XNOR U14052 ( .A(y[1089]), .B(x[1089]), .Z(n14064) );
  AND U14053 ( .A(n14066), .B(n14067), .Z(n14062) );
  XNOR U14054 ( .A(y[1090]), .B(x[1090]), .Z(n14067) );
  XNOR U14055 ( .A(y[1091]), .B(x[1091]), .Z(n14066) );
  AND U14056 ( .A(n14068), .B(n14069), .Z(n14052) );
  AND U14057 ( .A(n14070), .B(n14071), .Z(n14069) );
  AND U14058 ( .A(n14072), .B(n14073), .Z(n14071) );
  XNOR U14059 ( .A(y[1092]), .B(x[1092]), .Z(n14073) );
  XNOR U14060 ( .A(y[1093]), .B(x[1093]), .Z(n14072) );
  AND U14061 ( .A(n14074), .B(n14075), .Z(n14070) );
  XNOR U14062 ( .A(y[1094]), .B(x[1094]), .Z(n14075) );
  XNOR U14063 ( .A(y[1095]), .B(x[1095]), .Z(n14074) );
  AND U14064 ( .A(n14076), .B(n14077), .Z(n14068) );
  AND U14065 ( .A(n14078), .B(n14079), .Z(n14077) );
  XNOR U14066 ( .A(y[1096]), .B(x[1096]), .Z(n14079) );
  XNOR U14067 ( .A(y[1097]), .B(x[1097]), .Z(n14078) );
  AND U14068 ( .A(n14080), .B(n14081), .Z(n14076) );
  XNOR U14069 ( .A(y[1098]), .B(x[1098]), .Z(n14081) );
  XNOR U14070 ( .A(y[1099]), .B(x[1099]), .Z(n14080) );
  AND U14071 ( .A(n14082), .B(n14083), .Z(n14018) );
  AND U14072 ( .A(n14084), .B(n14085), .Z(n14083) );
  AND U14073 ( .A(n14086), .B(n14087), .Z(n14085) );
  AND U14074 ( .A(n14088), .B(n14089), .Z(n14087) );
  AND U14075 ( .A(n14090), .B(n14091), .Z(n14089) );
  XNOR U14076 ( .A(y[1100]), .B(x[1100]), .Z(n14091) );
  XNOR U14077 ( .A(y[1101]), .B(x[1101]), .Z(n14090) );
  AND U14078 ( .A(n14092), .B(n14093), .Z(n14088) );
  XNOR U14079 ( .A(y[1102]), .B(x[1102]), .Z(n14093) );
  XNOR U14080 ( .A(y[1103]), .B(x[1103]), .Z(n14092) );
  AND U14081 ( .A(n14094), .B(n14095), .Z(n14086) );
  AND U14082 ( .A(n14096), .B(n14097), .Z(n14095) );
  XNOR U14083 ( .A(y[1104]), .B(x[1104]), .Z(n14097) );
  XNOR U14084 ( .A(y[1105]), .B(x[1105]), .Z(n14096) );
  AND U14085 ( .A(n14098), .B(n14099), .Z(n14094) );
  XNOR U14086 ( .A(y[1106]), .B(x[1106]), .Z(n14099) );
  XNOR U14087 ( .A(y[1107]), .B(x[1107]), .Z(n14098) );
  AND U14088 ( .A(n14100), .B(n14101), .Z(n14084) );
  AND U14089 ( .A(n14102), .B(n14103), .Z(n14101) );
  AND U14090 ( .A(n14104), .B(n14105), .Z(n14103) );
  XNOR U14091 ( .A(y[1108]), .B(x[1108]), .Z(n14105) );
  XNOR U14092 ( .A(y[1109]), .B(x[1109]), .Z(n14104) );
  AND U14093 ( .A(n14106), .B(n14107), .Z(n14102) );
  XNOR U14094 ( .A(y[1110]), .B(x[1110]), .Z(n14107) );
  XNOR U14095 ( .A(y[1111]), .B(x[1111]), .Z(n14106) );
  AND U14096 ( .A(n14108), .B(n14109), .Z(n14100) );
  AND U14097 ( .A(n14110), .B(n14111), .Z(n14109) );
  XNOR U14098 ( .A(y[1112]), .B(x[1112]), .Z(n14111) );
  XNOR U14099 ( .A(y[1113]), .B(x[1113]), .Z(n14110) );
  AND U14100 ( .A(n14112), .B(n14113), .Z(n14108) );
  XNOR U14101 ( .A(y[1114]), .B(x[1114]), .Z(n14113) );
  XNOR U14102 ( .A(y[1115]), .B(x[1115]), .Z(n14112) );
  AND U14103 ( .A(n14114), .B(n14115), .Z(n14082) );
  AND U14104 ( .A(n14116), .B(n14117), .Z(n14115) );
  AND U14105 ( .A(n14118), .B(n14119), .Z(n14117) );
  AND U14106 ( .A(n14120), .B(n14121), .Z(n14119) );
  XNOR U14107 ( .A(y[1116]), .B(x[1116]), .Z(n14121) );
  XNOR U14108 ( .A(y[1117]), .B(x[1117]), .Z(n14120) );
  AND U14109 ( .A(n14122), .B(n14123), .Z(n14118) );
  XNOR U14110 ( .A(y[1118]), .B(x[1118]), .Z(n14123) );
  XNOR U14111 ( .A(y[1119]), .B(x[1119]), .Z(n14122) );
  AND U14112 ( .A(n14124), .B(n14125), .Z(n14116) );
  AND U14113 ( .A(n14126), .B(n14127), .Z(n14125) );
  XNOR U14114 ( .A(y[1120]), .B(x[1120]), .Z(n14127) );
  XNOR U14115 ( .A(y[1121]), .B(x[1121]), .Z(n14126) );
  AND U14116 ( .A(n14128), .B(n14129), .Z(n14124) );
  XNOR U14117 ( .A(y[1122]), .B(x[1122]), .Z(n14129) );
  XNOR U14118 ( .A(y[1123]), .B(x[1123]), .Z(n14128) );
  AND U14119 ( .A(n14130), .B(n14131), .Z(n14114) );
  AND U14120 ( .A(n14132), .B(n14133), .Z(n14131) );
  AND U14121 ( .A(n14134), .B(n14135), .Z(n14133) );
  XNOR U14122 ( .A(y[1124]), .B(x[1124]), .Z(n14135) );
  XNOR U14123 ( .A(y[1125]), .B(x[1125]), .Z(n14134) );
  AND U14124 ( .A(n14136), .B(n14137), .Z(n14132) );
  XNOR U14125 ( .A(y[1126]), .B(x[1126]), .Z(n14137) );
  XNOR U14126 ( .A(y[1127]), .B(x[1127]), .Z(n14136) );
  AND U14127 ( .A(n14138), .B(n14139), .Z(n14130) );
  AND U14128 ( .A(n14140), .B(n14141), .Z(n14139) );
  XNOR U14129 ( .A(y[1128]), .B(x[1128]), .Z(n14141) );
  XNOR U14130 ( .A(y[1129]), .B(x[1129]), .Z(n14140) );
  AND U14131 ( .A(n14142), .B(n14143), .Z(n14138) );
  XNOR U14132 ( .A(y[1130]), .B(x[1130]), .Z(n14143) );
  XNOR U14133 ( .A(y[1131]), .B(x[1131]), .Z(n14142) );
  AND U14134 ( .A(n14144), .B(n14145), .Z(n13888) );
  AND U14135 ( .A(n14146), .B(n14147), .Z(n14145) );
  AND U14136 ( .A(n14148), .B(n14149), .Z(n14147) );
  AND U14137 ( .A(n14150), .B(n14151), .Z(n14149) );
  AND U14138 ( .A(n14152), .B(n14153), .Z(n14151) );
  AND U14139 ( .A(n14154), .B(n14155), .Z(n14153) );
  AND U14140 ( .A(n14156), .B(n14157), .Z(n14155) );
  XNOR U14141 ( .A(y[1132]), .B(x[1132]), .Z(n14157) );
  XNOR U14142 ( .A(y[1133]), .B(x[1133]), .Z(n14156) );
  AND U14143 ( .A(n14158), .B(n14159), .Z(n14154) );
  XNOR U14144 ( .A(y[1134]), .B(x[1134]), .Z(n14159) );
  XNOR U14145 ( .A(y[1135]), .B(x[1135]), .Z(n14158) );
  AND U14146 ( .A(n14160), .B(n14161), .Z(n14152) );
  AND U14147 ( .A(n14162), .B(n14163), .Z(n14161) );
  XNOR U14148 ( .A(y[1136]), .B(x[1136]), .Z(n14163) );
  XNOR U14149 ( .A(y[1137]), .B(x[1137]), .Z(n14162) );
  AND U14150 ( .A(n14164), .B(n14165), .Z(n14160) );
  XNOR U14151 ( .A(y[1138]), .B(x[1138]), .Z(n14165) );
  XNOR U14152 ( .A(y[1139]), .B(x[1139]), .Z(n14164) );
  AND U14153 ( .A(n14166), .B(n14167), .Z(n14150) );
  AND U14154 ( .A(n14168), .B(n14169), .Z(n14167) );
  AND U14155 ( .A(n14170), .B(n14171), .Z(n14169) );
  XNOR U14156 ( .A(y[1140]), .B(x[1140]), .Z(n14171) );
  XNOR U14157 ( .A(y[1141]), .B(x[1141]), .Z(n14170) );
  AND U14158 ( .A(n14172), .B(n14173), .Z(n14168) );
  XNOR U14159 ( .A(y[1142]), .B(x[1142]), .Z(n14173) );
  XNOR U14160 ( .A(y[1143]), .B(x[1143]), .Z(n14172) );
  AND U14161 ( .A(n14174), .B(n14175), .Z(n14166) );
  AND U14162 ( .A(n14176), .B(n14177), .Z(n14175) );
  XNOR U14163 ( .A(y[1144]), .B(x[1144]), .Z(n14177) );
  XNOR U14164 ( .A(y[1145]), .B(x[1145]), .Z(n14176) );
  AND U14165 ( .A(n14178), .B(n14179), .Z(n14174) );
  XNOR U14166 ( .A(y[1146]), .B(x[1146]), .Z(n14179) );
  XNOR U14167 ( .A(y[1147]), .B(x[1147]), .Z(n14178) );
  AND U14168 ( .A(n14180), .B(n14181), .Z(n14148) );
  AND U14169 ( .A(n14182), .B(n14183), .Z(n14181) );
  AND U14170 ( .A(n14184), .B(n14185), .Z(n14183) );
  AND U14171 ( .A(n14186), .B(n14187), .Z(n14185) );
  XNOR U14172 ( .A(y[1148]), .B(x[1148]), .Z(n14187) );
  XNOR U14173 ( .A(y[1149]), .B(x[1149]), .Z(n14186) );
  AND U14174 ( .A(n14188), .B(n14189), .Z(n14184) );
  XNOR U14175 ( .A(y[1150]), .B(x[1150]), .Z(n14189) );
  XNOR U14176 ( .A(y[1151]), .B(x[1151]), .Z(n14188) );
  AND U14177 ( .A(n14190), .B(n14191), .Z(n14182) );
  AND U14178 ( .A(n14192), .B(n14193), .Z(n14191) );
  XNOR U14179 ( .A(y[1152]), .B(x[1152]), .Z(n14193) );
  XNOR U14180 ( .A(y[1153]), .B(x[1153]), .Z(n14192) );
  AND U14181 ( .A(n14194), .B(n14195), .Z(n14190) );
  XNOR U14182 ( .A(y[1154]), .B(x[1154]), .Z(n14195) );
  XNOR U14183 ( .A(y[1155]), .B(x[1155]), .Z(n14194) );
  AND U14184 ( .A(n14196), .B(n14197), .Z(n14180) );
  AND U14185 ( .A(n14198), .B(n14199), .Z(n14197) );
  AND U14186 ( .A(n14200), .B(n14201), .Z(n14199) );
  XNOR U14187 ( .A(y[1156]), .B(x[1156]), .Z(n14201) );
  XNOR U14188 ( .A(y[1157]), .B(x[1157]), .Z(n14200) );
  AND U14189 ( .A(n14202), .B(n14203), .Z(n14198) );
  XNOR U14190 ( .A(y[1158]), .B(x[1158]), .Z(n14203) );
  XNOR U14191 ( .A(y[1159]), .B(x[1159]), .Z(n14202) );
  AND U14192 ( .A(n14204), .B(n14205), .Z(n14196) );
  AND U14193 ( .A(n14206), .B(n14207), .Z(n14205) );
  XNOR U14194 ( .A(y[1160]), .B(x[1160]), .Z(n14207) );
  XNOR U14195 ( .A(y[1161]), .B(x[1161]), .Z(n14206) );
  AND U14196 ( .A(n14208), .B(n14209), .Z(n14204) );
  XNOR U14197 ( .A(y[1162]), .B(x[1162]), .Z(n14209) );
  XNOR U14198 ( .A(y[1163]), .B(x[1163]), .Z(n14208) );
  AND U14199 ( .A(n14210), .B(n14211), .Z(n14146) );
  AND U14200 ( .A(n14212), .B(n14213), .Z(n14211) );
  AND U14201 ( .A(n14214), .B(n14215), .Z(n14213) );
  AND U14202 ( .A(n14216), .B(n14217), .Z(n14215) );
  AND U14203 ( .A(n14218), .B(n14219), .Z(n14217) );
  XNOR U14204 ( .A(y[1164]), .B(x[1164]), .Z(n14219) );
  XNOR U14205 ( .A(y[1165]), .B(x[1165]), .Z(n14218) );
  AND U14206 ( .A(n14220), .B(n14221), .Z(n14216) );
  XNOR U14207 ( .A(y[1166]), .B(x[1166]), .Z(n14221) );
  XNOR U14208 ( .A(y[1167]), .B(x[1167]), .Z(n14220) );
  AND U14209 ( .A(n14222), .B(n14223), .Z(n14214) );
  AND U14210 ( .A(n14224), .B(n14225), .Z(n14223) );
  XNOR U14211 ( .A(y[1168]), .B(x[1168]), .Z(n14225) );
  XNOR U14212 ( .A(y[1169]), .B(x[1169]), .Z(n14224) );
  AND U14213 ( .A(n14226), .B(n14227), .Z(n14222) );
  XNOR U14214 ( .A(y[1170]), .B(x[1170]), .Z(n14227) );
  XNOR U14215 ( .A(y[1171]), .B(x[1171]), .Z(n14226) );
  AND U14216 ( .A(n14228), .B(n14229), .Z(n14212) );
  AND U14217 ( .A(n14230), .B(n14231), .Z(n14229) );
  AND U14218 ( .A(n14232), .B(n14233), .Z(n14231) );
  XNOR U14219 ( .A(y[1172]), .B(x[1172]), .Z(n14233) );
  XNOR U14220 ( .A(y[1173]), .B(x[1173]), .Z(n14232) );
  AND U14221 ( .A(n14234), .B(n14235), .Z(n14230) );
  XNOR U14222 ( .A(y[1174]), .B(x[1174]), .Z(n14235) );
  XNOR U14223 ( .A(y[1175]), .B(x[1175]), .Z(n14234) );
  AND U14224 ( .A(n14236), .B(n14237), .Z(n14228) );
  AND U14225 ( .A(n14238), .B(n14239), .Z(n14237) );
  XNOR U14226 ( .A(y[1176]), .B(x[1176]), .Z(n14239) );
  XNOR U14227 ( .A(y[1177]), .B(x[1177]), .Z(n14238) );
  AND U14228 ( .A(n14240), .B(n14241), .Z(n14236) );
  XNOR U14229 ( .A(y[1178]), .B(x[1178]), .Z(n14241) );
  XNOR U14230 ( .A(y[1179]), .B(x[1179]), .Z(n14240) );
  AND U14231 ( .A(n14242), .B(n14243), .Z(n14210) );
  AND U14232 ( .A(n14244), .B(n14245), .Z(n14243) );
  AND U14233 ( .A(n14246), .B(n14247), .Z(n14245) );
  AND U14234 ( .A(n14248), .B(n14249), .Z(n14247) );
  XNOR U14235 ( .A(y[1180]), .B(x[1180]), .Z(n14249) );
  XNOR U14236 ( .A(y[1181]), .B(x[1181]), .Z(n14248) );
  AND U14237 ( .A(n14250), .B(n14251), .Z(n14246) );
  XNOR U14238 ( .A(y[1182]), .B(x[1182]), .Z(n14251) );
  XNOR U14239 ( .A(y[1183]), .B(x[1183]), .Z(n14250) );
  AND U14240 ( .A(n14252), .B(n14253), .Z(n14244) );
  AND U14241 ( .A(n14254), .B(n14255), .Z(n14253) );
  XNOR U14242 ( .A(y[1184]), .B(x[1184]), .Z(n14255) );
  XNOR U14243 ( .A(y[1185]), .B(x[1185]), .Z(n14254) );
  AND U14244 ( .A(n14256), .B(n14257), .Z(n14252) );
  XNOR U14245 ( .A(y[1186]), .B(x[1186]), .Z(n14257) );
  XNOR U14246 ( .A(y[1187]), .B(x[1187]), .Z(n14256) );
  AND U14247 ( .A(n14258), .B(n14259), .Z(n14242) );
  AND U14248 ( .A(n14260), .B(n14261), .Z(n14259) );
  AND U14249 ( .A(n14262), .B(n14263), .Z(n14261) );
  XNOR U14250 ( .A(y[1188]), .B(x[1188]), .Z(n14263) );
  XNOR U14251 ( .A(y[1189]), .B(x[1189]), .Z(n14262) );
  AND U14252 ( .A(n14264), .B(n14265), .Z(n14260) );
  XNOR U14253 ( .A(y[1190]), .B(x[1190]), .Z(n14265) );
  XNOR U14254 ( .A(y[1191]), .B(x[1191]), .Z(n14264) );
  AND U14255 ( .A(n14266), .B(n14267), .Z(n14258) );
  AND U14256 ( .A(n14268), .B(n14269), .Z(n14267) );
  XNOR U14257 ( .A(y[1192]), .B(x[1192]), .Z(n14269) );
  XNOR U14258 ( .A(y[1193]), .B(x[1193]), .Z(n14268) );
  AND U14259 ( .A(n14270), .B(n14271), .Z(n14266) );
  XNOR U14260 ( .A(y[1194]), .B(x[1194]), .Z(n14271) );
  XNOR U14261 ( .A(y[1195]), .B(x[1195]), .Z(n14270) );
  AND U14262 ( .A(n14272), .B(n14273), .Z(n14144) );
  AND U14263 ( .A(n14274), .B(n14275), .Z(n14273) );
  AND U14264 ( .A(n14276), .B(n14277), .Z(n14275) );
  AND U14265 ( .A(n14278), .B(n14279), .Z(n14277) );
  AND U14266 ( .A(n14280), .B(n14281), .Z(n14279) );
  AND U14267 ( .A(n14282), .B(n14283), .Z(n14281) );
  XNOR U14268 ( .A(y[1196]), .B(x[1196]), .Z(n14283) );
  XNOR U14269 ( .A(y[1197]), .B(x[1197]), .Z(n14282) );
  AND U14270 ( .A(n14284), .B(n14285), .Z(n14280) );
  XNOR U14271 ( .A(y[1198]), .B(x[1198]), .Z(n14285) );
  XNOR U14272 ( .A(y[1199]), .B(x[1199]), .Z(n14284) );
  AND U14273 ( .A(n14286), .B(n14287), .Z(n14278) );
  AND U14274 ( .A(n14288), .B(n14289), .Z(n14287) );
  XNOR U14275 ( .A(y[1200]), .B(x[1200]), .Z(n14289) );
  XNOR U14276 ( .A(y[1201]), .B(x[1201]), .Z(n14288) );
  AND U14277 ( .A(n14290), .B(n14291), .Z(n14286) );
  XNOR U14278 ( .A(y[1202]), .B(x[1202]), .Z(n14291) );
  XNOR U14279 ( .A(y[1203]), .B(x[1203]), .Z(n14290) );
  AND U14280 ( .A(n14292), .B(n14293), .Z(n14276) );
  AND U14281 ( .A(n14294), .B(n14295), .Z(n14293) );
  AND U14282 ( .A(n14296), .B(n14297), .Z(n14295) );
  XNOR U14283 ( .A(y[1204]), .B(x[1204]), .Z(n14297) );
  XNOR U14284 ( .A(y[1205]), .B(x[1205]), .Z(n14296) );
  AND U14285 ( .A(n14298), .B(n14299), .Z(n14294) );
  XNOR U14286 ( .A(y[1206]), .B(x[1206]), .Z(n14299) );
  XNOR U14287 ( .A(y[1207]), .B(x[1207]), .Z(n14298) );
  AND U14288 ( .A(n14300), .B(n14301), .Z(n14292) );
  AND U14289 ( .A(n14302), .B(n14303), .Z(n14301) );
  XNOR U14290 ( .A(y[1208]), .B(x[1208]), .Z(n14303) );
  XNOR U14291 ( .A(y[1209]), .B(x[1209]), .Z(n14302) );
  AND U14292 ( .A(n14304), .B(n14305), .Z(n14300) );
  XNOR U14293 ( .A(y[1210]), .B(x[1210]), .Z(n14305) );
  XNOR U14294 ( .A(y[1211]), .B(x[1211]), .Z(n14304) );
  AND U14295 ( .A(n14306), .B(n14307), .Z(n14274) );
  AND U14296 ( .A(n14308), .B(n14309), .Z(n14307) );
  AND U14297 ( .A(n14310), .B(n14311), .Z(n14309) );
  AND U14298 ( .A(n14312), .B(n14313), .Z(n14311) );
  XNOR U14299 ( .A(y[1212]), .B(x[1212]), .Z(n14313) );
  XNOR U14300 ( .A(y[1213]), .B(x[1213]), .Z(n14312) );
  AND U14301 ( .A(n14314), .B(n14315), .Z(n14310) );
  XNOR U14302 ( .A(y[1214]), .B(x[1214]), .Z(n14315) );
  XNOR U14303 ( .A(y[1215]), .B(x[1215]), .Z(n14314) );
  AND U14304 ( .A(n14316), .B(n14317), .Z(n14308) );
  AND U14305 ( .A(n14318), .B(n14319), .Z(n14317) );
  XNOR U14306 ( .A(y[1216]), .B(x[1216]), .Z(n14319) );
  XNOR U14307 ( .A(y[1217]), .B(x[1217]), .Z(n14318) );
  AND U14308 ( .A(n14320), .B(n14321), .Z(n14316) );
  XNOR U14309 ( .A(y[1218]), .B(x[1218]), .Z(n14321) );
  XNOR U14310 ( .A(y[1219]), .B(x[1219]), .Z(n14320) );
  AND U14311 ( .A(n14322), .B(n14323), .Z(n14306) );
  AND U14312 ( .A(n14324), .B(n14325), .Z(n14323) );
  AND U14313 ( .A(n14326), .B(n14327), .Z(n14325) );
  XNOR U14314 ( .A(y[1220]), .B(x[1220]), .Z(n14327) );
  XNOR U14315 ( .A(y[1221]), .B(x[1221]), .Z(n14326) );
  AND U14316 ( .A(n14328), .B(n14329), .Z(n14324) );
  XNOR U14317 ( .A(y[1222]), .B(x[1222]), .Z(n14329) );
  XNOR U14318 ( .A(y[1223]), .B(x[1223]), .Z(n14328) );
  AND U14319 ( .A(n14330), .B(n14331), .Z(n14322) );
  AND U14320 ( .A(n14332), .B(n14333), .Z(n14331) );
  XNOR U14321 ( .A(y[1224]), .B(x[1224]), .Z(n14333) );
  XNOR U14322 ( .A(y[1225]), .B(x[1225]), .Z(n14332) );
  AND U14323 ( .A(n14334), .B(n14335), .Z(n14330) );
  XNOR U14324 ( .A(y[1226]), .B(x[1226]), .Z(n14335) );
  XNOR U14325 ( .A(y[1227]), .B(x[1227]), .Z(n14334) );
  AND U14326 ( .A(n14336), .B(n14337), .Z(n14272) );
  AND U14327 ( .A(n14338), .B(n14339), .Z(n14337) );
  AND U14328 ( .A(n14340), .B(n14341), .Z(n14339) );
  AND U14329 ( .A(n14342), .B(n14343), .Z(n14341) );
  AND U14330 ( .A(n14344), .B(n14345), .Z(n14343) );
  XNOR U14331 ( .A(y[1228]), .B(x[1228]), .Z(n14345) );
  XNOR U14332 ( .A(y[1229]), .B(x[1229]), .Z(n14344) );
  AND U14333 ( .A(n14346), .B(n14347), .Z(n14342) );
  XNOR U14334 ( .A(y[1230]), .B(x[1230]), .Z(n14347) );
  XNOR U14335 ( .A(y[1231]), .B(x[1231]), .Z(n14346) );
  AND U14336 ( .A(n14348), .B(n14349), .Z(n14340) );
  AND U14337 ( .A(n14350), .B(n14351), .Z(n14349) );
  XNOR U14338 ( .A(y[1232]), .B(x[1232]), .Z(n14351) );
  XNOR U14339 ( .A(y[1233]), .B(x[1233]), .Z(n14350) );
  AND U14340 ( .A(n14352), .B(n14353), .Z(n14348) );
  XNOR U14341 ( .A(y[1234]), .B(x[1234]), .Z(n14353) );
  XNOR U14342 ( .A(y[1235]), .B(x[1235]), .Z(n14352) );
  AND U14343 ( .A(n14354), .B(n14355), .Z(n14338) );
  AND U14344 ( .A(n14356), .B(n14357), .Z(n14355) );
  AND U14345 ( .A(n14358), .B(n14359), .Z(n14357) );
  XNOR U14346 ( .A(y[1236]), .B(x[1236]), .Z(n14359) );
  XNOR U14347 ( .A(y[1237]), .B(x[1237]), .Z(n14358) );
  AND U14348 ( .A(n14360), .B(n14361), .Z(n14356) );
  XNOR U14349 ( .A(y[1238]), .B(x[1238]), .Z(n14361) );
  XNOR U14350 ( .A(y[1239]), .B(x[1239]), .Z(n14360) );
  AND U14351 ( .A(n14362), .B(n14363), .Z(n14354) );
  AND U14352 ( .A(n14364), .B(n14365), .Z(n14363) );
  XNOR U14353 ( .A(y[1240]), .B(x[1240]), .Z(n14365) );
  XNOR U14354 ( .A(y[1241]), .B(x[1241]), .Z(n14364) );
  AND U14355 ( .A(n14366), .B(n14367), .Z(n14362) );
  XNOR U14356 ( .A(y[1242]), .B(x[1242]), .Z(n14367) );
  XNOR U14357 ( .A(y[1243]), .B(x[1243]), .Z(n14366) );
  AND U14358 ( .A(n14368), .B(n14369), .Z(n14336) );
  AND U14359 ( .A(n14370), .B(n14371), .Z(n14369) );
  AND U14360 ( .A(n14372), .B(n14373), .Z(n14371) );
  AND U14361 ( .A(n14374), .B(n14375), .Z(n14373) );
  XNOR U14362 ( .A(y[1244]), .B(x[1244]), .Z(n14375) );
  XNOR U14363 ( .A(y[1245]), .B(x[1245]), .Z(n14374) );
  AND U14364 ( .A(n14376), .B(n14377), .Z(n14372) );
  XNOR U14365 ( .A(y[1246]), .B(x[1246]), .Z(n14377) );
  XNOR U14366 ( .A(y[1247]), .B(x[1247]), .Z(n14376) );
  AND U14367 ( .A(n14378), .B(n14379), .Z(n14370) );
  AND U14368 ( .A(n14380), .B(n14381), .Z(n14379) );
  XNOR U14369 ( .A(y[1248]), .B(x[1248]), .Z(n14381) );
  XNOR U14370 ( .A(y[1249]), .B(x[1249]), .Z(n14380) );
  AND U14371 ( .A(n14382), .B(n14383), .Z(n14378) );
  XNOR U14372 ( .A(y[1250]), .B(x[1250]), .Z(n14383) );
  XNOR U14373 ( .A(y[1251]), .B(x[1251]), .Z(n14382) );
  AND U14374 ( .A(n14384), .B(n14385), .Z(n14368) );
  AND U14375 ( .A(n14386), .B(n14387), .Z(n14385) );
  AND U14376 ( .A(n14388), .B(n14389), .Z(n14387) );
  XNOR U14377 ( .A(y[1252]), .B(x[1252]), .Z(n14389) );
  XNOR U14378 ( .A(y[1253]), .B(x[1253]), .Z(n14388) );
  AND U14379 ( .A(n14390), .B(n14391), .Z(n14386) );
  XNOR U14380 ( .A(y[1254]), .B(x[1254]), .Z(n14391) );
  XNOR U14381 ( .A(y[1255]), .B(x[1255]), .Z(n14390) );
  AND U14382 ( .A(n14392), .B(n14393), .Z(n14384) );
  AND U14383 ( .A(n14394), .B(n14395), .Z(n14393) );
  XNOR U14384 ( .A(y[1256]), .B(x[1256]), .Z(n14395) );
  XNOR U14385 ( .A(y[1257]), .B(x[1257]), .Z(n14394) );
  AND U14386 ( .A(n14396), .B(n14397), .Z(n14392) );
  XNOR U14387 ( .A(y[1258]), .B(x[1258]), .Z(n14397) );
  XNOR U14388 ( .A(y[1259]), .B(x[1259]), .Z(n14396) );
  AND U14389 ( .A(n14398), .B(n14399), .Z(n8628) );
  XNOR U14390 ( .A(y[945]), .B(x[945]), .Z(n14399) );
  AND U14391 ( .A(n14400), .B(n14401), .Z(n14398) );
  XNOR U14392 ( .A(y[943]), .B(x[943]), .Z(n14401) );
  XNOR U14393 ( .A(y[944]), .B(x[944]), .Z(n14400) );
  AND U14394 ( .A(n14402), .B(n14403), .Z(n8626) );
  AND U14395 ( .A(n14404), .B(n14405), .Z(n14403) );
  XNOR U14396 ( .A(y[948]), .B(x[948]), .Z(n14405) );
  AND U14397 ( .A(n14406), .B(n14407), .Z(n14404) );
  XNOR U14398 ( .A(y[946]), .B(x[946]), .Z(n14407) );
  XNOR U14399 ( .A(y[947]), .B(x[947]), .Z(n14406) );
  AND U14400 ( .A(n14408), .B(n14409), .Z(n14402) );
  XNOR U14401 ( .A(y[949]), .B(x[949]), .Z(n14409) );
  XNOR U14402 ( .A(y[950]), .B(x[950]), .Z(n14408) );
  AND U14403 ( .A(n14410), .B(n14411), .Z(n8624) );
  AND U14404 ( .A(n14412), .B(n14413), .Z(n14411) );
  AND U14405 ( .A(n14414), .B(n14415), .Z(n14413) );
  XNOR U14406 ( .A(y[953]), .B(x[953]), .Z(n14415) );
  AND U14407 ( .A(n14416), .B(n14417), .Z(n14414) );
  XNOR U14408 ( .A(y[951]), .B(x[951]), .Z(n14417) );
  XNOR U14409 ( .A(y[952]), .B(x[952]), .Z(n14416) );
  AND U14410 ( .A(n14418), .B(n14419), .Z(n14412) );
  XNOR U14411 ( .A(y[954]), .B(x[954]), .Z(n14419) );
  XNOR U14412 ( .A(y[955]), .B(x[955]), .Z(n14418) );
  AND U14413 ( .A(n14420), .B(n14421), .Z(n14410) );
  AND U14414 ( .A(n14422), .B(n14423), .Z(n14421) );
  XNOR U14415 ( .A(y[398]), .B(x[398]), .Z(n14423) );
  AND U14416 ( .A(n14424), .B(n14425), .Z(n14422) );
  XNOR U14417 ( .A(y[956]), .B(x[956]), .Z(n14425) );
  XNOR U14418 ( .A(y[957]), .B(x[957]), .Z(n14424) );
  AND U14419 ( .A(n14426), .B(n14427), .Z(n14420) );
  XNOR U14420 ( .A(y[399]), .B(x[399]), .Z(n14427) );
  XNOR U14421 ( .A(y[400]), .B(x[400]), .Z(n14426) );
  AND U14422 ( .A(n14428), .B(n14429), .Z(n8622) );
  AND U14423 ( .A(n14430), .B(n14431), .Z(n14429) );
  AND U14424 ( .A(n14432), .B(n14433), .Z(n14431) );
  AND U14425 ( .A(n14434), .B(n14435), .Z(n14433) );
  XNOR U14426 ( .A(y[403]), .B(x[403]), .Z(n14435) );
  AND U14427 ( .A(n14436), .B(n14437), .Z(n14434) );
  XNOR U14428 ( .A(y[401]), .B(x[401]), .Z(n14437) );
  XNOR U14429 ( .A(y[402]), .B(x[402]), .Z(n14436) );
  AND U14430 ( .A(n14438), .B(n14439), .Z(n14432) );
  XNOR U14431 ( .A(y[406]), .B(x[406]), .Z(n14439) );
  AND U14432 ( .A(n14440), .B(n14441), .Z(n14438) );
  XNOR U14433 ( .A(y[404]), .B(x[404]), .Z(n14441) );
  XNOR U14434 ( .A(y[405]), .B(x[405]), .Z(n14440) );
  AND U14435 ( .A(n14442), .B(n14443), .Z(n14430) );
  AND U14436 ( .A(n14444), .B(n14445), .Z(n14443) );
  XNOR U14437 ( .A(y[409]), .B(x[409]), .Z(n14445) );
  AND U14438 ( .A(n14446), .B(n14447), .Z(n14444) );
  XNOR U14439 ( .A(y[407]), .B(x[407]), .Z(n14447) );
  XNOR U14440 ( .A(y[408]), .B(x[408]), .Z(n14446) );
  AND U14441 ( .A(n14448), .B(n14449), .Z(n14442) );
  XNOR U14442 ( .A(y[410]), .B(x[410]), .Z(n14449) );
  XNOR U14443 ( .A(y[411]), .B(x[411]), .Z(n14448) );
  AND U14444 ( .A(n14450), .B(n14451), .Z(n14428) );
  AND U14445 ( .A(n14452), .B(n14453), .Z(n14451) );
  AND U14446 ( .A(n14454), .B(n14455), .Z(n14453) );
  XNOR U14447 ( .A(y[414]), .B(x[414]), .Z(n14455) );
  AND U14448 ( .A(n14456), .B(n14457), .Z(n14454) );
  XNOR U14449 ( .A(y[412]), .B(x[412]), .Z(n14457) );
  XNOR U14450 ( .A(y[413]), .B(x[413]), .Z(n14456) );
  AND U14451 ( .A(n14458), .B(n14459), .Z(n14452) );
  XNOR U14452 ( .A(y[415]), .B(x[415]), .Z(n14459) );
  XNOR U14453 ( .A(y[416]), .B(x[416]), .Z(n14458) );
  AND U14454 ( .A(n14460), .B(n14461), .Z(n14450) );
  AND U14455 ( .A(n14462), .B(n14463), .Z(n14461) );
  XNOR U14456 ( .A(y[419]), .B(x[419]), .Z(n14463) );
  AND U14457 ( .A(n14464), .B(n14465), .Z(n14462) );
  XNOR U14458 ( .A(y[417]), .B(x[417]), .Z(n14465) );
  XNOR U14459 ( .A(y[418]), .B(x[418]), .Z(n14464) );
  AND U14460 ( .A(n14466), .B(n14467), .Z(n14460) );
  XNOR U14461 ( .A(y[420]), .B(x[420]), .Z(n14467) );
  XNOR U14462 ( .A(y[421]), .B(x[421]), .Z(n14466) );
  AND U14463 ( .A(n14468), .B(n14469), .Z(n8620) );
  AND U14464 ( .A(n14470), .B(n14471), .Z(n14469) );
  AND U14465 ( .A(n14472), .B(n14473), .Z(n14471) );
  AND U14466 ( .A(n14474), .B(n14475), .Z(n14473) );
  AND U14467 ( .A(n14476), .B(n14477), .Z(n14475) );
  XNOR U14468 ( .A(y[424]), .B(x[424]), .Z(n14477) );
  AND U14469 ( .A(n14478), .B(n14479), .Z(n14476) );
  XNOR U14470 ( .A(y[422]), .B(x[422]), .Z(n14479) );
  XNOR U14471 ( .A(y[423]), .B(x[423]), .Z(n14478) );
  AND U14472 ( .A(n14480), .B(n14481), .Z(n14474) );
  XNOR U14473 ( .A(y[427]), .B(x[427]), .Z(n14481) );
  AND U14474 ( .A(n14482), .B(n14483), .Z(n14480) );
  XNOR U14475 ( .A(y[425]), .B(x[425]), .Z(n14483) );
  XNOR U14476 ( .A(y[426]), .B(x[426]), .Z(n14482) );
  AND U14477 ( .A(n14484), .B(n14485), .Z(n14472) );
  AND U14478 ( .A(n14486), .B(n14487), .Z(n14485) );
  XNOR U14479 ( .A(y[430]), .B(x[430]), .Z(n14487) );
  AND U14480 ( .A(n14488), .B(n14489), .Z(n14486) );
  XNOR U14481 ( .A(y[428]), .B(x[428]), .Z(n14489) );
  XNOR U14482 ( .A(y[429]), .B(x[429]), .Z(n14488) );
  AND U14483 ( .A(n14490), .B(n14491), .Z(n14484) );
  XNOR U14484 ( .A(y[431]), .B(x[431]), .Z(n14491) );
  XNOR U14485 ( .A(y[432]), .B(x[432]), .Z(n14490) );
  AND U14486 ( .A(n14492), .B(n14493), .Z(n14470) );
  AND U14487 ( .A(n14494), .B(n14495), .Z(n14493) );
  AND U14488 ( .A(n14496), .B(n14497), .Z(n14495) );
  XNOR U14489 ( .A(y[435]), .B(x[435]), .Z(n14497) );
  AND U14490 ( .A(n14498), .B(n14499), .Z(n14496) );
  XNOR U14491 ( .A(y[433]), .B(x[433]), .Z(n14499) );
  XNOR U14492 ( .A(y[434]), .B(x[434]), .Z(n14498) );
  AND U14493 ( .A(n14500), .B(n14501), .Z(n14494) );
  XNOR U14494 ( .A(y[436]), .B(x[436]), .Z(n14501) );
  XNOR U14495 ( .A(y[437]), .B(x[437]), .Z(n14500) );
  AND U14496 ( .A(n14502), .B(n14503), .Z(n14492) );
  AND U14497 ( .A(n14504), .B(n14505), .Z(n14503) );
  XNOR U14498 ( .A(y[440]), .B(x[440]), .Z(n14505) );
  AND U14499 ( .A(n14506), .B(n14507), .Z(n14504) );
  XNOR U14500 ( .A(y[438]), .B(x[438]), .Z(n14507) );
  XNOR U14501 ( .A(y[439]), .B(x[439]), .Z(n14506) );
  AND U14502 ( .A(n14508), .B(n14509), .Z(n14502) );
  XNOR U14503 ( .A(y[441]), .B(x[441]), .Z(n14509) );
  XNOR U14504 ( .A(y[442]), .B(x[442]), .Z(n14508) );
  AND U14505 ( .A(n14510), .B(n14511), .Z(n14468) );
  AND U14506 ( .A(n14512), .B(n14513), .Z(n14511) );
  AND U14507 ( .A(n14514), .B(n14515), .Z(n14513) );
  AND U14508 ( .A(n14516), .B(n14517), .Z(n14515) );
  XNOR U14509 ( .A(y[445]), .B(x[445]), .Z(n14517) );
  AND U14510 ( .A(n14518), .B(n14519), .Z(n14516) );
  XNOR U14511 ( .A(y[443]), .B(x[443]), .Z(n14519) );
  XNOR U14512 ( .A(y[444]), .B(x[444]), .Z(n14518) );
  AND U14513 ( .A(n14520), .B(n14521), .Z(n14514) );
  XNOR U14514 ( .A(y[448]), .B(x[448]), .Z(n14521) );
  AND U14515 ( .A(n14522), .B(n14523), .Z(n14520) );
  XNOR U14516 ( .A(y[446]), .B(x[446]), .Z(n14523) );
  XNOR U14517 ( .A(y[447]), .B(x[447]), .Z(n14522) );
  AND U14518 ( .A(n14524), .B(n14525), .Z(n14512) );
  AND U14519 ( .A(n14526), .B(n14527), .Z(n14525) );
  XNOR U14520 ( .A(y[451]), .B(x[451]), .Z(n14527) );
  AND U14521 ( .A(n14528), .B(n14529), .Z(n14526) );
  XNOR U14522 ( .A(y[449]), .B(x[449]), .Z(n14529) );
  XNOR U14523 ( .A(y[450]), .B(x[450]), .Z(n14528) );
  AND U14524 ( .A(n14530), .B(n14531), .Z(n14524) );
  XNOR U14525 ( .A(y[452]), .B(x[452]), .Z(n14531) );
  XNOR U14526 ( .A(y[453]), .B(x[453]), .Z(n14530) );
  AND U14527 ( .A(n14532), .B(n14533), .Z(n14510) );
  AND U14528 ( .A(n14534), .B(n14535), .Z(n14533) );
  AND U14529 ( .A(n14536), .B(n14537), .Z(n14535) );
  XNOR U14530 ( .A(y[456]), .B(x[456]), .Z(n14537) );
  AND U14531 ( .A(n14538), .B(n14539), .Z(n14536) );
  XNOR U14532 ( .A(y[454]), .B(x[454]), .Z(n14539) );
  XNOR U14533 ( .A(y[455]), .B(x[455]), .Z(n14538) );
  AND U14534 ( .A(n14540), .B(n14541), .Z(n14534) );
  XNOR U14535 ( .A(y[457]), .B(x[457]), .Z(n14541) );
  XNOR U14536 ( .A(y[458]), .B(x[458]), .Z(n14540) );
  AND U14537 ( .A(n14542), .B(n14543), .Z(n14532) );
  AND U14538 ( .A(n14544), .B(n14545), .Z(n14543) );
  XNOR U14539 ( .A(y[461]), .B(x[461]), .Z(n14545) );
  AND U14540 ( .A(n14546), .B(n14547), .Z(n14544) );
  XNOR U14541 ( .A(y[459]), .B(x[459]), .Z(n14547) );
  XNOR U14542 ( .A(y[460]), .B(x[460]), .Z(n14546) );
  AND U14543 ( .A(n14548), .B(n14549), .Z(n14542) );
  XNOR U14544 ( .A(y[958]), .B(x[958]), .Z(n14549) );
  XNOR U14545 ( .A(y[959]), .B(x[959]), .Z(n14548) );
  AND U14546 ( .A(n14550), .B(n14551), .Z(n8618) );
  AND U14547 ( .A(n14552), .B(n14553), .Z(n14551) );
  AND U14548 ( .A(n14554), .B(n14555), .Z(n14553) );
  AND U14549 ( .A(n14556), .B(n14557), .Z(n14555) );
  AND U14550 ( .A(n14558), .B(n14559), .Z(n14557) );
  AND U14551 ( .A(n14560), .B(n14561), .Z(n14559) );
  XNOR U14552 ( .A(y[962]), .B(x[962]), .Z(n14561) );
  AND U14553 ( .A(n14562), .B(n14563), .Z(n14560) );
  XNOR U14554 ( .A(y[960]), .B(x[960]), .Z(n14563) );
  XNOR U14555 ( .A(y[961]), .B(x[961]), .Z(n14562) );
  AND U14556 ( .A(n14564), .B(n14565), .Z(n14558) );
  XNOR U14557 ( .A(y[965]), .B(x[965]), .Z(n14565) );
  AND U14558 ( .A(n14566), .B(n14567), .Z(n14564) );
  XNOR U14559 ( .A(y[963]), .B(x[963]), .Z(n14567) );
  XNOR U14560 ( .A(y[964]), .B(x[964]), .Z(n14566) );
  AND U14561 ( .A(n14568), .B(n14569), .Z(n14556) );
  AND U14562 ( .A(n14570), .B(n14571), .Z(n14569) );
  XNOR U14563 ( .A(y[968]), .B(x[968]), .Z(n14571) );
  AND U14564 ( .A(n14572), .B(n14573), .Z(n14570) );
  XNOR U14565 ( .A(y[966]), .B(x[966]), .Z(n14573) );
  XNOR U14566 ( .A(y[967]), .B(x[967]), .Z(n14572) );
  AND U14567 ( .A(n14574), .B(n14575), .Z(n14568) );
  XNOR U14568 ( .A(y[969]), .B(x[969]), .Z(n14575) );
  XNOR U14569 ( .A(y[970]), .B(x[970]), .Z(n14574) );
  AND U14570 ( .A(n14576), .B(n14577), .Z(n14554) );
  AND U14571 ( .A(n14578), .B(n14579), .Z(n14577) );
  AND U14572 ( .A(n14580), .B(n14581), .Z(n14579) );
  XNOR U14573 ( .A(y[1261]), .B(x[1261]), .Z(n14581) );
  AND U14574 ( .A(n14582), .B(n14583), .Z(n14580) );
  XNOR U14575 ( .A(y[971]), .B(x[971]), .Z(n14583) );
  XNOR U14576 ( .A(y[1260]), .B(x[1260]), .Z(n14582) );
  AND U14577 ( .A(n14584), .B(n14585), .Z(n14578) );
  XNOR U14578 ( .A(y[1262]), .B(x[1262]), .Z(n14585) );
  XNOR U14579 ( .A(y[1263]), .B(x[1263]), .Z(n14584) );
  AND U14580 ( .A(n14586), .B(n14587), .Z(n14576) );
  AND U14581 ( .A(n14588), .B(n14589), .Z(n14587) );
  XNOR U14582 ( .A(y[1266]), .B(x[1266]), .Z(n14589) );
  AND U14583 ( .A(n14590), .B(n14591), .Z(n14588) );
  XNOR U14584 ( .A(y[1264]), .B(x[1264]), .Z(n14591) );
  XNOR U14585 ( .A(y[1265]), .B(x[1265]), .Z(n14590) );
  AND U14586 ( .A(n14592), .B(n14593), .Z(n14586) );
  XNOR U14587 ( .A(y[1267]), .B(x[1267]), .Z(n14593) );
  XNOR U14588 ( .A(y[1268]), .B(x[1268]), .Z(n14592) );
  AND U14589 ( .A(n14594), .B(n14595), .Z(n14552) );
  AND U14590 ( .A(n14596), .B(n14597), .Z(n14595) );
  AND U14591 ( .A(n14598), .B(n14599), .Z(n14597) );
  AND U14592 ( .A(n14600), .B(n14601), .Z(n14599) );
  XNOR U14593 ( .A(y[1271]), .B(x[1271]), .Z(n14601) );
  AND U14594 ( .A(n14602), .B(n14603), .Z(n14600) );
  XNOR U14595 ( .A(y[1269]), .B(x[1269]), .Z(n14603) );
  XNOR U14596 ( .A(y[1270]), .B(x[1270]), .Z(n14602) );
  AND U14597 ( .A(n14604), .B(n14605), .Z(n14598) );
  XNOR U14598 ( .A(y[1274]), .B(x[1274]), .Z(n14605) );
  AND U14599 ( .A(n14606), .B(n14607), .Z(n14604) );
  XNOR U14600 ( .A(y[1272]), .B(x[1272]), .Z(n14607) );
  XNOR U14601 ( .A(y[1273]), .B(x[1273]), .Z(n14606) );
  AND U14602 ( .A(n14608), .B(n14609), .Z(n14596) );
  AND U14603 ( .A(n14610), .B(n14611), .Z(n14609) );
  XNOR U14604 ( .A(y[1277]), .B(x[1277]), .Z(n14611) );
  AND U14605 ( .A(n14612), .B(n14613), .Z(n14610) );
  XNOR U14606 ( .A(y[1275]), .B(x[1275]), .Z(n14613) );
  XNOR U14607 ( .A(y[1276]), .B(x[1276]), .Z(n14612) );
  AND U14608 ( .A(n14614), .B(n14615), .Z(n14608) );
  XNOR U14609 ( .A(y[1278]), .B(x[1278]), .Z(n14615) );
  XNOR U14610 ( .A(y[1279]), .B(x[1279]), .Z(n14614) );
  AND U14611 ( .A(n14616), .B(n14617), .Z(n14594) );
  AND U14612 ( .A(n14618), .B(n14619), .Z(n14617) );
  AND U14613 ( .A(n14620), .B(n14621), .Z(n14619) );
  XNOR U14614 ( .A(y[1282]), .B(x[1282]), .Z(n14621) );
  AND U14615 ( .A(n14622), .B(n14623), .Z(n14620) );
  XNOR U14616 ( .A(y[1280]), .B(x[1280]), .Z(n14623) );
  XNOR U14617 ( .A(y[1281]), .B(x[1281]), .Z(n14622) );
  AND U14618 ( .A(n14624), .B(n14625), .Z(n14618) );
  XNOR U14619 ( .A(y[1283]), .B(x[1283]), .Z(n14625) );
  XNOR U14620 ( .A(y[1284]), .B(x[1284]), .Z(n14624) );
  AND U14621 ( .A(n14626), .B(n14627), .Z(n14616) );
  AND U14622 ( .A(n14628), .B(n14629), .Z(n14627) );
  XNOR U14623 ( .A(y[1287]), .B(x[1287]), .Z(n14629) );
  AND U14624 ( .A(n14630), .B(n14631), .Z(n14628) );
  XNOR U14625 ( .A(y[1285]), .B(x[1285]), .Z(n14631) );
  XNOR U14626 ( .A(y[1286]), .B(x[1286]), .Z(n14630) );
  AND U14627 ( .A(n14632), .B(n14633), .Z(n14626) );
  XNOR U14628 ( .A(y[1288]), .B(x[1288]), .Z(n14633) );
  XNOR U14629 ( .A(y[1289]), .B(x[1289]), .Z(n14632) );
  AND U14630 ( .A(n14634), .B(n14635), .Z(n14550) );
  AND U14631 ( .A(n14636), .B(n14637), .Z(n14635) );
  AND U14632 ( .A(n14638), .B(n14639), .Z(n14637) );
  AND U14633 ( .A(n14640), .B(n14641), .Z(n14639) );
  AND U14634 ( .A(n14642), .B(n14643), .Z(n14641) );
  XNOR U14635 ( .A(y[1292]), .B(x[1292]), .Z(n14643) );
  AND U14636 ( .A(n14644), .B(n14645), .Z(n14642) );
  XNOR U14637 ( .A(y[1290]), .B(x[1290]), .Z(n14645) );
  XNOR U14638 ( .A(y[1291]), .B(x[1291]), .Z(n14644) );
  AND U14639 ( .A(n14646), .B(n14647), .Z(n14640) );
  XNOR U14640 ( .A(y[1295]), .B(x[1295]), .Z(n14647) );
  AND U14641 ( .A(n14648), .B(n14649), .Z(n14646) );
  XNOR U14642 ( .A(y[1293]), .B(x[1293]), .Z(n14649) );
  XNOR U14643 ( .A(y[1294]), .B(x[1294]), .Z(n14648) );
  AND U14644 ( .A(n14650), .B(n14651), .Z(n14638) );
  AND U14645 ( .A(n14652), .B(n14653), .Z(n14651) );
  XNOR U14646 ( .A(y[1298]), .B(x[1298]), .Z(n14653) );
  AND U14647 ( .A(n14654), .B(n14655), .Z(n14652) );
  XNOR U14648 ( .A(y[1296]), .B(x[1296]), .Z(n14655) );
  XNOR U14649 ( .A(y[1297]), .B(x[1297]), .Z(n14654) );
  AND U14650 ( .A(n14656), .B(n14657), .Z(n14650) );
  XNOR U14651 ( .A(y[1299]), .B(x[1299]), .Z(n14657) );
  XNOR U14652 ( .A(y[1300]), .B(x[1300]), .Z(n14656) );
  AND U14653 ( .A(n14658), .B(n14659), .Z(n14636) );
  AND U14654 ( .A(n14660), .B(n14661), .Z(n14659) );
  AND U14655 ( .A(n14662), .B(n14663), .Z(n14661) );
  XNOR U14656 ( .A(y[1303]), .B(x[1303]), .Z(n14663) );
  AND U14657 ( .A(n14664), .B(n14665), .Z(n14662) );
  XNOR U14658 ( .A(y[1301]), .B(x[1301]), .Z(n14665) );
  XNOR U14659 ( .A(y[1302]), .B(x[1302]), .Z(n14664) );
  AND U14660 ( .A(n14666), .B(n14667), .Z(n14660) );
  XNOR U14661 ( .A(y[1304]), .B(x[1304]), .Z(n14667) );
  XNOR U14662 ( .A(y[1305]), .B(x[1305]), .Z(n14666) );
  AND U14663 ( .A(n14668), .B(n14669), .Z(n14658) );
  AND U14664 ( .A(n14670), .B(n14671), .Z(n14669) );
  XNOR U14665 ( .A(y[1308]), .B(x[1308]), .Z(n14671) );
  AND U14666 ( .A(n14672), .B(n14673), .Z(n14670) );
  XNOR U14667 ( .A(y[1306]), .B(x[1306]), .Z(n14673) );
  XNOR U14668 ( .A(y[1307]), .B(x[1307]), .Z(n14672) );
  AND U14669 ( .A(n14674), .B(n14675), .Z(n14668) );
  XNOR U14670 ( .A(y[1309]), .B(x[1309]), .Z(n14675) );
  XNOR U14671 ( .A(y[1310]), .B(x[1310]), .Z(n14674) );
  AND U14672 ( .A(n14676), .B(n14677), .Z(n14634) );
  AND U14673 ( .A(n14678), .B(n14679), .Z(n14677) );
  AND U14674 ( .A(n14680), .B(n14681), .Z(n14679) );
  AND U14675 ( .A(n14682), .B(n14683), .Z(n14681) );
  XNOR U14676 ( .A(y[1313]), .B(x[1313]), .Z(n14683) );
  AND U14677 ( .A(n14684), .B(n14685), .Z(n14682) );
  XNOR U14678 ( .A(y[1311]), .B(x[1311]), .Z(n14685) );
  XNOR U14679 ( .A(y[1312]), .B(x[1312]), .Z(n14684) );
  AND U14680 ( .A(n14686), .B(n14687), .Z(n14680) );
  XNOR U14681 ( .A(y[1316]), .B(x[1316]), .Z(n14687) );
  AND U14682 ( .A(n14688), .B(n14689), .Z(n14686) );
  XNOR U14683 ( .A(y[1314]), .B(x[1314]), .Z(n14689) );
  XNOR U14684 ( .A(y[1315]), .B(x[1315]), .Z(n14688) );
  AND U14685 ( .A(n14690), .B(n14691), .Z(n14678) );
  AND U14686 ( .A(n14692), .B(n14693), .Z(n14691) );
  XNOR U14687 ( .A(y[1319]), .B(x[1319]), .Z(n14693) );
  AND U14688 ( .A(n14694), .B(n14695), .Z(n14692) );
  XNOR U14689 ( .A(y[1317]), .B(x[1317]), .Z(n14695) );
  XNOR U14690 ( .A(y[1318]), .B(x[1318]), .Z(n14694) );
  AND U14691 ( .A(n14696), .B(n14697), .Z(n14690) );
  XNOR U14692 ( .A(y[1320]), .B(x[1320]), .Z(n14697) );
  XNOR U14693 ( .A(y[1321]), .B(x[1321]), .Z(n14696) );
  AND U14694 ( .A(n14698), .B(n14699), .Z(n14676) );
  AND U14695 ( .A(n14700), .B(n14701), .Z(n14699) );
  AND U14696 ( .A(n14702), .B(n14703), .Z(n14701) );
  XNOR U14697 ( .A(y[1324]), .B(x[1324]), .Z(n14703) );
  AND U14698 ( .A(n14704), .B(n14705), .Z(n14702) );
  XNOR U14699 ( .A(y[1322]), .B(x[1322]), .Z(n14705) );
  XNOR U14700 ( .A(y[1323]), .B(x[1323]), .Z(n14704) );
  AND U14701 ( .A(n14706), .B(n14707), .Z(n14700) );
  XNOR U14702 ( .A(y[1325]), .B(x[1325]), .Z(n14707) );
  XNOR U14703 ( .A(y[1326]), .B(x[1326]), .Z(n14706) );
  AND U14704 ( .A(n14708), .B(n14709), .Z(n14698) );
  AND U14705 ( .A(n14710), .B(n14711), .Z(n14709) );
  XNOR U14706 ( .A(y[1329]), .B(x[1329]), .Z(n14711) );
  AND U14707 ( .A(n14712), .B(n14713), .Z(n14710) );
  XNOR U14708 ( .A(y[1327]), .B(x[1327]), .Z(n14713) );
  XNOR U14709 ( .A(y[1328]), .B(x[1328]), .Z(n14712) );
  AND U14710 ( .A(n14714), .B(n14715), .Z(n14708) );
  XNOR U14711 ( .A(y[1330]), .B(x[1330]), .Z(n14715) );
  XNOR U14712 ( .A(y[1331]), .B(x[1331]), .Z(n14714) );
  AND U14713 ( .A(n14716), .B(n14717), .Z(n8616) );
  AND U14714 ( .A(n14718), .B(n14719), .Z(n14717) );
  AND U14715 ( .A(n14720), .B(n14721), .Z(n14719) );
  AND U14716 ( .A(n14722), .B(n14723), .Z(n14721) );
  AND U14717 ( .A(n14724), .B(n14725), .Z(n14723) );
  AND U14718 ( .A(n14726), .B(n14727), .Z(n14725) );
  AND U14719 ( .A(n14728), .B(n14729), .Z(n14727) );
  XNOR U14720 ( .A(y[1334]), .B(x[1334]), .Z(n14729) );
  AND U14721 ( .A(n14730), .B(n14731), .Z(n14728) );
  XNOR U14722 ( .A(y[1332]), .B(x[1332]), .Z(n14731) );
  XNOR U14723 ( .A(y[1333]), .B(x[1333]), .Z(n14730) );
  AND U14724 ( .A(n14732), .B(n14733), .Z(n14726) );
  XNOR U14725 ( .A(y[1337]), .B(x[1337]), .Z(n14733) );
  AND U14726 ( .A(n14734), .B(n14735), .Z(n14732) );
  XNOR U14727 ( .A(y[1335]), .B(x[1335]), .Z(n14735) );
  XNOR U14728 ( .A(y[1336]), .B(x[1336]), .Z(n14734) );
  AND U14729 ( .A(n14736), .B(n14737), .Z(n14724) );
  AND U14730 ( .A(n14738), .B(n14739), .Z(n14737) );
  XNOR U14731 ( .A(y[1340]), .B(x[1340]), .Z(n14739) );
  AND U14732 ( .A(n14740), .B(n14741), .Z(n14738) );
  XNOR U14733 ( .A(y[1338]), .B(x[1338]), .Z(n14741) );
  XNOR U14734 ( .A(y[1339]), .B(x[1339]), .Z(n14740) );
  AND U14735 ( .A(n14742), .B(n14743), .Z(n14736) );
  XNOR U14736 ( .A(y[1341]), .B(x[1341]), .Z(n14743) );
  XNOR U14737 ( .A(y[1342]), .B(x[1342]), .Z(n14742) );
  AND U14738 ( .A(n14744), .B(n14745), .Z(n14722) );
  AND U14739 ( .A(n14746), .B(n14747), .Z(n14745) );
  AND U14740 ( .A(n14748), .B(n14749), .Z(n14747) );
  XNOR U14741 ( .A(y[1345]), .B(x[1345]), .Z(n14749) );
  AND U14742 ( .A(n14750), .B(n14751), .Z(n14748) );
  XNOR U14743 ( .A(y[1343]), .B(x[1343]), .Z(n14751) );
  XNOR U14744 ( .A(y[1344]), .B(x[1344]), .Z(n14750) );
  AND U14745 ( .A(n14752), .B(n14753), .Z(n14746) );
  XNOR U14746 ( .A(y[1346]), .B(x[1346]), .Z(n14753) );
  XNOR U14747 ( .A(y[1347]), .B(x[1347]), .Z(n14752) );
  AND U14748 ( .A(n14754), .B(n14755), .Z(n14744) );
  AND U14749 ( .A(n14756), .B(n14757), .Z(n14755) );
  XNOR U14750 ( .A(y[1350]), .B(x[1350]), .Z(n14757) );
  AND U14751 ( .A(n14758), .B(n14759), .Z(n14756) );
  XNOR U14752 ( .A(y[1348]), .B(x[1348]), .Z(n14759) );
  XNOR U14753 ( .A(y[1349]), .B(x[1349]), .Z(n14758) );
  AND U14754 ( .A(n14760), .B(n14761), .Z(n14754) );
  XNOR U14755 ( .A(y[1351]), .B(x[1351]), .Z(n14761) );
  XNOR U14756 ( .A(y[1352]), .B(x[1352]), .Z(n14760) );
  AND U14757 ( .A(n14762), .B(n14763), .Z(n14720) );
  AND U14758 ( .A(n14764), .B(n14765), .Z(n14763) );
  AND U14759 ( .A(n14766), .B(n14767), .Z(n14765) );
  AND U14760 ( .A(n14768), .B(n14769), .Z(n14767) );
  XNOR U14761 ( .A(y[1355]), .B(x[1355]), .Z(n14769) );
  AND U14762 ( .A(n14770), .B(n14771), .Z(n14768) );
  XNOR U14763 ( .A(y[1353]), .B(x[1353]), .Z(n14771) );
  XNOR U14764 ( .A(y[1354]), .B(x[1354]), .Z(n14770) );
  AND U14765 ( .A(n14772), .B(n14773), .Z(n14766) );
  XNOR U14766 ( .A(y[1358]), .B(x[1358]), .Z(n14773) );
  AND U14767 ( .A(n14774), .B(n14775), .Z(n14772) );
  XNOR U14768 ( .A(y[1356]), .B(x[1356]), .Z(n14775) );
  XNOR U14769 ( .A(y[1357]), .B(x[1357]), .Z(n14774) );
  AND U14770 ( .A(n14776), .B(n14777), .Z(n14764) );
  AND U14771 ( .A(n14778), .B(n14779), .Z(n14777) );
  XNOR U14772 ( .A(y[1361]), .B(x[1361]), .Z(n14779) );
  AND U14773 ( .A(n14780), .B(n14781), .Z(n14778) );
  XNOR U14774 ( .A(y[1359]), .B(x[1359]), .Z(n14781) );
  XNOR U14775 ( .A(y[1360]), .B(x[1360]), .Z(n14780) );
  AND U14776 ( .A(n14782), .B(n14783), .Z(n14776) );
  XNOR U14777 ( .A(y[1362]), .B(x[1362]), .Z(n14783) );
  XNOR U14778 ( .A(y[1363]), .B(x[1363]), .Z(n14782) );
  AND U14779 ( .A(n14784), .B(n14785), .Z(n14762) );
  AND U14780 ( .A(n14786), .B(n14787), .Z(n14785) );
  AND U14781 ( .A(n14788), .B(n14789), .Z(n14787) );
  XNOR U14782 ( .A(y[1366]), .B(x[1366]), .Z(n14789) );
  AND U14783 ( .A(n14790), .B(n14791), .Z(n14788) );
  XNOR U14784 ( .A(y[1364]), .B(x[1364]), .Z(n14791) );
  XNOR U14785 ( .A(y[1365]), .B(x[1365]), .Z(n14790) );
  AND U14786 ( .A(n14792), .B(n14793), .Z(n14786) );
  XNOR U14787 ( .A(y[1367]), .B(x[1367]), .Z(n14793) );
  XNOR U14788 ( .A(y[1368]), .B(x[1368]), .Z(n14792) );
  AND U14789 ( .A(n14794), .B(n14795), .Z(n14784) );
  AND U14790 ( .A(n14796), .B(n14797), .Z(n14795) );
  XNOR U14791 ( .A(y[1371]), .B(x[1371]), .Z(n14797) );
  AND U14792 ( .A(n14798), .B(n14799), .Z(n14796) );
  XNOR U14793 ( .A(y[1369]), .B(x[1369]), .Z(n14799) );
  XNOR U14794 ( .A(y[1370]), .B(x[1370]), .Z(n14798) );
  AND U14795 ( .A(n14800), .B(n14801), .Z(n14794) );
  XNOR U14796 ( .A(y[1372]), .B(x[1372]), .Z(n14801) );
  XNOR U14797 ( .A(y[1373]), .B(x[1373]), .Z(n14800) );
  AND U14798 ( .A(n14802), .B(n14803), .Z(n14718) );
  AND U14799 ( .A(n14804), .B(n14805), .Z(n14803) );
  AND U14800 ( .A(n14806), .B(n14807), .Z(n14805) );
  AND U14801 ( .A(n14808), .B(n14809), .Z(n14807) );
  AND U14802 ( .A(n14810), .B(n14811), .Z(n14809) );
  XNOR U14803 ( .A(y[1376]), .B(x[1376]), .Z(n14811) );
  AND U14804 ( .A(n14812), .B(n14813), .Z(n14810) );
  XNOR U14805 ( .A(y[1374]), .B(x[1374]), .Z(n14813) );
  XNOR U14806 ( .A(y[1375]), .B(x[1375]), .Z(n14812) );
  AND U14807 ( .A(n14814), .B(n14815), .Z(n14808) );
  XNOR U14808 ( .A(y[1379]), .B(x[1379]), .Z(n14815) );
  AND U14809 ( .A(n14816), .B(n14817), .Z(n14814) );
  XNOR U14810 ( .A(y[1377]), .B(x[1377]), .Z(n14817) );
  XNOR U14811 ( .A(y[1378]), .B(x[1378]), .Z(n14816) );
  AND U14812 ( .A(n14818), .B(n14819), .Z(n14806) );
  AND U14813 ( .A(n14820), .B(n14821), .Z(n14819) );
  XNOR U14814 ( .A(y[1382]), .B(x[1382]), .Z(n14821) );
  AND U14815 ( .A(n14822), .B(n14823), .Z(n14820) );
  XNOR U14816 ( .A(y[1380]), .B(x[1380]), .Z(n14823) );
  XNOR U14817 ( .A(y[1381]), .B(x[1381]), .Z(n14822) );
  AND U14818 ( .A(n14824), .B(n14825), .Z(n14818) );
  XNOR U14819 ( .A(y[1383]), .B(x[1383]), .Z(n14825) );
  XNOR U14820 ( .A(y[1384]), .B(x[1384]), .Z(n14824) );
  AND U14821 ( .A(n14826), .B(n14827), .Z(n14804) );
  AND U14822 ( .A(n14828), .B(n14829), .Z(n14827) );
  AND U14823 ( .A(n14830), .B(n14831), .Z(n14829) );
  XNOR U14824 ( .A(y[1387]), .B(x[1387]), .Z(n14831) );
  AND U14825 ( .A(n14832), .B(n14833), .Z(n14830) );
  XNOR U14826 ( .A(y[1385]), .B(x[1385]), .Z(n14833) );
  XNOR U14827 ( .A(y[1386]), .B(x[1386]), .Z(n14832) );
  AND U14828 ( .A(n14834), .B(n14835), .Z(n14828) );
  XNOR U14829 ( .A(y[1388]), .B(x[1388]), .Z(n14835) );
  XNOR U14830 ( .A(y[1389]), .B(x[1389]), .Z(n14834) );
  AND U14831 ( .A(n14836), .B(n14837), .Z(n14826) );
  AND U14832 ( .A(n14838), .B(n14839), .Z(n14837) );
  XNOR U14833 ( .A(y[1392]), .B(x[1392]), .Z(n14839) );
  AND U14834 ( .A(n14840), .B(n14841), .Z(n14838) );
  XNOR U14835 ( .A(y[1390]), .B(x[1390]), .Z(n14841) );
  XNOR U14836 ( .A(y[1391]), .B(x[1391]), .Z(n14840) );
  AND U14837 ( .A(n14842), .B(n14843), .Z(n14836) );
  XNOR U14838 ( .A(y[1393]), .B(x[1393]), .Z(n14843) );
  XNOR U14839 ( .A(y[1394]), .B(x[1394]), .Z(n14842) );
  AND U14840 ( .A(n14844), .B(n14845), .Z(n14802) );
  AND U14841 ( .A(n14846), .B(n14847), .Z(n14845) );
  AND U14842 ( .A(n14848), .B(n14849), .Z(n14847) );
  AND U14843 ( .A(n14850), .B(n14851), .Z(n14849) );
  XNOR U14844 ( .A(y[1397]), .B(x[1397]), .Z(n14851) );
  AND U14845 ( .A(n14852), .B(n14853), .Z(n14850) );
  XNOR U14846 ( .A(y[1395]), .B(x[1395]), .Z(n14853) );
  XNOR U14847 ( .A(y[1396]), .B(x[1396]), .Z(n14852) );
  AND U14848 ( .A(n14854), .B(n14855), .Z(n14848) );
  XNOR U14849 ( .A(y[1400]), .B(x[1400]), .Z(n14855) );
  AND U14850 ( .A(n14856), .B(n14857), .Z(n14854) );
  XNOR U14851 ( .A(y[1398]), .B(x[1398]), .Z(n14857) );
  XNOR U14852 ( .A(y[1399]), .B(x[1399]), .Z(n14856) );
  AND U14853 ( .A(n14858), .B(n14859), .Z(n14846) );
  AND U14854 ( .A(n14860), .B(n14861), .Z(n14859) );
  XNOR U14855 ( .A(y[1403]), .B(x[1403]), .Z(n14861) );
  AND U14856 ( .A(n14862), .B(n14863), .Z(n14860) );
  XNOR U14857 ( .A(y[1401]), .B(x[1401]), .Z(n14863) );
  XNOR U14858 ( .A(y[1402]), .B(x[1402]), .Z(n14862) );
  AND U14859 ( .A(n14864), .B(n14865), .Z(n14858) );
  XNOR U14860 ( .A(y[1404]), .B(x[1404]), .Z(n14865) );
  XNOR U14861 ( .A(y[1405]), .B(x[1405]), .Z(n14864) );
  AND U14862 ( .A(n14866), .B(n14867), .Z(n14844) );
  AND U14863 ( .A(n14868), .B(n14869), .Z(n14867) );
  AND U14864 ( .A(n14870), .B(n14871), .Z(n14869) );
  XNOR U14865 ( .A(y[1408]), .B(x[1408]), .Z(n14871) );
  AND U14866 ( .A(n14872), .B(n14873), .Z(n14870) );
  XNOR U14867 ( .A(y[1406]), .B(x[1406]), .Z(n14873) );
  XNOR U14868 ( .A(y[1407]), .B(x[1407]), .Z(n14872) );
  AND U14869 ( .A(n14874), .B(n14875), .Z(n14868) );
  XNOR U14870 ( .A(y[1409]), .B(x[1409]), .Z(n14875) );
  XNOR U14871 ( .A(y[1410]), .B(x[1410]), .Z(n14874) );
  AND U14872 ( .A(n14876), .B(n14877), .Z(n14866) );
  AND U14873 ( .A(n14878), .B(n14879), .Z(n14877) );
  XNOR U14874 ( .A(y[1413]), .B(x[1413]), .Z(n14879) );
  AND U14875 ( .A(n14880), .B(n14881), .Z(n14878) );
  XNOR U14876 ( .A(y[1411]), .B(x[1411]), .Z(n14881) );
  XNOR U14877 ( .A(y[1412]), .B(x[1412]), .Z(n14880) );
  AND U14878 ( .A(n14882), .B(n14883), .Z(n14876) );
  XNOR U14879 ( .A(y[1414]), .B(x[1414]), .Z(n14883) );
  XNOR U14880 ( .A(y[1415]), .B(x[1415]), .Z(n14882) );
  AND U14881 ( .A(n14884), .B(n14885), .Z(n14716) );
  AND U14882 ( .A(n14886), .B(n14887), .Z(n14885) );
  AND U14883 ( .A(n14888), .B(n14889), .Z(n14887) );
  AND U14884 ( .A(n14890), .B(n14891), .Z(n14889) );
  AND U14885 ( .A(n14892), .B(n14893), .Z(n14891) );
  AND U14886 ( .A(n14894), .B(n14895), .Z(n14893) );
  XNOR U14887 ( .A(y[1418]), .B(x[1418]), .Z(n14895) );
  AND U14888 ( .A(n14896), .B(n14897), .Z(n14894) );
  XNOR U14889 ( .A(y[1416]), .B(x[1416]), .Z(n14897) );
  XNOR U14890 ( .A(y[1417]), .B(x[1417]), .Z(n14896) );
  AND U14891 ( .A(n14898), .B(n14899), .Z(n14892) );
  XNOR U14892 ( .A(y[1421]), .B(x[1421]), .Z(n14899) );
  AND U14893 ( .A(n14900), .B(n14901), .Z(n14898) );
  XNOR U14894 ( .A(y[1419]), .B(x[1419]), .Z(n14901) );
  XNOR U14895 ( .A(y[1420]), .B(x[1420]), .Z(n14900) );
  AND U14896 ( .A(n14902), .B(n14903), .Z(n14890) );
  AND U14897 ( .A(n14904), .B(n14905), .Z(n14903) );
  XNOR U14898 ( .A(y[1424]), .B(x[1424]), .Z(n14905) );
  AND U14899 ( .A(n14906), .B(n14907), .Z(n14904) );
  XNOR U14900 ( .A(y[1422]), .B(x[1422]), .Z(n14907) );
  XNOR U14901 ( .A(y[1423]), .B(x[1423]), .Z(n14906) );
  AND U14902 ( .A(n14908), .B(n14909), .Z(n14902) );
  XNOR U14903 ( .A(y[1425]), .B(x[1425]), .Z(n14909) );
  XNOR U14904 ( .A(y[1426]), .B(x[1426]), .Z(n14908) );
  AND U14905 ( .A(n14910), .B(n14911), .Z(n14888) );
  AND U14906 ( .A(n14912), .B(n14913), .Z(n14911) );
  AND U14907 ( .A(n14914), .B(n14915), .Z(n14913) );
  XNOR U14908 ( .A(y[1429]), .B(x[1429]), .Z(n14915) );
  AND U14909 ( .A(n14916), .B(n14917), .Z(n14914) );
  XNOR U14910 ( .A(y[1427]), .B(x[1427]), .Z(n14917) );
  XNOR U14911 ( .A(y[1428]), .B(x[1428]), .Z(n14916) );
  AND U14912 ( .A(n14918), .B(n14919), .Z(n14912) );
  XNOR U14913 ( .A(y[1430]), .B(x[1430]), .Z(n14919) );
  XNOR U14914 ( .A(y[1431]), .B(x[1431]), .Z(n14918) );
  AND U14915 ( .A(n14920), .B(n14921), .Z(n14910) );
  AND U14916 ( .A(n14922), .B(n14923), .Z(n14921) );
  XNOR U14917 ( .A(y[1434]), .B(x[1434]), .Z(n14923) );
  AND U14918 ( .A(n14924), .B(n14925), .Z(n14922) );
  XNOR U14919 ( .A(y[1432]), .B(x[1432]), .Z(n14925) );
  XNOR U14920 ( .A(y[1433]), .B(x[1433]), .Z(n14924) );
  AND U14921 ( .A(n14926), .B(n14927), .Z(n14920) );
  XNOR U14922 ( .A(y[1435]), .B(x[1435]), .Z(n14927) );
  XNOR U14923 ( .A(y[1436]), .B(x[1436]), .Z(n14926) );
  AND U14924 ( .A(n14928), .B(n14929), .Z(n14886) );
  AND U14925 ( .A(n14930), .B(n14931), .Z(n14929) );
  AND U14926 ( .A(n14932), .B(n14933), .Z(n14931) );
  AND U14927 ( .A(n14934), .B(n14935), .Z(n14933) );
  XNOR U14928 ( .A(y[1439]), .B(x[1439]), .Z(n14935) );
  AND U14929 ( .A(n14936), .B(n14937), .Z(n14934) );
  XNOR U14930 ( .A(y[1437]), .B(x[1437]), .Z(n14937) );
  XNOR U14931 ( .A(y[1438]), .B(x[1438]), .Z(n14936) );
  AND U14932 ( .A(n14938), .B(n14939), .Z(n14932) );
  XNOR U14933 ( .A(y[1442]), .B(x[1442]), .Z(n14939) );
  AND U14934 ( .A(n14940), .B(n14941), .Z(n14938) );
  XNOR U14935 ( .A(y[1440]), .B(x[1440]), .Z(n14941) );
  XNOR U14936 ( .A(y[1441]), .B(x[1441]), .Z(n14940) );
  AND U14937 ( .A(n14942), .B(n14943), .Z(n14930) );
  AND U14938 ( .A(n14944), .B(n14945), .Z(n14943) );
  XNOR U14939 ( .A(y[1445]), .B(x[1445]), .Z(n14945) );
  AND U14940 ( .A(n14946), .B(n14947), .Z(n14944) );
  XNOR U14941 ( .A(y[1443]), .B(x[1443]), .Z(n14947) );
  XNOR U14942 ( .A(y[1444]), .B(x[1444]), .Z(n14946) );
  AND U14943 ( .A(n14948), .B(n14949), .Z(n14942) );
  XNOR U14944 ( .A(y[1446]), .B(x[1446]), .Z(n14949) );
  XNOR U14945 ( .A(y[1447]), .B(x[1447]), .Z(n14948) );
  AND U14946 ( .A(n14950), .B(n14951), .Z(n14928) );
  AND U14947 ( .A(n14952), .B(n14953), .Z(n14951) );
  AND U14948 ( .A(n14954), .B(n14955), .Z(n14953) );
  XNOR U14949 ( .A(y[1450]), .B(x[1450]), .Z(n14955) );
  AND U14950 ( .A(n14956), .B(n14957), .Z(n14954) );
  XNOR U14951 ( .A(y[1448]), .B(x[1448]), .Z(n14957) );
  XNOR U14952 ( .A(y[1449]), .B(x[1449]), .Z(n14956) );
  AND U14953 ( .A(n14958), .B(n14959), .Z(n14952) );
  XNOR U14954 ( .A(y[1451]), .B(x[1451]), .Z(n14959) );
  XNOR U14955 ( .A(y[1452]), .B(x[1452]), .Z(n14958) );
  AND U14956 ( .A(n14960), .B(n14961), .Z(n14950) );
  AND U14957 ( .A(n14962), .B(n14963), .Z(n14961) );
  XNOR U14958 ( .A(y[1455]), .B(x[1455]), .Z(n14963) );
  AND U14959 ( .A(n14964), .B(n14965), .Z(n14962) );
  XNOR U14960 ( .A(y[1453]), .B(x[1453]), .Z(n14965) );
  XNOR U14961 ( .A(y[1454]), .B(x[1454]), .Z(n14964) );
  AND U14962 ( .A(n14966), .B(n14967), .Z(n14960) );
  XNOR U14963 ( .A(y[1456]), .B(x[1456]), .Z(n14967) );
  XNOR U14964 ( .A(y[1457]), .B(x[1457]), .Z(n14966) );
  AND U14965 ( .A(n14968), .B(n14969), .Z(n14884) );
  AND U14966 ( .A(n14970), .B(n14971), .Z(n14969) );
  AND U14967 ( .A(n14972), .B(n14973), .Z(n14971) );
  AND U14968 ( .A(n14974), .B(n14975), .Z(n14973) );
  AND U14969 ( .A(n14976), .B(n14977), .Z(n14975) );
  XNOR U14970 ( .A(y[1460]), .B(x[1460]), .Z(n14977) );
  AND U14971 ( .A(n14978), .B(n14979), .Z(n14976) );
  XNOR U14972 ( .A(y[1458]), .B(x[1458]), .Z(n14979) );
  XNOR U14973 ( .A(y[1459]), .B(x[1459]), .Z(n14978) );
  AND U14974 ( .A(n14980), .B(n14981), .Z(n14974) );
  XNOR U14975 ( .A(y[1463]), .B(x[1463]), .Z(n14981) );
  AND U14976 ( .A(n14982), .B(n14983), .Z(n14980) );
  XNOR U14977 ( .A(y[1461]), .B(x[1461]), .Z(n14983) );
  XNOR U14978 ( .A(y[1462]), .B(x[1462]), .Z(n14982) );
  AND U14979 ( .A(n14984), .B(n14985), .Z(n14972) );
  AND U14980 ( .A(n14986), .B(n14987), .Z(n14985) );
  XNOR U14981 ( .A(y[1466]), .B(x[1466]), .Z(n14987) );
  AND U14982 ( .A(n14988), .B(n14989), .Z(n14986) );
  XNOR U14983 ( .A(y[1464]), .B(x[1464]), .Z(n14989) );
  XNOR U14984 ( .A(y[1465]), .B(x[1465]), .Z(n14988) );
  AND U14985 ( .A(n14990), .B(n14991), .Z(n14984) );
  XNOR U14986 ( .A(y[1467]), .B(x[1467]), .Z(n14991) );
  XNOR U14987 ( .A(y[1468]), .B(x[1468]), .Z(n14990) );
  AND U14988 ( .A(n14992), .B(n14993), .Z(n14970) );
  AND U14989 ( .A(n14994), .B(n14995), .Z(n14993) );
  AND U14990 ( .A(n14996), .B(n14997), .Z(n14995) );
  XNOR U14991 ( .A(y[1471]), .B(x[1471]), .Z(n14997) );
  AND U14992 ( .A(n14998), .B(n14999), .Z(n14996) );
  XNOR U14993 ( .A(y[1469]), .B(x[1469]), .Z(n14999) );
  XNOR U14994 ( .A(y[1470]), .B(x[1470]), .Z(n14998) );
  AND U14995 ( .A(n15000), .B(n15001), .Z(n14994) );
  XNOR U14996 ( .A(y[1472]), .B(x[1472]), .Z(n15001) );
  XNOR U14997 ( .A(y[1473]), .B(x[1473]), .Z(n15000) );
  AND U14998 ( .A(n15002), .B(n15003), .Z(n14992) );
  AND U14999 ( .A(n15004), .B(n15005), .Z(n15003) );
  XNOR U15000 ( .A(y[1476]), .B(x[1476]), .Z(n15005) );
  AND U15001 ( .A(n15006), .B(n15007), .Z(n15004) );
  XNOR U15002 ( .A(y[1474]), .B(x[1474]), .Z(n15007) );
  XNOR U15003 ( .A(y[1475]), .B(x[1475]), .Z(n15006) );
  AND U15004 ( .A(n15008), .B(n15009), .Z(n15002) );
  XNOR U15005 ( .A(y[1477]), .B(x[1477]), .Z(n15009) );
  XNOR U15006 ( .A(y[1478]), .B(x[1478]), .Z(n15008) );
  AND U15007 ( .A(n15010), .B(n15011), .Z(n14968) );
  AND U15008 ( .A(n15012), .B(n15013), .Z(n15011) );
  AND U15009 ( .A(n15014), .B(n15015), .Z(n15013) );
  AND U15010 ( .A(n15016), .B(n15017), .Z(n15015) );
  XNOR U15011 ( .A(y[1481]), .B(x[1481]), .Z(n15017) );
  AND U15012 ( .A(n15018), .B(n15019), .Z(n15016) );
  XNOR U15013 ( .A(y[1479]), .B(x[1479]), .Z(n15019) );
  XNOR U15014 ( .A(y[1480]), .B(x[1480]), .Z(n15018) );
  AND U15015 ( .A(n15020), .B(n15021), .Z(n15014) );
  XNOR U15016 ( .A(y[1484]), .B(x[1484]), .Z(n15021) );
  AND U15017 ( .A(n15022), .B(n15023), .Z(n15020) );
  XNOR U15018 ( .A(y[1482]), .B(x[1482]), .Z(n15023) );
  XNOR U15019 ( .A(y[1483]), .B(x[1483]), .Z(n15022) );
  AND U15020 ( .A(n15024), .B(n15025), .Z(n15012) );
  AND U15021 ( .A(n15026), .B(n15027), .Z(n15025) );
  XNOR U15022 ( .A(y[1487]), .B(x[1487]), .Z(n15027) );
  AND U15023 ( .A(n15028), .B(n15029), .Z(n15026) );
  XNOR U15024 ( .A(y[1485]), .B(x[1485]), .Z(n15029) );
  XNOR U15025 ( .A(y[1486]), .B(x[1486]), .Z(n15028) );
  AND U15026 ( .A(n15030), .B(n15031), .Z(n15024) );
  XNOR U15027 ( .A(y[1488]), .B(x[1488]), .Z(n15031) );
  XNOR U15028 ( .A(y[1489]), .B(x[1489]), .Z(n15030) );
  AND U15029 ( .A(n15032), .B(n15033), .Z(n15010) );
  AND U15030 ( .A(n15034), .B(n15035), .Z(n15033) );
  AND U15031 ( .A(n15036), .B(n15037), .Z(n15035) );
  XNOR U15032 ( .A(y[1492]), .B(x[1492]), .Z(n15037) );
  AND U15033 ( .A(n15038), .B(n15039), .Z(n15036) );
  XNOR U15034 ( .A(y[1490]), .B(x[1490]), .Z(n15039) );
  XNOR U15035 ( .A(y[1491]), .B(x[1491]), .Z(n15038) );
  AND U15036 ( .A(n15040), .B(n15041), .Z(n15034) );
  XNOR U15037 ( .A(y[1493]), .B(x[1493]), .Z(n15041) );
  XNOR U15038 ( .A(y[1494]), .B(x[1494]), .Z(n15040) );
  AND U15039 ( .A(n15042), .B(n15043), .Z(n15032) );
  AND U15040 ( .A(n15044), .B(n15045), .Z(n15043) );
  XNOR U15041 ( .A(y[1497]), .B(x[1497]), .Z(n15045) );
  AND U15042 ( .A(n15046), .B(n15047), .Z(n15044) );
  XNOR U15043 ( .A(y[1495]), .B(x[1495]), .Z(n15047) );
  XNOR U15044 ( .A(y[1496]), .B(x[1496]), .Z(n15046) );
  AND U15045 ( .A(n15048), .B(n15049), .Z(n15042) );
  XNOR U15046 ( .A(y[1498]), .B(x[1498]), .Z(n15049) );
  XNOR U15047 ( .A(y[1499]), .B(x[1499]), .Z(n15048) );
  AND U15048 ( .A(n15050), .B(n15051), .Z(n8214) );
  AND U15049 ( .A(n15052), .B(n15053), .Z(n15051) );
  AND U15050 ( .A(n15054), .B(n15055), .Z(n15053) );
  AND U15051 ( .A(n15056), .B(n15057), .Z(n15055) );
  AND U15052 ( .A(n15058), .B(n15059), .Z(n15057) );
  AND U15053 ( .A(n15060), .B(n15061), .Z(n15059) );
  AND U15054 ( .A(n15062), .B(n15063), .Z(n15061) );
  AND U15055 ( .A(n15064), .B(n15065), .Z(n15063) );
  AND U15056 ( .A(n15066), .B(n15067), .Z(n15065) );
  XNOR U15057 ( .A(y[462]), .B(x[462]), .Z(n15067) );
  XNOR U15058 ( .A(y[463]), .B(x[463]), .Z(n15066) );
  AND U15059 ( .A(n15068), .B(n15069), .Z(n15064) );
  XNOR U15060 ( .A(y[464]), .B(x[464]), .Z(n15069) );
  XNOR U15061 ( .A(y[465]), .B(x[465]), .Z(n15068) );
  AND U15062 ( .A(n15070), .B(n15071), .Z(n15062) );
  AND U15063 ( .A(n15072), .B(n15073), .Z(n15071) );
  XNOR U15064 ( .A(y[466]), .B(x[466]), .Z(n15073) );
  XNOR U15065 ( .A(y[467]), .B(x[467]), .Z(n15072) );
  AND U15066 ( .A(n15074), .B(n15075), .Z(n15070) );
  XNOR U15067 ( .A(y[468]), .B(x[468]), .Z(n15075) );
  XNOR U15068 ( .A(y[469]), .B(x[469]), .Z(n15074) );
  AND U15069 ( .A(n15076), .B(n15077), .Z(n15060) );
  AND U15070 ( .A(n15078), .B(n15079), .Z(n15077) );
  AND U15071 ( .A(n15080), .B(n15081), .Z(n15079) );
  XNOR U15072 ( .A(y[470]), .B(x[470]), .Z(n15081) );
  XNOR U15073 ( .A(y[471]), .B(x[471]), .Z(n15080) );
  AND U15074 ( .A(n15082), .B(n15083), .Z(n15078) );
  XNOR U15075 ( .A(y[472]), .B(x[472]), .Z(n15083) );
  XNOR U15076 ( .A(y[473]), .B(x[473]), .Z(n15082) );
  AND U15077 ( .A(n15084), .B(n15085), .Z(n15076) );
  AND U15078 ( .A(n15086), .B(n15087), .Z(n15085) );
  XNOR U15079 ( .A(y[474]), .B(x[474]), .Z(n15087) );
  XNOR U15080 ( .A(y[475]), .B(x[475]), .Z(n15086) );
  AND U15081 ( .A(n15088), .B(n15089), .Z(n15084) );
  XNOR U15082 ( .A(y[476]), .B(x[476]), .Z(n15089) );
  XNOR U15083 ( .A(y[477]), .B(x[477]), .Z(n15088) );
  AND U15084 ( .A(n15090), .B(n15091), .Z(n15058) );
  AND U15085 ( .A(n15092), .B(n15093), .Z(n15091) );
  AND U15086 ( .A(n15094), .B(n15095), .Z(n15093) );
  AND U15087 ( .A(n15096), .B(n15097), .Z(n15095) );
  XNOR U15088 ( .A(y[478]), .B(x[478]), .Z(n15097) );
  XNOR U15089 ( .A(y[479]), .B(x[479]), .Z(n15096) );
  AND U15090 ( .A(n15098), .B(n15099), .Z(n15094) );
  XNOR U15091 ( .A(y[480]), .B(x[480]), .Z(n15099) );
  XNOR U15092 ( .A(y[481]), .B(x[481]), .Z(n15098) );
  AND U15093 ( .A(n15100), .B(n15101), .Z(n15092) );
  AND U15094 ( .A(n15102), .B(n15103), .Z(n15101) );
  XNOR U15095 ( .A(y[482]), .B(x[482]), .Z(n15103) );
  XNOR U15096 ( .A(y[483]), .B(x[483]), .Z(n15102) );
  AND U15097 ( .A(n15104), .B(n15105), .Z(n15100) );
  XNOR U15098 ( .A(y[484]), .B(x[484]), .Z(n15105) );
  XNOR U15099 ( .A(y[485]), .B(x[485]), .Z(n15104) );
  AND U15100 ( .A(n15106), .B(n15107), .Z(n15090) );
  AND U15101 ( .A(n15108), .B(n15109), .Z(n15107) );
  AND U15102 ( .A(n15110), .B(n15111), .Z(n15109) );
  XNOR U15103 ( .A(y[486]), .B(x[486]), .Z(n15111) );
  XNOR U15104 ( .A(y[487]), .B(x[487]), .Z(n15110) );
  AND U15105 ( .A(n15112), .B(n15113), .Z(n15108) );
  XNOR U15106 ( .A(y[488]), .B(x[488]), .Z(n15113) );
  XNOR U15107 ( .A(y[489]), .B(x[489]), .Z(n15112) );
  AND U15108 ( .A(n15114), .B(n15115), .Z(n15106) );
  AND U15109 ( .A(n15116), .B(n15117), .Z(n15115) );
  XNOR U15110 ( .A(y[490]), .B(x[490]), .Z(n15117) );
  XNOR U15111 ( .A(y[491]), .B(x[491]), .Z(n15116) );
  AND U15112 ( .A(n15118), .B(n15119), .Z(n15114) );
  XNOR U15113 ( .A(y[492]), .B(x[492]), .Z(n15119) );
  XNOR U15114 ( .A(y[493]), .B(x[493]), .Z(n15118) );
  AND U15115 ( .A(n15120), .B(n15121), .Z(n15056) );
  AND U15116 ( .A(n15122), .B(n15123), .Z(n15121) );
  AND U15117 ( .A(n15124), .B(n15125), .Z(n15123) );
  AND U15118 ( .A(n15126), .B(n15127), .Z(n15125) );
  AND U15119 ( .A(n15128), .B(n15129), .Z(n15127) );
  XNOR U15120 ( .A(y[494]), .B(x[494]), .Z(n15129) );
  XNOR U15121 ( .A(y[495]), .B(x[495]), .Z(n15128) );
  AND U15122 ( .A(n15130), .B(n15131), .Z(n15126) );
  XNOR U15123 ( .A(y[496]), .B(x[496]), .Z(n15131) );
  XNOR U15124 ( .A(y[497]), .B(x[497]), .Z(n15130) );
  AND U15125 ( .A(n15132), .B(n15133), .Z(n15124) );
  AND U15126 ( .A(n15134), .B(n15135), .Z(n15133) );
  XNOR U15127 ( .A(y[498]), .B(x[498]), .Z(n15135) );
  XNOR U15128 ( .A(y[499]), .B(x[499]), .Z(n15134) );
  AND U15129 ( .A(n15136), .B(n15137), .Z(n15132) );
  XNOR U15130 ( .A(y[500]), .B(x[500]), .Z(n15137) );
  XNOR U15131 ( .A(y[501]), .B(x[501]), .Z(n15136) );
  AND U15132 ( .A(n15138), .B(n15139), .Z(n15122) );
  AND U15133 ( .A(n15140), .B(n15141), .Z(n15139) );
  AND U15134 ( .A(n15142), .B(n15143), .Z(n15141) );
  XNOR U15135 ( .A(y[502]), .B(x[502]), .Z(n15143) );
  XNOR U15136 ( .A(y[503]), .B(x[503]), .Z(n15142) );
  AND U15137 ( .A(n15144), .B(n15145), .Z(n15140) );
  XNOR U15138 ( .A(y[504]), .B(x[504]), .Z(n15145) );
  XNOR U15139 ( .A(y[505]), .B(x[505]), .Z(n15144) );
  AND U15140 ( .A(n15146), .B(n15147), .Z(n15138) );
  AND U15141 ( .A(n15148), .B(n15149), .Z(n15147) );
  XNOR U15142 ( .A(y[506]), .B(x[506]), .Z(n15149) );
  XNOR U15143 ( .A(y[507]), .B(x[507]), .Z(n15148) );
  AND U15144 ( .A(n15150), .B(n15151), .Z(n15146) );
  XNOR U15145 ( .A(y[508]), .B(x[508]), .Z(n15151) );
  XNOR U15146 ( .A(y[509]), .B(x[509]), .Z(n15150) );
  AND U15147 ( .A(n15152), .B(n15153), .Z(n15120) );
  AND U15148 ( .A(n15154), .B(n15155), .Z(n15153) );
  AND U15149 ( .A(n15156), .B(n15157), .Z(n15155) );
  AND U15150 ( .A(n15158), .B(n15159), .Z(n15157) );
  XNOR U15151 ( .A(y[510]), .B(x[510]), .Z(n15159) );
  XNOR U15152 ( .A(y[511]), .B(x[511]), .Z(n15158) );
  AND U15153 ( .A(n15160), .B(n15161), .Z(n15156) );
  XNOR U15154 ( .A(y[512]), .B(x[512]), .Z(n15161) );
  XNOR U15155 ( .A(y[513]), .B(x[513]), .Z(n15160) );
  AND U15156 ( .A(n15162), .B(n15163), .Z(n15154) );
  AND U15157 ( .A(n15164), .B(n15165), .Z(n15163) );
  XNOR U15158 ( .A(y[514]), .B(x[514]), .Z(n15165) );
  XNOR U15159 ( .A(y[515]), .B(x[515]), .Z(n15164) );
  AND U15160 ( .A(n15166), .B(n15167), .Z(n15162) );
  XNOR U15161 ( .A(y[516]), .B(x[516]), .Z(n15167) );
  XNOR U15162 ( .A(y[517]), .B(x[517]), .Z(n15166) );
  AND U15163 ( .A(n15168), .B(n15169), .Z(n15152) );
  AND U15164 ( .A(n15170), .B(n15171), .Z(n15169) );
  AND U15165 ( .A(n15172), .B(n15173), .Z(n15171) );
  XNOR U15166 ( .A(y[518]), .B(x[518]), .Z(n15173) );
  XNOR U15167 ( .A(y[519]), .B(x[519]), .Z(n15172) );
  AND U15168 ( .A(n15174), .B(n15175), .Z(n15170) );
  XNOR U15169 ( .A(y[520]), .B(x[520]), .Z(n15175) );
  XNOR U15170 ( .A(y[521]), .B(x[521]), .Z(n15174) );
  AND U15171 ( .A(n15176), .B(n15177), .Z(n15168) );
  AND U15172 ( .A(n15178), .B(n15179), .Z(n15177) );
  XNOR U15173 ( .A(y[522]), .B(x[522]), .Z(n15179) );
  XNOR U15174 ( .A(y[523]), .B(x[523]), .Z(n15178) );
  AND U15175 ( .A(n15180), .B(n15181), .Z(n15176) );
  XNOR U15176 ( .A(y[524]), .B(x[524]), .Z(n15181) );
  XNOR U15177 ( .A(y[527]), .B(x[527]), .Z(n15180) );
  AND U15178 ( .A(n15182), .B(n15183), .Z(n15054) );
  AND U15179 ( .A(n15184), .B(n15185), .Z(n15183) );
  AND U15180 ( .A(n15186), .B(n15187), .Z(n15185) );
  AND U15181 ( .A(n15188), .B(n15189), .Z(n15187) );
  AND U15182 ( .A(n15190), .B(n15191), .Z(n15189) );
  AND U15183 ( .A(n15192), .B(n15193), .Z(n15191) );
  XNOR U15184 ( .A(y[525]), .B(x[525]), .Z(n15193) );
  XNOR U15185 ( .A(y[526]), .B(x[526]), .Z(n15192) );
  AND U15186 ( .A(n15194), .B(n15195), .Z(n15190) );
  XNOR U15187 ( .A(y[528]), .B(x[528]), .Z(n15195) );
  XNOR U15188 ( .A(y[529]), .B(x[529]), .Z(n15194) );
  AND U15189 ( .A(n15196), .B(n15197), .Z(n15188) );
  AND U15190 ( .A(n15198), .B(n15199), .Z(n15197) );
  XNOR U15191 ( .A(y[530]), .B(x[530]), .Z(n15199) );
  XNOR U15192 ( .A(y[531]), .B(x[531]), .Z(n15198) );
  AND U15193 ( .A(n15200), .B(n15201), .Z(n15196) );
  XNOR U15194 ( .A(y[532]), .B(x[532]), .Z(n15201) );
  XNOR U15195 ( .A(y[533]), .B(x[533]), .Z(n15200) );
  AND U15196 ( .A(n15202), .B(n15203), .Z(n15186) );
  AND U15197 ( .A(n15204), .B(n15205), .Z(n15203) );
  AND U15198 ( .A(n15206), .B(n15207), .Z(n15205) );
  XNOR U15199 ( .A(y[534]), .B(x[534]), .Z(n15207) );
  XNOR U15200 ( .A(y[535]), .B(x[535]), .Z(n15206) );
  AND U15201 ( .A(n15208), .B(n15209), .Z(n15204) );
  XNOR U15202 ( .A(y[536]), .B(x[536]), .Z(n15209) );
  XNOR U15203 ( .A(y[537]), .B(x[537]), .Z(n15208) );
  AND U15204 ( .A(n15210), .B(n15211), .Z(n15202) );
  AND U15205 ( .A(n15212), .B(n15213), .Z(n15211) );
  XNOR U15206 ( .A(y[538]), .B(x[538]), .Z(n15213) );
  XNOR U15207 ( .A(y[539]), .B(x[539]), .Z(n15212) );
  AND U15208 ( .A(n15214), .B(n15215), .Z(n15210) );
  XNOR U15209 ( .A(y[540]), .B(x[540]), .Z(n15215) );
  XNOR U15210 ( .A(y[541]), .B(x[541]), .Z(n15214) );
  AND U15211 ( .A(n15216), .B(n15217), .Z(n15184) );
  AND U15212 ( .A(n15218), .B(n15219), .Z(n15217) );
  AND U15213 ( .A(n15220), .B(n15221), .Z(n15219) );
  AND U15214 ( .A(n15222), .B(n15223), .Z(n15221) );
  XNOR U15215 ( .A(y[542]), .B(x[542]), .Z(n15223) );
  XNOR U15216 ( .A(y[543]), .B(x[543]), .Z(n15222) );
  AND U15217 ( .A(n15224), .B(n15225), .Z(n15220) );
  XNOR U15218 ( .A(y[544]), .B(x[544]), .Z(n15225) );
  XNOR U15219 ( .A(y[545]), .B(x[545]), .Z(n15224) );
  AND U15220 ( .A(n15226), .B(n15227), .Z(n15218) );
  AND U15221 ( .A(n15228), .B(n15229), .Z(n15227) );
  XNOR U15222 ( .A(y[546]), .B(x[546]), .Z(n15229) );
  XNOR U15223 ( .A(y[547]), .B(x[547]), .Z(n15228) );
  AND U15224 ( .A(n15230), .B(n15231), .Z(n15226) );
  XNOR U15225 ( .A(y[548]), .B(x[548]), .Z(n15231) );
  XNOR U15226 ( .A(y[549]), .B(x[549]), .Z(n15230) );
  AND U15227 ( .A(n15232), .B(n15233), .Z(n15216) );
  AND U15228 ( .A(n15234), .B(n15235), .Z(n15233) );
  AND U15229 ( .A(n15236), .B(n15237), .Z(n15235) );
  XNOR U15230 ( .A(y[550]), .B(x[550]), .Z(n15237) );
  XNOR U15231 ( .A(y[551]), .B(x[551]), .Z(n15236) );
  AND U15232 ( .A(n15238), .B(n15239), .Z(n15234) );
  XNOR U15233 ( .A(y[552]), .B(x[552]), .Z(n15239) );
  XNOR U15234 ( .A(y[553]), .B(x[553]), .Z(n15238) );
  AND U15235 ( .A(n15240), .B(n15241), .Z(n15232) );
  AND U15236 ( .A(n15242), .B(n15243), .Z(n15241) );
  XNOR U15237 ( .A(y[554]), .B(x[554]), .Z(n15243) );
  XNOR U15238 ( .A(y[555]), .B(x[555]), .Z(n15242) );
  AND U15239 ( .A(n15244), .B(n15245), .Z(n15240) );
  XNOR U15240 ( .A(y[556]), .B(x[556]), .Z(n15245) );
  XNOR U15241 ( .A(y[557]), .B(x[557]), .Z(n15244) );
  AND U15242 ( .A(n15246), .B(n15247), .Z(n15182) );
  AND U15243 ( .A(n15248), .B(n15249), .Z(n15247) );
  AND U15244 ( .A(n15250), .B(n15251), .Z(n15249) );
  AND U15245 ( .A(n15252), .B(n15253), .Z(n15251) );
  AND U15246 ( .A(n15254), .B(n15255), .Z(n15253) );
  XNOR U15247 ( .A(y[558]), .B(x[558]), .Z(n15255) );
  XNOR U15248 ( .A(y[559]), .B(x[559]), .Z(n15254) );
  AND U15249 ( .A(n15256), .B(n15257), .Z(n15252) );
  XNOR U15250 ( .A(y[560]), .B(x[560]), .Z(n15257) );
  XNOR U15251 ( .A(y[561]), .B(x[561]), .Z(n15256) );
  AND U15252 ( .A(n15258), .B(n15259), .Z(n15250) );
  AND U15253 ( .A(n15260), .B(n15261), .Z(n15259) );
  XNOR U15254 ( .A(y[562]), .B(x[562]), .Z(n15261) );
  XNOR U15255 ( .A(y[563]), .B(x[563]), .Z(n15260) );
  AND U15256 ( .A(n15262), .B(n15263), .Z(n15258) );
  XNOR U15257 ( .A(y[564]), .B(x[564]), .Z(n15263) );
  XNOR U15258 ( .A(y[565]), .B(x[565]), .Z(n15262) );
  AND U15259 ( .A(n15264), .B(n15265), .Z(n15248) );
  AND U15260 ( .A(n15266), .B(n15267), .Z(n15265) );
  AND U15261 ( .A(n15268), .B(n15269), .Z(n15267) );
  XNOR U15262 ( .A(y[566]), .B(x[566]), .Z(n15269) );
  XNOR U15263 ( .A(y[567]), .B(x[567]), .Z(n15268) );
  AND U15264 ( .A(n15270), .B(n15271), .Z(n15266) );
  XNOR U15265 ( .A(y[568]), .B(x[568]), .Z(n15271) );
  XNOR U15266 ( .A(y[569]), .B(x[569]), .Z(n15270) );
  AND U15267 ( .A(n15272), .B(n15273), .Z(n15264) );
  AND U15268 ( .A(n15274), .B(n15275), .Z(n15273) );
  XNOR U15269 ( .A(y[570]), .B(x[570]), .Z(n15275) );
  XNOR U15270 ( .A(y[571]), .B(x[571]), .Z(n15274) );
  AND U15271 ( .A(n15276), .B(n15277), .Z(n15272) );
  XNOR U15272 ( .A(y[572]), .B(x[572]), .Z(n15277) );
  XNOR U15273 ( .A(y[573]), .B(x[573]), .Z(n15276) );
  AND U15274 ( .A(n15278), .B(n15279), .Z(n15246) );
  AND U15275 ( .A(n15280), .B(n15281), .Z(n15279) );
  AND U15276 ( .A(n15282), .B(n15283), .Z(n15281) );
  AND U15277 ( .A(n15284), .B(n15285), .Z(n15283) );
  XNOR U15278 ( .A(y[574]), .B(x[574]), .Z(n15285) );
  XNOR U15279 ( .A(y[575]), .B(x[575]), .Z(n15284) );
  AND U15280 ( .A(n15286), .B(n15287), .Z(n15282) );
  XNOR U15281 ( .A(y[576]), .B(x[576]), .Z(n15287) );
  XNOR U15282 ( .A(y[577]), .B(x[577]), .Z(n15286) );
  AND U15283 ( .A(n15288), .B(n15289), .Z(n15280) );
  AND U15284 ( .A(n15290), .B(n15291), .Z(n15289) );
  XNOR U15285 ( .A(y[578]), .B(x[578]), .Z(n15291) );
  XNOR U15286 ( .A(y[579]), .B(x[579]), .Z(n15290) );
  AND U15287 ( .A(n15292), .B(n15293), .Z(n15288) );
  XNOR U15288 ( .A(y[580]), .B(x[580]), .Z(n15293) );
  XNOR U15289 ( .A(y[581]), .B(x[581]), .Z(n15292) );
  AND U15290 ( .A(n15294), .B(n15295), .Z(n15278) );
  AND U15291 ( .A(n15296), .B(n15297), .Z(n15295) );
  AND U15292 ( .A(n15298), .B(n15299), .Z(n15297) );
  XNOR U15293 ( .A(y[582]), .B(x[582]), .Z(n15299) );
  XNOR U15294 ( .A(y[583]), .B(x[583]), .Z(n15298) );
  AND U15295 ( .A(n15300), .B(n15301), .Z(n15296) );
  XNOR U15296 ( .A(y[584]), .B(x[584]), .Z(n15301) );
  XNOR U15297 ( .A(y[585]), .B(x[585]), .Z(n15300) );
  AND U15298 ( .A(n15302), .B(n15303), .Z(n15294) );
  AND U15299 ( .A(n15304), .B(n15305), .Z(n15303) );
  XNOR U15300 ( .A(y[586]), .B(x[586]), .Z(n15305) );
  XNOR U15301 ( .A(y[587]), .B(x[587]), .Z(n15304) );
  AND U15302 ( .A(n15306), .B(n15307), .Z(n15302) );
  XNOR U15303 ( .A(y[588]), .B(x[588]), .Z(n15307) );
  XNOR U15304 ( .A(y[589]), .B(x[589]), .Z(n15306) );
  AND U15305 ( .A(n15308), .B(n15309), .Z(n15052) );
  AND U15306 ( .A(n15310), .B(n15311), .Z(n15309) );
  AND U15307 ( .A(n15312), .B(n15313), .Z(n15311) );
  AND U15308 ( .A(n15314), .B(n15315), .Z(n15313) );
  AND U15309 ( .A(n15316), .B(n15317), .Z(n15315) );
  AND U15310 ( .A(n15318), .B(n15319), .Z(n15317) );
  AND U15311 ( .A(n15320), .B(n15321), .Z(n15319) );
  XNOR U15312 ( .A(y[590]), .B(x[590]), .Z(n15321) );
  XNOR U15313 ( .A(y[591]), .B(x[591]), .Z(n15320) );
  AND U15314 ( .A(n15322), .B(n15323), .Z(n15318) );
  XNOR U15315 ( .A(y[592]), .B(x[592]), .Z(n15323) );
  XNOR U15316 ( .A(y[593]), .B(x[593]), .Z(n15322) );
  AND U15317 ( .A(n15324), .B(n15325), .Z(n15316) );
  AND U15318 ( .A(n15326), .B(n15327), .Z(n15325) );
  XNOR U15319 ( .A(y[594]), .B(x[594]), .Z(n15327) );
  XNOR U15320 ( .A(y[595]), .B(x[595]), .Z(n15326) );
  AND U15321 ( .A(n15328), .B(n15329), .Z(n15324) );
  XNOR U15322 ( .A(y[596]), .B(x[596]), .Z(n15329) );
  XNOR U15323 ( .A(y[597]), .B(x[597]), .Z(n15328) );
  AND U15324 ( .A(n15330), .B(n15331), .Z(n15314) );
  AND U15325 ( .A(n15332), .B(n15333), .Z(n15331) );
  AND U15326 ( .A(n15334), .B(n15335), .Z(n15333) );
  XNOR U15327 ( .A(y[598]), .B(x[598]), .Z(n15335) );
  XNOR U15328 ( .A(y[599]), .B(x[599]), .Z(n15334) );
  AND U15329 ( .A(n15336), .B(n15337), .Z(n15332) );
  XNOR U15330 ( .A(y[600]), .B(x[600]), .Z(n15337) );
  XNOR U15331 ( .A(y[601]), .B(x[601]), .Z(n15336) );
  AND U15332 ( .A(n15338), .B(n15339), .Z(n15330) );
  AND U15333 ( .A(n15340), .B(n15341), .Z(n15339) );
  XNOR U15334 ( .A(y[602]), .B(x[602]), .Z(n15341) );
  XNOR U15335 ( .A(y[603]), .B(x[603]), .Z(n15340) );
  AND U15336 ( .A(n15342), .B(n15343), .Z(n15338) );
  XNOR U15337 ( .A(y[604]), .B(x[604]), .Z(n15343) );
  XNOR U15338 ( .A(y[605]), .B(x[605]), .Z(n15342) );
  AND U15339 ( .A(n15344), .B(n15345), .Z(n15312) );
  AND U15340 ( .A(n15346), .B(n15347), .Z(n15345) );
  AND U15341 ( .A(n15348), .B(n15349), .Z(n15347) );
  AND U15342 ( .A(n15350), .B(n15351), .Z(n15349) );
  XNOR U15343 ( .A(y[606]), .B(x[606]), .Z(n15351) );
  XNOR U15344 ( .A(y[607]), .B(x[607]), .Z(n15350) );
  AND U15345 ( .A(n15352), .B(n15353), .Z(n15348) );
  XNOR U15346 ( .A(y[608]), .B(x[608]), .Z(n15353) );
  XNOR U15347 ( .A(y[609]), .B(x[609]), .Z(n15352) );
  AND U15348 ( .A(n15354), .B(n15355), .Z(n15346) );
  AND U15349 ( .A(n15356), .B(n15357), .Z(n15355) );
  XNOR U15350 ( .A(y[610]), .B(x[610]), .Z(n15357) );
  XNOR U15351 ( .A(y[611]), .B(x[611]), .Z(n15356) );
  AND U15352 ( .A(n15358), .B(n15359), .Z(n15354) );
  XNOR U15353 ( .A(y[612]), .B(x[612]), .Z(n15359) );
  XNOR U15354 ( .A(y[613]), .B(x[613]), .Z(n15358) );
  AND U15355 ( .A(n15360), .B(n15361), .Z(n15344) );
  AND U15356 ( .A(n15362), .B(n15363), .Z(n15361) );
  AND U15357 ( .A(n15364), .B(n15365), .Z(n15363) );
  XNOR U15358 ( .A(y[614]), .B(x[614]), .Z(n15365) );
  XNOR U15359 ( .A(y[615]), .B(x[615]), .Z(n15364) );
  AND U15360 ( .A(n15366), .B(n15367), .Z(n15362) );
  XNOR U15361 ( .A(y[616]), .B(x[616]), .Z(n15367) );
  XNOR U15362 ( .A(y[617]), .B(x[617]), .Z(n15366) );
  AND U15363 ( .A(n15368), .B(n15369), .Z(n15360) );
  AND U15364 ( .A(n15370), .B(n15371), .Z(n15369) );
  XNOR U15365 ( .A(y[618]), .B(x[618]), .Z(n15371) );
  XNOR U15366 ( .A(y[619]), .B(x[619]), .Z(n15370) );
  AND U15367 ( .A(n15372), .B(n15373), .Z(n15368) );
  XNOR U15368 ( .A(y[620]), .B(x[620]), .Z(n15373) );
  XNOR U15369 ( .A(y[621]), .B(x[621]), .Z(n15372) );
  AND U15370 ( .A(n15374), .B(n15375), .Z(n15310) );
  AND U15371 ( .A(n15376), .B(n15377), .Z(n15375) );
  AND U15372 ( .A(n15378), .B(n15379), .Z(n15377) );
  AND U15373 ( .A(n15380), .B(n15381), .Z(n15379) );
  AND U15374 ( .A(n15382), .B(n15383), .Z(n15381) );
  XNOR U15375 ( .A(y[622]), .B(x[622]), .Z(n15383) );
  XNOR U15376 ( .A(y[623]), .B(x[623]), .Z(n15382) );
  AND U15377 ( .A(n15384), .B(n15385), .Z(n15380) );
  XNOR U15378 ( .A(y[624]), .B(x[624]), .Z(n15385) );
  XNOR U15379 ( .A(y[625]), .B(x[625]), .Z(n15384) );
  AND U15380 ( .A(n15386), .B(n15387), .Z(n15378) );
  AND U15381 ( .A(n15388), .B(n15389), .Z(n15387) );
  XNOR U15382 ( .A(y[626]), .B(x[626]), .Z(n15389) );
  XNOR U15383 ( .A(y[627]), .B(x[627]), .Z(n15388) );
  AND U15384 ( .A(n15390), .B(n15391), .Z(n15386) );
  XNOR U15385 ( .A(y[628]), .B(x[628]), .Z(n15391) );
  XNOR U15386 ( .A(y[629]), .B(x[629]), .Z(n15390) );
  AND U15387 ( .A(n15392), .B(n15393), .Z(n15376) );
  AND U15388 ( .A(n15394), .B(n15395), .Z(n15393) );
  AND U15389 ( .A(n15396), .B(n15397), .Z(n15395) );
  XNOR U15390 ( .A(y[630]), .B(x[630]), .Z(n15397) );
  XNOR U15391 ( .A(y[631]), .B(x[631]), .Z(n15396) );
  AND U15392 ( .A(n15398), .B(n15399), .Z(n15394) );
  XNOR U15393 ( .A(y[632]), .B(x[632]), .Z(n15399) );
  XNOR U15394 ( .A(y[633]), .B(x[633]), .Z(n15398) );
  AND U15395 ( .A(n15400), .B(n15401), .Z(n15392) );
  AND U15396 ( .A(n15402), .B(n15403), .Z(n15401) );
  XNOR U15397 ( .A(y[634]), .B(x[634]), .Z(n15403) );
  XNOR U15398 ( .A(y[635]), .B(x[635]), .Z(n15402) );
  AND U15399 ( .A(n15404), .B(n15405), .Z(n15400) );
  XNOR U15400 ( .A(y[636]), .B(x[636]), .Z(n15405) );
  XNOR U15401 ( .A(y[637]), .B(x[637]), .Z(n15404) );
  AND U15402 ( .A(n15406), .B(n15407), .Z(n15374) );
  AND U15403 ( .A(n15408), .B(n15409), .Z(n15407) );
  AND U15404 ( .A(n15410), .B(n15411), .Z(n15409) );
  AND U15405 ( .A(n15412), .B(n15413), .Z(n15411) );
  XNOR U15406 ( .A(y[638]), .B(x[638]), .Z(n15413) );
  XNOR U15407 ( .A(y[639]), .B(x[639]), .Z(n15412) );
  AND U15408 ( .A(n15414), .B(n15415), .Z(n15410) );
  XNOR U15409 ( .A(y[640]), .B(x[640]), .Z(n15415) );
  XNOR U15410 ( .A(y[641]), .B(x[641]), .Z(n15414) );
  AND U15411 ( .A(n15416), .B(n15417), .Z(n15408) );
  AND U15412 ( .A(n15418), .B(n15419), .Z(n15417) );
  XNOR U15413 ( .A(y[642]), .B(x[642]), .Z(n15419) );
  XNOR U15414 ( .A(y[643]), .B(x[643]), .Z(n15418) );
  AND U15415 ( .A(n15420), .B(n15421), .Z(n15416) );
  XNOR U15416 ( .A(y[644]), .B(x[644]), .Z(n15421) );
  XNOR U15417 ( .A(y[645]), .B(x[645]), .Z(n15420) );
  AND U15418 ( .A(n15422), .B(n15423), .Z(n15406) );
  AND U15419 ( .A(n15424), .B(n15425), .Z(n15423) );
  AND U15420 ( .A(n15426), .B(n15427), .Z(n15425) );
  XNOR U15421 ( .A(y[646]), .B(x[646]), .Z(n15427) );
  XNOR U15422 ( .A(y[647]), .B(x[647]), .Z(n15426) );
  AND U15423 ( .A(n15428), .B(n15429), .Z(n15424) );
  XNOR U15424 ( .A(y[648]), .B(x[648]), .Z(n15429) );
  XNOR U15425 ( .A(y[649]), .B(x[649]), .Z(n15428) );
  AND U15426 ( .A(n15430), .B(n15431), .Z(n15422) );
  AND U15427 ( .A(n15432), .B(n15433), .Z(n15431) );
  XNOR U15428 ( .A(y[650]), .B(x[650]), .Z(n15433) );
  XNOR U15429 ( .A(y[651]), .B(x[651]), .Z(n15432) );
  AND U15430 ( .A(n15434), .B(n15435), .Z(n15430) );
  XNOR U15431 ( .A(y[652]), .B(x[652]), .Z(n15435) );
  XNOR U15432 ( .A(y[653]), .B(x[653]), .Z(n15434) );
  AND U15433 ( .A(n15436), .B(n15437), .Z(n15308) );
  AND U15434 ( .A(n15438), .B(n15439), .Z(n15437) );
  AND U15435 ( .A(n15440), .B(n15441), .Z(n15439) );
  AND U15436 ( .A(n15442), .B(n15443), .Z(n15441) );
  AND U15437 ( .A(n15444), .B(n15445), .Z(n15443) );
  AND U15438 ( .A(n15446), .B(n15447), .Z(n15445) );
  XNOR U15439 ( .A(y[654]), .B(x[654]), .Z(n15447) );
  XNOR U15440 ( .A(y[655]), .B(x[655]), .Z(n15446) );
  AND U15441 ( .A(n15448), .B(n15449), .Z(n15444) );
  XNOR U15442 ( .A(y[656]), .B(x[656]), .Z(n15449) );
  XNOR U15443 ( .A(y[657]), .B(x[657]), .Z(n15448) );
  AND U15444 ( .A(n15450), .B(n15451), .Z(n15442) );
  AND U15445 ( .A(n15452), .B(n15453), .Z(n15451) );
  XNOR U15446 ( .A(y[658]), .B(x[658]), .Z(n15453) );
  XNOR U15447 ( .A(y[659]), .B(x[659]), .Z(n15452) );
  AND U15448 ( .A(n15454), .B(n15455), .Z(n15450) );
  XNOR U15449 ( .A(y[660]), .B(x[660]), .Z(n15455) );
  XNOR U15450 ( .A(y[661]), .B(x[661]), .Z(n15454) );
  AND U15451 ( .A(n15456), .B(n15457), .Z(n15440) );
  AND U15452 ( .A(n15458), .B(n15459), .Z(n15457) );
  AND U15453 ( .A(n15460), .B(n15461), .Z(n15459) );
  XNOR U15454 ( .A(y[662]), .B(x[662]), .Z(n15461) );
  XNOR U15455 ( .A(y[663]), .B(x[663]), .Z(n15460) );
  AND U15456 ( .A(n15462), .B(n15463), .Z(n15458) );
  XNOR U15457 ( .A(y[664]), .B(x[664]), .Z(n15463) );
  XNOR U15458 ( .A(y[665]), .B(x[665]), .Z(n15462) );
  AND U15459 ( .A(n15464), .B(n15465), .Z(n15456) );
  AND U15460 ( .A(n15466), .B(n15467), .Z(n15465) );
  XNOR U15461 ( .A(y[666]), .B(x[666]), .Z(n15467) );
  XNOR U15462 ( .A(y[667]), .B(x[667]), .Z(n15466) );
  AND U15463 ( .A(n15468), .B(n15469), .Z(n15464) );
  XNOR U15464 ( .A(y[668]), .B(x[668]), .Z(n15469) );
  XNOR U15465 ( .A(y[669]), .B(x[669]), .Z(n15468) );
  AND U15466 ( .A(n15470), .B(n15471), .Z(n15438) );
  AND U15467 ( .A(n15472), .B(n15473), .Z(n15471) );
  AND U15468 ( .A(n15474), .B(n15475), .Z(n15473) );
  AND U15469 ( .A(n15476), .B(n15477), .Z(n15475) );
  XNOR U15470 ( .A(y[670]), .B(x[670]), .Z(n15477) );
  XNOR U15471 ( .A(y[671]), .B(x[671]), .Z(n15476) );
  AND U15472 ( .A(n15478), .B(n15479), .Z(n15474) );
  XNOR U15473 ( .A(y[672]), .B(x[672]), .Z(n15479) );
  XNOR U15474 ( .A(y[673]), .B(x[673]), .Z(n15478) );
  AND U15475 ( .A(n15480), .B(n15481), .Z(n15472) );
  AND U15476 ( .A(n15482), .B(n15483), .Z(n15481) );
  XNOR U15477 ( .A(y[674]), .B(x[674]), .Z(n15483) );
  XNOR U15478 ( .A(y[675]), .B(x[675]), .Z(n15482) );
  AND U15479 ( .A(n15484), .B(n15485), .Z(n15480) );
  XNOR U15480 ( .A(y[676]), .B(x[676]), .Z(n15485) );
  XNOR U15481 ( .A(y[677]), .B(x[677]), .Z(n15484) );
  AND U15482 ( .A(n15486), .B(n15487), .Z(n15470) );
  AND U15483 ( .A(n15488), .B(n15489), .Z(n15487) );
  AND U15484 ( .A(n15490), .B(n15491), .Z(n15489) );
  XNOR U15485 ( .A(y[678]), .B(x[678]), .Z(n15491) );
  XNOR U15486 ( .A(y[679]), .B(x[679]), .Z(n15490) );
  AND U15487 ( .A(n15492), .B(n15493), .Z(n15488) );
  XNOR U15488 ( .A(y[680]), .B(x[680]), .Z(n15493) );
  XNOR U15489 ( .A(y[681]), .B(x[681]), .Z(n15492) );
  AND U15490 ( .A(n15494), .B(n15495), .Z(n15486) );
  AND U15491 ( .A(n15496), .B(n15497), .Z(n15495) );
  XNOR U15492 ( .A(y[682]), .B(x[682]), .Z(n15497) );
  XNOR U15493 ( .A(y[683]), .B(x[683]), .Z(n15496) );
  AND U15494 ( .A(n15498), .B(n15499), .Z(n15494) );
  XNOR U15495 ( .A(y[684]), .B(x[684]), .Z(n15499) );
  XNOR U15496 ( .A(y[685]), .B(x[685]), .Z(n15498) );
  AND U15497 ( .A(n15500), .B(n15501), .Z(n15436) );
  AND U15498 ( .A(n15502), .B(n15503), .Z(n15501) );
  AND U15499 ( .A(n15504), .B(n15505), .Z(n15503) );
  AND U15500 ( .A(n15506), .B(n15507), .Z(n15505) );
  AND U15501 ( .A(n15508), .B(n15509), .Z(n15507) );
  XNOR U15502 ( .A(y[686]), .B(x[686]), .Z(n15509) );
  XNOR U15503 ( .A(y[687]), .B(x[687]), .Z(n15508) );
  AND U15504 ( .A(n15510), .B(n15511), .Z(n15506) );
  XNOR U15505 ( .A(y[688]), .B(x[688]), .Z(n15511) );
  XNOR U15506 ( .A(y[689]), .B(x[689]), .Z(n15510) );
  AND U15507 ( .A(n15512), .B(n15513), .Z(n15504) );
  AND U15508 ( .A(n15514), .B(n15515), .Z(n15513) );
  XNOR U15509 ( .A(y[690]), .B(x[690]), .Z(n15515) );
  XNOR U15510 ( .A(y[691]), .B(x[691]), .Z(n15514) );
  AND U15511 ( .A(n15516), .B(n15517), .Z(n15512) );
  XNOR U15512 ( .A(y[692]), .B(x[692]), .Z(n15517) );
  XNOR U15513 ( .A(y[693]), .B(x[693]), .Z(n15516) );
  AND U15514 ( .A(n15518), .B(n15519), .Z(n15502) );
  AND U15515 ( .A(n15520), .B(n15521), .Z(n15519) );
  AND U15516 ( .A(n15522), .B(n15523), .Z(n15521) );
  XNOR U15517 ( .A(y[694]), .B(x[694]), .Z(n15523) );
  XNOR U15518 ( .A(y[695]), .B(x[695]), .Z(n15522) );
  AND U15519 ( .A(n15524), .B(n15525), .Z(n15520) );
  XNOR U15520 ( .A(y[696]), .B(x[696]), .Z(n15525) );
  XNOR U15521 ( .A(y[697]), .B(x[697]), .Z(n15524) );
  AND U15522 ( .A(n15526), .B(n15527), .Z(n15518) );
  AND U15523 ( .A(n15528), .B(n15529), .Z(n15527) );
  XNOR U15524 ( .A(y[698]), .B(x[698]), .Z(n15529) );
  XNOR U15525 ( .A(y[699]), .B(x[699]), .Z(n15528) );
  AND U15526 ( .A(n15530), .B(n15531), .Z(n15526) );
  XNOR U15527 ( .A(y[700]), .B(x[700]), .Z(n15531) );
  XNOR U15528 ( .A(y[701]), .B(x[701]), .Z(n15530) );
  AND U15529 ( .A(n15532), .B(n15533), .Z(n15500) );
  AND U15530 ( .A(n15534), .B(n15535), .Z(n15533) );
  AND U15531 ( .A(n15536), .B(n15537), .Z(n15535) );
  AND U15532 ( .A(n15538), .B(n15539), .Z(n15537) );
  XNOR U15533 ( .A(y[702]), .B(x[702]), .Z(n15539) );
  XNOR U15534 ( .A(y[703]), .B(x[703]), .Z(n15538) );
  AND U15535 ( .A(n15540), .B(n15541), .Z(n15536) );
  XNOR U15536 ( .A(y[704]), .B(x[704]), .Z(n15541) );
  XNOR U15537 ( .A(y[705]), .B(x[705]), .Z(n15540) );
  AND U15538 ( .A(n15542), .B(n15543), .Z(n15534) );
  AND U15539 ( .A(n15544), .B(n15545), .Z(n15543) );
  XNOR U15540 ( .A(y[706]), .B(x[706]), .Z(n15545) );
  XNOR U15541 ( .A(y[707]), .B(x[707]), .Z(n15544) );
  AND U15542 ( .A(n15546), .B(n15547), .Z(n15542) );
  XNOR U15543 ( .A(y[708]), .B(x[708]), .Z(n15547) );
  XNOR U15544 ( .A(y[709]), .B(x[709]), .Z(n15546) );
  AND U15545 ( .A(n15548), .B(n15549), .Z(n15532) );
  AND U15546 ( .A(n15550), .B(n15551), .Z(n15549) );
  AND U15547 ( .A(n15552), .B(n15553), .Z(n15551) );
  XNOR U15548 ( .A(y[710]), .B(x[710]), .Z(n15553) );
  XNOR U15549 ( .A(y[711]), .B(x[711]), .Z(n15552) );
  AND U15550 ( .A(n15554), .B(n15555), .Z(n15550) );
  XNOR U15551 ( .A(y[712]), .B(x[712]), .Z(n15555) );
  XNOR U15552 ( .A(y[713]), .B(x[713]), .Z(n15554) );
  AND U15553 ( .A(n15556), .B(n15557), .Z(n15548) );
  AND U15554 ( .A(n15558), .B(n15559), .Z(n15557) );
  XNOR U15555 ( .A(y[714]), .B(x[714]), .Z(n15559) );
  XNOR U15556 ( .A(y[715]), .B(x[715]), .Z(n15558) );
  AND U15557 ( .A(n15560), .B(n15561), .Z(n15556) );
  XNOR U15558 ( .A(y[716]), .B(x[716]), .Z(n15561) );
  XNOR U15559 ( .A(y[717]), .B(x[717]), .Z(n15560) );
  XNOR U15560 ( .A(y[350]), .B(x[350]), .Z(n15050) );
  AND U15561 ( .A(n15562), .B(n15563), .Z(n8212) );
  XNOR U15562 ( .A(y[353]), .B(x[353]), .Z(n15563) );
  AND U15563 ( .A(n15564), .B(n15565), .Z(n15562) );
  XNOR U15564 ( .A(y[351]), .B(x[351]), .Z(n15565) );
  XNOR U15565 ( .A(y[352]), .B(x[352]), .Z(n15564) );
  AND U15566 ( .A(n15566), .B(n15567), .Z(n8210) );
  AND U15567 ( .A(n15568), .B(n15569), .Z(n15567) );
  AND U15568 ( .A(n15570), .B(n15571), .Z(n15569) );
  XNOR U15569 ( .A(y[356]), .B(x[356]), .Z(n15571) );
  XNOR U15570 ( .A(y[354]), .B(x[354]), .Z(n15570) );
  AND U15571 ( .A(n15572), .B(n15573), .Z(n15568) );
  XNOR U15572 ( .A(y[355]), .B(x[355]), .Z(n15573) );
  XNOR U15573 ( .A(y[359]), .B(x[359]), .Z(n15572) );
  AND U15574 ( .A(n15574), .B(n15575), .Z(n15566) );
  XNOR U15575 ( .A(y[362]), .B(x[362]), .Z(n15575) );
  AND U15576 ( .A(n15576), .B(n15577), .Z(n15574) );
  XNOR U15577 ( .A(y[357]), .B(x[357]), .Z(n15577) );
  XNOR U15578 ( .A(y[358]), .B(x[358]), .Z(n15576) );
  AND U15579 ( .A(n15578), .B(n15579), .Z(n8208) );
  AND U15580 ( .A(n15580), .B(n15581), .Z(n15579) );
  AND U15581 ( .A(n15582), .B(n15583), .Z(n15581) );
  AND U15582 ( .A(n15584), .B(n15585), .Z(n15583) );
  XNOR U15583 ( .A(y[360]), .B(x[360]), .Z(n15585) );
  XNOR U15584 ( .A(y[361]), .B(x[361]), .Z(n15584) );
  AND U15585 ( .A(n15586), .B(n15587), .Z(n15582) );
  XNOR U15586 ( .A(y[365]), .B(x[365]), .Z(n15587) );
  XNOR U15587 ( .A(y[363]), .B(x[363]), .Z(n15586) );
  AND U15588 ( .A(n15588), .B(n15589), .Z(n15580) );
  XNOR U15589 ( .A(y[366]), .B(x[366]), .Z(n15589) );
  AND U15590 ( .A(n15590), .B(n15591), .Z(n15588) );
  XNOR U15591 ( .A(y[364]), .B(x[364]), .Z(n15591) );
  XNOR U15592 ( .A(y[368]), .B(x[368]), .Z(n15590) );
  AND U15593 ( .A(n15592), .B(n15593), .Z(n15578) );
  AND U15594 ( .A(n15594), .B(n15595), .Z(n15593) );
  XNOR U15595 ( .A(y[369]), .B(x[369]), .Z(n15595) );
  AND U15596 ( .A(n15596), .B(n15597), .Z(n15594) );
  XNOR U15597 ( .A(y[367]), .B(x[367]), .Z(n15597) );
  XNOR U15598 ( .A(y[371]), .B(x[371]), .Z(n15596) );
  AND U15599 ( .A(n15598), .B(n15599), .Z(n15592) );
  XNOR U15600 ( .A(y[372]), .B(x[372]), .Z(n15599) );
  AND U15601 ( .A(n15600), .B(n15601), .Z(n15598) );
  XNOR U15602 ( .A(y[370]), .B(x[370]), .Z(n15601) );
  XNOR U15603 ( .A(y[374]), .B(x[374]), .Z(n15600) );
  AND U15604 ( .A(n15602), .B(n15603), .Z(n8206) );
  AND U15605 ( .A(n15604), .B(n15605), .Z(n15603) );
  AND U15606 ( .A(n15606), .B(n15607), .Z(n15605) );
  AND U15607 ( .A(n15608), .B(n15609), .Z(n15607) );
  AND U15608 ( .A(n15610), .B(n15611), .Z(n15609) );
  XNOR U15609 ( .A(y[373]), .B(x[373]), .Z(n15611) );
  XNOR U15610 ( .A(y[300]), .B(x[300]), .Z(n15610) );
  AND U15611 ( .A(n15612), .B(n15613), .Z(n15608) );
  XNOR U15612 ( .A(y[301]), .B(x[301]), .Z(n15613) );
  XNOR U15613 ( .A(y[302]), .B(x[302]), .Z(n15612) );
  AND U15614 ( .A(n15614), .B(n15615), .Z(n15606) );
  XNOR U15615 ( .A(y[304]), .B(x[304]), .Z(n15615) );
  AND U15616 ( .A(n15616), .B(n15617), .Z(n15614) );
  XNOR U15617 ( .A(y[303]), .B(x[303]), .Z(n15617) );
  XNOR U15618 ( .A(y[306]), .B(x[306]), .Z(n15616) );
  AND U15619 ( .A(n15618), .B(n15619), .Z(n15604) );
  AND U15620 ( .A(n15620), .B(n15621), .Z(n15619) );
  AND U15621 ( .A(n15622), .B(n15623), .Z(n15621) );
  XNOR U15622 ( .A(y[305]), .B(x[305]), .Z(n15623) );
  XNOR U15623 ( .A(y[309]), .B(x[309]), .Z(n15622) );
  AND U15624 ( .A(n15624), .B(n15625), .Z(n15620) );
  XNOR U15625 ( .A(y[307]), .B(x[307]), .Z(n15625) );
  XNOR U15626 ( .A(y[308]), .B(x[308]), .Z(n15624) );
  AND U15627 ( .A(n15626), .B(n15627), .Z(n15618) );
  XNOR U15628 ( .A(y[311]), .B(x[311]), .Z(n15627) );
  AND U15629 ( .A(n15628), .B(n15629), .Z(n15626) );
  XNOR U15630 ( .A(y[312]), .B(x[312]), .Z(n15629) );
  XNOR U15631 ( .A(y[310]), .B(x[310]), .Z(n15628) );
  AND U15632 ( .A(n15630), .B(n15631), .Z(n15602) );
  AND U15633 ( .A(n15632), .B(n15633), .Z(n15631) );
  AND U15634 ( .A(n15634), .B(n15635), .Z(n15633) );
  AND U15635 ( .A(n15636), .B(n15637), .Z(n15635) );
  XNOR U15636 ( .A(y[315]), .B(x[315]), .Z(n15637) );
  XNOR U15637 ( .A(y[313]), .B(x[313]), .Z(n15636) );
  AND U15638 ( .A(n15638), .B(n15639), .Z(n15634) );
  XNOR U15639 ( .A(y[314]), .B(x[314]), .Z(n15639) );
  XNOR U15640 ( .A(y[318]), .B(x[318]), .Z(n15638) );
  AND U15641 ( .A(n15640), .B(n15641), .Z(n15632) );
  XNOR U15642 ( .A(y[321]), .B(x[321]), .Z(n15641) );
  AND U15643 ( .A(n15642), .B(n15643), .Z(n15640) );
  XNOR U15644 ( .A(y[316]), .B(x[316]), .Z(n15643) );
  XNOR U15645 ( .A(y[317]), .B(x[317]), .Z(n15642) );
  AND U15646 ( .A(n15644), .B(n15645), .Z(n15630) );
  AND U15647 ( .A(n15646), .B(n15647), .Z(n15645) );
  XNOR U15648 ( .A(y[324]), .B(x[324]), .Z(n15647) );
  AND U15649 ( .A(n15648), .B(n15649), .Z(n15646) );
  XNOR U15650 ( .A(y[319]), .B(x[319]), .Z(n15649) );
  XNOR U15651 ( .A(y[320]), .B(x[320]), .Z(n15648) );
  AND U15652 ( .A(n15650), .B(n15651), .Z(n15644) );
  XNOR U15653 ( .A(y[325]), .B(x[325]), .Z(n15651) );
  AND U15654 ( .A(n15652), .B(n15653), .Z(n15650) );
  XNOR U15655 ( .A(y[322]), .B(x[322]), .Z(n15653) );
  XNOR U15656 ( .A(y[323]), .B(x[323]), .Z(n15652) );
  AND U15657 ( .A(n15654), .B(n15655), .Z(n8204) );
  AND U15658 ( .A(n15656), .B(n15657), .Z(n15655) );
  AND U15659 ( .A(n15658), .B(n15659), .Z(n15657) );
  AND U15660 ( .A(n15660), .B(n15661), .Z(n15659) );
  AND U15661 ( .A(n15662), .B(n15663), .Z(n15661) );
  AND U15662 ( .A(n15664), .B(n15665), .Z(n15663) );
  XNOR U15663 ( .A(y[326]), .B(x[326]), .Z(n15665) );
  XNOR U15664 ( .A(y[327]), .B(x[327]), .Z(n15664) );
  AND U15665 ( .A(n15666), .B(n15667), .Z(n15662) );
  XNOR U15666 ( .A(y[328]), .B(x[328]), .Z(n15667) );
  XNOR U15667 ( .A(y[331]), .B(x[331]), .Z(n15666) );
  AND U15668 ( .A(n15668), .B(n15669), .Z(n15660) );
  XNOR U15669 ( .A(y[334]), .B(x[334]), .Z(n15669) );
  AND U15670 ( .A(n15670), .B(n15671), .Z(n15668) );
  XNOR U15671 ( .A(y[329]), .B(x[329]), .Z(n15671) );
  XNOR U15672 ( .A(y[330]), .B(x[330]), .Z(n15670) );
  AND U15673 ( .A(n15672), .B(n15673), .Z(n15658) );
  AND U15674 ( .A(n15674), .B(n15675), .Z(n15673) );
  AND U15675 ( .A(n15676), .B(n15677), .Z(n15675) );
  XNOR U15676 ( .A(y[332]), .B(x[332]), .Z(n15677) );
  XNOR U15677 ( .A(y[333]), .B(x[333]), .Z(n15676) );
  AND U15678 ( .A(n15678), .B(n15679), .Z(n15674) );
  XNOR U15679 ( .A(y[337]), .B(x[337]), .Z(n15679) );
  XNOR U15680 ( .A(y[335]), .B(x[335]), .Z(n15678) );
  AND U15681 ( .A(n15680), .B(n15681), .Z(n15672) );
  XNOR U15682 ( .A(y[338]), .B(x[338]), .Z(n15681) );
  AND U15683 ( .A(n15682), .B(n15683), .Z(n15680) );
  XNOR U15684 ( .A(y[336]), .B(x[336]), .Z(n15683) );
  XNOR U15685 ( .A(y[340]), .B(x[340]), .Z(n15682) );
  AND U15686 ( .A(n15684), .B(n15685), .Z(n15656) );
  AND U15687 ( .A(n15686), .B(n15687), .Z(n15685) );
  AND U15688 ( .A(n15688), .B(n15689), .Z(n15687) );
  AND U15689 ( .A(n15690), .B(n15691), .Z(n15689) );
  XNOR U15690 ( .A(y[339]), .B(x[339]), .Z(n15691) );
  XNOR U15691 ( .A(y[343]), .B(x[343]), .Z(n15690) );
  AND U15692 ( .A(n15692), .B(n15693), .Z(n15688) );
  XNOR U15693 ( .A(y[341]), .B(x[341]), .Z(n15693) );
  XNOR U15694 ( .A(y[342]), .B(x[342]), .Z(n15692) );
  AND U15695 ( .A(n15694), .B(n15695), .Z(n15686) );
  XNOR U15696 ( .A(y[345]), .B(x[345]), .Z(n15695) );
  AND U15697 ( .A(n15696), .B(n15697), .Z(n15694) );
  XNOR U15698 ( .A(y[346]), .B(x[346]), .Z(n15697) );
  XNOR U15699 ( .A(y[344]), .B(x[344]), .Z(n15696) );
  AND U15700 ( .A(n15698), .B(n15699), .Z(n15684) );
  AND U15701 ( .A(n15700), .B(n15701), .Z(n15699) );
  XNOR U15702 ( .A(y[348]), .B(x[348]), .Z(n15701) );
  AND U15703 ( .A(n15702), .B(n15703), .Z(n15700) );
  XNOR U15704 ( .A(y[349]), .B(x[349]), .Z(n15703) );
  XNOR U15705 ( .A(y[347]), .B(x[347]), .Z(n15702) );
  AND U15706 ( .A(n15704), .B(n15705), .Z(n15698) );
  XNOR U15707 ( .A(y[202]), .B(x[202]), .Z(n15705) );
  AND U15708 ( .A(n15706), .B(n15707), .Z(n15704) );
  XNOR U15709 ( .A(y[200]), .B(x[200]), .Z(n15707) );
  XNOR U15710 ( .A(y[201]), .B(x[201]), .Z(n15706) );
  AND U15711 ( .A(n15708), .B(n15709), .Z(n15654) );
  AND U15712 ( .A(n15710), .B(n15711), .Z(n15709) );
  AND U15713 ( .A(n15712), .B(n15713), .Z(n15711) );
  AND U15714 ( .A(n15714), .B(n15715), .Z(n15713) );
  AND U15715 ( .A(n15716), .B(n15717), .Z(n15715) );
  XNOR U15716 ( .A(y[203]), .B(x[203]), .Z(n15717) );
  XNOR U15717 ( .A(y[206]), .B(x[206]), .Z(n15716) );
  AND U15718 ( .A(n15718), .B(n15719), .Z(n15714) );
  XNOR U15719 ( .A(y[204]), .B(x[204]), .Z(n15719) );
  XNOR U15720 ( .A(y[205]), .B(x[205]), .Z(n15718) );
  AND U15721 ( .A(n15720), .B(n15721), .Z(n15712) );
  XNOR U15722 ( .A(y[208]), .B(x[208]), .Z(n15721) );
  AND U15723 ( .A(n15722), .B(n15723), .Z(n15720) );
  XNOR U15724 ( .A(y[209]), .B(x[209]), .Z(n15723) );
  XNOR U15725 ( .A(y[207]), .B(x[207]), .Z(n15722) );
  AND U15726 ( .A(n15724), .B(n15725), .Z(n15710) );
  AND U15727 ( .A(n15726), .B(n15727), .Z(n15725) );
  XNOR U15728 ( .A(y[211]), .B(x[211]), .Z(n15727) );
  AND U15729 ( .A(n15728), .B(n15729), .Z(n15726) );
  XNOR U15730 ( .A(y[212]), .B(x[212]), .Z(n15729) );
  XNOR U15731 ( .A(y[210]), .B(x[210]), .Z(n15728) );
  AND U15732 ( .A(n15730), .B(n15731), .Z(n15724) );
  XNOR U15733 ( .A(y[214]), .B(x[214]), .Z(n15731) );
  AND U15734 ( .A(n15732), .B(n15733), .Z(n15730) );
  XNOR U15735 ( .A(y[215]), .B(x[215]), .Z(n15733) );
  XNOR U15736 ( .A(y[213]), .B(x[213]), .Z(n15732) );
  AND U15737 ( .A(n15734), .B(n15735), .Z(n15708) );
  AND U15738 ( .A(n15736), .B(n15737), .Z(n15735) );
  AND U15739 ( .A(n15738), .B(n15739), .Z(n15737) );
  AND U15740 ( .A(n15740), .B(n15741), .Z(n15739) );
  XNOR U15741 ( .A(y[218]), .B(x[218]), .Z(n15741) );
  XNOR U15742 ( .A(y[216]), .B(x[216]), .Z(n15740) );
  AND U15743 ( .A(n15742), .B(n15743), .Z(n15738) );
  XNOR U15744 ( .A(y[217]), .B(x[217]), .Z(n15743) );
  XNOR U15745 ( .A(y[221]), .B(x[221]), .Z(n15742) );
  AND U15746 ( .A(n15744), .B(n15745), .Z(n15736) );
  XNOR U15747 ( .A(y[224]), .B(x[224]), .Z(n15745) );
  AND U15748 ( .A(n15746), .B(n15747), .Z(n15744) );
  XNOR U15749 ( .A(y[219]), .B(x[219]), .Z(n15747) );
  XNOR U15750 ( .A(y[220]), .B(x[220]), .Z(n15746) );
  AND U15751 ( .A(n15748), .B(n15749), .Z(n15734) );
  AND U15752 ( .A(n15750), .B(n15751), .Z(n15749) );
  XNOR U15753 ( .A(y[225]), .B(x[225]), .Z(n15751) );
  AND U15754 ( .A(n15752), .B(n15753), .Z(n15750) );
  XNOR U15755 ( .A(y[222]), .B(x[222]), .Z(n15753) );
  XNOR U15756 ( .A(y[223]), .B(x[223]), .Z(n15752) );
  AND U15757 ( .A(n15754), .B(n15755), .Z(n15748) );
  XNOR U15758 ( .A(y[228]), .B(x[228]), .Z(n15755) );
  AND U15759 ( .A(n15756), .B(n15757), .Z(n15754) );
  XNOR U15760 ( .A(y[226]), .B(x[226]), .Z(n15757) );
  XNOR U15761 ( .A(y[227]), .B(x[227]), .Z(n15756) );
  AND U15762 ( .A(n15758), .B(n15759), .Z(n8202) );
  AND U15763 ( .A(n15760), .B(n15761), .Z(n15759) );
  AND U15764 ( .A(n15762), .B(n15763), .Z(n15761) );
  AND U15765 ( .A(n15764), .B(n15765), .Z(n15763) );
  AND U15766 ( .A(n15766), .B(n15767), .Z(n15765) );
  AND U15767 ( .A(n15768), .B(n15769), .Z(n15767) );
  AND U15768 ( .A(n15770), .B(n15771), .Z(n15769) );
  XNOR U15769 ( .A(y[231]), .B(x[231]), .Z(n15771) );
  XNOR U15770 ( .A(y[229]), .B(x[229]), .Z(n15770) );
  AND U15771 ( .A(n15772), .B(n15773), .Z(n15768) );
  XNOR U15772 ( .A(y[230]), .B(x[230]), .Z(n15773) );
  XNOR U15773 ( .A(y[234]), .B(x[234]), .Z(n15772) );
  AND U15774 ( .A(n15774), .B(n15775), .Z(n15766) );
  XNOR U15775 ( .A(y[237]), .B(x[237]), .Z(n15775) );
  AND U15776 ( .A(n15776), .B(n15777), .Z(n15774) );
  XNOR U15777 ( .A(y[232]), .B(x[232]), .Z(n15777) );
  XNOR U15778 ( .A(y[233]), .B(x[233]), .Z(n15776) );
  AND U15779 ( .A(n15778), .B(n15779), .Z(n15764) );
  AND U15780 ( .A(n15780), .B(n15781), .Z(n15779) );
  AND U15781 ( .A(n15782), .B(n15783), .Z(n15781) );
  XNOR U15782 ( .A(y[235]), .B(x[235]), .Z(n15783) );
  XNOR U15783 ( .A(y[236]), .B(x[236]), .Z(n15782) );
  AND U15784 ( .A(n15784), .B(n15785), .Z(n15780) );
  XNOR U15785 ( .A(y[240]), .B(x[240]), .Z(n15785) );
  XNOR U15786 ( .A(y[238]), .B(x[238]), .Z(n15784) );
  AND U15787 ( .A(n15786), .B(n15787), .Z(n15778) );
  XNOR U15788 ( .A(y[241]), .B(x[241]), .Z(n15787) );
  AND U15789 ( .A(n15788), .B(n15789), .Z(n15786) );
  XNOR U15790 ( .A(y[239]), .B(x[239]), .Z(n15789) );
  XNOR U15791 ( .A(y[243]), .B(x[243]), .Z(n15788) );
  AND U15792 ( .A(n15790), .B(n15791), .Z(n15762) );
  AND U15793 ( .A(n15792), .B(n15793), .Z(n15791) );
  AND U15794 ( .A(n15794), .B(n15795), .Z(n15793) );
  AND U15795 ( .A(n15796), .B(n15797), .Z(n15795) );
  XNOR U15796 ( .A(y[242]), .B(x[242]), .Z(n15797) );
  XNOR U15797 ( .A(y[246]), .B(x[246]), .Z(n15796) );
  AND U15798 ( .A(n15798), .B(n15799), .Z(n15794) );
  XNOR U15799 ( .A(y[244]), .B(x[244]), .Z(n15799) );
  XNOR U15800 ( .A(y[245]), .B(x[245]), .Z(n15798) );
  AND U15801 ( .A(n15800), .B(n15801), .Z(n15792) );
  XNOR U15802 ( .A(y[248]), .B(x[248]), .Z(n15801) );
  AND U15803 ( .A(n15802), .B(n15803), .Z(n15800) );
  XNOR U15804 ( .A(y[249]), .B(x[249]), .Z(n15803) );
  XNOR U15805 ( .A(y[247]), .B(x[247]), .Z(n15802) );
  AND U15806 ( .A(n15804), .B(n15805), .Z(n15790) );
  AND U15807 ( .A(n15806), .B(n15807), .Z(n15805) );
  XNOR U15808 ( .A(y[252]), .B(x[252]), .Z(n15807) );
  AND U15809 ( .A(n15808), .B(n15809), .Z(n15806) );
  XNOR U15810 ( .A(y[250]), .B(x[250]), .Z(n15809) );
  XNOR U15811 ( .A(y[251]), .B(x[251]), .Z(n15808) );
  AND U15812 ( .A(n15810), .B(n15811), .Z(n15804) );
  XNOR U15813 ( .A(y[254]), .B(x[254]), .Z(n15811) );
  AND U15814 ( .A(n15812), .B(n15813), .Z(n15810) );
  XNOR U15815 ( .A(y[253]), .B(x[253]), .Z(n15813) );
  XNOR U15816 ( .A(y[256]), .B(x[256]), .Z(n15812) );
  AND U15817 ( .A(n15814), .B(n15815), .Z(n15760) );
  AND U15818 ( .A(n15816), .B(n15817), .Z(n15815) );
  AND U15819 ( .A(n15818), .B(n15819), .Z(n15817) );
  AND U15820 ( .A(n15820), .B(n15821), .Z(n15819) );
  AND U15821 ( .A(n15822), .B(n15823), .Z(n15821) );
  XNOR U15822 ( .A(y[255]), .B(x[255]), .Z(n15823) );
  XNOR U15823 ( .A(y[259]), .B(x[259]), .Z(n15822) );
  AND U15824 ( .A(n15824), .B(n15825), .Z(n15820) );
  XNOR U15825 ( .A(y[257]), .B(x[257]), .Z(n15825) );
  XNOR U15826 ( .A(y[258]), .B(x[258]), .Z(n15824) );
  AND U15827 ( .A(n15826), .B(n15827), .Z(n15818) );
  XNOR U15828 ( .A(y[261]), .B(x[261]), .Z(n15827) );
  AND U15829 ( .A(n15828), .B(n15829), .Z(n15826) );
  XNOR U15830 ( .A(y[262]), .B(x[262]), .Z(n15829) );
  XNOR U15831 ( .A(y[260]), .B(x[260]), .Z(n15828) );
  AND U15832 ( .A(n15830), .B(n15831), .Z(n15816) );
  AND U15833 ( .A(n15832), .B(n15833), .Z(n15831) );
  XNOR U15834 ( .A(y[264]), .B(x[264]), .Z(n15833) );
  AND U15835 ( .A(n15834), .B(n15835), .Z(n15832) );
  XNOR U15836 ( .A(y[265]), .B(x[265]), .Z(n15835) );
  XNOR U15837 ( .A(y[263]), .B(x[263]), .Z(n15834) );
  AND U15838 ( .A(n15836), .B(n15837), .Z(n15830) );
  XNOR U15839 ( .A(y[267]), .B(x[267]), .Z(n15837) );
  AND U15840 ( .A(n15838), .B(n15839), .Z(n15836) );
  XNOR U15841 ( .A(y[268]), .B(x[268]), .Z(n15839) );
  XNOR U15842 ( .A(y[266]), .B(x[266]), .Z(n15838) );
  AND U15843 ( .A(n15840), .B(n15841), .Z(n15814) );
  AND U15844 ( .A(n15842), .B(n15843), .Z(n15841) );
  AND U15845 ( .A(n15844), .B(n15845), .Z(n15843) );
  AND U15846 ( .A(n15846), .B(n15847), .Z(n15845) );
  XNOR U15847 ( .A(y[271]), .B(x[271]), .Z(n15847) );
  XNOR U15848 ( .A(y[269]), .B(x[269]), .Z(n15846) );
  AND U15849 ( .A(n15848), .B(n15849), .Z(n15844) );
  XNOR U15850 ( .A(y[270]), .B(x[270]), .Z(n15849) );
  XNOR U15851 ( .A(y[274]), .B(x[274]), .Z(n15848) );
  AND U15852 ( .A(n15850), .B(n15851), .Z(n15842) );
  XNOR U15853 ( .A(y[275]), .B(x[275]), .Z(n15851) );
  AND U15854 ( .A(n15852), .B(n15853), .Z(n15850) );
  XNOR U15855 ( .A(y[272]), .B(x[272]), .Z(n15853) );
  XNOR U15856 ( .A(y[273]), .B(x[273]), .Z(n15852) );
  AND U15857 ( .A(n15854), .B(n15855), .Z(n15840) );
  AND U15858 ( .A(n15856), .B(n15857), .Z(n15855) );
  XNOR U15859 ( .A(y[278]), .B(x[278]), .Z(n15857) );
  AND U15860 ( .A(n15858), .B(n15859), .Z(n15856) );
  XNOR U15861 ( .A(y[276]), .B(x[276]), .Z(n15859) );
  XNOR U15862 ( .A(y[277]), .B(x[277]), .Z(n15858) );
  AND U15863 ( .A(n15860), .B(n15861), .Z(n15854) );
  XNOR U15864 ( .A(y[280]), .B(x[280]), .Z(n15861) );
  AND U15865 ( .A(n15862), .B(n15863), .Z(n15860) );
  XNOR U15866 ( .A(y[281]), .B(x[281]), .Z(n15863) );
  XNOR U15867 ( .A(y[279]), .B(x[279]), .Z(n15862) );
  AND U15868 ( .A(n15864), .B(n15865), .Z(n15758) );
  AND U15869 ( .A(n15866), .B(n15867), .Z(n15865) );
  AND U15870 ( .A(n15868), .B(n15869), .Z(n15867) );
  AND U15871 ( .A(n15870), .B(n15871), .Z(n15869) );
  AND U15872 ( .A(n15872), .B(n15873), .Z(n15871) );
  AND U15873 ( .A(n15874), .B(n15875), .Z(n15873) );
  XNOR U15874 ( .A(y[284]), .B(x[284]), .Z(n15875) );
  XNOR U15875 ( .A(y[282]), .B(x[282]), .Z(n15874) );
  AND U15876 ( .A(n15876), .B(n15877), .Z(n15872) );
  XNOR U15877 ( .A(y[283]), .B(x[283]), .Z(n15877) );
  XNOR U15878 ( .A(y[287]), .B(x[287]), .Z(n15876) );
  AND U15879 ( .A(n15878), .B(n15879), .Z(n15870) );
  XNOR U15880 ( .A(y[290]), .B(x[290]), .Z(n15879) );
  AND U15881 ( .A(n15880), .B(n15881), .Z(n15878) );
  XNOR U15882 ( .A(y[285]), .B(x[285]), .Z(n15881) );
  XNOR U15883 ( .A(y[286]), .B(x[286]), .Z(n15880) );
  AND U15884 ( .A(n15882), .B(n15883), .Z(n15868) );
  AND U15885 ( .A(n15884), .B(n15885), .Z(n15883) );
  AND U15886 ( .A(n15886), .B(n15887), .Z(n15885) );
  XNOR U15887 ( .A(y[288]), .B(x[288]), .Z(n15887) );
  XNOR U15888 ( .A(y[289]), .B(x[289]), .Z(n15886) );
  AND U15889 ( .A(n15888), .B(n15889), .Z(n15884) );
  XNOR U15890 ( .A(y[293]), .B(x[293]), .Z(n15889) );
  XNOR U15891 ( .A(y[291]), .B(x[291]), .Z(n15888) );
  AND U15892 ( .A(n15890), .B(n15891), .Z(n15882) );
  XNOR U15893 ( .A(y[294]), .B(x[294]), .Z(n15891) );
  AND U15894 ( .A(n15892), .B(n15893), .Z(n15890) );
  XNOR U15895 ( .A(y[292]), .B(x[292]), .Z(n15893) );
  XNOR U15896 ( .A(y[296]), .B(x[296]), .Z(n15892) );
  AND U15897 ( .A(n15894), .B(n15895), .Z(n15866) );
  AND U15898 ( .A(n15896), .B(n15897), .Z(n15895) );
  AND U15899 ( .A(n15898), .B(n15899), .Z(n15897) );
  AND U15900 ( .A(n15900), .B(n15901), .Z(n15899) );
  XNOR U15901 ( .A(y[295]), .B(x[295]), .Z(n15901) );
  XNOR U15902 ( .A(y[299]), .B(x[299]), .Z(n15900) );
  AND U15903 ( .A(n15902), .B(n15903), .Z(n15898) );
  XNOR U15904 ( .A(y[297]), .B(x[297]), .Z(n15903) );
  XNOR U15905 ( .A(y[298]), .B(x[298]), .Z(n15902) );
  AND U15906 ( .A(n15904), .B(n15905), .Z(n15896) );
  XNOR U15907 ( .A(y[376]), .B(x[376]), .Z(n15905) );
  AND U15908 ( .A(n15906), .B(n15907), .Z(n15904) );
  XNOR U15909 ( .A(y[377]), .B(x[377]), .Z(n15907) );
  XNOR U15910 ( .A(y[375]), .B(x[375]), .Z(n15906) );
  AND U15911 ( .A(n15908), .B(n15909), .Z(n15894) );
  AND U15912 ( .A(n15910), .B(n15911), .Z(n15909) );
  XNOR U15913 ( .A(y[379]), .B(x[379]), .Z(n15911) );
  AND U15914 ( .A(n15912), .B(n15913), .Z(n15910) );
  XNOR U15915 ( .A(y[380]), .B(x[380]), .Z(n15913) );
  XNOR U15916 ( .A(y[378]), .B(x[378]), .Z(n15912) );
  AND U15917 ( .A(n15914), .B(n15915), .Z(n15908) );
  XNOR U15918 ( .A(y[382]), .B(x[382]), .Z(n15915) );
  AND U15919 ( .A(n15916), .B(n15917), .Z(n15914) );
  XNOR U15920 ( .A(y[383]), .B(x[383]), .Z(n15917) );
  XNOR U15921 ( .A(y[381]), .B(x[381]), .Z(n15916) );
  AND U15922 ( .A(n15918), .B(n15919), .Z(n15864) );
  AND U15923 ( .A(n15920), .B(n15921), .Z(n15919) );
  AND U15924 ( .A(n15922), .B(n15923), .Z(n15921) );
  AND U15925 ( .A(n15924), .B(n15925), .Z(n15923) );
  AND U15926 ( .A(n15926), .B(n15927), .Z(n15925) );
  XNOR U15927 ( .A(y[386]), .B(x[386]), .Z(n15927) );
  XNOR U15928 ( .A(y[384]), .B(x[384]), .Z(n15926) );
  AND U15929 ( .A(n15928), .B(n15929), .Z(n15924) );
  XNOR U15930 ( .A(y[385]), .B(x[385]), .Z(n15929) );
  XNOR U15931 ( .A(y[389]), .B(x[389]), .Z(n15928) );
  AND U15932 ( .A(n15930), .B(n15931), .Z(n15922) );
  XNOR U15933 ( .A(y[392]), .B(x[392]), .Z(n15931) );
  AND U15934 ( .A(n15932), .B(n15933), .Z(n15930) );
  XNOR U15935 ( .A(y[387]), .B(x[387]), .Z(n15933) );
  XNOR U15936 ( .A(y[388]), .B(x[388]), .Z(n15932) );
  AND U15937 ( .A(n15934), .B(n15935), .Z(n15920) );
  AND U15938 ( .A(n15936), .B(n15937), .Z(n15935) );
  XNOR U15939 ( .A(y[395]), .B(x[395]), .Z(n15937) );
  AND U15940 ( .A(n15938), .B(n15939), .Z(n15936) );
  XNOR U15941 ( .A(y[390]), .B(x[390]), .Z(n15939) );
  XNOR U15942 ( .A(y[391]), .B(x[391]), .Z(n15938) );
  AND U15943 ( .A(n15940), .B(n15941), .Z(n15934) );
  XNOR U15944 ( .A(y[718]), .B(x[718]), .Z(n15941) );
  AND U15945 ( .A(n15942), .B(n15943), .Z(n15940) );
  XNOR U15946 ( .A(y[393]), .B(x[393]), .Z(n15943) );
  XNOR U15947 ( .A(y[394]), .B(x[394]), .Z(n15942) );
  AND U15948 ( .A(n15944), .B(n15945), .Z(n15918) );
  AND U15949 ( .A(n15946), .B(n15947), .Z(n15945) );
  AND U15950 ( .A(n15948), .B(n15949), .Z(n15947) );
  AND U15951 ( .A(n15950), .B(n15951), .Z(n15949) );
  XNOR U15952 ( .A(y[719]), .B(x[719]), .Z(n15951) );
  XNOR U15953 ( .A(y[720]), .B(x[720]), .Z(n15950) );
  AND U15954 ( .A(n15952), .B(n15953), .Z(n15948) );
  XNOR U15955 ( .A(y[721]), .B(x[721]), .Z(n15953) );
  XNOR U15956 ( .A(y[722]), .B(x[722]), .Z(n15952) );
  AND U15957 ( .A(n15954), .B(n15955), .Z(n15946) );
  XNOR U15958 ( .A(y[725]), .B(x[725]), .Z(n15955) );
  AND U15959 ( .A(n15956), .B(n15957), .Z(n15954) );
  XNOR U15960 ( .A(y[723]), .B(x[723]), .Z(n15957) );
  XNOR U15961 ( .A(y[724]), .B(x[724]), .Z(n15956) );
  AND U15962 ( .A(n15958), .B(n15959), .Z(n15944) );
  AND U15963 ( .A(n15960), .B(n15961), .Z(n15959) );
  XNOR U15964 ( .A(y[728]), .B(x[728]), .Z(n15961) );
  AND U15965 ( .A(n15962), .B(n15963), .Z(n15960) );
  XNOR U15966 ( .A(y[726]), .B(x[726]), .Z(n15963) );
  XNOR U15967 ( .A(y[727]), .B(x[727]), .Z(n15962) );
  AND U15968 ( .A(n15964), .B(n15965), .Z(n15958) );
  XNOR U15969 ( .A(y[731]), .B(x[731]), .Z(n15965) );
  AND U15970 ( .A(n15966), .B(n15967), .Z(n15964) );
  XNOR U15971 ( .A(y[729]), .B(x[729]), .Z(n15967) );
  XNOR U15972 ( .A(y[730]), .B(x[730]), .Z(n15966) );
  AND U15973 ( .A(n15968), .B(n15969), .Z(n8200) );
  AND U15974 ( .A(n15970), .B(n15971), .Z(n15969) );
  AND U15975 ( .A(n15972), .B(n15973), .Z(n15971) );
  AND U15976 ( .A(n15974), .B(n15975), .Z(n15973) );
  AND U15977 ( .A(n15976), .B(n15977), .Z(n15975) );
  AND U15978 ( .A(n15978), .B(n15979), .Z(n15977) );
  AND U15979 ( .A(n15980), .B(n15981), .Z(n15979) );
  AND U15980 ( .A(n15982), .B(n15983), .Z(n15981) );
  XNOR U15981 ( .A(y[732]), .B(x[732]), .Z(n15983) );
  XNOR U15982 ( .A(y[733]), .B(x[733]), .Z(n15982) );
  AND U15983 ( .A(n15984), .B(n15985), .Z(n15980) );
  XNOR U15984 ( .A(y[734]), .B(x[734]), .Z(n15985) );
  XNOR U15985 ( .A(y[735]), .B(x[735]), .Z(n15984) );
  AND U15986 ( .A(n15986), .B(n15987), .Z(n15978) );
  XNOR U15987 ( .A(y[738]), .B(x[738]), .Z(n15987) );
  AND U15988 ( .A(n15988), .B(n15989), .Z(n15986) );
  XNOR U15989 ( .A(y[736]), .B(x[736]), .Z(n15989) );
  XNOR U15990 ( .A(y[737]), .B(x[737]), .Z(n15988) );
  AND U15991 ( .A(n15990), .B(n15991), .Z(n15976) );
  AND U15992 ( .A(n15992), .B(n15993), .Z(n15991) );
  AND U15993 ( .A(n15994), .B(n15995), .Z(n15993) );
  XNOR U15994 ( .A(y[739]), .B(x[739]), .Z(n15995) );
  XNOR U15995 ( .A(y[740]), .B(x[740]), .Z(n15994) );
  AND U15996 ( .A(n15996), .B(n15997), .Z(n15992) );
  XNOR U15997 ( .A(y[741]), .B(x[741]), .Z(n15997) );
  XNOR U15998 ( .A(y[742]), .B(x[742]), .Z(n15996) );
  AND U15999 ( .A(n15998), .B(n15999), .Z(n15990) );
  XNOR U16000 ( .A(y[745]), .B(x[745]), .Z(n15999) );
  AND U16001 ( .A(n16000), .B(n16001), .Z(n15998) );
  XNOR U16002 ( .A(y[743]), .B(x[743]), .Z(n16001) );
  XNOR U16003 ( .A(y[744]), .B(x[744]), .Z(n16000) );
  AND U16004 ( .A(n16002), .B(n16003), .Z(n15974) );
  AND U16005 ( .A(n16004), .B(n16005), .Z(n16003) );
  AND U16006 ( .A(n16006), .B(n16007), .Z(n16005) );
  AND U16007 ( .A(n16008), .B(n16009), .Z(n16007) );
  XNOR U16008 ( .A(y[746]), .B(x[746]), .Z(n16009) );
  XNOR U16009 ( .A(y[747]), .B(x[747]), .Z(n16008) );
  AND U16010 ( .A(n16010), .B(n16011), .Z(n16006) );
  XNOR U16011 ( .A(y[748]), .B(x[748]), .Z(n16011) );
  XNOR U16012 ( .A(y[749]), .B(x[749]), .Z(n16010) );
  AND U16013 ( .A(n16012), .B(n16013), .Z(n16004) );
  XNOR U16014 ( .A(y[752]), .B(x[752]), .Z(n16013) );
  AND U16015 ( .A(n16014), .B(n16015), .Z(n16012) );
  XNOR U16016 ( .A(y[750]), .B(x[750]), .Z(n16015) );
  XNOR U16017 ( .A(y[751]), .B(x[751]), .Z(n16014) );
  AND U16018 ( .A(n16016), .B(n16017), .Z(n16002) );
  AND U16019 ( .A(n16018), .B(n16019), .Z(n16017) );
  XNOR U16020 ( .A(y[755]), .B(x[755]), .Z(n16019) );
  AND U16021 ( .A(n16020), .B(n16021), .Z(n16018) );
  XNOR U16022 ( .A(y[753]), .B(x[753]), .Z(n16021) );
  XNOR U16023 ( .A(y[754]), .B(x[754]), .Z(n16020) );
  AND U16024 ( .A(n16022), .B(n16023), .Z(n16016) );
  XNOR U16025 ( .A(y[758]), .B(x[758]), .Z(n16023) );
  AND U16026 ( .A(n16024), .B(n16025), .Z(n16022) );
  XNOR U16027 ( .A(y[756]), .B(x[756]), .Z(n16025) );
  XNOR U16028 ( .A(y[757]), .B(x[757]), .Z(n16024) );
  AND U16029 ( .A(n16026), .B(n16027), .Z(n15972) );
  AND U16030 ( .A(n16028), .B(n16029), .Z(n16027) );
  AND U16031 ( .A(n16030), .B(n16031), .Z(n16029) );
  AND U16032 ( .A(n16032), .B(n16033), .Z(n16031) );
  AND U16033 ( .A(n16034), .B(n16035), .Z(n16033) );
  XNOR U16034 ( .A(y[759]), .B(x[759]), .Z(n16035) );
  XNOR U16035 ( .A(y[760]), .B(x[760]), .Z(n16034) );
  AND U16036 ( .A(n16036), .B(n16037), .Z(n16032) );
  XNOR U16037 ( .A(y[761]), .B(x[761]), .Z(n16037) );
  XNOR U16038 ( .A(y[762]), .B(x[762]), .Z(n16036) );
  AND U16039 ( .A(n16038), .B(n16039), .Z(n16030) );
  XNOR U16040 ( .A(y[765]), .B(x[765]), .Z(n16039) );
  AND U16041 ( .A(n16040), .B(n16041), .Z(n16038) );
  XNOR U16042 ( .A(y[763]), .B(x[763]), .Z(n16041) );
  XNOR U16043 ( .A(y[764]), .B(x[764]), .Z(n16040) );
  AND U16044 ( .A(n16042), .B(n16043), .Z(n16028) );
  AND U16045 ( .A(n16044), .B(n16045), .Z(n16043) );
  XNOR U16046 ( .A(y[768]), .B(x[768]), .Z(n16045) );
  AND U16047 ( .A(n16046), .B(n16047), .Z(n16044) );
  XNOR U16048 ( .A(y[766]), .B(x[766]), .Z(n16047) );
  XNOR U16049 ( .A(y[767]), .B(x[767]), .Z(n16046) );
  AND U16050 ( .A(n16048), .B(n16049), .Z(n16042) );
  XNOR U16051 ( .A(y[771]), .B(x[771]), .Z(n16049) );
  AND U16052 ( .A(n16050), .B(n16051), .Z(n16048) );
  XNOR U16053 ( .A(y[769]), .B(x[769]), .Z(n16051) );
  XNOR U16054 ( .A(y[770]), .B(x[770]), .Z(n16050) );
  AND U16055 ( .A(n16052), .B(n16053), .Z(n16026) );
  AND U16056 ( .A(n16054), .B(n16055), .Z(n16053) );
  AND U16057 ( .A(n16056), .B(n16057), .Z(n16055) );
  AND U16058 ( .A(n16058), .B(n16059), .Z(n16057) );
  XNOR U16059 ( .A(y[772]), .B(x[772]), .Z(n16059) );
  XNOR U16060 ( .A(y[773]), .B(x[773]), .Z(n16058) );
  AND U16061 ( .A(n16060), .B(n16061), .Z(n16056) );
  XNOR U16062 ( .A(y[774]), .B(x[774]), .Z(n16061) );
  XNOR U16063 ( .A(y[775]), .B(x[775]), .Z(n16060) );
  AND U16064 ( .A(n16062), .B(n16063), .Z(n16054) );
  XNOR U16065 ( .A(y[778]), .B(x[778]), .Z(n16063) );
  AND U16066 ( .A(n16064), .B(n16065), .Z(n16062) );
  XNOR U16067 ( .A(y[776]), .B(x[776]), .Z(n16065) );
  XNOR U16068 ( .A(y[777]), .B(x[777]), .Z(n16064) );
  AND U16069 ( .A(n16066), .B(n16067), .Z(n16052) );
  AND U16070 ( .A(n16068), .B(n16069), .Z(n16067) );
  XNOR U16071 ( .A(y[781]), .B(x[781]), .Z(n16069) );
  AND U16072 ( .A(n16070), .B(n16071), .Z(n16068) );
  XNOR U16073 ( .A(y[779]), .B(x[779]), .Z(n16071) );
  XNOR U16074 ( .A(y[780]), .B(x[780]), .Z(n16070) );
  AND U16075 ( .A(n16072), .B(n16073), .Z(n16066) );
  XNOR U16076 ( .A(y[784]), .B(x[784]), .Z(n16073) );
  AND U16077 ( .A(n16074), .B(n16075), .Z(n16072) );
  XNOR U16078 ( .A(y[782]), .B(x[782]), .Z(n16075) );
  XNOR U16079 ( .A(y[783]), .B(x[783]), .Z(n16074) );
  AND U16080 ( .A(n16076), .B(n16077), .Z(n15970) );
  AND U16081 ( .A(n16078), .B(n16079), .Z(n16077) );
  AND U16082 ( .A(n16080), .B(n16081), .Z(n16079) );
  AND U16083 ( .A(n16082), .B(n16083), .Z(n16081) );
  AND U16084 ( .A(n16084), .B(n16085), .Z(n16083) );
  AND U16085 ( .A(n16086), .B(n16087), .Z(n16085) );
  XNOR U16086 ( .A(y[785]), .B(x[785]), .Z(n16087) );
  XNOR U16087 ( .A(y[786]), .B(x[786]), .Z(n16086) );
  AND U16088 ( .A(n16088), .B(n16089), .Z(n16084) );
  XNOR U16089 ( .A(y[787]), .B(x[787]), .Z(n16089) );
  XNOR U16090 ( .A(y[788]), .B(x[788]), .Z(n16088) );
  AND U16091 ( .A(n16090), .B(n16091), .Z(n16082) );
  XNOR U16092 ( .A(y[791]), .B(x[791]), .Z(n16091) );
  AND U16093 ( .A(n16092), .B(n16093), .Z(n16090) );
  XNOR U16094 ( .A(y[789]), .B(x[789]), .Z(n16093) );
  XNOR U16095 ( .A(y[790]), .B(x[790]), .Z(n16092) );
  AND U16096 ( .A(n16094), .B(n16095), .Z(n16080) );
  AND U16097 ( .A(n16096), .B(n16097), .Z(n16095) );
  AND U16098 ( .A(n16098), .B(n16099), .Z(n16097) );
  XNOR U16099 ( .A(y[792]), .B(x[792]), .Z(n16099) );
  XNOR U16100 ( .A(y[793]), .B(x[793]), .Z(n16098) );
  AND U16101 ( .A(n16100), .B(n16101), .Z(n16096) );
  XNOR U16102 ( .A(y[794]), .B(x[794]), .Z(n16101) );
  XNOR U16103 ( .A(y[795]), .B(x[795]), .Z(n16100) );
  AND U16104 ( .A(n16102), .B(n16103), .Z(n16094) );
  XNOR U16105 ( .A(y[798]), .B(x[798]), .Z(n16103) );
  AND U16106 ( .A(n16104), .B(n16105), .Z(n16102) );
  XNOR U16107 ( .A(y[796]), .B(x[796]), .Z(n16105) );
  XNOR U16108 ( .A(y[797]), .B(x[797]), .Z(n16104) );
  AND U16109 ( .A(n16106), .B(n16107), .Z(n16078) );
  AND U16110 ( .A(n16108), .B(n16109), .Z(n16107) );
  AND U16111 ( .A(n16110), .B(n16111), .Z(n16109) );
  AND U16112 ( .A(n16112), .B(n16113), .Z(n16111) );
  XNOR U16113 ( .A(y[799]), .B(x[799]), .Z(n16113) );
  XNOR U16114 ( .A(y[800]), .B(x[800]), .Z(n16112) );
  AND U16115 ( .A(n16114), .B(n16115), .Z(n16110) );
  XNOR U16116 ( .A(y[801]), .B(x[801]), .Z(n16115) );
  XNOR U16117 ( .A(y[802]), .B(x[802]), .Z(n16114) );
  AND U16118 ( .A(n16116), .B(n16117), .Z(n16108) );
  XNOR U16119 ( .A(y[805]), .B(x[805]), .Z(n16117) );
  AND U16120 ( .A(n16118), .B(n16119), .Z(n16116) );
  XNOR U16121 ( .A(y[803]), .B(x[803]), .Z(n16119) );
  XNOR U16122 ( .A(y[804]), .B(x[804]), .Z(n16118) );
  AND U16123 ( .A(n16120), .B(n16121), .Z(n16106) );
  AND U16124 ( .A(n16122), .B(n16123), .Z(n16121) );
  XNOR U16125 ( .A(y[808]), .B(x[808]), .Z(n16123) );
  AND U16126 ( .A(n16124), .B(n16125), .Z(n16122) );
  XNOR U16127 ( .A(y[806]), .B(x[806]), .Z(n16125) );
  XNOR U16128 ( .A(y[807]), .B(x[807]), .Z(n16124) );
  AND U16129 ( .A(n16126), .B(n16127), .Z(n16120) );
  XNOR U16130 ( .A(y[811]), .B(x[811]), .Z(n16127) );
  AND U16131 ( .A(n16128), .B(n16129), .Z(n16126) );
  XNOR U16132 ( .A(y[809]), .B(x[809]), .Z(n16129) );
  XNOR U16133 ( .A(y[810]), .B(x[810]), .Z(n16128) );
  AND U16134 ( .A(n16130), .B(n16131), .Z(n16076) );
  AND U16135 ( .A(n16132), .B(n16133), .Z(n16131) );
  AND U16136 ( .A(n16134), .B(n16135), .Z(n16133) );
  AND U16137 ( .A(n16136), .B(n16137), .Z(n16135) );
  AND U16138 ( .A(n16138), .B(n16139), .Z(n16137) );
  XNOR U16139 ( .A(y[812]), .B(x[812]), .Z(n16139) );
  XNOR U16140 ( .A(y[813]), .B(x[813]), .Z(n16138) );
  AND U16141 ( .A(n16140), .B(n16141), .Z(n16136) );
  XNOR U16142 ( .A(y[814]), .B(x[814]), .Z(n16141) );
  XNOR U16143 ( .A(y[815]), .B(x[815]), .Z(n16140) );
  AND U16144 ( .A(n16142), .B(n16143), .Z(n16134) );
  XNOR U16145 ( .A(y[818]), .B(x[818]), .Z(n16143) );
  AND U16146 ( .A(n16144), .B(n16145), .Z(n16142) );
  XNOR U16147 ( .A(y[816]), .B(x[816]), .Z(n16145) );
  XNOR U16148 ( .A(y[817]), .B(x[817]), .Z(n16144) );
  AND U16149 ( .A(n16146), .B(n16147), .Z(n16132) );
  AND U16150 ( .A(n16148), .B(n16149), .Z(n16147) );
  XNOR U16151 ( .A(y[821]), .B(x[821]), .Z(n16149) );
  AND U16152 ( .A(n16150), .B(n16151), .Z(n16148) );
  XNOR U16153 ( .A(y[819]), .B(x[819]), .Z(n16151) );
  XNOR U16154 ( .A(y[820]), .B(x[820]), .Z(n16150) );
  AND U16155 ( .A(n16152), .B(n16153), .Z(n16146) );
  XNOR U16156 ( .A(y[824]), .B(x[824]), .Z(n16153) );
  AND U16157 ( .A(n16154), .B(n16155), .Z(n16152) );
  XNOR U16158 ( .A(y[822]), .B(x[822]), .Z(n16155) );
  XNOR U16159 ( .A(y[823]), .B(x[823]), .Z(n16154) );
  AND U16160 ( .A(n16156), .B(n16157), .Z(n16130) );
  AND U16161 ( .A(n16158), .B(n16159), .Z(n16157) );
  AND U16162 ( .A(n16160), .B(n16161), .Z(n16159) );
  AND U16163 ( .A(n16162), .B(n16163), .Z(n16161) );
  XNOR U16164 ( .A(y[825]), .B(x[825]), .Z(n16163) );
  XNOR U16165 ( .A(y[826]), .B(x[826]), .Z(n16162) );
  AND U16166 ( .A(n16164), .B(n16165), .Z(n16160) );
  XNOR U16167 ( .A(y[827]), .B(x[827]), .Z(n16165) );
  XNOR U16168 ( .A(y[828]), .B(x[828]), .Z(n16164) );
  AND U16169 ( .A(n16166), .B(n16167), .Z(n16158) );
  XNOR U16170 ( .A(y[831]), .B(x[831]), .Z(n16167) );
  AND U16171 ( .A(n16168), .B(n16169), .Z(n16166) );
  XNOR U16172 ( .A(y[829]), .B(x[829]), .Z(n16169) );
  XNOR U16173 ( .A(y[830]), .B(x[830]), .Z(n16168) );
  AND U16174 ( .A(n16170), .B(n16171), .Z(n16156) );
  AND U16175 ( .A(n16172), .B(n16173), .Z(n16171) );
  XNOR U16176 ( .A(y[834]), .B(x[834]), .Z(n16173) );
  AND U16177 ( .A(n16174), .B(n16175), .Z(n16172) );
  XNOR U16178 ( .A(y[832]), .B(x[832]), .Z(n16175) );
  XNOR U16179 ( .A(y[833]), .B(x[833]), .Z(n16174) );
  AND U16180 ( .A(n16176), .B(n16177), .Z(n16170) );
  XNOR U16181 ( .A(y[837]), .B(x[837]), .Z(n16177) );
  AND U16182 ( .A(n16178), .B(n16179), .Z(n16176) );
  XNOR U16183 ( .A(y[835]), .B(x[835]), .Z(n16179) );
  XNOR U16184 ( .A(y[836]), .B(x[836]), .Z(n16178) );
  AND U16185 ( .A(n16180), .B(n16181), .Z(n15968) );
  AND U16186 ( .A(n16182), .B(n16183), .Z(n16181) );
  AND U16187 ( .A(n16184), .B(n16185), .Z(n16183) );
  AND U16188 ( .A(n16186), .B(n16187), .Z(n16185) );
  AND U16189 ( .A(n16188), .B(n16189), .Z(n16187) );
  AND U16190 ( .A(n16190), .B(n16191), .Z(n16189) );
  AND U16191 ( .A(n16192), .B(n16193), .Z(n16191) );
  XNOR U16192 ( .A(y[838]), .B(x[838]), .Z(n16193) );
  XNOR U16193 ( .A(y[839]), .B(x[839]), .Z(n16192) );
  AND U16194 ( .A(n16194), .B(n16195), .Z(n16190) );
  XNOR U16195 ( .A(y[840]), .B(x[840]), .Z(n16195) );
  XNOR U16196 ( .A(y[841]), .B(x[841]), .Z(n16194) );
  AND U16197 ( .A(n16196), .B(n16197), .Z(n16188) );
  XNOR U16198 ( .A(y[844]), .B(x[844]), .Z(n16197) );
  AND U16199 ( .A(n16198), .B(n16199), .Z(n16196) );
  XNOR U16200 ( .A(y[842]), .B(x[842]), .Z(n16199) );
  XNOR U16201 ( .A(y[843]), .B(x[843]), .Z(n16198) );
  AND U16202 ( .A(n16200), .B(n16201), .Z(n16186) );
  AND U16203 ( .A(n16202), .B(n16203), .Z(n16201) );
  AND U16204 ( .A(n16204), .B(n16205), .Z(n16203) );
  XNOR U16205 ( .A(y[845]), .B(x[845]), .Z(n16205) );
  XNOR U16206 ( .A(y[846]), .B(x[846]), .Z(n16204) );
  AND U16207 ( .A(n16206), .B(n16207), .Z(n16202) );
  XNOR U16208 ( .A(y[847]), .B(x[847]), .Z(n16207) );
  XNOR U16209 ( .A(y[848]), .B(x[848]), .Z(n16206) );
  AND U16210 ( .A(n16208), .B(n16209), .Z(n16200) );
  XNOR U16211 ( .A(y[851]), .B(x[851]), .Z(n16209) );
  AND U16212 ( .A(n16210), .B(n16211), .Z(n16208) );
  XNOR U16213 ( .A(y[849]), .B(x[849]), .Z(n16211) );
  XNOR U16214 ( .A(y[850]), .B(x[850]), .Z(n16210) );
  AND U16215 ( .A(n16212), .B(n16213), .Z(n16184) );
  AND U16216 ( .A(n16214), .B(n16215), .Z(n16213) );
  AND U16217 ( .A(n16216), .B(n16217), .Z(n16215) );
  AND U16218 ( .A(n16218), .B(n16219), .Z(n16217) );
  XNOR U16219 ( .A(y[852]), .B(x[852]), .Z(n16219) );
  XNOR U16220 ( .A(y[853]), .B(x[853]), .Z(n16218) );
  AND U16221 ( .A(n16220), .B(n16221), .Z(n16216) );
  XNOR U16222 ( .A(y[854]), .B(x[854]), .Z(n16221) );
  XNOR U16223 ( .A(y[855]), .B(x[855]), .Z(n16220) );
  AND U16224 ( .A(n16222), .B(n16223), .Z(n16214) );
  XNOR U16225 ( .A(y[858]), .B(x[858]), .Z(n16223) );
  AND U16226 ( .A(n16224), .B(n16225), .Z(n16222) );
  XNOR U16227 ( .A(y[856]), .B(x[856]), .Z(n16225) );
  XNOR U16228 ( .A(y[857]), .B(x[857]), .Z(n16224) );
  AND U16229 ( .A(n16226), .B(n16227), .Z(n16212) );
  AND U16230 ( .A(n16228), .B(n16229), .Z(n16227) );
  XNOR U16231 ( .A(y[861]), .B(x[861]), .Z(n16229) );
  AND U16232 ( .A(n16230), .B(n16231), .Z(n16228) );
  XNOR U16233 ( .A(y[859]), .B(x[859]), .Z(n16231) );
  XNOR U16234 ( .A(y[860]), .B(x[860]), .Z(n16230) );
  AND U16235 ( .A(n16232), .B(n16233), .Z(n16226) );
  XNOR U16236 ( .A(y[864]), .B(x[864]), .Z(n16233) );
  AND U16237 ( .A(n16234), .B(n16235), .Z(n16232) );
  XNOR U16238 ( .A(y[862]), .B(x[862]), .Z(n16235) );
  XNOR U16239 ( .A(y[863]), .B(x[863]), .Z(n16234) );
  AND U16240 ( .A(n16236), .B(n16237), .Z(n16182) );
  AND U16241 ( .A(n16238), .B(n16239), .Z(n16237) );
  AND U16242 ( .A(n16240), .B(n16241), .Z(n16239) );
  AND U16243 ( .A(n16242), .B(n16243), .Z(n16241) );
  AND U16244 ( .A(n16244), .B(n16245), .Z(n16243) );
  XNOR U16245 ( .A(y[865]), .B(x[865]), .Z(n16245) );
  XNOR U16246 ( .A(y[866]), .B(x[866]), .Z(n16244) );
  AND U16247 ( .A(n16246), .B(n16247), .Z(n16242) );
  XNOR U16248 ( .A(y[867]), .B(x[867]), .Z(n16247) );
  XNOR U16249 ( .A(y[868]), .B(x[868]), .Z(n16246) );
  AND U16250 ( .A(n16248), .B(n16249), .Z(n16240) );
  XNOR U16251 ( .A(y[871]), .B(x[871]), .Z(n16249) );
  AND U16252 ( .A(n16250), .B(n16251), .Z(n16248) );
  XNOR U16253 ( .A(y[869]), .B(x[869]), .Z(n16251) );
  XNOR U16254 ( .A(y[870]), .B(x[870]), .Z(n16250) );
  AND U16255 ( .A(n16252), .B(n16253), .Z(n16238) );
  AND U16256 ( .A(n16254), .B(n16255), .Z(n16253) );
  XNOR U16257 ( .A(y[874]), .B(x[874]), .Z(n16255) );
  AND U16258 ( .A(n16256), .B(n16257), .Z(n16254) );
  XNOR U16259 ( .A(y[872]), .B(x[872]), .Z(n16257) );
  XNOR U16260 ( .A(y[873]), .B(x[873]), .Z(n16256) );
  AND U16261 ( .A(n16258), .B(n16259), .Z(n16252) );
  XNOR U16262 ( .A(y[877]), .B(x[877]), .Z(n16259) );
  AND U16263 ( .A(n16260), .B(n16261), .Z(n16258) );
  XNOR U16264 ( .A(y[875]), .B(x[875]), .Z(n16261) );
  XNOR U16265 ( .A(y[876]), .B(x[876]), .Z(n16260) );
  AND U16266 ( .A(n16262), .B(n16263), .Z(n16236) );
  AND U16267 ( .A(n16264), .B(n16265), .Z(n16263) );
  AND U16268 ( .A(n16266), .B(n16267), .Z(n16265) );
  AND U16269 ( .A(n16268), .B(n16269), .Z(n16267) );
  XNOR U16270 ( .A(y[878]), .B(x[878]), .Z(n16269) );
  XNOR U16271 ( .A(y[879]), .B(x[879]), .Z(n16268) );
  AND U16272 ( .A(n16270), .B(n16271), .Z(n16266) );
  XNOR U16273 ( .A(y[880]), .B(x[880]), .Z(n16271) );
  XNOR U16274 ( .A(y[881]), .B(x[881]), .Z(n16270) );
  AND U16275 ( .A(n16272), .B(n16273), .Z(n16264) );
  XNOR U16276 ( .A(y[884]), .B(x[884]), .Z(n16273) );
  AND U16277 ( .A(n16274), .B(n16275), .Z(n16272) );
  XNOR U16278 ( .A(y[882]), .B(x[882]), .Z(n16275) );
  XNOR U16279 ( .A(y[883]), .B(x[883]), .Z(n16274) );
  AND U16280 ( .A(n16276), .B(n16277), .Z(n16262) );
  AND U16281 ( .A(n16278), .B(n16279), .Z(n16277) );
  XNOR U16282 ( .A(y[887]), .B(x[887]), .Z(n16279) );
  AND U16283 ( .A(n16280), .B(n16281), .Z(n16278) );
  XNOR U16284 ( .A(y[885]), .B(x[885]), .Z(n16281) );
  XNOR U16285 ( .A(y[886]), .B(x[886]), .Z(n16280) );
  AND U16286 ( .A(n16282), .B(n16283), .Z(n16276) );
  XNOR U16287 ( .A(y[890]), .B(x[890]), .Z(n16283) );
  AND U16288 ( .A(n16284), .B(n16285), .Z(n16282) );
  XNOR U16289 ( .A(y[888]), .B(x[888]), .Z(n16285) );
  XNOR U16290 ( .A(y[889]), .B(x[889]), .Z(n16284) );
  AND U16291 ( .A(n16286), .B(n16287), .Z(n16180) );
  AND U16292 ( .A(n16288), .B(n16289), .Z(n16287) );
  AND U16293 ( .A(n16290), .B(n16291), .Z(n16289) );
  AND U16294 ( .A(n16292), .B(n16293), .Z(n16291) );
  AND U16295 ( .A(n16294), .B(n16295), .Z(n16293) );
  AND U16296 ( .A(n16296), .B(n16297), .Z(n16295) );
  XNOR U16297 ( .A(y[891]), .B(x[891]), .Z(n16297) );
  XNOR U16298 ( .A(y[892]), .B(x[892]), .Z(n16296) );
  AND U16299 ( .A(n16298), .B(n16299), .Z(n16294) );
  XNOR U16300 ( .A(y[893]), .B(x[893]), .Z(n16299) );
  XNOR U16301 ( .A(y[894]), .B(x[894]), .Z(n16298) );
  AND U16302 ( .A(n16300), .B(n16301), .Z(n16292) );
  XNOR U16303 ( .A(y[897]), .B(x[897]), .Z(n16301) );
  AND U16304 ( .A(n16302), .B(n16303), .Z(n16300) );
  XNOR U16305 ( .A(y[895]), .B(x[895]), .Z(n16303) );
  XNOR U16306 ( .A(y[896]), .B(x[896]), .Z(n16302) );
  AND U16307 ( .A(n16304), .B(n16305), .Z(n16290) );
  AND U16308 ( .A(n16306), .B(n16307), .Z(n16305) );
  AND U16309 ( .A(n16308), .B(n16309), .Z(n16307) );
  XNOR U16310 ( .A(y[898]), .B(x[898]), .Z(n16309) );
  XNOR U16311 ( .A(y[899]), .B(x[899]), .Z(n16308) );
  AND U16312 ( .A(n16310), .B(n16311), .Z(n16306) );
  XNOR U16313 ( .A(y[900]), .B(x[900]), .Z(n16311) );
  XNOR U16314 ( .A(y[901]), .B(x[901]), .Z(n16310) );
  AND U16315 ( .A(n16312), .B(n16313), .Z(n16304) );
  XNOR U16316 ( .A(y[904]), .B(x[904]), .Z(n16313) );
  AND U16317 ( .A(n16314), .B(n16315), .Z(n16312) );
  XNOR U16318 ( .A(y[902]), .B(x[902]), .Z(n16315) );
  XNOR U16319 ( .A(y[903]), .B(x[903]), .Z(n16314) );
  AND U16320 ( .A(n16316), .B(n16317), .Z(n16288) );
  AND U16321 ( .A(n16318), .B(n16319), .Z(n16317) );
  AND U16322 ( .A(n16320), .B(n16321), .Z(n16319) );
  AND U16323 ( .A(n16322), .B(n16323), .Z(n16321) );
  XNOR U16324 ( .A(y[905]), .B(x[905]), .Z(n16323) );
  XNOR U16325 ( .A(y[906]), .B(x[906]), .Z(n16322) );
  AND U16326 ( .A(n16324), .B(n16325), .Z(n16320) );
  XNOR U16327 ( .A(y[907]), .B(x[907]), .Z(n16325) );
  XNOR U16328 ( .A(y[908]), .B(x[908]), .Z(n16324) );
  AND U16329 ( .A(n16326), .B(n16327), .Z(n16318) );
  XNOR U16330 ( .A(y[911]), .B(x[911]), .Z(n16327) );
  AND U16331 ( .A(n16328), .B(n16329), .Z(n16326) );
  XNOR U16332 ( .A(y[909]), .B(x[909]), .Z(n16329) );
  XNOR U16333 ( .A(y[910]), .B(x[910]), .Z(n16328) );
  AND U16334 ( .A(n16330), .B(n16331), .Z(n16316) );
  AND U16335 ( .A(n16332), .B(n16333), .Z(n16331) );
  XNOR U16336 ( .A(y[914]), .B(x[914]), .Z(n16333) );
  AND U16337 ( .A(n16334), .B(n16335), .Z(n16332) );
  XNOR U16338 ( .A(y[912]), .B(x[912]), .Z(n16335) );
  XNOR U16339 ( .A(y[913]), .B(x[913]), .Z(n16334) );
  AND U16340 ( .A(n16336), .B(n16337), .Z(n16330) );
  XNOR U16341 ( .A(y[917]), .B(x[917]), .Z(n16337) );
  AND U16342 ( .A(n16338), .B(n16339), .Z(n16336) );
  XNOR U16343 ( .A(y[915]), .B(x[915]), .Z(n16339) );
  XNOR U16344 ( .A(y[916]), .B(x[916]), .Z(n16338) );
  AND U16345 ( .A(n16340), .B(n16341), .Z(n16286) );
  AND U16346 ( .A(n16342), .B(n16343), .Z(n16341) );
  AND U16347 ( .A(n16344), .B(n16345), .Z(n16343) );
  AND U16348 ( .A(n16346), .B(n16347), .Z(n16345) );
  AND U16349 ( .A(n16348), .B(n16349), .Z(n16347) );
  XNOR U16350 ( .A(y[918]), .B(x[918]), .Z(n16349) );
  XNOR U16351 ( .A(y[919]), .B(x[919]), .Z(n16348) );
  AND U16352 ( .A(n16350), .B(n16351), .Z(n16346) );
  XNOR U16353 ( .A(y[920]), .B(x[920]), .Z(n16351) );
  XNOR U16354 ( .A(y[921]), .B(x[921]), .Z(n16350) );
  AND U16355 ( .A(n16352), .B(n16353), .Z(n16344) );
  XNOR U16356 ( .A(y[924]), .B(x[924]), .Z(n16353) );
  AND U16357 ( .A(n16354), .B(n16355), .Z(n16352) );
  XNOR U16358 ( .A(y[922]), .B(x[922]), .Z(n16355) );
  XNOR U16359 ( .A(y[923]), .B(x[923]), .Z(n16354) );
  AND U16360 ( .A(n16356), .B(n16357), .Z(n16342) );
  AND U16361 ( .A(n16358), .B(n16359), .Z(n16357) );
  XNOR U16362 ( .A(y[927]), .B(x[927]), .Z(n16359) );
  AND U16363 ( .A(n16360), .B(n16361), .Z(n16358) );
  XNOR U16364 ( .A(y[925]), .B(x[925]), .Z(n16361) );
  XNOR U16365 ( .A(y[926]), .B(x[926]), .Z(n16360) );
  AND U16366 ( .A(n16362), .B(n16363), .Z(n16356) );
  XNOR U16367 ( .A(y[930]), .B(x[930]), .Z(n16363) );
  AND U16368 ( .A(n16364), .B(n16365), .Z(n16362) );
  XNOR U16369 ( .A(y[928]), .B(x[928]), .Z(n16365) );
  XNOR U16370 ( .A(y[929]), .B(x[929]), .Z(n16364) );
  AND U16371 ( .A(n16366), .B(n16367), .Z(n16340) );
  AND U16372 ( .A(n16368), .B(n16369), .Z(n16367) );
  AND U16373 ( .A(n16370), .B(n16371), .Z(n16369) );
  AND U16374 ( .A(n16372), .B(n16373), .Z(n16371) );
  XNOR U16375 ( .A(y[931]), .B(x[931]), .Z(n16373) );
  XNOR U16376 ( .A(y[932]), .B(x[932]), .Z(n16372) );
  AND U16377 ( .A(n16374), .B(n16375), .Z(n16370) );
  XNOR U16378 ( .A(y[933]), .B(x[933]), .Z(n16375) );
  XNOR U16379 ( .A(y[934]), .B(x[934]), .Z(n16374) );
  AND U16380 ( .A(n16376), .B(n16377), .Z(n16368) );
  XNOR U16381 ( .A(y[937]), .B(x[937]), .Z(n16377) );
  AND U16382 ( .A(n16378), .B(n16379), .Z(n16376) );
  XNOR U16383 ( .A(y[935]), .B(x[935]), .Z(n16379) );
  XNOR U16384 ( .A(y[936]), .B(x[936]), .Z(n16378) );
  AND U16385 ( .A(n16380), .B(n16381), .Z(n16366) );
  AND U16386 ( .A(n16382), .B(n16383), .Z(n16381) );
  XNOR U16387 ( .A(y[940]), .B(x[940]), .Z(n16383) );
  AND U16388 ( .A(n16384), .B(n16385), .Z(n16382) );
  XNOR U16389 ( .A(y[938]), .B(x[938]), .Z(n16385) );
  XNOR U16390 ( .A(y[939]), .B(x[939]), .Z(n16384) );
  AND U16391 ( .A(n16386), .B(n16387), .Z(n16380) );
  XNOR U16392 ( .A(y[397]), .B(x[397]), .Z(n16387) );
  AND U16393 ( .A(n16388), .B(n16389), .Z(n16386) );
  XNOR U16394 ( .A(y[941]), .B(x[941]), .Z(n16389) );
  XNOR U16395 ( .A(y[396]), .B(x[396]), .Z(n16388) );
  IV U16396 ( .A(ebreg), .Z(e) );
endmodule

