
module sum_N256_CC32 ( clk, rst, a, b, c );
  input [7:0] a;
  input [7:0] b;
  output [7:0] c;
  input clk, rst;
  wire   N18, N19, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N19), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N18), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[7]  ( .D(n32), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n31), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n30), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n29), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n28), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n27), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n26), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n25), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NANDN U35 ( .A(n64), .B(n65), .Z(n33) );
  NANDN U36 ( .A(n98), .B(n97), .Z(n34) );
  AND U37 ( .A(n33), .B(n34), .Z(n35) );
  OR U38 ( .A(n66), .B(n35), .Z(n36) );
  NAND U39 ( .A(n102), .B(n103), .Z(n37) );
  AND U40 ( .A(n36), .B(n37), .Z(n67) );
  XOR U41 ( .A(n55), .B(n54), .Z(n87) );
  AND U42 ( .A(b[7]), .B(a[7]), .Z(n72) );
  AND U43 ( .A(a[5]), .B(b[5]), .Z(n66) );
  AND U44 ( .A(a[4]), .B(b[4]), .Z(n64) );
  XNOR U45 ( .A(a[1]), .B(b[1]), .Z(n40) );
  XNOR U46 ( .A(carry_on[1]), .B(n40), .Z(n78) );
  NAND U47 ( .A(a[0]), .B(b[0]), .Z(n39) );
  XOR U48 ( .A(a[0]), .B(b[0]), .Z(n73) );
  NAND U49 ( .A(n73), .B(carry_on[0]), .Z(n38) );
  NAND U50 ( .A(n39), .B(n38), .Z(n77) );
  NAND U51 ( .A(n78), .B(n77), .Z(n42) );
  ANDN U52 ( .B(carry_on[1]), .A(n40), .Z(n43) );
  ANDN U53 ( .B(n42), .A(n43), .Z(n41) );
  NAND U54 ( .A(a[1]), .B(b[1]), .Z(n44) );
  NAND U55 ( .A(n41), .B(n44), .Z(n48) );
  XNOR U56 ( .A(n44), .B(n42), .Z(n46) );
  NAND U57 ( .A(n44), .B(n43), .Z(n45) );
  NAND U58 ( .A(n46), .B(n45), .Z(n83) );
  XNOR U59 ( .A(a[2]), .B(b[2]), .Z(n82) );
  NAND U60 ( .A(n83), .B(n82), .Z(n47) );
  NAND U61 ( .A(n48), .B(n47), .Z(n54) );
  NAND U62 ( .A(a[2]), .B(b[2]), .Z(n55) );
  AND U63 ( .A(n54), .B(n55), .Z(n50) );
  XOR U64 ( .A(a[3]), .B(b[3]), .Z(n88) );
  ANDN U65 ( .B(n87), .A(n88), .Z(n49) );
  OR U66 ( .A(n50), .B(n49), .Z(n51) );
  AND U67 ( .A(a[3]), .B(b[3]), .Z(n53) );
  ANDN U68 ( .B(n51), .A(n53), .Z(n60) );
  NOR U69 ( .A(n55), .B(n54), .Z(n52) );
  XNOR U70 ( .A(n53), .B(n52), .Z(n58) );
  XOR U71 ( .A(n55), .B(n54), .Z(n56) );
  NAND U72 ( .A(n56), .B(n88), .Z(n57) );
  NAND U73 ( .A(n58), .B(n57), .Z(n93) );
  XNOR U74 ( .A(a[4]), .B(b[4]), .Z(n92) );
  NAND U75 ( .A(n93), .B(n92), .Z(n59) );
  NANDN U76 ( .A(n60), .B(n59), .Z(n65) );
  ANDN U77 ( .B(n64), .A(n65), .Z(n61) );
  XNOR U78 ( .A(n66), .B(n61), .Z(n63) );
  XOR U79 ( .A(a[5]), .B(b[5]), .Z(n98) );
  XNOR U80 ( .A(n64), .B(n65), .Z(n97) );
  NAND U81 ( .A(n98), .B(n97), .Z(n62) );
  NAND U82 ( .A(n63), .B(n62), .Z(n103) );
  XNOR U83 ( .A(a[6]), .B(b[6]), .Z(n102) );
  NAND U84 ( .A(a[6]), .B(b[6]), .Z(n68) );
  ANDN U85 ( .B(n67), .A(n68), .Z(n71) );
  XNOR U86 ( .A(n72), .B(n71), .Z(n70) );
  XNOR U87 ( .A(n68), .B(n67), .Z(n107) );
  XOR U88 ( .A(b[7]), .B(a[7]), .Z(n108) );
  NAND U89 ( .A(n107), .B(n108), .Z(n69) );
  NAND U90 ( .A(n70), .B(n69), .Z(N18) );
  AND U91 ( .A(n72), .B(n71), .Z(N19) );
  NAND U93 ( .A(c[0]), .B(rst), .Z(n76) );
  XOR U94 ( .A(n73), .B(carry_on[0]), .Z(n74) );
  NANDN U95 ( .A(rst), .B(n74), .Z(n75) );
  NAND U96 ( .A(n76), .B(n75), .Z(n25) );
  NAND U97 ( .A(c[1]), .B(rst), .Z(n81) );
  XOR U98 ( .A(n78), .B(n77), .Z(n79) );
  NANDN U99 ( .A(rst), .B(n79), .Z(n80) );
  NAND U100 ( .A(n81), .B(n80), .Z(n26) );
  NAND U101 ( .A(c[2]), .B(rst), .Z(n86) );
  XNOR U102 ( .A(n83), .B(n82), .Z(n84) );
  NANDN U103 ( .A(rst), .B(n84), .Z(n85) );
  NAND U104 ( .A(n86), .B(n85), .Z(n27) );
  NAND U105 ( .A(c[3]), .B(rst), .Z(n91) );
  XOR U106 ( .A(n88), .B(n87), .Z(n89) );
  NANDN U107 ( .A(rst), .B(n89), .Z(n90) );
  NAND U108 ( .A(n91), .B(n90), .Z(n28) );
  NAND U109 ( .A(c[4]), .B(rst), .Z(n96) );
  XNOR U110 ( .A(n93), .B(n92), .Z(n94) );
  NANDN U111 ( .A(rst), .B(n94), .Z(n95) );
  NAND U112 ( .A(n96), .B(n95), .Z(n29) );
  NAND U113 ( .A(c[5]), .B(rst), .Z(n101) );
  XOR U114 ( .A(n98), .B(n97), .Z(n99) );
  NANDN U115 ( .A(rst), .B(n99), .Z(n100) );
  NAND U116 ( .A(n101), .B(n100), .Z(n30) );
  NAND U117 ( .A(c[6]), .B(rst), .Z(n106) );
  XNOR U118 ( .A(n103), .B(n102), .Z(n104) );
  NANDN U119 ( .A(rst), .B(n104), .Z(n105) );
  NAND U120 ( .A(n106), .B(n105), .Z(n31) );
  NAND U121 ( .A(c[7]), .B(rst), .Z(n111) );
  XOR U122 ( .A(n108), .B(n107), .Z(n109) );
  NANDN U123 ( .A(rst), .B(n109), .Z(n110) );
  NAND U124 ( .A(n111), .B(n110), .Z(n32) );
endmodule

