
module sum_N1024_CC2 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, \ADD_/c[511] , \ADD_/c[510] , \ADD_/c[509] ,
         \ADD_/c[508] , \ADD_/c[507] , \ADD_/c[506] , \ADD_/c[505] ,
         \ADD_/c[504] , \ADD_/c[503] , \ADD_/c[502] , \ADD_/c[501] ,
         \ADD_/c[500] , \ADD_/c[499] , \ADD_/c[498] , \ADD_/c[497] ,
         \ADD_/c[496] , \ADD_/c[495] , \ADD_/c[494] , \ADD_/c[493] ,
         \ADD_/c[492] , \ADD_/c[491] , \ADD_/c[490] , \ADD_/c[489] ,
         \ADD_/c[488] , \ADD_/c[487] , \ADD_/c[486] , \ADD_/c[485] ,
         \ADD_/c[484] , \ADD_/c[483] , \ADD_/c[482] , \ADD_/c[481] ,
         \ADD_/c[480] , \ADD_/c[479] , \ADD_/c[478] , \ADD_/c[477] ,
         \ADD_/c[476] , \ADD_/c[475] , \ADD_/c[474] , \ADD_/c[473] ,
         \ADD_/c[472] , \ADD_/c[471] , \ADD_/c[470] , \ADD_/c[469] ,
         \ADD_/c[468] , \ADD_/c[467] , \ADD_/c[466] , \ADD_/c[465] ,
         \ADD_/c[464] , \ADD_/c[463] , \ADD_/c[462] , \ADD_/c[461] ,
         \ADD_/c[460] , \ADD_/c[459] , \ADD_/c[458] , \ADD_/c[457] ,
         \ADD_/c[456] , \ADD_/c[455] , \ADD_/c[454] , \ADD_/c[453] ,
         \ADD_/c[452] , \ADD_/c[451] , \ADD_/c[450] , \ADD_/c[449] ,
         \ADD_/c[448] , \ADD_/c[447] , \ADD_/c[446] , \ADD_/c[445] ,
         \ADD_/c[444] , \ADD_/c[443] , \ADD_/c[442] , \ADD_/c[441] ,
         \ADD_/c[440] , \ADD_/c[439] , \ADD_/c[438] , \ADD_/c[437] ,
         \ADD_/c[436] , \ADD_/c[435] , \ADD_/c[434] , \ADD_/c[433] ,
         \ADD_/c[432] , \ADD_/c[431] , \ADD_/c[430] , \ADD_/c[429] ,
         \ADD_/c[428] , \ADD_/c[427] , \ADD_/c[426] , \ADD_/c[425] ,
         \ADD_/c[424] , \ADD_/c[423] , \ADD_/c[422] , \ADD_/c[421] ,
         \ADD_/c[420] , \ADD_/c[419] , \ADD_/c[418] , \ADD_/c[417] ,
         \ADD_/c[416] , \ADD_/c[415] , \ADD_/c[414] , \ADD_/c[413] ,
         \ADD_/c[412] , \ADD_/c[411] , \ADD_/c[410] , \ADD_/c[409] ,
         \ADD_/c[408] , \ADD_/c[407] , \ADD_/c[406] , \ADD_/c[405] ,
         \ADD_/c[404] , \ADD_/c[403] , \ADD_/c[402] , \ADD_/c[401] ,
         \ADD_/c[400] , \ADD_/c[399] , \ADD_/c[398] , \ADD_/c[397] ,
         \ADD_/c[396] , \ADD_/c[395] , \ADD_/c[394] , \ADD_/c[393] ,
         \ADD_/c[392] , \ADD_/c[391] , \ADD_/c[390] , \ADD_/c[389] ,
         \ADD_/c[388] , \ADD_/c[387] , \ADD_/c[386] , \ADD_/c[385] ,
         \ADD_/c[384] , \ADD_/c[383] , \ADD_/c[382] , \ADD_/c[381] ,
         \ADD_/c[380] , \ADD_/c[379] , \ADD_/c[378] , \ADD_/c[377] ,
         \ADD_/c[376] , \ADD_/c[375] , \ADD_/c[374] , \ADD_/c[373] ,
         \ADD_/c[372] , \ADD_/c[371] , \ADD_/c[370] , \ADD_/c[369] ,
         \ADD_/c[368] , \ADD_/c[367] , \ADD_/c[366] , \ADD_/c[365] ,
         \ADD_/c[364] , \ADD_/c[363] , \ADD_/c[362] , \ADD_/c[361] ,
         \ADD_/c[360] , \ADD_/c[359] , \ADD_/c[358] , \ADD_/c[357] ,
         \ADD_/c[356] , \ADD_/c[355] , \ADD_/c[354] , \ADD_/c[353] ,
         \ADD_/c[352] , \ADD_/c[351] , \ADD_/c[350] , \ADD_/c[349] ,
         \ADD_/c[348] , \ADD_/c[347] , \ADD_/c[346] , \ADD_/c[345] ,
         \ADD_/c[344] , \ADD_/c[343] , \ADD_/c[342] , \ADD_/c[341] ,
         \ADD_/c[340] , \ADD_/c[339] , \ADD_/c[338] , \ADD_/c[337] ,
         \ADD_/c[336] , \ADD_/c[335] , \ADD_/c[334] , \ADD_/c[333] ,
         \ADD_/c[332] , \ADD_/c[331] , \ADD_/c[330] , \ADD_/c[329] ,
         \ADD_/c[328] , \ADD_/c[327] , \ADD_/c[326] , \ADD_/c[325] ,
         \ADD_/c[324] , \ADD_/c[323] , \ADD_/c[322] , \ADD_/c[321] ,
         \ADD_/c[320] , \ADD_/c[319] , \ADD_/c[318] , \ADD_/c[317] ,
         \ADD_/c[316] , \ADD_/c[315] , \ADD_/c[314] , \ADD_/c[313] ,
         \ADD_/c[312] , \ADD_/c[311] , \ADD_/c[310] , \ADD_/c[309] ,
         \ADD_/c[308] , \ADD_/c[307] , \ADD_/c[306] , \ADD_/c[305] ,
         \ADD_/c[304] , \ADD_/c[303] , \ADD_/c[302] , \ADD_/c[301] ,
         \ADD_/c[300] , \ADD_/c[299] , \ADD_/c[298] , \ADD_/c[297] ,
         \ADD_/c[296] , \ADD_/c[295] , \ADD_/c[294] , \ADD_/c[293] ,
         \ADD_/c[292] , \ADD_/c[291] , \ADD_/c[290] , \ADD_/c[289] ,
         \ADD_/c[288] , \ADD_/c[287] , \ADD_/c[286] , \ADD_/c[285] ,
         \ADD_/c[284] , \ADD_/c[283] , \ADD_/c[282] , \ADD_/c[281] ,
         \ADD_/c[280] , \ADD_/c[279] , \ADD_/c[278] , \ADD_/c[277] ,
         \ADD_/c[276] , \ADD_/c[275] , \ADD_/c[274] , \ADD_/c[273] ,
         \ADD_/c[272] , \ADD_/c[271] , \ADD_/c[270] , \ADD_/c[269] ,
         \ADD_/c[268] , \ADD_/c[267] , \ADD_/c[266] , \ADD_/c[265] ,
         \ADD_/c[264] , \ADD_/c[263] , \ADD_/c[262] , \ADD_/c[261] ,
         \ADD_/c[260] , \ADD_/c[259] , \ADD_/c[258] , \ADD_/c[257] ,
         \ADD_/c[256] , \ADD_/c[255] , \ADD_/c[254] , \ADD_/c[253] ,
         \ADD_/c[252] , \ADD_/c[251] , \ADD_/c[250] , \ADD_/c[249] ,
         \ADD_/c[248] , \ADD_/c[247] , \ADD_/c[246] , \ADD_/c[245] ,
         \ADD_/c[244] , \ADD_/c[243] , \ADD_/c[242] , \ADD_/c[241] ,
         \ADD_/c[240] , \ADD_/c[239] , \ADD_/c[238] , \ADD_/c[237] ,
         \ADD_/c[236] , \ADD_/c[235] , \ADD_/c[234] , \ADD_/c[233] ,
         \ADD_/c[232] , \ADD_/c[231] , \ADD_/c[230] , \ADD_/c[229] ,
         \ADD_/c[228] , \ADD_/c[227] , \ADD_/c[226] , \ADD_/c[225] ,
         \ADD_/c[224] , \ADD_/c[223] , \ADD_/c[222] , \ADD_/c[221] ,
         \ADD_/c[220] , \ADD_/c[219] , \ADD_/c[218] , \ADD_/c[217] ,
         \ADD_/c[216] , \ADD_/c[215] , \ADD_/c[214] , \ADD_/c[213] ,
         \ADD_/c[212] , \ADD_/c[211] , \ADD_/c[210] , \ADD_/c[209] ,
         \ADD_/c[208] , \ADD_/c[207] , \ADD_/c[206] , \ADD_/c[205] ,
         \ADD_/c[204] , \ADD_/c[203] , \ADD_/c[202] , \ADD_/c[201] ,
         \ADD_/c[200] , \ADD_/c[199] , \ADD_/c[198] , \ADD_/c[197] ,
         \ADD_/c[196] , \ADD_/c[195] , \ADD_/c[194] , \ADD_/c[193] ,
         \ADD_/c[192] , \ADD_/c[191] , \ADD_/c[190] , \ADD_/c[189] ,
         \ADD_/c[188] , \ADD_/c[187] , \ADD_/c[186] , \ADD_/c[185] ,
         \ADD_/c[184] , \ADD_/c[183] , \ADD_/c[182] , \ADD_/c[181] ,
         \ADD_/c[180] , \ADD_/c[179] , \ADD_/c[178] , \ADD_/c[177] ,
         \ADD_/c[176] , \ADD_/c[175] , \ADD_/c[174] , \ADD_/c[173] ,
         \ADD_/c[172] , \ADD_/c[171] , \ADD_/c[170] , \ADD_/c[169] ,
         \ADD_/c[168] , \ADD_/c[167] , \ADD_/c[166] , \ADD_/c[165] ,
         \ADD_/c[164] , \ADD_/c[163] , \ADD_/c[162] , \ADD_/c[161] ,
         \ADD_/c[160] , \ADD_/c[159] , \ADD_/c[158] , \ADD_/c[157] ,
         \ADD_/c[156] , \ADD_/c[155] , \ADD_/c[154] , \ADD_/c[153] ,
         \ADD_/c[152] , \ADD_/c[151] , \ADD_/c[150] , \ADD_/c[149] ,
         \ADD_/c[148] , \ADD_/c[147] , \ADD_/c[146] , \ADD_/c[145] ,
         \ADD_/c[144] , \ADD_/c[143] , \ADD_/c[142] , \ADD_/c[141] ,
         \ADD_/c[140] , \ADD_/c[139] , \ADD_/c[138] , \ADD_/c[137] ,
         \ADD_/c[136] , \ADD_/c[135] , \ADD_/c[134] , \ADD_/c[133] ,
         \ADD_/c[132] , \ADD_/c[131] , \ADD_/c[130] , \ADD_/c[129] ,
         \ADD_/c[128] , \ADD_/c[127] , \ADD_/c[126] , \ADD_/c[125] ,
         \ADD_/c[124] , \ADD_/c[123] , \ADD_/c[122] , \ADD_/c[121] ,
         \ADD_/c[120] , \ADD_/c[119] , \ADD_/c[118] , \ADD_/c[117] ,
         \ADD_/c[116] , \ADD_/c[115] , \ADD_/c[114] , \ADD_/c[113] ,
         \ADD_/c[112] , \ADD_/c[111] , \ADD_/c[110] , \ADD_/c[109] ,
         \ADD_/c[108] , \ADD_/c[107] , \ADD_/c[106] , \ADD_/c[105] ,
         \ADD_/c[104] , \ADD_/c[103] , \ADD_/c[102] , \ADD_/c[101] ,
         \ADD_/c[100] , \ADD_/c[99] , \ADD_/c[98] , \ADD_/c[97] , \ADD_/c[96] ,
         \ADD_/c[95] , \ADD_/c[94] , \ADD_/c[93] , \ADD_/c[92] , \ADD_/c[91] ,
         \ADD_/c[90] , \ADD_/c[89] , \ADD_/c[88] , \ADD_/c[87] , \ADD_/c[86] ,
         \ADD_/c[85] , \ADD_/c[84] , \ADD_/c[83] , \ADD_/c[82] , \ADD_/c[81] ,
         \ADD_/c[80] , \ADD_/c[79] , \ADD_/c[78] , \ADD_/c[77] , \ADD_/c[76] ,
         \ADD_/c[75] , \ADD_/c[74] , \ADD_/c[73] , \ADD_/c[72] , \ADD_/c[71] ,
         \ADD_/c[70] , \ADD_/c[69] , \ADD_/c[68] , \ADD_/c[67] , \ADD_/c[66] ,
         \ADD_/c[65] , \ADD_/c[64] , \ADD_/c[63] , \ADD_/c[62] , \ADD_/c[61] ,
         \ADD_/c[60] , \ADD_/c[59] , \ADD_/c[58] , \ADD_/c[57] , \ADD_/c[56] ,
         \ADD_/c[55] , \ADD_/c[54] , \ADD_/c[53] , \ADD_/c[52] , \ADD_/c[51] ,
         \ADD_/c[50] , \ADD_/c[49] , \ADD_/c[48] , \ADD_/c[47] , \ADD_/c[46] ,
         \ADD_/c[45] , \ADD_/c[44] , \ADD_/c[43] , \ADD_/c[42] , \ADD_/c[41] ,
         \ADD_/c[40] , \ADD_/c[39] , \ADD_/c[38] , \ADD_/c[37] , \ADD_/c[36] ,
         \ADD_/c[35] , \ADD_/c[34] , \ADD_/c[33] , \ADD_/c[32] , \ADD_/c[31] ,
         \ADD_/c[30] , \ADD_/c[29] , \ADD_/c[28] , \ADD_/c[27] , \ADD_/c[26] ,
         \ADD_/c[25] , \ADD_/c[24] , \ADD_/c[23] , \ADD_/c[22] , \ADD_/c[21] ,
         \ADD_/c[20] , \ADD_/c[19] , \ADD_/c[18] , \ADD_/c[17] , \ADD_/c[16] ,
         \ADD_/c[15] , \ADD_/c[14] , \ADD_/c[13] , \ADD_/c[12] , \ADD_/c[11] ,
         \ADD_/c[10] , \ADD_/c[9] , \ADD_/c[8] , \ADD_/c[7] , \ADD_/c[6] ,
         \ADD_/c[5] , \ADD_/c[4] , \ADD_/c[3] , \ADD_/c[2] , \ADD_/c[1] ,
         \ADD_/FAINST[0].FA_/n3 , \ADD_/FAINST[0].FA_/n2 ,
         \ADD_/FAINST[0].FA_/n1 , \ADD_/FAINST[511].FA_/n3 ,
         \ADD_/FAINST[511].FA_/n2 , \ADD_/FAINST[511].FA_/n1 ,
         \ADD_/FAINST[510].FA_/n3 , \ADD_/FAINST[510].FA_/n2 ,
         \ADD_/FAINST[510].FA_/n1 , \ADD_/FAINST[509].FA_/n3 ,
         \ADD_/FAINST[509].FA_/n2 , \ADD_/FAINST[509].FA_/n1 ,
         \ADD_/FAINST[508].FA_/n3 , \ADD_/FAINST[508].FA_/n2 ,
         \ADD_/FAINST[508].FA_/n1 , \ADD_/FAINST[507].FA_/n3 ,
         \ADD_/FAINST[507].FA_/n2 , \ADD_/FAINST[507].FA_/n1 ,
         \ADD_/FAINST[506].FA_/n3 , \ADD_/FAINST[506].FA_/n2 ,
         \ADD_/FAINST[506].FA_/n1 , \ADD_/FAINST[505].FA_/n3 ,
         \ADD_/FAINST[505].FA_/n2 , \ADD_/FAINST[505].FA_/n1 ,
         \ADD_/FAINST[504].FA_/n3 , \ADD_/FAINST[504].FA_/n2 ,
         \ADD_/FAINST[504].FA_/n1 , \ADD_/FAINST[503].FA_/n3 ,
         \ADD_/FAINST[503].FA_/n2 , \ADD_/FAINST[503].FA_/n1 ,
         \ADD_/FAINST[502].FA_/n3 , \ADD_/FAINST[502].FA_/n2 ,
         \ADD_/FAINST[502].FA_/n1 , \ADD_/FAINST[501].FA_/n3 ,
         \ADD_/FAINST[501].FA_/n2 , \ADD_/FAINST[501].FA_/n1 ,
         \ADD_/FAINST[500].FA_/n3 , \ADD_/FAINST[500].FA_/n2 ,
         \ADD_/FAINST[500].FA_/n1 , \ADD_/FAINST[499].FA_/n3 ,
         \ADD_/FAINST[499].FA_/n2 , \ADD_/FAINST[499].FA_/n1 ,
         \ADD_/FAINST[498].FA_/n3 , \ADD_/FAINST[498].FA_/n2 ,
         \ADD_/FAINST[498].FA_/n1 , \ADD_/FAINST[497].FA_/n3 ,
         \ADD_/FAINST[497].FA_/n2 , \ADD_/FAINST[497].FA_/n1 ,
         \ADD_/FAINST[496].FA_/n3 , \ADD_/FAINST[496].FA_/n2 ,
         \ADD_/FAINST[496].FA_/n1 , \ADD_/FAINST[495].FA_/n3 ,
         \ADD_/FAINST[495].FA_/n2 , \ADD_/FAINST[495].FA_/n1 ,
         \ADD_/FAINST[494].FA_/n3 , \ADD_/FAINST[494].FA_/n2 ,
         \ADD_/FAINST[494].FA_/n1 , \ADD_/FAINST[493].FA_/n3 ,
         \ADD_/FAINST[493].FA_/n2 , \ADD_/FAINST[493].FA_/n1 ,
         \ADD_/FAINST[492].FA_/n3 , \ADD_/FAINST[492].FA_/n2 ,
         \ADD_/FAINST[492].FA_/n1 , \ADD_/FAINST[491].FA_/n3 ,
         \ADD_/FAINST[491].FA_/n2 , \ADD_/FAINST[491].FA_/n1 ,
         \ADD_/FAINST[490].FA_/n3 , \ADD_/FAINST[490].FA_/n2 ,
         \ADD_/FAINST[490].FA_/n1 , \ADD_/FAINST[489].FA_/n3 ,
         \ADD_/FAINST[489].FA_/n2 , \ADD_/FAINST[489].FA_/n1 ,
         \ADD_/FAINST[488].FA_/n3 , \ADD_/FAINST[488].FA_/n2 ,
         \ADD_/FAINST[488].FA_/n1 , \ADD_/FAINST[487].FA_/n3 ,
         \ADD_/FAINST[487].FA_/n2 , \ADD_/FAINST[487].FA_/n1 ,
         \ADD_/FAINST[486].FA_/n3 , \ADD_/FAINST[486].FA_/n2 ,
         \ADD_/FAINST[486].FA_/n1 , \ADD_/FAINST[485].FA_/n3 ,
         \ADD_/FAINST[485].FA_/n2 , \ADD_/FAINST[485].FA_/n1 ,
         \ADD_/FAINST[484].FA_/n3 , \ADD_/FAINST[484].FA_/n2 ,
         \ADD_/FAINST[484].FA_/n1 , \ADD_/FAINST[483].FA_/n3 ,
         \ADD_/FAINST[483].FA_/n2 , \ADD_/FAINST[483].FA_/n1 ,
         \ADD_/FAINST[482].FA_/n3 , \ADD_/FAINST[482].FA_/n2 ,
         \ADD_/FAINST[482].FA_/n1 , \ADD_/FAINST[481].FA_/n3 ,
         \ADD_/FAINST[481].FA_/n2 , \ADD_/FAINST[481].FA_/n1 ,
         \ADD_/FAINST[480].FA_/n3 , \ADD_/FAINST[480].FA_/n2 ,
         \ADD_/FAINST[480].FA_/n1 , \ADD_/FAINST[479].FA_/n3 ,
         \ADD_/FAINST[479].FA_/n2 , \ADD_/FAINST[479].FA_/n1 ,
         \ADD_/FAINST[478].FA_/n3 , \ADD_/FAINST[478].FA_/n2 ,
         \ADD_/FAINST[478].FA_/n1 , \ADD_/FAINST[477].FA_/n3 ,
         \ADD_/FAINST[477].FA_/n2 , \ADD_/FAINST[477].FA_/n1 ,
         \ADD_/FAINST[476].FA_/n3 , \ADD_/FAINST[476].FA_/n2 ,
         \ADD_/FAINST[476].FA_/n1 , \ADD_/FAINST[475].FA_/n3 ,
         \ADD_/FAINST[475].FA_/n2 , \ADD_/FAINST[475].FA_/n1 ,
         \ADD_/FAINST[474].FA_/n3 , \ADD_/FAINST[474].FA_/n2 ,
         \ADD_/FAINST[474].FA_/n1 , \ADD_/FAINST[473].FA_/n3 ,
         \ADD_/FAINST[473].FA_/n2 , \ADD_/FAINST[473].FA_/n1 ,
         \ADD_/FAINST[472].FA_/n3 , \ADD_/FAINST[472].FA_/n2 ,
         \ADD_/FAINST[472].FA_/n1 , \ADD_/FAINST[471].FA_/n3 ,
         \ADD_/FAINST[471].FA_/n2 , \ADD_/FAINST[471].FA_/n1 ,
         \ADD_/FAINST[470].FA_/n3 , \ADD_/FAINST[470].FA_/n2 ,
         \ADD_/FAINST[470].FA_/n1 , \ADD_/FAINST[469].FA_/n3 ,
         \ADD_/FAINST[469].FA_/n2 , \ADD_/FAINST[469].FA_/n1 ,
         \ADD_/FAINST[468].FA_/n3 , \ADD_/FAINST[468].FA_/n2 ,
         \ADD_/FAINST[468].FA_/n1 , \ADD_/FAINST[467].FA_/n3 ,
         \ADD_/FAINST[467].FA_/n2 , \ADD_/FAINST[467].FA_/n1 ,
         \ADD_/FAINST[466].FA_/n3 , \ADD_/FAINST[466].FA_/n2 ,
         \ADD_/FAINST[466].FA_/n1 , \ADD_/FAINST[465].FA_/n3 ,
         \ADD_/FAINST[465].FA_/n2 , \ADD_/FAINST[465].FA_/n1 ,
         \ADD_/FAINST[464].FA_/n3 , \ADD_/FAINST[464].FA_/n2 ,
         \ADD_/FAINST[464].FA_/n1 , \ADD_/FAINST[463].FA_/n3 ,
         \ADD_/FAINST[463].FA_/n2 , \ADD_/FAINST[463].FA_/n1 ,
         \ADD_/FAINST[462].FA_/n3 , \ADD_/FAINST[462].FA_/n2 ,
         \ADD_/FAINST[462].FA_/n1 , \ADD_/FAINST[461].FA_/n3 ,
         \ADD_/FAINST[461].FA_/n2 , \ADD_/FAINST[461].FA_/n1 ,
         \ADD_/FAINST[460].FA_/n3 , \ADD_/FAINST[460].FA_/n2 ,
         \ADD_/FAINST[460].FA_/n1 , \ADD_/FAINST[459].FA_/n3 ,
         \ADD_/FAINST[459].FA_/n2 , \ADD_/FAINST[459].FA_/n1 ,
         \ADD_/FAINST[458].FA_/n3 , \ADD_/FAINST[458].FA_/n2 ,
         \ADD_/FAINST[458].FA_/n1 , \ADD_/FAINST[457].FA_/n3 ,
         \ADD_/FAINST[457].FA_/n2 , \ADD_/FAINST[457].FA_/n1 ,
         \ADD_/FAINST[456].FA_/n3 , \ADD_/FAINST[456].FA_/n2 ,
         \ADD_/FAINST[456].FA_/n1 , \ADD_/FAINST[455].FA_/n3 ,
         \ADD_/FAINST[455].FA_/n2 , \ADD_/FAINST[455].FA_/n1 ,
         \ADD_/FAINST[454].FA_/n3 , \ADD_/FAINST[454].FA_/n2 ,
         \ADD_/FAINST[454].FA_/n1 , \ADD_/FAINST[453].FA_/n3 ,
         \ADD_/FAINST[453].FA_/n2 , \ADD_/FAINST[453].FA_/n1 ,
         \ADD_/FAINST[452].FA_/n3 , \ADD_/FAINST[452].FA_/n2 ,
         \ADD_/FAINST[452].FA_/n1 , \ADD_/FAINST[451].FA_/n3 ,
         \ADD_/FAINST[451].FA_/n2 , \ADD_/FAINST[451].FA_/n1 ,
         \ADD_/FAINST[450].FA_/n3 , \ADD_/FAINST[450].FA_/n2 ,
         \ADD_/FAINST[450].FA_/n1 , \ADD_/FAINST[449].FA_/n3 ,
         \ADD_/FAINST[449].FA_/n2 , \ADD_/FAINST[449].FA_/n1 ,
         \ADD_/FAINST[448].FA_/n3 , \ADD_/FAINST[448].FA_/n2 ,
         \ADD_/FAINST[448].FA_/n1 , \ADD_/FAINST[447].FA_/n3 ,
         \ADD_/FAINST[447].FA_/n2 , \ADD_/FAINST[447].FA_/n1 ,
         \ADD_/FAINST[446].FA_/n3 , \ADD_/FAINST[446].FA_/n2 ,
         \ADD_/FAINST[446].FA_/n1 , \ADD_/FAINST[445].FA_/n3 ,
         \ADD_/FAINST[445].FA_/n2 , \ADD_/FAINST[445].FA_/n1 ,
         \ADD_/FAINST[444].FA_/n3 , \ADD_/FAINST[444].FA_/n2 ,
         \ADD_/FAINST[444].FA_/n1 , \ADD_/FAINST[443].FA_/n3 ,
         \ADD_/FAINST[443].FA_/n2 , \ADD_/FAINST[443].FA_/n1 ,
         \ADD_/FAINST[442].FA_/n3 , \ADD_/FAINST[442].FA_/n2 ,
         \ADD_/FAINST[442].FA_/n1 , \ADD_/FAINST[441].FA_/n3 ,
         \ADD_/FAINST[441].FA_/n2 , \ADD_/FAINST[441].FA_/n1 ,
         \ADD_/FAINST[440].FA_/n3 , \ADD_/FAINST[440].FA_/n2 ,
         \ADD_/FAINST[440].FA_/n1 , \ADD_/FAINST[439].FA_/n3 ,
         \ADD_/FAINST[439].FA_/n2 , \ADD_/FAINST[439].FA_/n1 ,
         \ADD_/FAINST[438].FA_/n3 , \ADD_/FAINST[438].FA_/n2 ,
         \ADD_/FAINST[438].FA_/n1 , \ADD_/FAINST[437].FA_/n3 ,
         \ADD_/FAINST[437].FA_/n2 , \ADD_/FAINST[437].FA_/n1 ,
         \ADD_/FAINST[436].FA_/n3 , \ADD_/FAINST[436].FA_/n2 ,
         \ADD_/FAINST[436].FA_/n1 , \ADD_/FAINST[435].FA_/n3 ,
         \ADD_/FAINST[435].FA_/n2 , \ADD_/FAINST[435].FA_/n1 ,
         \ADD_/FAINST[434].FA_/n3 , \ADD_/FAINST[434].FA_/n2 ,
         \ADD_/FAINST[434].FA_/n1 , \ADD_/FAINST[433].FA_/n3 ,
         \ADD_/FAINST[433].FA_/n2 , \ADD_/FAINST[433].FA_/n1 ,
         \ADD_/FAINST[432].FA_/n3 , \ADD_/FAINST[432].FA_/n2 ,
         \ADD_/FAINST[432].FA_/n1 , \ADD_/FAINST[431].FA_/n3 ,
         \ADD_/FAINST[431].FA_/n2 , \ADD_/FAINST[431].FA_/n1 ,
         \ADD_/FAINST[430].FA_/n3 , \ADD_/FAINST[430].FA_/n2 ,
         \ADD_/FAINST[430].FA_/n1 , \ADD_/FAINST[429].FA_/n3 ,
         \ADD_/FAINST[429].FA_/n2 , \ADD_/FAINST[429].FA_/n1 ,
         \ADD_/FAINST[428].FA_/n3 , \ADD_/FAINST[428].FA_/n2 ,
         \ADD_/FAINST[428].FA_/n1 , \ADD_/FAINST[427].FA_/n3 ,
         \ADD_/FAINST[427].FA_/n2 , \ADD_/FAINST[427].FA_/n1 ,
         \ADD_/FAINST[426].FA_/n3 , \ADD_/FAINST[426].FA_/n2 ,
         \ADD_/FAINST[426].FA_/n1 , \ADD_/FAINST[425].FA_/n3 ,
         \ADD_/FAINST[425].FA_/n2 , \ADD_/FAINST[425].FA_/n1 ,
         \ADD_/FAINST[424].FA_/n3 , \ADD_/FAINST[424].FA_/n2 ,
         \ADD_/FAINST[424].FA_/n1 , \ADD_/FAINST[423].FA_/n3 ,
         \ADD_/FAINST[423].FA_/n2 , \ADD_/FAINST[423].FA_/n1 ,
         \ADD_/FAINST[422].FA_/n3 , \ADD_/FAINST[422].FA_/n2 ,
         \ADD_/FAINST[422].FA_/n1 , \ADD_/FAINST[421].FA_/n3 ,
         \ADD_/FAINST[421].FA_/n2 , \ADD_/FAINST[421].FA_/n1 ,
         \ADD_/FAINST[420].FA_/n3 , \ADD_/FAINST[420].FA_/n2 ,
         \ADD_/FAINST[420].FA_/n1 , \ADD_/FAINST[419].FA_/n3 ,
         \ADD_/FAINST[419].FA_/n2 , \ADD_/FAINST[419].FA_/n1 ,
         \ADD_/FAINST[418].FA_/n3 , \ADD_/FAINST[418].FA_/n2 ,
         \ADD_/FAINST[418].FA_/n1 , \ADD_/FAINST[417].FA_/n3 ,
         \ADD_/FAINST[417].FA_/n2 , \ADD_/FAINST[417].FA_/n1 ,
         \ADD_/FAINST[416].FA_/n3 , \ADD_/FAINST[416].FA_/n2 ,
         \ADD_/FAINST[416].FA_/n1 , \ADD_/FAINST[415].FA_/n3 ,
         \ADD_/FAINST[415].FA_/n2 , \ADD_/FAINST[415].FA_/n1 ,
         \ADD_/FAINST[414].FA_/n3 , \ADD_/FAINST[414].FA_/n2 ,
         \ADD_/FAINST[414].FA_/n1 , \ADD_/FAINST[413].FA_/n3 ,
         \ADD_/FAINST[413].FA_/n2 , \ADD_/FAINST[413].FA_/n1 ,
         \ADD_/FAINST[412].FA_/n3 , \ADD_/FAINST[412].FA_/n2 ,
         \ADD_/FAINST[412].FA_/n1 , \ADD_/FAINST[411].FA_/n3 ,
         \ADD_/FAINST[411].FA_/n2 , \ADD_/FAINST[411].FA_/n1 ,
         \ADD_/FAINST[410].FA_/n3 , \ADD_/FAINST[410].FA_/n2 ,
         \ADD_/FAINST[410].FA_/n1 , \ADD_/FAINST[409].FA_/n3 ,
         \ADD_/FAINST[409].FA_/n2 , \ADD_/FAINST[409].FA_/n1 ,
         \ADD_/FAINST[408].FA_/n3 , \ADD_/FAINST[408].FA_/n2 ,
         \ADD_/FAINST[408].FA_/n1 , \ADD_/FAINST[407].FA_/n3 ,
         \ADD_/FAINST[407].FA_/n2 , \ADD_/FAINST[407].FA_/n1 ,
         \ADD_/FAINST[406].FA_/n3 , \ADD_/FAINST[406].FA_/n2 ,
         \ADD_/FAINST[406].FA_/n1 , \ADD_/FAINST[405].FA_/n3 ,
         \ADD_/FAINST[405].FA_/n2 , \ADD_/FAINST[405].FA_/n1 ,
         \ADD_/FAINST[404].FA_/n3 , \ADD_/FAINST[404].FA_/n2 ,
         \ADD_/FAINST[404].FA_/n1 , \ADD_/FAINST[403].FA_/n3 ,
         \ADD_/FAINST[403].FA_/n2 , \ADD_/FAINST[403].FA_/n1 ,
         \ADD_/FAINST[402].FA_/n3 , \ADD_/FAINST[402].FA_/n2 ,
         \ADD_/FAINST[402].FA_/n1 , \ADD_/FAINST[401].FA_/n3 ,
         \ADD_/FAINST[401].FA_/n2 , \ADD_/FAINST[401].FA_/n1 ,
         \ADD_/FAINST[400].FA_/n3 , \ADD_/FAINST[400].FA_/n2 ,
         \ADD_/FAINST[400].FA_/n1 , \ADD_/FAINST[399].FA_/n3 ,
         \ADD_/FAINST[399].FA_/n2 , \ADD_/FAINST[399].FA_/n1 ,
         \ADD_/FAINST[398].FA_/n3 , \ADD_/FAINST[398].FA_/n2 ,
         \ADD_/FAINST[398].FA_/n1 , \ADD_/FAINST[397].FA_/n3 ,
         \ADD_/FAINST[397].FA_/n2 , \ADD_/FAINST[397].FA_/n1 ,
         \ADD_/FAINST[396].FA_/n3 , \ADD_/FAINST[396].FA_/n2 ,
         \ADD_/FAINST[396].FA_/n1 , \ADD_/FAINST[395].FA_/n3 ,
         \ADD_/FAINST[395].FA_/n2 , \ADD_/FAINST[395].FA_/n1 ,
         \ADD_/FAINST[394].FA_/n3 , \ADD_/FAINST[394].FA_/n2 ,
         \ADD_/FAINST[394].FA_/n1 , \ADD_/FAINST[393].FA_/n3 ,
         \ADD_/FAINST[393].FA_/n2 , \ADD_/FAINST[393].FA_/n1 ,
         \ADD_/FAINST[392].FA_/n3 , \ADD_/FAINST[392].FA_/n2 ,
         \ADD_/FAINST[392].FA_/n1 , \ADD_/FAINST[391].FA_/n3 ,
         \ADD_/FAINST[391].FA_/n2 , \ADD_/FAINST[391].FA_/n1 ,
         \ADD_/FAINST[390].FA_/n3 , \ADD_/FAINST[390].FA_/n2 ,
         \ADD_/FAINST[390].FA_/n1 , \ADD_/FAINST[389].FA_/n3 ,
         \ADD_/FAINST[389].FA_/n2 , \ADD_/FAINST[389].FA_/n1 ,
         \ADD_/FAINST[388].FA_/n3 , \ADD_/FAINST[388].FA_/n2 ,
         \ADD_/FAINST[388].FA_/n1 , \ADD_/FAINST[387].FA_/n3 ,
         \ADD_/FAINST[387].FA_/n2 , \ADD_/FAINST[387].FA_/n1 ,
         \ADD_/FAINST[386].FA_/n3 , \ADD_/FAINST[386].FA_/n2 ,
         \ADD_/FAINST[386].FA_/n1 , \ADD_/FAINST[385].FA_/n3 ,
         \ADD_/FAINST[385].FA_/n2 , \ADD_/FAINST[385].FA_/n1 ,
         \ADD_/FAINST[384].FA_/n3 , \ADD_/FAINST[384].FA_/n2 ,
         \ADD_/FAINST[384].FA_/n1 , \ADD_/FAINST[383].FA_/n3 ,
         \ADD_/FAINST[383].FA_/n2 , \ADD_/FAINST[383].FA_/n1 ,
         \ADD_/FAINST[382].FA_/n3 , \ADD_/FAINST[382].FA_/n2 ,
         \ADD_/FAINST[382].FA_/n1 , \ADD_/FAINST[381].FA_/n3 ,
         \ADD_/FAINST[381].FA_/n2 , \ADD_/FAINST[381].FA_/n1 ,
         \ADD_/FAINST[380].FA_/n3 , \ADD_/FAINST[380].FA_/n2 ,
         \ADD_/FAINST[380].FA_/n1 , \ADD_/FAINST[379].FA_/n3 ,
         \ADD_/FAINST[379].FA_/n2 , \ADD_/FAINST[379].FA_/n1 ,
         \ADD_/FAINST[378].FA_/n3 , \ADD_/FAINST[378].FA_/n2 ,
         \ADD_/FAINST[378].FA_/n1 , \ADD_/FAINST[377].FA_/n3 ,
         \ADD_/FAINST[377].FA_/n2 , \ADD_/FAINST[377].FA_/n1 ,
         \ADD_/FAINST[376].FA_/n3 , \ADD_/FAINST[376].FA_/n2 ,
         \ADD_/FAINST[376].FA_/n1 , \ADD_/FAINST[375].FA_/n3 ,
         \ADD_/FAINST[375].FA_/n2 , \ADD_/FAINST[375].FA_/n1 ,
         \ADD_/FAINST[374].FA_/n3 , \ADD_/FAINST[374].FA_/n2 ,
         \ADD_/FAINST[374].FA_/n1 , \ADD_/FAINST[373].FA_/n3 ,
         \ADD_/FAINST[373].FA_/n2 , \ADD_/FAINST[373].FA_/n1 ,
         \ADD_/FAINST[372].FA_/n3 , \ADD_/FAINST[372].FA_/n2 ,
         \ADD_/FAINST[372].FA_/n1 , \ADD_/FAINST[371].FA_/n3 ,
         \ADD_/FAINST[371].FA_/n2 , \ADD_/FAINST[371].FA_/n1 ,
         \ADD_/FAINST[370].FA_/n3 , \ADD_/FAINST[370].FA_/n2 ,
         \ADD_/FAINST[370].FA_/n1 , \ADD_/FAINST[369].FA_/n3 ,
         \ADD_/FAINST[369].FA_/n2 , \ADD_/FAINST[369].FA_/n1 ,
         \ADD_/FAINST[368].FA_/n3 , \ADD_/FAINST[368].FA_/n2 ,
         \ADD_/FAINST[368].FA_/n1 , \ADD_/FAINST[367].FA_/n3 ,
         \ADD_/FAINST[367].FA_/n2 , \ADD_/FAINST[367].FA_/n1 ,
         \ADD_/FAINST[366].FA_/n3 , \ADD_/FAINST[366].FA_/n2 ,
         \ADD_/FAINST[366].FA_/n1 , \ADD_/FAINST[365].FA_/n3 ,
         \ADD_/FAINST[365].FA_/n2 , \ADD_/FAINST[365].FA_/n1 ,
         \ADD_/FAINST[364].FA_/n3 , \ADD_/FAINST[364].FA_/n2 ,
         \ADD_/FAINST[364].FA_/n1 , \ADD_/FAINST[363].FA_/n3 ,
         \ADD_/FAINST[363].FA_/n2 , \ADD_/FAINST[363].FA_/n1 ,
         \ADD_/FAINST[362].FA_/n3 , \ADD_/FAINST[362].FA_/n2 ,
         \ADD_/FAINST[362].FA_/n1 , \ADD_/FAINST[361].FA_/n3 ,
         \ADD_/FAINST[361].FA_/n2 , \ADD_/FAINST[361].FA_/n1 ,
         \ADD_/FAINST[360].FA_/n3 , \ADD_/FAINST[360].FA_/n2 ,
         \ADD_/FAINST[360].FA_/n1 , \ADD_/FAINST[359].FA_/n3 ,
         \ADD_/FAINST[359].FA_/n2 , \ADD_/FAINST[359].FA_/n1 ,
         \ADD_/FAINST[358].FA_/n3 , \ADD_/FAINST[358].FA_/n2 ,
         \ADD_/FAINST[358].FA_/n1 , \ADD_/FAINST[357].FA_/n3 ,
         \ADD_/FAINST[357].FA_/n2 , \ADD_/FAINST[357].FA_/n1 ,
         \ADD_/FAINST[356].FA_/n3 , \ADD_/FAINST[356].FA_/n2 ,
         \ADD_/FAINST[356].FA_/n1 , \ADD_/FAINST[355].FA_/n3 ,
         \ADD_/FAINST[355].FA_/n2 , \ADD_/FAINST[355].FA_/n1 ,
         \ADD_/FAINST[354].FA_/n3 , \ADD_/FAINST[354].FA_/n2 ,
         \ADD_/FAINST[354].FA_/n1 , \ADD_/FAINST[353].FA_/n3 ,
         \ADD_/FAINST[353].FA_/n2 , \ADD_/FAINST[353].FA_/n1 ,
         \ADD_/FAINST[352].FA_/n3 , \ADD_/FAINST[352].FA_/n2 ,
         \ADD_/FAINST[352].FA_/n1 , \ADD_/FAINST[351].FA_/n3 ,
         \ADD_/FAINST[351].FA_/n2 , \ADD_/FAINST[351].FA_/n1 ,
         \ADD_/FAINST[350].FA_/n3 , \ADD_/FAINST[350].FA_/n2 ,
         \ADD_/FAINST[350].FA_/n1 , \ADD_/FAINST[349].FA_/n3 ,
         \ADD_/FAINST[349].FA_/n2 , \ADD_/FAINST[349].FA_/n1 ,
         \ADD_/FAINST[348].FA_/n3 , \ADD_/FAINST[348].FA_/n2 ,
         \ADD_/FAINST[348].FA_/n1 , \ADD_/FAINST[347].FA_/n3 ,
         \ADD_/FAINST[347].FA_/n2 , \ADD_/FAINST[347].FA_/n1 ,
         \ADD_/FAINST[346].FA_/n3 , \ADD_/FAINST[346].FA_/n2 ,
         \ADD_/FAINST[346].FA_/n1 , \ADD_/FAINST[345].FA_/n3 ,
         \ADD_/FAINST[345].FA_/n2 , \ADD_/FAINST[345].FA_/n1 ,
         \ADD_/FAINST[344].FA_/n3 , \ADD_/FAINST[344].FA_/n2 ,
         \ADD_/FAINST[344].FA_/n1 , \ADD_/FAINST[343].FA_/n3 ,
         \ADD_/FAINST[343].FA_/n2 , \ADD_/FAINST[343].FA_/n1 ,
         \ADD_/FAINST[342].FA_/n3 , \ADD_/FAINST[342].FA_/n2 ,
         \ADD_/FAINST[342].FA_/n1 , \ADD_/FAINST[341].FA_/n3 ,
         \ADD_/FAINST[341].FA_/n2 , \ADD_/FAINST[341].FA_/n1 ,
         \ADD_/FAINST[340].FA_/n3 , \ADD_/FAINST[340].FA_/n2 ,
         \ADD_/FAINST[340].FA_/n1 , \ADD_/FAINST[339].FA_/n3 ,
         \ADD_/FAINST[339].FA_/n2 , \ADD_/FAINST[339].FA_/n1 ,
         \ADD_/FAINST[338].FA_/n3 , \ADD_/FAINST[338].FA_/n2 ,
         \ADD_/FAINST[338].FA_/n1 , \ADD_/FAINST[337].FA_/n3 ,
         \ADD_/FAINST[337].FA_/n2 , \ADD_/FAINST[337].FA_/n1 ,
         \ADD_/FAINST[336].FA_/n3 , \ADD_/FAINST[336].FA_/n2 ,
         \ADD_/FAINST[336].FA_/n1 , \ADD_/FAINST[335].FA_/n3 ,
         \ADD_/FAINST[335].FA_/n2 , \ADD_/FAINST[335].FA_/n1 ,
         \ADD_/FAINST[334].FA_/n3 , \ADD_/FAINST[334].FA_/n2 ,
         \ADD_/FAINST[334].FA_/n1 , \ADD_/FAINST[333].FA_/n3 ,
         \ADD_/FAINST[333].FA_/n2 , \ADD_/FAINST[333].FA_/n1 ,
         \ADD_/FAINST[332].FA_/n3 , \ADD_/FAINST[332].FA_/n2 ,
         \ADD_/FAINST[332].FA_/n1 , \ADD_/FAINST[331].FA_/n3 ,
         \ADD_/FAINST[331].FA_/n2 , \ADD_/FAINST[331].FA_/n1 ,
         \ADD_/FAINST[330].FA_/n3 , \ADD_/FAINST[330].FA_/n2 ,
         \ADD_/FAINST[330].FA_/n1 , \ADD_/FAINST[329].FA_/n3 ,
         \ADD_/FAINST[329].FA_/n2 , \ADD_/FAINST[329].FA_/n1 ,
         \ADD_/FAINST[328].FA_/n3 , \ADD_/FAINST[328].FA_/n2 ,
         \ADD_/FAINST[328].FA_/n1 , \ADD_/FAINST[327].FA_/n3 ,
         \ADD_/FAINST[327].FA_/n2 , \ADD_/FAINST[327].FA_/n1 ,
         \ADD_/FAINST[326].FA_/n3 , \ADD_/FAINST[326].FA_/n2 ,
         \ADD_/FAINST[326].FA_/n1 , \ADD_/FAINST[325].FA_/n3 ,
         \ADD_/FAINST[325].FA_/n2 , \ADD_/FAINST[325].FA_/n1 ,
         \ADD_/FAINST[324].FA_/n3 , \ADD_/FAINST[324].FA_/n2 ,
         \ADD_/FAINST[324].FA_/n1 , \ADD_/FAINST[323].FA_/n3 ,
         \ADD_/FAINST[323].FA_/n2 , \ADD_/FAINST[323].FA_/n1 ,
         \ADD_/FAINST[322].FA_/n3 , \ADD_/FAINST[322].FA_/n2 ,
         \ADD_/FAINST[322].FA_/n1 , \ADD_/FAINST[321].FA_/n3 ,
         \ADD_/FAINST[321].FA_/n2 , \ADD_/FAINST[321].FA_/n1 ,
         \ADD_/FAINST[320].FA_/n3 , \ADD_/FAINST[320].FA_/n2 ,
         \ADD_/FAINST[320].FA_/n1 , \ADD_/FAINST[319].FA_/n3 ,
         \ADD_/FAINST[319].FA_/n2 , \ADD_/FAINST[319].FA_/n1 ,
         \ADD_/FAINST[318].FA_/n3 , \ADD_/FAINST[318].FA_/n2 ,
         \ADD_/FAINST[318].FA_/n1 , \ADD_/FAINST[317].FA_/n3 ,
         \ADD_/FAINST[317].FA_/n2 , \ADD_/FAINST[317].FA_/n1 ,
         \ADD_/FAINST[316].FA_/n3 , \ADD_/FAINST[316].FA_/n2 ,
         \ADD_/FAINST[316].FA_/n1 , \ADD_/FAINST[315].FA_/n3 ,
         \ADD_/FAINST[315].FA_/n2 , \ADD_/FAINST[315].FA_/n1 ,
         \ADD_/FAINST[314].FA_/n3 , \ADD_/FAINST[314].FA_/n2 ,
         \ADD_/FAINST[314].FA_/n1 , \ADD_/FAINST[313].FA_/n3 ,
         \ADD_/FAINST[313].FA_/n2 , \ADD_/FAINST[313].FA_/n1 ,
         \ADD_/FAINST[312].FA_/n3 , \ADD_/FAINST[312].FA_/n2 ,
         \ADD_/FAINST[312].FA_/n1 , \ADD_/FAINST[311].FA_/n3 ,
         \ADD_/FAINST[311].FA_/n2 , \ADD_/FAINST[311].FA_/n1 ,
         \ADD_/FAINST[310].FA_/n3 , \ADD_/FAINST[310].FA_/n2 ,
         \ADD_/FAINST[310].FA_/n1 , \ADD_/FAINST[309].FA_/n3 ,
         \ADD_/FAINST[309].FA_/n2 , \ADD_/FAINST[309].FA_/n1 ,
         \ADD_/FAINST[308].FA_/n3 , \ADD_/FAINST[308].FA_/n2 ,
         \ADD_/FAINST[308].FA_/n1 , \ADD_/FAINST[307].FA_/n3 ,
         \ADD_/FAINST[307].FA_/n2 , \ADD_/FAINST[307].FA_/n1 ,
         \ADD_/FAINST[306].FA_/n3 , \ADD_/FAINST[306].FA_/n2 ,
         \ADD_/FAINST[306].FA_/n1 , \ADD_/FAINST[305].FA_/n3 ,
         \ADD_/FAINST[305].FA_/n2 , \ADD_/FAINST[305].FA_/n1 ,
         \ADD_/FAINST[304].FA_/n3 , \ADD_/FAINST[304].FA_/n2 ,
         \ADD_/FAINST[304].FA_/n1 , \ADD_/FAINST[303].FA_/n3 ,
         \ADD_/FAINST[303].FA_/n2 , \ADD_/FAINST[303].FA_/n1 ,
         \ADD_/FAINST[302].FA_/n3 , \ADD_/FAINST[302].FA_/n2 ,
         \ADD_/FAINST[302].FA_/n1 , \ADD_/FAINST[301].FA_/n3 ,
         \ADD_/FAINST[301].FA_/n2 , \ADD_/FAINST[301].FA_/n1 ,
         \ADD_/FAINST[300].FA_/n3 , \ADD_/FAINST[300].FA_/n2 ,
         \ADD_/FAINST[300].FA_/n1 , \ADD_/FAINST[299].FA_/n3 ,
         \ADD_/FAINST[299].FA_/n2 , \ADD_/FAINST[299].FA_/n1 ,
         \ADD_/FAINST[298].FA_/n3 , \ADD_/FAINST[298].FA_/n2 ,
         \ADD_/FAINST[298].FA_/n1 , \ADD_/FAINST[297].FA_/n3 ,
         \ADD_/FAINST[297].FA_/n2 , \ADD_/FAINST[297].FA_/n1 ,
         \ADD_/FAINST[296].FA_/n3 , \ADD_/FAINST[296].FA_/n2 ,
         \ADD_/FAINST[296].FA_/n1 , \ADD_/FAINST[295].FA_/n3 ,
         \ADD_/FAINST[295].FA_/n2 , \ADD_/FAINST[295].FA_/n1 ,
         \ADD_/FAINST[294].FA_/n3 , \ADD_/FAINST[294].FA_/n2 ,
         \ADD_/FAINST[294].FA_/n1 , \ADD_/FAINST[293].FA_/n3 ,
         \ADD_/FAINST[293].FA_/n2 , \ADD_/FAINST[293].FA_/n1 ,
         \ADD_/FAINST[292].FA_/n3 , \ADD_/FAINST[292].FA_/n2 ,
         \ADD_/FAINST[292].FA_/n1 , \ADD_/FAINST[291].FA_/n3 ,
         \ADD_/FAINST[291].FA_/n2 , \ADD_/FAINST[291].FA_/n1 ,
         \ADD_/FAINST[290].FA_/n3 , \ADD_/FAINST[290].FA_/n2 ,
         \ADD_/FAINST[290].FA_/n1 , \ADD_/FAINST[289].FA_/n3 ,
         \ADD_/FAINST[289].FA_/n2 , \ADD_/FAINST[289].FA_/n1 ,
         \ADD_/FAINST[288].FA_/n3 , \ADD_/FAINST[288].FA_/n2 ,
         \ADD_/FAINST[288].FA_/n1 , \ADD_/FAINST[287].FA_/n3 ,
         \ADD_/FAINST[287].FA_/n2 , \ADD_/FAINST[287].FA_/n1 ,
         \ADD_/FAINST[286].FA_/n3 , \ADD_/FAINST[286].FA_/n2 ,
         \ADD_/FAINST[286].FA_/n1 , \ADD_/FAINST[285].FA_/n3 ,
         \ADD_/FAINST[285].FA_/n2 , \ADD_/FAINST[285].FA_/n1 ,
         \ADD_/FAINST[284].FA_/n3 , \ADD_/FAINST[284].FA_/n2 ,
         \ADD_/FAINST[284].FA_/n1 , \ADD_/FAINST[283].FA_/n3 ,
         \ADD_/FAINST[283].FA_/n2 , \ADD_/FAINST[283].FA_/n1 ,
         \ADD_/FAINST[282].FA_/n3 , \ADD_/FAINST[282].FA_/n2 ,
         \ADD_/FAINST[282].FA_/n1 , \ADD_/FAINST[281].FA_/n3 ,
         \ADD_/FAINST[281].FA_/n2 , \ADD_/FAINST[281].FA_/n1 ,
         \ADD_/FAINST[280].FA_/n3 , \ADD_/FAINST[280].FA_/n2 ,
         \ADD_/FAINST[280].FA_/n1 , \ADD_/FAINST[279].FA_/n3 ,
         \ADD_/FAINST[279].FA_/n2 , \ADD_/FAINST[279].FA_/n1 ,
         \ADD_/FAINST[278].FA_/n3 , \ADD_/FAINST[278].FA_/n2 ,
         \ADD_/FAINST[278].FA_/n1 , \ADD_/FAINST[277].FA_/n3 ,
         \ADD_/FAINST[277].FA_/n2 , \ADD_/FAINST[277].FA_/n1 ,
         \ADD_/FAINST[276].FA_/n3 , \ADD_/FAINST[276].FA_/n2 ,
         \ADD_/FAINST[276].FA_/n1 , \ADD_/FAINST[275].FA_/n3 ,
         \ADD_/FAINST[275].FA_/n2 , \ADD_/FAINST[275].FA_/n1 ,
         \ADD_/FAINST[274].FA_/n3 , \ADD_/FAINST[274].FA_/n2 ,
         \ADD_/FAINST[274].FA_/n1 , \ADD_/FAINST[273].FA_/n3 ,
         \ADD_/FAINST[273].FA_/n2 , \ADD_/FAINST[273].FA_/n1 ,
         \ADD_/FAINST[272].FA_/n3 , \ADD_/FAINST[272].FA_/n2 ,
         \ADD_/FAINST[272].FA_/n1 , \ADD_/FAINST[271].FA_/n3 ,
         \ADD_/FAINST[271].FA_/n2 , \ADD_/FAINST[271].FA_/n1 ,
         \ADD_/FAINST[270].FA_/n3 , \ADD_/FAINST[270].FA_/n2 ,
         \ADD_/FAINST[270].FA_/n1 , \ADD_/FAINST[269].FA_/n3 ,
         \ADD_/FAINST[269].FA_/n2 , \ADD_/FAINST[269].FA_/n1 ,
         \ADD_/FAINST[268].FA_/n3 , \ADD_/FAINST[268].FA_/n2 ,
         \ADD_/FAINST[268].FA_/n1 , \ADD_/FAINST[267].FA_/n3 ,
         \ADD_/FAINST[267].FA_/n2 , \ADD_/FAINST[267].FA_/n1 ,
         \ADD_/FAINST[266].FA_/n3 , \ADD_/FAINST[266].FA_/n2 ,
         \ADD_/FAINST[266].FA_/n1 , \ADD_/FAINST[265].FA_/n3 ,
         \ADD_/FAINST[265].FA_/n2 , \ADD_/FAINST[265].FA_/n1 ,
         \ADD_/FAINST[264].FA_/n3 , \ADD_/FAINST[264].FA_/n2 ,
         \ADD_/FAINST[264].FA_/n1 , \ADD_/FAINST[263].FA_/n3 ,
         \ADD_/FAINST[263].FA_/n2 , \ADD_/FAINST[263].FA_/n1 ,
         \ADD_/FAINST[262].FA_/n3 , \ADD_/FAINST[262].FA_/n2 ,
         \ADD_/FAINST[262].FA_/n1 , \ADD_/FAINST[261].FA_/n3 ,
         \ADD_/FAINST[261].FA_/n2 , \ADD_/FAINST[261].FA_/n1 ,
         \ADD_/FAINST[260].FA_/n3 , \ADD_/FAINST[260].FA_/n2 ,
         \ADD_/FAINST[260].FA_/n1 , \ADD_/FAINST[259].FA_/n3 ,
         \ADD_/FAINST[259].FA_/n2 , \ADD_/FAINST[259].FA_/n1 ,
         \ADD_/FAINST[258].FA_/n3 , \ADD_/FAINST[258].FA_/n2 ,
         \ADD_/FAINST[258].FA_/n1 , \ADD_/FAINST[257].FA_/n3 ,
         \ADD_/FAINST[257].FA_/n2 , \ADD_/FAINST[257].FA_/n1 ,
         \ADD_/FAINST[256].FA_/n3 , \ADD_/FAINST[256].FA_/n2 ,
         \ADD_/FAINST[256].FA_/n1 , \ADD_/FAINST[255].FA_/n3 ,
         \ADD_/FAINST[255].FA_/n2 , \ADD_/FAINST[255].FA_/n1 ,
         \ADD_/FAINST[254].FA_/n3 , \ADD_/FAINST[254].FA_/n2 ,
         \ADD_/FAINST[254].FA_/n1 , \ADD_/FAINST[253].FA_/n3 ,
         \ADD_/FAINST[253].FA_/n2 , \ADD_/FAINST[253].FA_/n1 ,
         \ADD_/FAINST[252].FA_/n3 , \ADD_/FAINST[252].FA_/n2 ,
         \ADD_/FAINST[252].FA_/n1 , \ADD_/FAINST[251].FA_/n3 ,
         \ADD_/FAINST[251].FA_/n2 , \ADD_/FAINST[251].FA_/n1 ,
         \ADD_/FAINST[250].FA_/n3 , \ADD_/FAINST[250].FA_/n2 ,
         \ADD_/FAINST[250].FA_/n1 , \ADD_/FAINST[249].FA_/n3 ,
         \ADD_/FAINST[249].FA_/n2 , \ADD_/FAINST[249].FA_/n1 ,
         \ADD_/FAINST[248].FA_/n3 , \ADD_/FAINST[248].FA_/n2 ,
         \ADD_/FAINST[248].FA_/n1 , \ADD_/FAINST[247].FA_/n3 ,
         \ADD_/FAINST[247].FA_/n2 , \ADD_/FAINST[247].FA_/n1 ,
         \ADD_/FAINST[246].FA_/n3 , \ADD_/FAINST[246].FA_/n2 ,
         \ADD_/FAINST[246].FA_/n1 , \ADD_/FAINST[245].FA_/n3 ,
         \ADD_/FAINST[245].FA_/n2 , \ADD_/FAINST[245].FA_/n1 ,
         \ADD_/FAINST[244].FA_/n3 , \ADD_/FAINST[244].FA_/n2 ,
         \ADD_/FAINST[244].FA_/n1 , \ADD_/FAINST[243].FA_/n3 ,
         \ADD_/FAINST[243].FA_/n2 , \ADD_/FAINST[243].FA_/n1 ,
         \ADD_/FAINST[242].FA_/n3 , \ADD_/FAINST[242].FA_/n2 ,
         \ADD_/FAINST[242].FA_/n1 , \ADD_/FAINST[241].FA_/n3 ,
         \ADD_/FAINST[241].FA_/n2 , \ADD_/FAINST[241].FA_/n1 ,
         \ADD_/FAINST[240].FA_/n3 , \ADD_/FAINST[240].FA_/n2 ,
         \ADD_/FAINST[240].FA_/n1 , \ADD_/FAINST[239].FA_/n3 ,
         \ADD_/FAINST[239].FA_/n2 , \ADD_/FAINST[239].FA_/n1 ,
         \ADD_/FAINST[238].FA_/n3 , \ADD_/FAINST[238].FA_/n2 ,
         \ADD_/FAINST[238].FA_/n1 , \ADD_/FAINST[237].FA_/n3 ,
         \ADD_/FAINST[237].FA_/n2 , \ADD_/FAINST[237].FA_/n1 ,
         \ADD_/FAINST[236].FA_/n3 , \ADD_/FAINST[236].FA_/n2 ,
         \ADD_/FAINST[236].FA_/n1 , \ADD_/FAINST[235].FA_/n3 ,
         \ADD_/FAINST[235].FA_/n2 , \ADD_/FAINST[235].FA_/n1 ,
         \ADD_/FAINST[234].FA_/n3 , \ADD_/FAINST[234].FA_/n2 ,
         \ADD_/FAINST[234].FA_/n1 , \ADD_/FAINST[233].FA_/n3 ,
         \ADD_/FAINST[233].FA_/n2 , \ADD_/FAINST[233].FA_/n1 ,
         \ADD_/FAINST[232].FA_/n3 , \ADD_/FAINST[232].FA_/n2 ,
         \ADD_/FAINST[232].FA_/n1 , \ADD_/FAINST[231].FA_/n3 ,
         \ADD_/FAINST[231].FA_/n2 , \ADD_/FAINST[231].FA_/n1 ,
         \ADD_/FAINST[230].FA_/n3 , \ADD_/FAINST[230].FA_/n2 ,
         \ADD_/FAINST[230].FA_/n1 , \ADD_/FAINST[229].FA_/n3 ,
         \ADD_/FAINST[229].FA_/n2 , \ADD_/FAINST[229].FA_/n1 ,
         \ADD_/FAINST[228].FA_/n3 , \ADD_/FAINST[228].FA_/n2 ,
         \ADD_/FAINST[228].FA_/n1 , \ADD_/FAINST[227].FA_/n3 ,
         \ADD_/FAINST[227].FA_/n2 , \ADD_/FAINST[227].FA_/n1 ,
         \ADD_/FAINST[226].FA_/n3 , \ADD_/FAINST[226].FA_/n2 ,
         \ADD_/FAINST[226].FA_/n1 , \ADD_/FAINST[225].FA_/n3 ,
         \ADD_/FAINST[225].FA_/n2 , \ADD_/FAINST[225].FA_/n1 ,
         \ADD_/FAINST[224].FA_/n3 , \ADD_/FAINST[224].FA_/n2 ,
         \ADD_/FAINST[224].FA_/n1 , \ADD_/FAINST[223].FA_/n3 ,
         \ADD_/FAINST[223].FA_/n2 , \ADD_/FAINST[223].FA_/n1 ,
         \ADD_/FAINST[222].FA_/n3 , \ADD_/FAINST[222].FA_/n2 ,
         \ADD_/FAINST[222].FA_/n1 , \ADD_/FAINST[221].FA_/n3 ,
         \ADD_/FAINST[221].FA_/n2 , \ADD_/FAINST[221].FA_/n1 ,
         \ADD_/FAINST[220].FA_/n3 , \ADD_/FAINST[220].FA_/n2 ,
         \ADD_/FAINST[220].FA_/n1 , \ADD_/FAINST[219].FA_/n3 ,
         \ADD_/FAINST[219].FA_/n2 , \ADD_/FAINST[219].FA_/n1 ,
         \ADD_/FAINST[218].FA_/n3 , \ADD_/FAINST[218].FA_/n2 ,
         \ADD_/FAINST[218].FA_/n1 , \ADD_/FAINST[217].FA_/n3 ,
         \ADD_/FAINST[217].FA_/n2 , \ADD_/FAINST[217].FA_/n1 ,
         \ADD_/FAINST[216].FA_/n3 , \ADD_/FAINST[216].FA_/n2 ,
         \ADD_/FAINST[216].FA_/n1 , \ADD_/FAINST[215].FA_/n3 ,
         \ADD_/FAINST[215].FA_/n2 , \ADD_/FAINST[215].FA_/n1 ,
         \ADD_/FAINST[214].FA_/n3 , \ADD_/FAINST[214].FA_/n2 ,
         \ADD_/FAINST[214].FA_/n1 , \ADD_/FAINST[213].FA_/n3 ,
         \ADD_/FAINST[213].FA_/n2 , \ADD_/FAINST[213].FA_/n1 ,
         \ADD_/FAINST[212].FA_/n3 , \ADD_/FAINST[212].FA_/n2 ,
         \ADD_/FAINST[212].FA_/n1 , \ADD_/FAINST[211].FA_/n3 ,
         \ADD_/FAINST[211].FA_/n2 , \ADD_/FAINST[211].FA_/n1 ,
         \ADD_/FAINST[210].FA_/n3 , \ADD_/FAINST[210].FA_/n2 ,
         \ADD_/FAINST[210].FA_/n1 , \ADD_/FAINST[209].FA_/n3 ,
         \ADD_/FAINST[209].FA_/n2 , \ADD_/FAINST[209].FA_/n1 ,
         \ADD_/FAINST[208].FA_/n3 , \ADD_/FAINST[208].FA_/n2 ,
         \ADD_/FAINST[208].FA_/n1 , \ADD_/FAINST[207].FA_/n3 ,
         \ADD_/FAINST[207].FA_/n2 , \ADD_/FAINST[207].FA_/n1 ,
         \ADD_/FAINST[206].FA_/n3 , \ADD_/FAINST[206].FA_/n2 ,
         \ADD_/FAINST[206].FA_/n1 , \ADD_/FAINST[205].FA_/n3 ,
         \ADD_/FAINST[205].FA_/n2 , \ADD_/FAINST[205].FA_/n1 ,
         \ADD_/FAINST[204].FA_/n3 , \ADD_/FAINST[204].FA_/n2 ,
         \ADD_/FAINST[204].FA_/n1 , \ADD_/FAINST[203].FA_/n3 ,
         \ADD_/FAINST[203].FA_/n2 , \ADD_/FAINST[203].FA_/n1 ,
         \ADD_/FAINST[202].FA_/n3 , \ADD_/FAINST[202].FA_/n2 ,
         \ADD_/FAINST[202].FA_/n1 , \ADD_/FAINST[201].FA_/n3 ,
         \ADD_/FAINST[201].FA_/n2 , \ADD_/FAINST[201].FA_/n1 ,
         \ADD_/FAINST[200].FA_/n3 , \ADD_/FAINST[200].FA_/n2 ,
         \ADD_/FAINST[200].FA_/n1 , \ADD_/FAINST[199].FA_/n3 ,
         \ADD_/FAINST[199].FA_/n2 , \ADD_/FAINST[199].FA_/n1 ,
         \ADD_/FAINST[198].FA_/n3 , \ADD_/FAINST[198].FA_/n2 ,
         \ADD_/FAINST[198].FA_/n1 , \ADD_/FAINST[197].FA_/n3 ,
         \ADD_/FAINST[197].FA_/n2 , \ADD_/FAINST[197].FA_/n1 ,
         \ADD_/FAINST[196].FA_/n3 , \ADD_/FAINST[196].FA_/n2 ,
         \ADD_/FAINST[196].FA_/n1 , \ADD_/FAINST[195].FA_/n3 ,
         \ADD_/FAINST[195].FA_/n2 , \ADD_/FAINST[195].FA_/n1 ,
         \ADD_/FAINST[194].FA_/n3 , \ADD_/FAINST[194].FA_/n2 ,
         \ADD_/FAINST[194].FA_/n1 , \ADD_/FAINST[193].FA_/n3 ,
         \ADD_/FAINST[193].FA_/n2 , \ADD_/FAINST[193].FA_/n1 ,
         \ADD_/FAINST[192].FA_/n3 , \ADD_/FAINST[192].FA_/n2 ,
         \ADD_/FAINST[192].FA_/n1 , \ADD_/FAINST[191].FA_/n3 ,
         \ADD_/FAINST[191].FA_/n2 , \ADD_/FAINST[191].FA_/n1 ,
         \ADD_/FAINST[190].FA_/n3 , \ADD_/FAINST[190].FA_/n2 ,
         \ADD_/FAINST[190].FA_/n1 , \ADD_/FAINST[189].FA_/n3 ,
         \ADD_/FAINST[189].FA_/n2 , \ADD_/FAINST[189].FA_/n1 ,
         \ADD_/FAINST[188].FA_/n3 , \ADD_/FAINST[188].FA_/n2 ,
         \ADD_/FAINST[188].FA_/n1 , \ADD_/FAINST[187].FA_/n3 ,
         \ADD_/FAINST[187].FA_/n2 , \ADD_/FAINST[187].FA_/n1 ,
         \ADD_/FAINST[186].FA_/n3 , \ADD_/FAINST[186].FA_/n2 ,
         \ADD_/FAINST[186].FA_/n1 , \ADD_/FAINST[185].FA_/n3 ,
         \ADD_/FAINST[185].FA_/n2 , \ADD_/FAINST[185].FA_/n1 ,
         \ADD_/FAINST[184].FA_/n3 , \ADD_/FAINST[184].FA_/n2 ,
         \ADD_/FAINST[184].FA_/n1 , \ADD_/FAINST[183].FA_/n3 ,
         \ADD_/FAINST[183].FA_/n2 , \ADD_/FAINST[183].FA_/n1 ,
         \ADD_/FAINST[182].FA_/n3 , \ADD_/FAINST[182].FA_/n2 ,
         \ADD_/FAINST[182].FA_/n1 , \ADD_/FAINST[181].FA_/n3 ,
         \ADD_/FAINST[181].FA_/n2 , \ADD_/FAINST[181].FA_/n1 ,
         \ADD_/FAINST[180].FA_/n3 , \ADD_/FAINST[180].FA_/n2 ,
         \ADD_/FAINST[180].FA_/n1 , \ADD_/FAINST[179].FA_/n3 ,
         \ADD_/FAINST[179].FA_/n2 , \ADD_/FAINST[179].FA_/n1 ,
         \ADD_/FAINST[178].FA_/n3 , \ADD_/FAINST[178].FA_/n2 ,
         \ADD_/FAINST[178].FA_/n1 , \ADD_/FAINST[177].FA_/n3 ,
         \ADD_/FAINST[177].FA_/n2 , \ADD_/FAINST[177].FA_/n1 ,
         \ADD_/FAINST[176].FA_/n3 , \ADD_/FAINST[176].FA_/n2 ,
         \ADD_/FAINST[176].FA_/n1 , \ADD_/FAINST[175].FA_/n3 ,
         \ADD_/FAINST[175].FA_/n2 , \ADD_/FAINST[175].FA_/n1 ,
         \ADD_/FAINST[174].FA_/n3 , \ADD_/FAINST[174].FA_/n2 ,
         \ADD_/FAINST[174].FA_/n1 , \ADD_/FAINST[173].FA_/n3 ,
         \ADD_/FAINST[173].FA_/n2 , \ADD_/FAINST[173].FA_/n1 ,
         \ADD_/FAINST[172].FA_/n3 , \ADD_/FAINST[172].FA_/n2 ,
         \ADD_/FAINST[172].FA_/n1 , \ADD_/FAINST[171].FA_/n3 ,
         \ADD_/FAINST[171].FA_/n2 , \ADD_/FAINST[171].FA_/n1 ,
         \ADD_/FAINST[170].FA_/n3 , \ADD_/FAINST[170].FA_/n2 ,
         \ADD_/FAINST[170].FA_/n1 , \ADD_/FAINST[169].FA_/n3 ,
         \ADD_/FAINST[169].FA_/n2 , \ADD_/FAINST[169].FA_/n1 ,
         \ADD_/FAINST[168].FA_/n3 , \ADD_/FAINST[168].FA_/n2 ,
         \ADD_/FAINST[168].FA_/n1 , \ADD_/FAINST[167].FA_/n3 ,
         \ADD_/FAINST[167].FA_/n2 , \ADD_/FAINST[167].FA_/n1 ,
         \ADD_/FAINST[166].FA_/n3 , \ADD_/FAINST[166].FA_/n2 ,
         \ADD_/FAINST[166].FA_/n1 , \ADD_/FAINST[165].FA_/n3 ,
         \ADD_/FAINST[165].FA_/n2 , \ADD_/FAINST[165].FA_/n1 ,
         \ADD_/FAINST[164].FA_/n3 , \ADD_/FAINST[164].FA_/n2 ,
         \ADD_/FAINST[164].FA_/n1 , \ADD_/FAINST[163].FA_/n3 ,
         \ADD_/FAINST[163].FA_/n2 , \ADD_/FAINST[163].FA_/n1 ,
         \ADD_/FAINST[162].FA_/n3 , \ADD_/FAINST[162].FA_/n2 ,
         \ADD_/FAINST[162].FA_/n1 , \ADD_/FAINST[161].FA_/n3 ,
         \ADD_/FAINST[161].FA_/n2 , \ADD_/FAINST[161].FA_/n1 ,
         \ADD_/FAINST[160].FA_/n3 , \ADD_/FAINST[160].FA_/n2 ,
         \ADD_/FAINST[160].FA_/n1 , \ADD_/FAINST[159].FA_/n3 ,
         \ADD_/FAINST[159].FA_/n2 , \ADD_/FAINST[159].FA_/n1 ,
         \ADD_/FAINST[158].FA_/n3 , \ADD_/FAINST[158].FA_/n2 ,
         \ADD_/FAINST[158].FA_/n1 , \ADD_/FAINST[157].FA_/n3 ,
         \ADD_/FAINST[157].FA_/n2 , \ADD_/FAINST[157].FA_/n1 ,
         \ADD_/FAINST[156].FA_/n3 , \ADD_/FAINST[156].FA_/n2 ,
         \ADD_/FAINST[156].FA_/n1 , \ADD_/FAINST[155].FA_/n3 ,
         \ADD_/FAINST[155].FA_/n2 , \ADD_/FAINST[155].FA_/n1 ,
         \ADD_/FAINST[154].FA_/n3 , \ADD_/FAINST[154].FA_/n2 ,
         \ADD_/FAINST[154].FA_/n1 , \ADD_/FAINST[153].FA_/n3 ,
         \ADD_/FAINST[153].FA_/n2 , \ADD_/FAINST[153].FA_/n1 ,
         \ADD_/FAINST[152].FA_/n3 , \ADD_/FAINST[152].FA_/n2 ,
         \ADD_/FAINST[152].FA_/n1 , \ADD_/FAINST[151].FA_/n3 ,
         \ADD_/FAINST[151].FA_/n2 , \ADD_/FAINST[151].FA_/n1 ,
         \ADD_/FAINST[150].FA_/n3 , \ADD_/FAINST[150].FA_/n2 ,
         \ADD_/FAINST[150].FA_/n1 , \ADD_/FAINST[149].FA_/n3 ,
         \ADD_/FAINST[149].FA_/n2 , \ADD_/FAINST[149].FA_/n1 ,
         \ADD_/FAINST[148].FA_/n3 , \ADD_/FAINST[148].FA_/n2 ,
         \ADD_/FAINST[148].FA_/n1 , \ADD_/FAINST[147].FA_/n3 ,
         \ADD_/FAINST[147].FA_/n2 , \ADD_/FAINST[147].FA_/n1 ,
         \ADD_/FAINST[146].FA_/n3 , \ADD_/FAINST[146].FA_/n2 ,
         \ADD_/FAINST[146].FA_/n1 , \ADD_/FAINST[145].FA_/n3 ,
         \ADD_/FAINST[145].FA_/n2 , \ADD_/FAINST[145].FA_/n1 ,
         \ADD_/FAINST[144].FA_/n3 , \ADD_/FAINST[144].FA_/n2 ,
         \ADD_/FAINST[144].FA_/n1 , \ADD_/FAINST[143].FA_/n3 ,
         \ADD_/FAINST[143].FA_/n2 , \ADD_/FAINST[143].FA_/n1 ,
         \ADD_/FAINST[142].FA_/n3 , \ADD_/FAINST[142].FA_/n2 ,
         \ADD_/FAINST[142].FA_/n1 , \ADD_/FAINST[141].FA_/n3 ,
         \ADD_/FAINST[141].FA_/n2 , \ADD_/FAINST[141].FA_/n1 ,
         \ADD_/FAINST[140].FA_/n3 , \ADD_/FAINST[140].FA_/n2 ,
         \ADD_/FAINST[140].FA_/n1 , \ADD_/FAINST[139].FA_/n3 ,
         \ADD_/FAINST[139].FA_/n2 , \ADD_/FAINST[139].FA_/n1 ,
         \ADD_/FAINST[138].FA_/n3 , \ADD_/FAINST[138].FA_/n2 ,
         \ADD_/FAINST[138].FA_/n1 , \ADD_/FAINST[137].FA_/n3 ,
         \ADD_/FAINST[137].FA_/n2 , \ADD_/FAINST[137].FA_/n1 ,
         \ADD_/FAINST[136].FA_/n3 , \ADD_/FAINST[136].FA_/n2 ,
         \ADD_/FAINST[136].FA_/n1 , \ADD_/FAINST[135].FA_/n3 ,
         \ADD_/FAINST[135].FA_/n2 , \ADD_/FAINST[135].FA_/n1 ,
         \ADD_/FAINST[134].FA_/n3 , \ADD_/FAINST[134].FA_/n2 ,
         \ADD_/FAINST[134].FA_/n1 , \ADD_/FAINST[133].FA_/n3 ,
         \ADD_/FAINST[133].FA_/n2 , \ADD_/FAINST[133].FA_/n1 ,
         \ADD_/FAINST[132].FA_/n3 , \ADD_/FAINST[132].FA_/n2 ,
         \ADD_/FAINST[132].FA_/n1 , \ADD_/FAINST[131].FA_/n3 ,
         \ADD_/FAINST[131].FA_/n2 , \ADD_/FAINST[131].FA_/n1 ,
         \ADD_/FAINST[130].FA_/n3 , \ADD_/FAINST[130].FA_/n2 ,
         \ADD_/FAINST[130].FA_/n1 , \ADD_/FAINST[129].FA_/n3 ,
         \ADD_/FAINST[129].FA_/n2 , \ADD_/FAINST[129].FA_/n1 ,
         \ADD_/FAINST[128].FA_/n3 , \ADD_/FAINST[128].FA_/n2 ,
         \ADD_/FAINST[128].FA_/n1 , \ADD_/FAINST[127].FA_/n3 ,
         \ADD_/FAINST[127].FA_/n2 , \ADD_/FAINST[127].FA_/n1 ,
         \ADD_/FAINST[126].FA_/n3 , \ADD_/FAINST[126].FA_/n2 ,
         \ADD_/FAINST[126].FA_/n1 , \ADD_/FAINST[125].FA_/n3 ,
         \ADD_/FAINST[125].FA_/n2 , \ADD_/FAINST[125].FA_/n1 ,
         \ADD_/FAINST[124].FA_/n3 , \ADD_/FAINST[124].FA_/n2 ,
         \ADD_/FAINST[124].FA_/n1 , \ADD_/FAINST[123].FA_/n3 ,
         \ADD_/FAINST[123].FA_/n2 , \ADD_/FAINST[123].FA_/n1 ,
         \ADD_/FAINST[122].FA_/n3 , \ADD_/FAINST[122].FA_/n2 ,
         \ADD_/FAINST[122].FA_/n1 , \ADD_/FAINST[121].FA_/n3 ,
         \ADD_/FAINST[121].FA_/n2 , \ADD_/FAINST[121].FA_/n1 ,
         \ADD_/FAINST[120].FA_/n3 , \ADD_/FAINST[120].FA_/n2 ,
         \ADD_/FAINST[120].FA_/n1 , \ADD_/FAINST[119].FA_/n3 ,
         \ADD_/FAINST[119].FA_/n2 , \ADD_/FAINST[119].FA_/n1 ,
         \ADD_/FAINST[118].FA_/n3 , \ADD_/FAINST[118].FA_/n2 ,
         \ADD_/FAINST[118].FA_/n1 , \ADD_/FAINST[117].FA_/n3 ,
         \ADD_/FAINST[117].FA_/n2 , \ADD_/FAINST[117].FA_/n1 ,
         \ADD_/FAINST[116].FA_/n3 , \ADD_/FAINST[116].FA_/n2 ,
         \ADD_/FAINST[116].FA_/n1 , \ADD_/FAINST[115].FA_/n3 ,
         \ADD_/FAINST[115].FA_/n2 , \ADD_/FAINST[115].FA_/n1 ,
         \ADD_/FAINST[114].FA_/n3 , \ADD_/FAINST[114].FA_/n2 ,
         \ADD_/FAINST[114].FA_/n1 , \ADD_/FAINST[113].FA_/n3 ,
         \ADD_/FAINST[113].FA_/n2 , \ADD_/FAINST[113].FA_/n1 ,
         \ADD_/FAINST[112].FA_/n3 , \ADD_/FAINST[112].FA_/n2 ,
         \ADD_/FAINST[112].FA_/n1 , \ADD_/FAINST[111].FA_/n3 ,
         \ADD_/FAINST[111].FA_/n2 , \ADD_/FAINST[111].FA_/n1 ,
         \ADD_/FAINST[110].FA_/n3 , \ADD_/FAINST[110].FA_/n2 ,
         \ADD_/FAINST[110].FA_/n1 , \ADD_/FAINST[109].FA_/n3 ,
         \ADD_/FAINST[109].FA_/n2 , \ADD_/FAINST[109].FA_/n1 ,
         \ADD_/FAINST[108].FA_/n3 , \ADD_/FAINST[108].FA_/n2 ,
         \ADD_/FAINST[108].FA_/n1 , \ADD_/FAINST[107].FA_/n3 ,
         \ADD_/FAINST[107].FA_/n2 , \ADD_/FAINST[107].FA_/n1 ,
         \ADD_/FAINST[106].FA_/n3 , \ADD_/FAINST[106].FA_/n2 ,
         \ADD_/FAINST[106].FA_/n1 , \ADD_/FAINST[105].FA_/n3 ,
         \ADD_/FAINST[105].FA_/n2 , \ADD_/FAINST[105].FA_/n1 ,
         \ADD_/FAINST[104].FA_/n3 , \ADD_/FAINST[104].FA_/n2 ,
         \ADD_/FAINST[104].FA_/n1 , \ADD_/FAINST[103].FA_/n3 ,
         \ADD_/FAINST[103].FA_/n2 , \ADD_/FAINST[103].FA_/n1 ,
         \ADD_/FAINST[102].FA_/n3 , \ADD_/FAINST[102].FA_/n2 ,
         \ADD_/FAINST[102].FA_/n1 , \ADD_/FAINST[101].FA_/n3 ,
         \ADD_/FAINST[101].FA_/n2 , \ADD_/FAINST[101].FA_/n1 ,
         \ADD_/FAINST[100].FA_/n3 , \ADD_/FAINST[100].FA_/n2 ,
         \ADD_/FAINST[100].FA_/n1 , \ADD_/FAINST[99].FA_/n3 ,
         \ADD_/FAINST[99].FA_/n2 , \ADD_/FAINST[99].FA_/n1 ,
         \ADD_/FAINST[98].FA_/n3 , \ADD_/FAINST[98].FA_/n2 ,
         \ADD_/FAINST[98].FA_/n1 , \ADD_/FAINST[97].FA_/n3 ,
         \ADD_/FAINST[97].FA_/n2 , \ADD_/FAINST[97].FA_/n1 ,
         \ADD_/FAINST[96].FA_/n3 , \ADD_/FAINST[96].FA_/n2 ,
         \ADD_/FAINST[96].FA_/n1 , \ADD_/FAINST[95].FA_/n3 ,
         \ADD_/FAINST[95].FA_/n2 , \ADD_/FAINST[95].FA_/n1 ,
         \ADD_/FAINST[94].FA_/n3 , \ADD_/FAINST[94].FA_/n2 ,
         \ADD_/FAINST[94].FA_/n1 , \ADD_/FAINST[93].FA_/n3 ,
         \ADD_/FAINST[93].FA_/n2 , \ADD_/FAINST[93].FA_/n1 ,
         \ADD_/FAINST[92].FA_/n3 , \ADD_/FAINST[92].FA_/n2 ,
         \ADD_/FAINST[92].FA_/n1 , \ADD_/FAINST[91].FA_/n3 ,
         \ADD_/FAINST[91].FA_/n2 , \ADD_/FAINST[91].FA_/n1 ,
         \ADD_/FAINST[90].FA_/n3 , \ADD_/FAINST[90].FA_/n2 ,
         \ADD_/FAINST[90].FA_/n1 , \ADD_/FAINST[89].FA_/n3 ,
         \ADD_/FAINST[89].FA_/n2 , \ADD_/FAINST[89].FA_/n1 ,
         \ADD_/FAINST[88].FA_/n3 , \ADD_/FAINST[88].FA_/n2 ,
         \ADD_/FAINST[88].FA_/n1 , \ADD_/FAINST[87].FA_/n3 ,
         \ADD_/FAINST[87].FA_/n2 , \ADD_/FAINST[87].FA_/n1 ,
         \ADD_/FAINST[86].FA_/n3 , \ADD_/FAINST[86].FA_/n2 ,
         \ADD_/FAINST[86].FA_/n1 , \ADD_/FAINST[85].FA_/n3 ,
         \ADD_/FAINST[85].FA_/n2 , \ADD_/FAINST[85].FA_/n1 ,
         \ADD_/FAINST[84].FA_/n3 , \ADD_/FAINST[84].FA_/n2 ,
         \ADD_/FAINST[84].FA_/n1 , \ADD_/FAINST[83].FA_/n3 ,
         \ADD_/FAINST[83].FA_/n2 , \ADD_/FAINST[83].FA_/n1 ,
         \ADD_/FAINST[82].FA_/n3 , \ADD_/FAINST[82].FA_/n2 ,
         \ADD_/FAINST[82].FA_/n1 , \ADD_/FAINST[81].FA_/n3 ,
         \ADD_/FAINST[81].FA_/n2 , \ADD_/FAINST[81].FA_/n1 ,
         \ADD_/FAINST[80].FA_/n3 , \ADD_/FAINST[80].FA_/n2 ,
         \ADD_/FAINST[80].FA_/n1 , \ADD_/FAINST[79].FA_/n3 ,
         \ADD_/FAINST[79].FA_/n2 , \ADD_/FAINST[79].FA_/n1 ,
         \ADD_/FAINST[78].FA_/n3 , \ADD_/FAINST[78].FA_/n2 ,
         \ADD_/FAINST[78].FA_/n1 , \ADD_/FAINST[77].FA_/n3 ,
         \ADD_/FAINST[77].FA_/n2 , \ADD_/FAINST[77].FA_/n1 ,
         \ADD_/FAINST[76].FA_/n3 , \ADD_/FAINST[76].FA_/n2 ,
         \ADD_/FAINST[76].FA_/n1 , \ADD_/FAINST[75].FA_/n3 ,
         \ADD_/FAINST[75].FA_/n2 , \ADD_/FAINST[75].FA_/n1 ,
         \ADD_/FAINST[74].FA_/n3 , \ADD_/FAINST[74].FA_/n2 ,
         \ADD_/FAINST[74].FA_/n1 , \ADD_/FAINST[73].FA_/n3 ,
         \ADD_/FAINST[73].FA_/n2 , \ADD_/FAINST[73].FA_/n1 ,
         \ADD_/FAINST[72].FA_/n3 , \ADD_/FAINST[72].FA_/n2 ,
         \ADD_/FAINST[72].FA_/n1 , \ADD_/FAINST[71].FA_/n3 ,
         \ADD_/FAINST[71].FA_/n2 , \ADD_/FAINST[71].FA_/n1 ,
         \ADD_/FAINST[70].FA_/n3 , \ADD_/FAINST[70].FA_/n2 ,
         \ADD_/FAINST[70].FA_/n1 , \ADD_/FAINST[69].FA_/n3 ,
         \ADD_/FAINST[69].FA_/n2 , \ADD_/FAINST[69].FA_/n1 ,
         \ADD_/FAINST[68].FA_/n3 , \ADD_/FAINST[68].FA_/n2 ,
         \ADD_/FAINST[68].FA_/n1 , \ADD_/FAINST[67].FA_/n3 ,
         \ADD_/FAINST[67].FA_/n2 , \ADD_/FAINST[67].FA_/n1 ,
         \ADD_/FAINST[66].FA_/n3 , \ADD_/FAINST[66].FA_/n2 ,
         \ADD_/FAINST[66].FA_/n1 , \ADD_/FAINST[65].FA_/n3 ,
         \ADD_/FAINST[65].FA_/n2 , \ADD_/FAINST[65].FA_/n1 ,
         \ADD_/FAINST[64].FA_/n3 , \ADD_/FAINST[64].FA_/n2 ,
         \ADD_/FAINST[64].FA_/n1 , \ADD_/FAINST[63].FA_/n3 ,
         \ADD_/FAINST[63].FA_/n2 , \ADD_/FAINST[63].FA_/n1 ,
         \ADD_/FAINST[62].FA_/n3 , \ADD_/FAINST[62].FA_/n2 ,
         \ADD_/FAINST[62].FA_/n1 , \ADD_/FAINST[61].FA_/n3 ,
         \ADD_/FAINST[61].FA_/n2 , \ADD_/FAINST[61].FA_/n1 ,
         \ADD_/FAINST[60].FA_/n3 , \ADD_/FAINST[60].FA_/n2 ,
         \ADD_/FAINST[60].FA_/n1 , \ADD_/FAINST[59].FA_/n3 ,
         \ADD_/FAINST[59].FA_/n2 , \ADD_/FAINST[59].FA_/n1 ,
         \ADD_/FAINST[58].FA_/n3 , \ADD_/FAINST[58].FA_/n2 ,
         \ADD_/FAINST[58].FA_/n1 , \ADD_/FAINST[57].FA_/n3 ,
         \ADD_/FAINST[57].FA_/n2 , \ADD_/FAINST[57].FA_/n1 ,
         \ADD_/FAINST[56].FA_/n3 , \ADD_/FAINST[56].FA_/n2 ,
         \ADD_/FAINST[56].FA_/n1 , \ADD_/FAINST[55].FA_/n3 ,
         \ADD_/FAINST[55].FA_/n2 , \ADD_/FAINST[55].FA_/n1 ,
         \ADD_/FAINST[54].FA_/n3 , \ADD_/FAINST[54].FA_/n2 ,
         \ADD_/FAINST[54].FA_/n1 , \ADD_/FAINST[53].FA_/n3 ,
         \ADD_/FAINST[53].FA_/n2 , \ADD_/FAINST[53].FA_/n1 ,
         \ADD_/FAINST[52].FA_/n3 , \ADD_/FAINST[52].FA_/n2 ,
         \ADD_/FAINST[52].FA_/n1 , \ADD_/FAINST[51].FA_/n3 ,
         \ADD_/FAINST[51].FA_/n2 , \ADD_/FAINST[51].FA_/n1 ,
         \ADD_/FAINST[50].FA_/n3 , \ADD_/FAINST[50].FA_/n2 ,
         \ADD_/FAINST[50].FA_/n1 , \ADD_/FAINST[49].FA_/n3 ,
         \ADD_/FAINST[49].FA_/n2 , \ADD_/FAINST[49].FA_/n1 ,
         \ADD_/FAINST[48].FA_/n3 , \ADD_/FAINST[48].FA_/n2 ,
         \ADD_/FAINST[48].FA_/n1 , \ADD_/FAINST[47].FA_/n3 ,
         \ADD_/FAINST[47].FA_/n2 , \ADD_/FAINST[47].FA_/n1 ,
         \ADD_/FAINST[46].FA_/n3 , \ADD_/FAINST[46].FA_/n2 ,
         \ADD_/FAINST[46].FA_/n1 , \ADD_/FAINST[45].FA_/n3 ,
         \ADD_/FAINST[45].FA_/n2 , \ADD_/FAINST[45].FA_/n1 ,
         \ADD_/FAINST[44].FA_/n3 , \ADD_/FAINST[44].FA_/n2 ,
         \ADD_/FAINST[44].FA_/n1 , \ADD_/FAINST[43].FA_/n3 ,
         \ADD_/FAINST[43].FA_/n2 , \ADD_/FAINST[43].FA_/n1 ,
         \ADD_/FAINST[42].FA_/n3 , \ADD_/FAINST[42].FA_/n2 ,
         \ADD_/FAINST[42].FA_/n1 , \ADD_/FAINST[41].FA_/n3 ,
         \ADD_/FAINST[41].FA_/n2 , \ADD_/FAINST[41].FA_/n1 ,
         \ADD_/FAINST[40].FA_/n3 , \ADD_/FAINST[40].FA_/n2 ,
         \ADD_/FAINST[40].FA_/n1 , \ADD_/FAINST[39].FA_/n3 ,
         \ADD_/FAINST[39].FA_/n2 , \ADD_/FAINST[39].FA_/n1 ,
         \ADD_/FAINST[38].FA_/n3 , \ADD_/FAINST[38].FA_/n2 ,
         \ADD_/FAINST[38].FA_/n1 , \ADD_/FAINST[37].FA_/n3 ,
         \ADD_/FAINST[37].FA_/n2 , \ADD_/FAINST[37].FA_/n1 ,
         \ADD_/FAINST[36].FA_/n3 , \ADD_/FAINST[36].FA_/n2 ,
         \ADD_/FAINST[36].FA_/n1 , \ADD_/FAINST[35].FA_/n3 ,
         \ADD_/FAINST[35].FA_/n2 , \ADD_/FAINST[35].FA_/n1 ,
         \ADD_/FAINST[34].FA_/n3 , \ADD_/FAINST[34].FA_/n2 ,
         \ADD_/FAINST[34].FA_/n1 , \ADD_/FAINST[33].FA_/n3 ,
         \ADD_/FAINST[33].FA_/n2 , \ADD_/FAINST[33].FA_/n1 ,
         \ADD_/FAINST[32].FA_/n3 , \ADD_/FAINST[32].FA_/n2 ,
         \ADD_/FAINST[32].FA_/n1 , \ADD_/FAINST[31].FA_/n3 ,
         \ADD_/FAINST[31].FA_/n2 , \ADD_/FAINST[31].FA_/n1 ,
         \ADD_/FAINST[30].FA_/n3 , \ADD_/FAINST[30].FA_/n2 ,
         \ADD_/FAINST[30].FA_/n1 , \ADD_/FAINST[29].FA_/n3 ,
         \ADD_/FAINST[29].FA_/n2 , \ADD_/FAINST[29].FA_/n1 ,
         \ADD_/FAINST[28].FA_/n3 , \ADD_/FAINST[28].FA_/n2 ,
         \ADD_/FAINST[28].FA_/n1 , \ADD_/FAINST[27].FA_/n3 ,
         \ADD_/FAINST[27].FA_/n2 , \ADD_/FAINST[27].FA_/n1 ,
         \ADD_/FAINST[26].FA_/n3 , \ADD_/FAINST[26].FA_/n2 ,
         \ADD_/FAINST[26].FA_/n1 , \ADD_/FAINST[25].FA_/n3 ,
         \ADD_/FAINST[25].FA_/n2 , \ADD_/FAINST[25].FA_/n1 ,
         \ADD_/FAINST[24].FA_/n3 , \ADD_/FAINST[24].FA_/n2 ,
         \ADD_/FAINST[24].FA_/n1 , \ADD_/FAINST[23].FA_/n3 ,
         \ADD_/FAINST[23].FA_/n2 , \ADD_/FAINST[23].FA_/n1 ,
         \ADD_/FAINST[22].FA_/n3 , \ADD_/FAINST[22].FA_/n2 ,
         \ADD_/FAINST[22].FA_/n1 , \ADD_/FAINST[21].FA_/n3 ,
         \ADD_/FAINST[21].FA_/n2 , \ADD_/FAINST[21].FA_/n1 ,
         \ADD_/FAINST[20].FA_/n3 , \ADD_/FAINST[20].FA_/n2 ,
         \ADD_/FAINST[20].FA_/n1 , \ADD_/FAINST[19].FA_/n3 ,
         \ADD_/FAINST[19].FA_/n2 , \ADD_/FAINST[19].FA_/n1 ,
         \ADD_/FAINST[18].FA_/n3 , \ADD_/FAINST[18].FA_/n2 ,
         \ADD_/FAINST[18].FA_/n1 , \ADD_/FAINST[17].FA_/n3 ,
         \ADD_/FAINST[17].FA_/n2 , \ADD_/FAINST[17].FA_/n1 ,
         \ADD_/FAINST[16].FA_/n3 , \ADD_/FAINST[16].FA_/n2 ,
         \ADD_/FAINST[16].FA_/n1 , \ADD_/FAINST[15].FA_/n3 ,
         \ADD_/FAINST[15].FA_/n2 , \ADD_/FAINST[15].FA_/n1 ,
         \ADD_/FAINST[14].FA_/n3 , \ADD_/FAINST[14].FA_/n2 ,
         \ADD_/FAINST[14].FA_/n1 , \ADD_/FAINST[13].FA_/n3 ,
         \ADD_/FAINST[13].FA_/n2 , \ADD_/FAINST[13].FA_/n1 ,
         \ADD_/FAINST[12].FA_/n3 , \ADD_/FAINST[12].FA_/n2 ,
         \ADD_/FAINST[12].FA_/n1 , \ADD_/FAINST[11].FA_/n3 ,
         \ADD_/FAINST[11].FA_/n2 , \ADD_/FAINST[11].FA_/n1 ,
         \ADD_/FAINST[10].FA_/n3 , \ADD_/FAINST[10].FA_/n2 ,
         \ADD_/FAINST[10].FA_/n1 , \ADD_/FAINST[9].FA_/n3 ,
         \ADD_/FAINST[9].FA_/n2 , \ADD_/FAINST[9].FA_/n1 ,
         \ADD_/FAINST[8].FA_/n3 , \ADD_/FAINST[8].FA_/n2 ,
         \ADD_/FAINST[8].FA_/n1 , \ADD_/FAINST[7].FA_/n3 ,
         \ADD_/FAINST[7].FA_/n2 , \ADD_/FAINST[7].FA_/n1 ,
         \ADD_/FAINST[6].FA_/n3 , \ADD_/FAINST[6].FA_/n2 ,
         \ADD_/FAINST[6].FA_/n1 , \ADD_/FAINST[5].FA_/n3 ,
         \ADD_/FAINST[5].FA_/n2 , \ADD_/FAINST[5].FA_/n1 ,
         \ADD_/FAINST[4].FA_/n3 , \ADD_/FAINST[4].FA_/n2 ,
         \ADD_/FAINST[4].FA_/n1 , \ADD_/FAINST[3].FA_/n3 ,
         \ADD_/FAINST[3].FA_/n2 , \ADD_/FAINST[3].FA_/n1 ,
         \ADD_/FAINST[2].FA_/n3 , \ADD_/FAINST[2].FA_/n2 ,
         \ADD_/FAINST[2].FA_/n1 , \ADD_/FAINST[1].FA_/n3 ,
         \ADD_/FAINST[1].FA_/n2 , \ADD_/FAINST[1].FA_/n1 ;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR \ADD_/FAINST[0].FA_/U5  ( .A(\ADD_/FAINST[0].FA_/n3 ), .B(carry_on), .Z(
        \ADD_/c[1] ) );
  XOR \ADD_/FAINST[0].FA_/U4  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(b[0]), .Z(c[0]) );
  AND \ADD_/FAINST[0].FA_/U3  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(
        \ADD_/FAINST[0].FA_/n2 ), .Z(\ADD_/FAINST[0].FA_/n3 ) );
  XOR \ADD_/FAINST[0].FA_/U2  ( .A(b[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n2 ) );
  XOR \ADD_/FAINST[0].FA_/U1  ( .A(a[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n1 ) );
  XOR \ADD_/FAINST[511].FA_/U5  ( .A(\ADD_/FAINST[511].FA_/n3 ), .B(
        \ADD_/c[511] ), .Z(carry_on_d) );
  XOR \ADD_/FAINST[511].FA_/U4  ( .A(\ADD_/FAINST[511].FA_/n1 ), .B(b[511]), 
        .Z(c[511]) );
  AND \ADD_/FAINST[511].FA_/U3  ( .A(\ADD_/FAINST[511].FA_/n1 ), .B(
        \ADD_/FAINST[511].FA_/n2 ), .Z(\ADD_/FAINST[511].FA_/n3 ) );
  XOR \ADD_/FAINST[511].FA_/U2  ( .A(b[511]), .B(\ADD_/c[511] ), .Z(
        \ADD_/FAINST[511].FA_/n2 ) );
  XOR \ADD_/FAINST[511].FA_/U1  ( .A(a[511]), .B(\ADD_/c[511] ), .Z(
        \ADD_/FAINST[511].FA_/n1 ) );
  XOR \ADD_/FAINST[510].FA_/U5  ( .A(\ADD_/FAINST[510].FA_/n3 ), .B(
        \ADD_/c[510] ), .Z(\ADD_/c[511] ) );
  XOR \ADD_/FAINST[510].FA_/U4  ( .A(\ADD_/FAINST[510].FA_/n1 ), .B(b[510]), 
        .Z(c[510]) );
  AND \ADD_/FAINST[510].FA_/U3  ( .A(\ADD_/FAINST[510].FA_/n1 ), .B(
        \ADD_/FAINST[510].FA_/n2 ), .Z(\ADD_/FAINST[510].FA_/n3 ) );
  XOR \ADD_/FAINST[510].FA_/U2  ( .A(b[510]), .B(\ADD_/c[510] ), .Z(
        \ADD_/FAINST[510].FA_/n2 ) );
  XOR \ADD_/FAINST[510].FA_/U1  ( .A(a[510]), .B(\ADD_/c[510] ), .Z(
        \ADD_/FAINST[510].FA_/n1 ) );
  XOR \ADD_/FAINST[509].FA_/U5  ( .A(\ADD_/FAINST[509].FA_/n3 ), .B(
        \ADD_/c[509] ), .Z(\ADD_/c[510] ) );
  XOR \ADD_/FAINST[509].FA_/U4  ( .A(\ADD_/FAINST[509].FA_/n1 ), .B(b[509]), 
        .Z(c[509]) );
  AND \ADD_/FAINST[509].FA_/U3  ( .A(\ADD_/FAINST[509].FA_/n1 ), .B(
        \ADD_/FAINST[509].FA_/n2 ), .Z(\ADD_/FAINST[509].FA_/n3 ) );
  XOR \ADD_/FAINST[509].FA_/U2  ( .A(b[509]), .B(\ADD_/c[509] ), .Z(
        \ADD_/FAINST[509].FA_/n2 ) );
  XOR \ADD_/FAINST[509].FA_/U1  ( .A(a[509]), .B(\ADD_/c[509] ), .Z(
        \ADD_/FAINST[509].FA_/n1 ) );
  XOR \ADD_/FAINST[508].FA_/U5  ( .A(\ADD_/FAINST[508].FA_/n3 ), .B(
        \ADD_/c[508] ), .Z(\ADD_/c[509] ) );
  XOR \ADD_/FAINST[508].FA_/U4  ( .A(\ADD_/FAINST[508].FA_/n1 ), .B(b[508]), 
        .Z(c[508]) );
  AND \ADD_/FAINST[508].FA_/U3  ( .A(\ADD_/FAINST[508].FA_/n1 ), .B(
        \ADD_/FAINST[508].FA_/n2 ), .Z(\ADD_/FAINST[508].FA_/n3 ) );
  XOR \ADD_/FAINST[508].FA_/U2  ( .A(b[508]), .B(\ADD_/c[508] ), .Z(
        \ADD_/FAINST[508].FA_/n2 ) );
  XOR \ADD_/FAINST[508].FA_/U1  ( .A(a[508]), .B(\ADD_/c[508] ), .Z(
        \ADD_/FAINST[508].FA_/n1 ) );
  XOR \ADD_/FAINST[507].FA_/U5  ( .A(\ADD_/FAINST[507].FA_/n3 ), .B(
        \ADD_/c[507] ), .Z(\ADD_/c[508] ) );
  XOR \ADD_/FAINST[507].FA_/U4  ( .A(\ADD_/FAINST[507].FA_/n1 ), .B(b[507]), 
        .Z(c[507]) );
  AND \ADD_/FAINST[507].FA_/U3  ( .A(\ADD_/FAINST[507].FA_/n1 ), .B(
        \ADD_/FAINST[507].FA_/n2 ), .Z(\ADD_/FAINST[507].FA_/n3 ) );
  XOR \ADD_/FAINST[507].FA_/U2  ( .A(b[507]), .B(\ADD_/c[507] ), .Z(
        \ADD_/FAINST[507].FA_/n2 ) );
  XOR \ADD_/FAINST[507].FA_/U1  ( .A(a[507]), .B(\ADD_/c[507] ), .Z(
        \ADD_/FAINST[507].FA_/n1 ) );
  XOR \ADD_/FAINST[506].FA_/U5  ( .A(\ADD_/FAINST[506].FA_/n3 ), .B(
        \ADD_/c[506] ), .Z(\ADD_/c[507] ) );
  XOR \ADD_/FAINST[506].FA_/U4  ( .A(\ADD_/FAINST[506].FA_/n1 ), .B(b[506]), 
        .Z(c[506]) );
  AND \ADD_/FAINST[506].FA_/U3  ( .A(\ADD_/FAINST[506].FA_/n1 ), .B(
        \ADD_/FAINST[506].FA_/n2 ), .Z(\ADD_/FAINST[506].FA_/n3 ) );
  XOR \ADD_/FAINST[506].FA_/U2  ( .A(b[506]), .B(\ADD_/c[506] ), .Z(
        \ADD_/FAINST[506].FA_/n2 ) );
  XOR \ADD_/FAINST[506].FA_/U1  ( .A(a[506]), .B(\ADD_/c[506] ), .Z(
        \ADD_/FAINST[506].FA_/n1 ) );
  XOR \ADD_/FAINST[505].FA_/U5  ( .A(\ADD_/FAINST[505].FA_/n3 ), .B(
        \ADD_/c[505] ), .Z(\ADD_/c[506] ) );
  XOR \ADD_/FAINST[505].FA_/U4  ( .A(\ADD_/FAINST[505].FA_/n1 ), .B(b[505]), 
        .Z(c[505]) );
  AND \ADD_/FAINST[505].FA_/U3  ( .A(\ADD_/FAINST[505].FA_/n1 ), .B(
        \ADD_/FAINST[505].FA_/n2 ), .Z(\ADD_/FAINST[505].FA_/n3 ) );
  XOR \ADD_/FAINST[505].FA_/U2  ( .A(b[505]), .B(\ADD_/c[505] ), .Z(
        \ADD_/FAINST[505].FA_/n2 ) );
  XOR \ADD_/FAINST[505].FA_/U1  ( .A(a[505]), .B(\ADD_/c[505] ), .Z(
        \ADD_/FAINST[505].FA_/n1 ) );
  XOR \ADD_/FAINST[504].FA_/U5  ( .A(\ADD_/FAINST[504].FA_/n3 ), .B(
        \ADD_/c[504] ), .Z(\ADD_/c[505] ) );
  XOR \ADD_/FAINST[504].FA_/U4  ( .A(\ADD_/FAINST[504].FA_/n1 ), .B(b[504]), 
        .Z(c[504]) );
  AND \ADD_/FAINST[504].FA_/U3  ( .A(\ADD_/FAINST[504].FA_/n1 ), .B(
        \ADD_/FAINST[504].FA_/n2 ), .Z(\ADD_/FAINST[504].FA_/n3 ) );
  XOR \ADD_/FAINST[504].FA_/U2  ( .A(b[504]), .B(\ADD_/c[504] ), .Z(
        \ADD_/FAINST[504].FA_/n2 ) );
  XOR \ADD_/FAINST[504].FA_/U1  ( .A(a[504]), .B(\ADD_/c[504] ), .Z(
        \ADD_/FAINST[504].FA_/n1 ) );
  XOR \ADD_/FAINST[503].FA_/U5  ( .A(\ADD_/FAINST[503].FA_/n3 ), .B(
        \ADD_/c[503] ), .Z(\ADD_/c[504] ) );
  XOR \ADD_/FAINST[503].FA_/U4  ( .A(\ADD_/FAINST[503].FA_/n1 ), .B(b[503]), 
        .Z(c[503]) );
  AND \ADD_/FAINST[503].FA_/U3  ( .A(\ADD_/FAINST[503].FA_/n1 ), .B(
        \ADD_/FAINST[503].FA_/n2 ), .Z(\ADD_/FAINST[503].FA_/n3 ) );
  XOR \ADD_/FAINST[503].FA_/U2  ( .A(b[503]), .B(\ADD_/c[503] ), .Z(
        \ADD_/FAINST[503].FA_/n2 ) );
  XOR \ADD_/FAINST[503].FA_/U1  ( .A(a[503]), .B(\ADD_/c[503] ), .Z(
        \ADD_/FAINST[503].FA_/n1 ) );
  XOR \ADD_/FAINST[502].FA_/U5  ( .A(\ADD_/FAINST[502].FA_/n3 ), .B(
        \ADD_/c[502] ), .Z(\ADD_/c[503] ) );
  XOR \ADD_/FAINST[502].FA_/U4  ( .A(\ADD_/FAINST[502].FA_/n1 ), .B(b[502]), 
        .Z(c[502]) );
  AND \ADD_/FAINST[502].FA_/U3  ( .A(\ADD_/FAINST[502].FA_/n1 ), .B(
        \ADD_/FAINST[502].FA_/n2 ), .Z(\ADD_/FAINST[502].FA_/n3 ) );
  XOR \ADD_/FAINST[502].FA_/U2  ( .A(b[502]), .B(\ADD_/c[502] ), .Z(
        \ADD_/FAINST[502].FA_/n2 ) );
  XOR \ADD_/FAINST[502].FA_/U1  ( .A(a[502]), .B(\ADD_/c[502] ), .Z(
        \ADD_/FAINST[502].FA_/n1 ) );
  XOR \ADD_/FAINST[501].FA_/U5  ( .A(\ADD_/FAINST[501].FA_/n3 ), .B(
        \ADD_/c[501] ), .Z(\ADD_/c[502] ) );
  XOR \ADD_/FAINST[501].FA_/U4  ( .A(\ADD_/FAINST[501].FA_/n1 ), .B(b[501]), 
        .Z(c[501]) );
  AND \ADD_/FAINST[501].FA_/U3  ( .A(\ADD_/FAINST[501].FA_/n1 ), .B(
        \ADD_/FAINST[501].FA_/n2 ), .Z(\ADD_/FAINST[501].FA_/n3 ) );
  XOR \ADD_/FAINST[501].FA_/U2  ( .A(b[501]), .B(\ADD_/c[501] ), .Z(
        \ADD_/FAINST[501].FA_/n2 ) );
  XOR \ADD_/FAINST[501].FA_/U1  ( .A(a[501]), .B(\ADD_/c[501] ), .Z(
        \ADD_/FAINST[501].FA_/n1 ) );
  XOR \ADD_/FAINST[500].FA_/U5  ( .A(\ADD_/FAINST[500].FA_/n3 ), .B(
        \ADD_/c[500] ), .Z(\ADD_/c[501] ) );
  XOR \ADD_/FAINST[500].FA_/U4  ( .A(\ADD_/FAINST[500].FA_/n1 ), .B(b[500]), 
        .Z(c[500]) );
  AND \ADD_/FAINST[500].FA_/U3  ( .A(\ADD_/FAINST[500].FA_/n1 ), .B(
        \ADD_/FAINST[500].FA_/n2 ), .Z(\ADD_/FAINST[500].FA_/n3 ) );
  XOR \ADD_/FAINST[500].FA_/U2  ( .A(b[500]), .B(\ADD_/c[500] ), .Z(
        \ADD_/FAINST[500].FA_/n2 ) );
  XOR \ADD_/FAINST[500].FA_/U1  ( .A(a[500]), .B(\ADD_/c[500] ), .Z(
        \ADD_/FAINST[500].FA_/n1 ) );
  XOR \ADD_/FAINST[499].FA_/U5  ( .A(\ADD_/FAINST[499].FA_/n3 ), .B(
        \ADD_/c[499] ), .Z(\ADD_/c[500] ) );
  XOR \ADD_/FAINST[499].FA_/U4  ( .A(\ADD_/FAINST[499].FA_/n1 ), .B(b[499]), 
        .Z(c[499]) );
  AND \ADD_/FAINST[499].FA_/U3  ( .A(\ADD_/FAINST[499].FA_/n1 ), .B(
        \ADD_/FAINST[499].FA_/n2 ), .Z(\ADD_/FAINST[499].FA_/n3 ) );
  XOR \ADD_/FAINST[499].FA_/U2  ( .A(b[499]), .B(\ADD_/c[499] ), .Z(
        \ADD_/FAINST[499].FA_/n2 ) );
  XOR \ADD_/FAINST[499].FA_/U1  ( .A(a[499]), .B(\ADD_/c[499] ), .Z(
        \ADD_/FAINST[499].FA_/n1 ) );
  XOR \ADD_/FAINST[498].FA_/U5  ( .A(\ADD_/FAINST[498].FA_/n3 ), .B(
        \ADD_/c[498] ), .Z(\ADD_/c[499] ) );
  XOR \ADD_/FAINST[498].FA_/U4  ( .A(\ADD_/FAINST[498].FA_/n1 ), .B(b[498]), 
        .Z(c[498]) );
  AND \ADD_/FAINST[498].FA_/U3  ( .A(\ADD_/FAINST[498].FA_/n1 ), .B(
        \ADD_/FAINST[498].FA_/n2 ), .Z(\ADD_/FAINST[498].FA_/n3 ) );
  XOR \ADD_/FAINST[498].FA_/U2  ( .A(b[498]), .B(\ADD_/c[498] ), .Z(
        \ADD_/FAINST[498].FA_/n2 ) );
  XOR \ADD_/FAINST[498].FA_/U1  ( .A(a[498]), .B(\ADD_/c[498] ), .Z(
        \ADD_/FAINST[498].FA_/n1 ) );
  XOR \ADD_/FAINST[497].FA_/U5  ( .A(\ADD_/FAINST[497].FA_/n3 ), .B(
        \ADD_/c[497] ), .Z(\ADD_/c[498] ) );
  XOR \ADD_/FAINST[497].FA_/U4  ( .A(\ADD_/FAINST[497].FA_/n1 ), .B(b[497]), 
        .Z(c[497]) );
  AND \ADD_/FAINST[497].FA_/U3  ( .A(\ADD_/FAINST[497].FA_/n1 ), .B(
        \ADD_/FAINST[497].FA_/n2 ), .Z(\ADD_/FAINST[497].FA_/n3 ) );
  XOR \ADD_/FAINST[497].FA_/U2  ( .A(b[497]), .B(\ADD_/c[497] ), .Z(
        \ADD_/FAINST[497].FA_/n2 ) );
  XOR \ADD_/FAINST[497].FA_/U1  ( .A(a[497]), .B(\ADD_/c[497] ), .Z(
        \ADD_/FAINST[497].FA_/n1 ) );
  XOR \ADD_/FAINST[496].FA_/U5  ( .A(\ADD_/FAINST[496].FA_/n3 ), .B(
        \ADD_/c[496] ), .Z(\ADD_/c[497] ) );
  XOR \ADD_/FAINST[496].FA_/U4  ( .A(\ADD_/FAINST[496].FA_/n1 ), .B(b[496]), 
        .Z(c[496]) );
  AND \ADD_/FAINST[496].FA_/U3  ( .A(\ADD_/FAINST[496].FA_/n1 ), .B(
        \ADD_/FAINST[496].FA_/n2 ), .Z(\ADD_/FAINST[496].FA_/n3 ) );
  XOR \ADD_/FAINST[496].FA_/U2  ( .A(b[496]), .B(\ADD_/c[496] ), .Z(
        \ADD_/FAINST[496].FA_/n2 ) );
  XOR \ADD_/FAINST[496].FA_/U1  ( .A(a[496]), .B(\ADD_/c[496] ), .Z(
        \ADD_/FAINST[496].FA_/n1 ) );
  XOR \ADD_/FAINST[495].FA_/U5  ( .A(\ADD_/FAINST[495].FA_/n3 ), .B(
        \ADD_/c[495] ), .Z(\ADD_/c[496] ) );
  XOR \ADD_/FAINST[495].FA_/U4  ( .A(\ADD_/FAINST[495].FA_/n1 ), .B(b[495]), 
        .Z(c[495]) );
  AND \ADD_/FAINST[495].FA_/U3  ( .A(\ADD_/FAINST[495].FA_/n1 ), .B(
        \ADD_/FAINST[495].FA_/n2 ), .Z(\ADD_/FAINST[495].FA_/n3 ) );
  XOR \ADD_/FAINST[495].FA_/U2  ( .A(b[495]), .B(\ADD_/c[495] ), .Z(
        \ADD_/FAINST[495].FA_/n2 ) );
  XOR \ADD_/FAINST[495].FA_/U1  ( .A(a[495]), .B(\ADD_/c[495] ), .Z(
        \ADD_/FAINST[495].FA_/n1 ) );
  XOR \ADD_/FAINST[494].FA_/U5  ( .A(\ADD_/FAINST[494].FA_/n3 ), .B(
        \ADD_/c[494] ), .Z(\ADD_/c[495] ) );
  XOR \ADD_/FAINST[494].FA_/U4  ( .A(\ADD_/FAINST[494].FA_/n1 ), .B(b[494]), 
        .Z(c[494]) );
  AND \ADD_/FAINST[494].FA_/U3  ( .A(\ADD_/FAINST[494].FA_/n1 ), .B(
        \ADD_/FAINST[494].FA_/n2 ), .Z(\ADD_/FAINST[494].FA_/n3 ) );
  XOR \ADD_/FAINST[494].FA_/U2  ( .A(b[494]), .B(\ADD_/c[494] ), .Z(
        \ADD_/FAINST[494].FA_/n2 ) );
  XOR \ADD_/FAINST[494].FA_/U1  ( .A(a[494]), .B(\ADD_/c[494] ), .Z(
        \ADD_/FAINST[494].FA_/n1 ) );
  XOR \ADD_/FAINST[493].FA_/U5  ( .A(\ADD_/FAINST[493].FA_/n3 ), .B(
        \ADD_/c[493] ), .Z(\ADD_/c[494] ) );
  XOR \ADD_/FAINST[493].FA_/U4  ( .A(\ADD_/FAINST[493].FA_/n1 ), .B(b[493]), 
        .Z(c[493]) );
  AND \ADD_/FAINST[493].FA_/U3  ( .A(\ADD_/FAINST[493].FA_/n1 ), .B(
        \ADD_/FAINST[493].FA_/n2 ), .Z(\ADD_/FAINST[493].FA_/n3 ) );
  XOR \ADD_/FAINST[493].FA_/U2  ( .A(b[493]), .B(\ADD_/c[493] ), .Z(
        \ADD_/FAINST[493].FA_/n2 ) );
  XOR \ADD_/FAINST[493].FA_/U1  ( .A(a[493]), .B(\ADD_/c[493] ), .Z(
        \ADD_/FAINST[493].FA_/n1 ) );
  XOR \ADD_/FAINST[492].FA_/U5  ( .A(\ADD_/FAINST[492].FA_/n3 ), .B(
        \ADD_/c[492] ), .Z(\ADD_/c[493] ) );
  XOR \ADD_/FAINST[492].FA_/U4  ( .A(\ADD_/FAINST[492].FA_/n1 ), .B(b[492]), 
        .Z(c[492]) );
  AND \ADD_/FAINST[492].FA_/U3  ( .A(\ADD_/FAINST[492].FA_/n1 ), .B(
        \ADD_/FAINST[492].FA_/n2 ), .Z(\ADD_/FAINST[492].FA_/n3 ) );
  XOR \ADD_/FAINST[492].FA_/U2  ( .A(b[492]), .B(\ADD_/c[492] ), .Z(
        \ADD_/FAINST[492].FA_/n2 ) );
  XOR \ADD_/FAINST[492].FA_/U1  ( .A(a[492]), .B(\ADD_/c[492] ), .Z(
        \ADD_/FAINST[492].FA_/n1 ) );
  XOR \ADD_/FAINST[491].FA_/U5  ( .A(\ADD_/FAINST[491].FA_/n3 ), .B(
        \ADD_/c[491] ), .Z(\ADD_/c[492] ) );
  XOR \ADD_/FAINST[491].FA_/U4  ( .A(\ADD_/FAINST[491].FA_/n1 ), .B(b[491]), 
        .Z(c[491]) );
  AND \ADD_/FAINST[491].FA_/U3  ( .A(\ADD_/FAINST[491].FA_/n1 ), .B(
        \ADD_/FAINST[491].FA_/n2 ), .Z(\ADD_/FAINST[491].FA_/n3 ) );
  XOR \ADD_/FAINST[491].FA_/U2  ( .A(b[491]), .B(\ADD_/c[491] ), .Z(
        \ADD_/FAINST[491].FA_/n2 ) );
  XOR \ADD_/FAINST[491].FA_/U1  ( .A(a[491]), .B(\ADD_/c[491] ), .Z(
        \ADD_/FAINST[491].FA_/n1 ) );
  XOR \ADD_/FAINST[490].FA_/U5  ( .A(\ADD_/FAINST[490].FA_/n3 ), .B(
        \ADD_/c[490] ), .Z(\ADD_/c[491] ) );
  XOR \ADD_/FAINST[490].FA_/U4  ( .A(\ADD_/FAINST[490].FA_/n1 ), .B(b[490]), 
        .Z(c[490]) );
  AND \ADD_/FAINST[490].FA_/U3  ( .A(\ADD_/FAINST[490].FA_/n1 ), .B(
        \ADD_/FAINST[490].FA_/n2 ), .Z(\ADD_/FAINST[490].FA_/n3 ) );
  XOR \ADD_/FAINST[490].FA_/U2  ( .A(b[490]), .B(\ADD_/c[490] ), .Z(
        \ADD_/FAINST[490].FA_/n2 ) );
  XOR \ADD_/FAINST[490].FA_/U1  ( .A(a[490]), .B(\ADD_/c[490] ), .Z(
        \ADD_/FAINST[490].FA_/n1 ) );
  XOR \ADD_/FAINST[489].FA_/U5  ( .A(\ADD_/FAINST[489].FA_/n3 ), .B(
        \ADD_/c[489] ), .Z(\ADD_/c[490] ) );
  XOR \ADD_/FAINST[489].FA_/U4  ( .A(\ADD_/FAINST[489].FA_/n1 ), .B(b[489]), 
        .Z(c[489]) );
  AND \ADD_/FAINST[489].FA_/U3  ( .A(\ADD_/FAINST[489].FA_/n1 ), .B(
        \ADD_/FAINST[489].FA_/n2 ), .Z(\ADD_/FAINST[489].FA_/n3 ) );
  XOR \ADD_/FAINST[489].FA_/U2  ( .A(b[489]), .B(\ADD_/c[489] ), .Z(
        \ADD_/FAINST[489].FA_/n2 ) );
  XOR \ADD_/FAINST[489].FA_/U1  ( .A(a[489]), .B(\ADD_/c[489] ), .Z(
        \ADD_/FAINST[489].FA_/n1 ) );
  XOR \ADD_/FAINST[488].FA_/U5  ( .A(\ADD_/FAINST[488].FA_/n3 ), .B(
        \ADD_/c[488] ), .Z(\ADD_/c[489] ) );
  XOR \ADD_/FAINST[488].FA_/U4  ( .A(\ADD_/FAINST[488].FA_/n1 ), .B(b[488]), 
        .Z(c[488]) );
  AND \ADD_/FAINST[488].FA_/U3  ( .A(\ADD_/FAINST[488].FA_/n1 ), .B(
        \ADD_/FAINST[488].FA_/n2 ), .Z(\ADD_/FAINST[488].FA_/n3 ) );
  XOR \ADD_/FAINST[488].FA_/U2  ( .A(b[488]), .B(\ADD_/c[488] ), .Z(
        \ADD_/FAINST[488].FA_/n2 ) );
  XOR \ADD_/FAINST[488].FA_/U1  ( .A(a[488]), .B(\ADD_/c[488] ), .Z(
        \ADD_/FAINST[488].FA_/n1 ) );
  XOR \ADD_/FAINST[487].FA_/U5  ( .A(\ADD_/FAINST[487].FA_/n3 ), .B(
        \ADD_/c[487] ), .Z(\ADD_/c[488] ) );
  XOR \ADD_/FAINST[487].FA_/U4  ( .A(\ADD_/FAINST[487].FA_/n1 ), .B(b[487]), 
        .Z(c[487]) );
  AND \ADD_/FAINST[487].FA_/U3  ( .A(\ADD_/FAINST[487].FA_/n1 ), .B(
        \ADD_/FAINST[487].FA_/n2 ), .Z(\ADD_/FAINST[487].FA_/n3 ) );
  XOR \ADD_/FAINST[487].FA_/U2  ( .A(b[487]), .B(\ADD_/c[487] ), .Z(
        \ADD_/FAINST[487].FA_/n2 ) );
  XOR \ADD_/FAINST[487].FA_/U1  ( .A(a[487]), .B(\ADD_/c[487] ), .Z(
        \ADD_/FAINST[487].FA_/n1 ) );
  XOR \ADD_/FAINST[486].FA_/U5  ( .A(\ADD_/FAINST[486].FA_/n3 ), .B(
        \ADD_/c[486] ), .Z(\ADD_/c[487] ) );
  XOR \ADD_/FAINST[486].FA_/U4  ( .A(\ADD_/FAINST[486].FA_/n1 ), .B(b[486]), 
        .Z(c[486]) );
  AND \ADD_/FAINST[486].FA_/U3  ( .A(\ADD_/FAINST[486].FA_/n1 ), .B(
        \ADD_/FAINST[486].FA_/n2 ), .Z(\ADD_/FAINST[486].FA_/n3 ) );
  XOR \ADD_/FAINST[486].FA_/U2  ( .A(b[486]), .B(\ADD_/c[486] ), .Z(
        \ADD_/FAINST[486].FA_/n2 ) );
  XOR \ADD_/FAINST[486].FA_/U1  ( .A(a[486]), .B(\ADD_/c[486] ), .Z(
        \ADD_/FAINST[486].FA_/n1 ) );
  XOR \ADD_/FAINST[485].FA_/U5  ( .A(\ADD_/FAINST[485].FA_/n3 ), .B(
        \ADD_/c[485] ), .Z(\ADD_/c[486] ) );
  XOR \ADD_/FAINST[485].FA_/U4  ( .A(\ADD_/FAINST[485].FA_/n1 ), .B(b[485]), 
        .Z(c[485]) );
  AND \ADD_/FAINST[485].FA_/U3  ( .A(\ADD_/FAINST[485].FA_/n1 ), .B(
        \ADD_/FAINST[485].FA_/n2 ), .Z(\ADD_/FAINST[485].FA_/n3 ) );
  XOR \ADD_/FAINST[485].FA_/U2  ( .A(b[485]), .B(\ADD_/c[485] ), .Z(
        \ADD_/FAINST[485].FA_/n2 ) );
  XOR \ADD_/FAINST[485].FA_/U1  ( .A(a[485]), .B(\ADD_/c[485] ), .Z(
        \ADD_/FAINST[485].FA_/n1 ) );
  XOR \ADD_/FAINST[484].FA_/U5  ( .A(\ADD_/FAINST[484].FA_/n3 ), .B(
        \ADD_/c[484] ), .Z(\ADD_/c[485] ) );
  XOR \ADD_/FAINST[484].FA_/U4  ( .A(\ADD_/FAINST[484].FA_/n1 ), .B(b[484]), 
        .Z(c[484]) );
  AND \ADD_/FAINST[484].FA_/U3  ( .A(\ADD_/FAINST[484].FA_/n1 ), .B(
        \ADD_/FAINST[484].FA_/n2 ), .Z(\ADD_/FAINST[484].FA_/n3 ) );
  XOR \ADD_/FAINST[484].FA_/U2  ( .A(b[484]), .B(\ADD_/c[484] ), .Z(
        \ADD_/FAINST[484].FA_/n2 ) );
  XOR \ADD_/FAINST[484].FA_/U1  ( .A(a[484]), .B(\ADD_/c[484] ), .Z(
        \ADD_/FAINST[484].FA_/n1 ) );
  XOR \ADD_/FAINST[483].FA_/U5  ( .A(\ADD_/FAINST[483].FA_/n3 ), .B(
        \ADD_/c[483] ), .Z(\ADD_/c[484] ) );
  XOR \ADD_/FAINST[483].FA_/U4  ( .A(\ADD_/FAINST[483].FA_/n1 ), .B(b[483]), 
        .Z(c[483]) );
  AND \ADD_/FAINST[483].FA_/U3  ( .A(\ADD_/FAINST[483].FA_/n1 ), .B(
        \ADD_/FAINST[483].FA_/n2 ), .Z(\ADD_/FAINST[483].FA_/n3 ) );
  XOR \ADD_/FAINST[483].FA_/U2  ( .A(b[483]), .B(\ADD_/c[483] ), .Z(
        \ADD_/FAINST[483].FA_/n2 ) );
  XOR \ADD_/FAINST[483].FA_/U1  ( .A(a[483]), .B(\ADD_/c[483] ), .Z(
        \ADD_/FAINST[483].FA_/n1 ) );
  XOR \ADD_/FAINST[482].FA_/U5  ( .A(\ADD_/FAINST[482].FA_/n3 ), .B(
        \ADD_/c[482] ), .Z(\ADD_/c[483] ) );
  XOR \ADD_/FAINST[482].FA_/U4  ( .A(\ADD_/FAINST[482].FA_/n1 ), .B(b[482]), 
        .Z(c[482]) );
  AND \ADD_/FAINST[482].FA_/U3  ( .A(\ADD_/FAINST[482].FA_/n1 ), .B(
        \ADD_/FAINST[482].FA_/n2 ), .Z(\ADD_/FAINST[482].FA_/n3 ) );
  XOR \ADD_/FAINST[482].FA_/U2  ( .A(b[482]), .B(\ADD_/c[482] ), .Z(
        \ADD_/FAINST[482].FA_/n2 ) );
  XOR \ADD_/FAINST[482].FA_/U1  ( .A(a[482]), .B(\ADD_/c[482] ), .Z(
        \ADD_/FAINST[482].FA_/n1 ) );
  XOR \ADD_/FAINST[481].FA_/U5  ( .A(\ADD_/FAINST[481].FA_/n3 ), .B(
        \ADD_/c[481] ), .Z(\ADD_/c[482] ) );
  XOR \ADD_/FAINST[481].FA_/U4  ( .A(\ADD_/FAINST[481].FA_/n1 ), .B(b[481]), 
        .Z(c[481]) );
  AND \ADD_/FAINST[481].FA_/U3  ( .A(\ADD_/FAINST[481].FA_/n1 ), .B(
        \ADD_/FAINST[481].FA_/n2 ), .Z(\ADD_/FAINST[481].FA_/n3 ) );
  XOR \ADD_/FAINST[481].FA_/U2  ( .A(b[481]), .B(\ADD_/c[481] ), .Z(
        \ADD_/FAINST[481].FA_/n2 ) );
  XOR \ADD_/FAINST[481].FA_/U1  ( .A(a[481]), .B(\ADD_/c[481] ), .Z(
        \ADD_/FAINST[481].FA_/n1 ) );
  XOR \ADD_/FAINST[480].FA_/U5  ( .A(\ADD_/FAINST[480].FA_/n3 ), .B(
        \ADD_/c[480] ), .Z(\ADD_/c[481] ) );
  XOR \ADD_/FAINST[480].FA_/U4  ( .A(\ADD_/FAINST[480].FA_/n1 ), .B(b[480]), 
        .Z(c[480]) );
  AND \ADD_/FAINST[480].FA_/U3  ( .A(\ADD_/FAINST[480].FA_/n1 ), .B(
        \ADD_/FAINST[480].FA_/n2 ), .Z(\ADD_/FAINST[480].FA_/n3 ) );
  XOR \ADD_/FAINST[480].FA_/U2  ( .A(b[480]), .B(\ADD_/c[480] ), .Z(
        \ADD_/FAINST[480].FA_/n2 ) );
  XOR \ADD_/FAINST[480].FA_/U1  ( .A(a[480]), .B(\ADD_/c[480] ), .Z(
        \ADD_/FAINST[480].FA_/n1 ) );
  XOR \ADD_/FAINST[479].FA_/U5  ( .A(\ADD_/FAINST[479].FA_/n3 ), .B(
        \ADD_/c[479] ), .Z(\ADD_/c[480] ) );
  XOR \ADD_/FAINST[479].FA_/U4  ( .A(\ADD_/FAINST[479].FA_/n1 ), .B(b[479]), 
        .Z(c[479]) );
  AND \ADD_/FAINST[479].FA_/U3  ( .A(\ADD_/FAINST[479].FA_/n1 ), .B(
        \ADD_/FAINST[479].FA_/n2 ), .Z(\ADD_/FAINST[479].FA_/n3 ) );
  XOR \ADD_/FAINST[479].FA_/U2  ( .A(b[479]), .B(\ADD_/c[479] ), .Z(
        \ADD_/FAINST[479].FA_/n2 ) );
  XOR \ADD_/FAINST[479].FA_/U1  ( .A(a[479]), .B(\ADD_/c[479] ), .Z(
        \ADD_/FAINST[479].FA_/n1 ) );
  XOR \ADD_/FAINST[478].FA_/U5  ( .A(\ADD_/FAINST[478].FA_/n3 ), .B(
        \ADD_/c[478] ), .Z(\ADD_/c[479] ) );
  XOR \ADD_/FAINST[478].FA_/U4  ( .A(\ADD_/FAINST[478].FA_/n1 ), .B(b[478]), 
        .Z(c[478]) );
  AND \ADD_/FAINST[478].FA_/U3  ( .A(\ADD_/FAINST[478].FA_/n1 ), .B(
        \ADD_/FAINST[478].FA_/n2 ), .Z(\ADD_/FAINST[478].FA_/n3 ) );
  XOR \ADD_/FAINST[478].FA_/U2  ( .A(b[478]), .B(\ADD_/c[478] ), .Z(
        \ADD_/FAINST[478].FA_/n2 ) );
  XOR \ADD_/FAINST[478].FA_/U1  ( .A(a[478]), .B(\ADD_/c[478] ), .Z(
        \ADD_/FAINST[478].FA_/n1 ) );
  XOR \ADD_/FAINST[477].FA_/U5  ( .A(\ADD_/FAINST[477].FA_/n3 ), .B(
        \ADD_/c[477] ), .Z(\ADD_/c[478] ) );
  XOR \ADD_/FAINST[477].FA_/U4  ( .A(\ADD_/FAINST[477].FA_/n1 ), .B(b[477]), 
        .Z(c[477]) );
  AND \ADD_/FAINST[477].FA_/U3  ( .A(\ADD_/FAINST[477].FA_/n1 ), .B(
        \ADD_/FAINST[477].FA_/n2 ), .Z(\ADD_/FAINST[477].FA_/n3 ) );
  XOR \ADD_/FAINST[477].FA_/U2  ( .A(b[477]), .B(\ADD_/c[477] ), .Z(
        \ADD_/FAINST[477].FA_/n2 ) );
  XOR \ADD_/FAINST[477].FA_/U1  ( .A(a[477]), .B(\ADD_/c[477] ), .Z(
        \ADD_/FAINST[477].FA_/n1 ) );
  XOR \ADD_/FAINST[476].FA_/U5  ( .A(\ADD_/FAINST[476].FA_/n3 ), .B(
        \ADD_/c[476] ), .Z(\ADD_/c[477] ) );
  XOR \ADD_/FAINST[476].FA_/U4  ( .A(\ADD_/FAINST[476].FA_/n1 ), .B(b[476]), 
        .Z(c[476]) );
  AND \ADD_/FAINST[476].FA_/U3  ( .A(\ADD_/FAINST[476].FA_/n1 ), .B(
        \ADD_/FAINST[476].FA_/n2 ), .Z(\ADD_/FAINST[476].FA_/n3 ) );
  XOR \ADD_/FAINST[476].FA_/U2  ( .A(b[476]), .B(\ADD_/c[476] ), .Z(
        \ADD_/FAINST[476].FA_/n2 ) );
  XOR \ADD_/FAINST[476].FA_/U1  ( .A(a[476]), .B(\ADD_/c[476] ), .Z(
        \ADD_/FAINST[476].FA_/n1 ) );
  XOR \ADD_/FAINST[475].FA_/U5  ( .A(\ADD_/FAINST[475].FA_/n3 ), .B(
        \ADD_/c[475] ), .Z(\ADD_/c[476] ) );
  XOR \ADD_/FAINST[475].FA_/U4  ( .A(\ADD_/FAINST[475].FA_/n1 ), .B(b[475]), 
        .Z(c[475]) );
  AND \ADD_/FAINST[475].FA_/U3  ( .A(\ADD_/FAINST[475].FA_/n1 ), .B(
        \ADD_/FAINST[475].FA_/n2 ), .Z(\ADD_/FAINST[475].FA_/n3 ) );
  XOR \ADD_/FAINST[475].FA_/U2  ( .A(b[475]), .B(\ADD_/c[475] ), .Z(
        \ADD_/FAINST[475].FA_/n2 ) );
  XOR \ADD_/FAINST[475].FA_/U1  ( .A(a[475]), .B(\ADD_/c[475] ), .Z(
        \ADD_/FAINST[475].FA_/n1 ) );
  XOR \ADD_/FAINST[474].FA_/U5  ( .A(\ADD_/FAINST[474].FA_/n3 ), .B(
        \ADD_/c[474] ), .Z(\ADD_/c[475] ) );
  XOR \ADD_/FAINST[474].FA_/U4  ( .A(\ADD_/FAINST[474].FA_/n1 ), .B(b[474]), 
        .Z(c[474]) );
  AND \ADD_/FAINST[474].FA_/U3  ( .A(\ADD_/FAINST[474].FA_/n1 ), .B(
        \ADD_/FAINST[474].FA_/n2 ), .Z(\ADD_/FAINST[474].FA_/n3 ) );
  XOR \ADD_/FAINST[474].FA_/U2  ( .A(b[474]), .B(\ADD_/c[474] ), .Z(
        \ADD_/FAINST[474].FA_/n2 ) );
  XOR \ADD_/FAINST[474].FA_/U1  ( .A(a[474]), .B(\ADD_/c[474] ), .Z(
        \ADD_/FAINST[474].FA_/n1 ) );
  XOR \ADD_/FAINST[473].FA_/U5  ( .A(\ADD_/FAINST[473].FA_/n3 ), .B(
        \ADD_/c[473] ), .Z(\ADD_/c[474] ) );
  XOR \ADD_/FAINST[473].FA_/U4  ( .A(\ADD_/FAINST[473].FA_/n1 ), .B(b[473]), 
        .Z(c[473]) );
  AND \ADD_/FAINST[473].FA_/U3  ( .A(\ADD_/FAINST[473].FA_/n1 ), .B(
        \ADD_/FAINST[473].FA_/n2 ), .Z(\ADD_/FAINST[473].FA_/n3 ) );
  XOR \ADD_/FAINST[473].FA_/U2  ( .A(b[473]), .B(\ADD_/c[473] ), .Z(
        \ADD_/FAINST[473].FA_/n2 ) );
  XOR \ADD_/FAINST[473].FA_/U1  ( .A(a[473]), .B(\ADD_/c[473] ), .Z(
        \ADD_/FAINST[473].FA_/n1 ) );
  XOR \ADD_/FAINST[472].FA_/U5  ( .A(\ADD_/FAINST[472].FA_/n3 ), .B(
        \ADD_/c[472] ), .Z(\ADD_/c[473] ) );
  XOR \ADD_/FAINST[472].FA_/U4  ( .A(\ADD_/FAINST[472].FA_/n1 ), .B(b[472]), 
        .Z(c[472]) );
  AND \ADD_/FAINST[472].FA_/U3  ( .A(\ADD_/FAINST[472].FA_/n1 ), .B(
        \ADD_/FAINST[472].FA_/n2 ), .Z(\ADD_/FAINST[472].FA_/n3 ) );
  XOR \ADD_/FAINST[472].FA_/U2  ( .A(b[472]), .B(\ADD_/c[472] ), .Z(
        \ADD_/FAINST[472].FA_/n2 ) );
  XOR \ADD_/FAINST[472].FA_/U1  ( .A(a[472]), .B(\ADD_/c[472] ), .Z(
        \ADD_/FAINST[472].FA_/n1 ) );
  XOR \ADD_/FAINST[471].FA_/U5  ( .A(\ADD_/FAINST[471].FA_/n3 ), .B(
        \ADD_/c[471] ), .Z(\ADD_/c[472] ) );
  XOR \ADD_/FAINST[471].FA_/U4  ( .A(\ADD_/FAINST[471].FA_/n1 ), .B(b[471]), 
        .Z(c[471]) );
  AND \ADD_/FAINST[471].FA_/U3  ( .A(\ADD_/FAINST[471].FA_/n1 ), .B(
        \ADD_/FAINST[471].FA_/n2 ), .Z(\ADD_/FAINST[471].FA_/n3 ) );
  XOR \ADD_/FAINST[471].FA_/U2  ( .A(b[471]), .B(\ADD_/c[471] ), .Z(
        \ADD_/FAINST[471].FA_/n2 ) );
  XOR \ADD_/FAINST[471].FA_/U1  ( .A(a[471]), .B(\ADD_/c[471] ), .Z(
        \ADD_/FAINST[471].FA_/n1 ) );
  XOR \ADD_/FAINST[470].FA_/U5  ( .A(\ADD_/FAINST[470].FA_/n3 ), .B(
        \ADD_/c[470] ), .Z(\ADD_/c[471] ) );
  XOR \ADD_/FAINST[470].FA_/U4  ( .A(\ADD_/FAINST[470].FA_/n1 ), .B(b[470]), 
        .Z(c[470]) );
  AND \ADD_/FAINST[470].FA_/U3  ( .A(\ADD_/FAINST[470].FA_/n1 ), .B(
        \ADD_/FAINST[470].FA_/n2 ), .Z(\ADD_/FAINST[470].FA_/n3 ) );
  XOR \ADD_/FAINST[470].FA_/U2  ( .A(b[470]), .B(\ADD_/c[470] ), .Z(
        \ADD_/FAINST[470].FA_/n2 ) );
  XOR \ADD_/FAINST[470].FA_/U1  ( .A(a[470]), .B(\ADD_/c[470] ), .Z(
        \ADD_/FAINST[470].FA_/n1 ) );
  XOR \ADD_/FAINST[469].FA_/U5  ( .A(\ADD_/FAINST[469].FA_/n3 ), .B(
        \ADD_/c[469] ), .Z(\ADD_/c[470] ) );
  XOR \ADD_/FAINST[469].FA_/U4  ( .A(\ADD_/FAINST[469].FA_/n1 ), .B(b[469]), 
        .Z(c[469]) );
  AND \ADD_/FAINST[469].FA_/U3  ( .A(\ADD_/FAINST[469].FA_/n1 ), .B(
        \ADD_/FAINST[469].FA_/n2 ), .Z(\ADD_/FAINST[469].FA_/n3 ) );
  XOR \ADD_/FAINST[469].FA_/U2  ( .A(b[469]), .B(\ADD_/c[469] ), .Z(
        \ADD_/FAINST[469].FA_/n2 ) );
  XOR \ADD_/FAINST[469].FA_/U1  ( .A(a[469]), .B(\ADD_/c[469] ), .Z(
        \ADD_/FAINST[469].FA_/n1 ) );
  XOR \ADD_/FAINST[468].FA_/U5  ( .A(\ADD_/FAINST[468].FA_/n3 ), .B(
        \ADD_/c[468] ), .Z(\ADD_/c[469] ) );
  XOR \ADD_/FAINST[468].FA_/U4  ( .A(\ADD_/FAINST[468].FA_/n1 ), .B(b[468]), 
        .Z(c[468]) );
  AND \ADD_/FAINST[468].FA_/U3  ( .A(\ADD_/FAINST[468].FA_/n1 ), .B(
        \ADD_/FAINST[468].FA_/n2 ), .Z(\ADD_/FAINST[468].FA_/n3 ) );
  XOR \ADD_/FAINST[468].FA_/U2  ( .A(b[468]), .B(\ADD_/c[468] ), .Z(
        \ADD_/FAINST[468].FA_/n2 ) );
  XOR \ADD_/FAINST[468].FA_/U1  ( .A(a[468]), .B(\ADD_/c[468] ), .Z(
        \ADD_/FAINST[468].FA_/n1 ) );
  XOR \ADD_/FAINST[467].FA_/U5  ( .A(\ADD_/FAINST[467].FA_/n3 ), .B(
        \ADD_/c[467] ), .Z(\ADD_/c[468] ) );
  XOR \ADD_/FAINST[467].FA_/U4  ( .A(\ADD_/FAINST[467].FA_/n1 ), .B(b[467]), 
        .Z(c[467]) );
  AND \ADD_/FAINST[467].FA_/U3  ( .A(\ADD_/FAINST[467].FA_/n1 ), .B(
        \ADD_/FAINST[467].FA_/n2 ), .Z(\ADD_/FAINST[467].FA_/n3 ) );
  XOR \ADD_/FAINST[467].FA_/U2  ( .A(b[467]), .B(\ADD_/c[467] ), .Z(
        \ADD_/FAINST[467].FA_/n2 ) );
  XOR \ADD_/FAINST[467].FA_/U1  ( .A(a[467]), .B(\ADD_/c[467] ), .Z(
        \ADD_/FAINST[467].FA_/n1 ) );
  XOR \ADD_/FAINST[466].FA_/U5  ( .A(\ADD_/FAINST[466].FA_/n3 ), .B(
        \ADD_/c[466] ), .Z(\ADD_/c[467] ) );
  XOR \ADD_/FAINST[466].FA_/U4  ( .A(\ADD_/FAINST[466].FA_/n1 ), .B(b[466]), 
        .Z(c[466]) );
  AND \ADD_/FAINST[466].FA_/U3  ( .A(\ADD_/FAINST[466].FA_/n1 ), .B(
        \ADD_/FAINST[466].FA_/n2 ), .Z(\ADD_/FAINST[466].FA_/n3 ) );
  XOR \ADD_/FAINST[466].FA_/U2  ( .A(b[466]), .B(\ADD_/c[466] ), .Z(
        \ADD_/FAINST[466].FA_/n2 ) );
  XOR \ADD_/FAINST[466].FA_/U1  ( .A(a[466]), .B(\ADD_/c[466] ), .Z(
        \ADD_/FAINST[466].FA_/n1 ) );
  XOR \ADD_/FAINST[465].FA_/U5  ( .A(\ADD_/FAINST[465].FA_/n3 ), .B(
        \ADD_/c[465] ), .Z(\ADD_/c[466] ) );
  XOR \ADD_/FAINST[465].FA_/U4  ( .A(\ADD_/FAINST[465].FA_/n1 ), .B(b[465]), 
        .Z(c[465]) );
  AND \ADD_/FAINST[465].FA_/U3  ( .A(\ADD_/FAINST[465].FA_/n1 ), .B(
        \ADD_/FAINST[465].FA_/n2 ), .Z(\ADD_/FAINST[465].FA_/n3 ) );
  XOR \ADD_/FAINST[465].FA_/U2  ( .A(b[465]), .B(\ADD_/c[465] ), .Z(
        \ADD_/FAINST[465].FA_/n2 ) );
  XOR \ADD_/FAINST[465].FA_/U1  ( .A(a[465]), .B(\ADD_/c[465] ), .Z(
        \ADD_/FAINST[465].FA_/n1 ) );
  XOR \ADD_/FAINST[464].FA_/U5  ( .A(\ADD_/FAINST[464].FA_/n3 ), .B(
        \ADD_/c[464] ), .Z(\ADD_/c[465] ) );
  XOR \ADD_/FAINST[464].FA_/U4  ( .A(\ADD_/FAINST[464].FA_/n1 ), .B(b[464]), 
        .Z(c[464]) );
  AND \ADD_/FAINST[464].FA_/U3  ( .A(\ADD_/FAINST[464].FA_/n1 ), .B(
        \ADD_/FAINST[464].FA_/n2 ), .Z(\ADD_/FAINST[464].FA_/n3 ) );
  XOR \ADD_/FAINST[464].FA_/U2  ( .A(b[464]), .B(\ADD_/c[464] ), .Z(
        \ADD_/FAINST[464].FA_/n2 ) );
  XOR \ADD_/FAINST[464].FA_/U1  ( .A(a[464]), .B(\ADD_/c[464] ), .Z(
        \ADD_/FAINST[464].FA_/n1 ) );
  XOR \ADD_/FAINST[463].FA_/U5  ( .A(\ADD_/FAINST[463].FA_/n3 ), .B(
        \ADD_/c[463] ), .Z(\ADD_/c[464] ) );
  XOR \ADD_/FAINST[463].FA_/U4  ( .A(\ADD_/FAINST[463].FA_/n1 ), .B(b[463]), 
        .Z(c[463]) );
  AND \ADD_/FAINST[463].FA_/U3  ( .A(\ADD_/FAINST[463].FA_/n1 ), .B(
        \ADD_/FAINST[463].FA_/n2 ), .Z(\ADD_/FAINST[463].FA_/n3 ) );
  XOR \ADD_/FAINST[463].FA_/U2  ( .A(b[463]), .B(\ADD_/c[463] ), .Z(
        \ADD_/FAINST[463].FA_/n2 ) );
  XOR \ADD_/FAINST[463].FA_/U1  ( .A(a[463]), .B(\ADD_/c[463] ), .Z(
        \ADD_/FAINST[463].FA_/n1 ) );
  XOR \ADD_/FAINST[462].FA_/U5  ( .A(\ADD_/FAINST[462].FA_/n3 ), .B(
        \ADD_/c[462] ), .Z(\ADD_/c[463] ) );
  XOR \ADD_/FAINST[462].FA_/U4  ( .A(\ADD_/FAINST[462].FA_/n1 ), .B(b[462]), 
        .Z(c[462]) );
  AND \ADD_/FAINST[462].FA_/U3  ( .A(\ADD_/FAINST[462].FA_/n1 ), .B(
        \ADD_/FAINST[462].FA_/n2 ), .Z(\ADD_/FAINST[462].FA_/n3 ) );
  XOR \ADD_/FAINST[462].FA_/U2  ( .A(b[462]), .B(\ADD_/c[462] ), .Z(
        \ADD_/FAINST[462].FA_/n2 ) );
  XOR \ADD_/FAINST[462].FA_/U1  ( .A(a[462]), .B(\ADD_/c[462] ), .Z(
        \ADD_/FAINST[462].FA_/n1 ) );
  XOR \ADD_/FAINST[461].FA_/U5  ( .A(\ADD_/FAINST[461].FA_/n3 ), .B(
        \ADD_/c[461] ), .Z(\ADD_/c[462] ) );
  XOR \ADD_/FAINST[461].FA_/U4  ( .A(\ADD_/FAINST[461].FA_/n1 ), .B(b[461]), 
        .Z(c[461]) );
  AND \ADD_/FAINST[461].FA_/U3  ( .A(\ADD_/FAINST[461].FA_/n1 ), .B(
        \ADD_/FAINST[461].FA_/n2 ), .Z(\ADD_/FAINST[461].FA_/n3 ) );
  XOR \ADD_/FAINST[461].FA_/U2  ( .A(b[461]), .B(\ADD_/c[461] ), .Z(
        \ADD_/FAINST[461].FA_/n2 ) );
  XOR \ADD_/FAINST[461].FA_/U1  ( .A(a[461]), .B(\ADD_/c[461] ), .Z(
        \ADD_/FAINST[461].FA_/n1 ) );
  XOR \ADD_/FAINST[460].FA_/U5  ( .A(\ADD_/FAINST[460].FA_/n3 ), .B(
        \ADD_/c[460] ), .Z(\ADD_/c[461] ) );
  XOR \ADD_/FAINST[460].FA_/U4  ( .A(\ADD_/FAINST[460].FA_/n1 ), .B(b[460]), 
        .Z(c[460]) );
  AND \ADD_/FAINST[460].FA_/U3  ( .A(\ADD_/FAINST[460].FA_/n1 ), .B(
        \ADD_/FAINST[460].FA_/n2 ), .Z(\ADD_/FAINST[460].FA_/n3 ) );
  XOR \ADD_/FAINST[460].FA_/U2  ( .A(b[460]), .B(\ADD_/c[460] ), .Z(
        \ADD_/FAINST[460].FA_/n2 ) );
  XOR \ADD_/FAINST[460].FA_/U1  ( .A(a[460]), .B(\ADD_/c[460] ), .Z(
        \ADD_/FAINST[460].FA_/n1 ) );
  XOR \ADD_/FAINST[459].FA_/U5  ( .A(\ADD_/FAINST[459].FA_/n3 ), .B(
        \ADD_/c[459] ), .Z(\ADD_/c[460] ) );
  XOR \ADD_/FAINST[459].FA_/U4  ( .A(\ADD_/FAINST[459].FA_/n1 ), .B(b[459]), 
        .Z(c[459]) );
  AND \ADD_/FAINST[459].FA_/U3  ( .A(\ADD_/FAINST[459].FA_/n1 ), .B(
        \ADD_/FAINST[459].FA_/n2 ), .Z(\ADD_/FAINST[459].FA_/n3 ) );
  XOR \ADD_/FAINST[459].FA_/U2  ( .A(b[459]), .B(\ADD_/c[459] ), .Z(
        \ADD_/FAINST[459].FA_/n2 ) );
  XOR \ADD_/FAINST[459].FA_/U1  ( .A(a[459]), .B(\ADD_/c[459] ), .Z(
        \ADD_/FAINST[459].FA_/n1 ) );
  XOR \ADD_/FAINST[458].FA_/U5  ( .A(\ADD_/FAINST[458].FA_/n3 ), .B(
        \ADD_/c[458] ), .Z(\ADD_/c[459] ) );
  XOR \ADD_/FAINST[458].FA_/U4  ( .A(\ADD_/FAINST[458].FA_/n1 ), .B(b[458]), 
        .Z(c[458]) );
  AND \ADD_/FAINST[458].FA_/U3  ( .A(\ADD_/FAINST[458].FA_/n1 ), .B(
        \ADD_/FAINST[458].FA_/n2 ), .Z(\ADD_/FAINST[458].FA_/n3 ) );
  XOR \ADD_/FAINST[458].FA_/U2  ( .A(b[458]), .B(\ADD_/c[458] ), .Z(
        \ADD_/FAINST[458].FA_/n2 ) );
  XOR \ADD_/FAINST[458].FA_/U1  ( .A(a[458]), .B(\ADD_/c[458] ), .Z(
        \ADD_/FAINST[458].FA_/n1 ) );
  XOR \ADD_/FAINST[457].FA_/U5  ( .A(\ADD_/FAINST[457].FA_/n3 ), .B(
        \ADD_/c[457] ), .Z(\ADD_/c[458] ) );
  XOR \ADD_/FAINST[457].FA_/U4  ( .A(\ADD_/FAINST[457].FA_/n1 ), .B(b[457]), 
        .Z(c[457]) );
  AND \ADD_/FAINST[457].FA_/U3  ( .A(\ADD_/FAINST[457].FA_/n1 ), .B(
        \ADD_/FAINST[457].FA_/n2 ), .Z(\ADD_/FAINST[457].FA_/n3 ) );
  XOR \ADD_/FAINST[457].FA_/U2  ( .A(b[457]), .B(\ADD_/c[457] ), .Z(
        \ADD_/FAINST[457].FA_/n2 ) );
  XOR \ADD_/FAINST[457].FA_/U1  ( .A(a[457]), .B(\ADD_/c[457] ), .Z(
        \ADD_/FAINST[457].FA_/n1 ) );
  XOR \ADD_/FAINST[456].FA_/U5  ( .A(\ADD_/FAINST[456].FA_/n3 ), .B(
        \ADD_/c[456] ), .Z(\ADD_/c[457] ) );
  XOR \ADD_/FAINST[456].FA_/U4  ( .A(\ADD_/FAINST[456].FA_/n1 ), .B(b[456]), 
        .Z(c[456]) );
  AND \ADD_/FAINST[456].FA_/U3  ( .A(\ADD_/FAINST[456].FA_/n1 ), .B(
        \ADD_/FAINST[456].FA_/n2 ), .Z(\ADD_/FAINST[456].FA_/n3 ) );
  XOR \ADD_/FAINST[456].FA_/U2  ( .A(b[456]), .B(\ADD_/c[456] ), .Z(
        \ADD_/FAINST[456].FA_/n2 ) );
  XOR \ADD_/FAINST[456].FA_/U1  ( .A(a[456]), .B(\ADD_/c[456] ), .Z(
        \ADD_/FAINST[456].FA_/n1 ) );
  XOR \ADD_/FAINST[455].FA_/U5  ( .A(\ADD_/FAINST[455].FA_/n3 ), .B(
        \ADD_/c[455] ), .Z(\ADD_/c[456] ) );
  XOR \ADD_/FAINST[455].FA_/U4  ( .A(\ADD_/FAINST[455].FA_/n1 ), .B(b[455]), 
        .Z(c[455]) );
  AND \ADD_/FAINST[455].FA_/U3  ( .A(\ADD_/FAINST[455].FA_/n1 ), .B(
        \ADD_/FAINST[455].FA_/n2 ), .Z(\ADD_/FAINST[455].FA_/n3 ) );
  XOR \ADD_/FAINST[455].FA_/U2  ( .A(b[455]), .B(\ADD_/c[455] ), .Z(
        \ADD_/FAINST[455].FA_/n2 ) );
  XOR \ADD_/FAINST[455].FA_/U1  ( .A(a[455]), .B(\ADD_/c[455] ), .Z(
        \ADD_/FAINST[455].FA_/n1 ) );
  XOR \ADD_/FAINST[454].FA_/U5  ( .A(\ADD_/FAINST[454].FA_/n3 ), .B(
        \ADD_/c[454] ), .Z(\ADD_/c[455] ) );
  XOR \ADD_/FAINST[454].FA_/U4  ( .A(\ADD_/FAINST[454].FA_/n1 ), .B(b[454]), 
        .Z(c[454]) );
  AND \ADD_/FAINST[454].FA_/U3  ( .A(\ADD_/FAINST[454].FA_/n1 ), .B(
        \ADD_/FAINST[454].FA_/n2 ), .Z(\ADD_/FAINST[454].FA_/n3 ) );
  XOR \ADD_/FAINST[454].FA_/U2  ( .A(b[454]), .B(\ADD_/c[454] ), .Z(
        \ADD_/FAINST[454].FA_/n2 ) );
  XOR \ADD_/FAINST[454].FA_/U1  ( .A(a[454]), .B(\ADD_/c[454] ), .Z(
        \ADD_/FAINST[454].FA_/n1 ) );
  XOR \ADD_/FAINST[453].FA_/U5  ( .A(\ADD_/FAINST[453].FA_/n3 ), .B(
        \ADD_/c[453] ), .Z(\ADD_/c[454] ) );
  XOR \ADD_/FAINST[453].FA_/U4  ( .A(\ADD_/FAINST[453].FA_/n1 ), .B(b[453]), 
        .Z(c[453]) );
  AND \ADD_/FAINST[453].FA_/U3  ( .A(\ADD_/FAINST[453].FA_/n1 ), .B(
        \ADD_/FAINST[453].FA_/n2 ), .Z(\ADD_/FAINST[453].FA_/n3 ) );
  XOR \ADD_/FAINST[453].FA_/U2  ( .A(b[453]), .B(\ADD_/c[453] ), .Z(
        \ADD_/FAINST[453].FA_/n2 ) );
  XOR \ADD_/FAINST[453].FA_/U1  ( .A(a[453]), .B(\ADD_/c[453] ), .Z(
        \ADD_/FAINST[453].FA_/n1 ) );
  XOR \ADD_/FAINST[452].FA_/U5  ( .A(\ADD_/FAINST[452].FA_/n3 ), .B(
        \ADD_/c[452] ), .Z(\ADD_/c[453] ) );
  XOR \ADD_/FAINST[452].FA_/U4  ( .A(\ADD_/FAINST[452].FA_/n1 ), .B(b[452]), 
        .Z(c[452]) );
  AND \ADD_/FAINST[452].FA_/U3  ( .A(\ADD_/FAINST[452].FA_/n1 ), .B(
        \ADD_/FAINST[452].FA_/n2 ), .Z(\ADD_/FAINST[452].FA_/n3 ) );
  XOR \ADD_/FAINST[452].FA_/U2  ( .A(b[452]), .B(\ADD_/c[452] ), .Z(
        \ADD_/FAINST[452].FA_/n2 ) );
  XOR \ADD_/FAINST[452].FA_/U1  ( .A(a[452]), .B(\ADD_/c[452] ), .Z(
        \ADD_/FAINST[452].FA_/n1 ) );
  XOR \ADD_/FAINST[451].FA_/U5  ( .A(\ADD_/FAINST[451].FA_/n3 ), .B(
        \ADD_/c[451] ), .Z(\ADD_/c[452] ) );
  XOR \ADD_/FAINST[451].FA_/U4  ( .A(\ADD_/FAINST[451].FA_/n1 ), .B(b[451]), 
        .Z(c[451]) );
  AND \ADD_/FAINST[451].FA_/U3  ( .A(\ADD_/FAINST[451].FA_/n1 ), .B(
        \ADD_/FAINST[451].FA_/n2 ), .Z(\ADD_/FAINST[451].FA_/n3 ) );
  XOR \ADD_/FAINST[451].FA_/U2  ( .A(b[451]), .B(\ADD_/c[451] ), .Z(
        \ADD_/FAINST[451].FA_/n2 ) );
  XOR \ADD_/FAINST[451].FA_/U1  ( .A(a[451]), .B(\ADD_/c[451] ), .Z(
        \ADD_/FAINST[451].FA_/n1 ) );
  XOR \ADD_/FAINST[450].FA_/U5  ( .A(\ADD_/FAINST[450].FA_/n3 ), .B(
        \ADD_/c[450] ), .Z(\ADD_/c[451] ) );
  XOR \ADD_/FAINST[450].FA_/U4  ( .A(\ADD_/FAINST[450].FA_/n1 ), .B(b[450]), 
        .Z(c[450]) );
  AND \ADD_/FAINST[450].FA_/U3  ( .A(\ADD_/FAINST[450].FA_/n1 ), .B(
        \ADD_/FAINST[450].FA_/n2 ), .Z(\ADD_/FAINST[450].FA_/n3 ) );
  XOR \ADD_/FAINST[450].FA_/U2  ( .A(b[450]), .B(\ADD_/c[450] ), .Z(
        \ADD_/FAINST[450].FA_/n2 ) );
  XOR \ADD_/FAINST[450].FA_/U1  ( .A(a[450]), .B(\ADD_/c[450] ), .Z(
        \ADD_/FAINST[450].FA_/n1 ) );
  XOR \ADD_/FAINST[449].FA_/U5  ( .A(\ADD_/FAINST[449].FA_/n3 ), .B(
        \ADD_/c[449] ), .Z(\ADD_/c[450] ) );
  XOR \ADD_/FAINST[449].FA_/U4  ( .A(\ADD_/FAINST[449].FA_/n1 ), .B(b[449]), 
        .Z(c[449]) );
  AND \ADD_/FAINST[449].FA_/U3  ( .A(\ADD_/FAINST[449].FA_/n1 ), .B(
        \ADD_/FAINST[449].FA_/n2 ), .Z(\ADD_/FAINST[449].FA_/n3 ) );
  XOR \ADD_/FAINST[449].FA_/U2  ( .A(b[449]), .B(\ADD_/c[449] ), .Z(
        \ADD_/FAINST[449].FA_/n2 ) );
  XOR \ADD_/FAINST[449].FA_/U1  ( .A(a[449]), .B(\ADD_/c[449] ), .Z(
        \ADD_/FAINST[449].FA_/n1 ) );
  XOR \ADD_/FAINST[448].FA_/U5  ( .A(\ADD_/FAINST[448].FA_/n3 ), .B(
        \ADD_/c[448] ), .Z(\ADD_/c[449] ) );
  XOR \ADD_/FAINST[448].FA_/U4  ( .A(\ADD_/FAINST[448].FA_/n1 ), .B(b[448]), 
        .Z(c[448]) );
  AND \ADD_/FAINST[448].FA_/U3  ( .A(\ADD_/FAINST[448].FA_/n1 ), .B(
        \ADD_/FAINST[448].FA_/n2 ), .Z(\ADD_/FAINST[448].FA_/n3 ) );
  XOR \ADD_/FAINST[448].FA_/U2  ( .A(b[448]), .B(\ADD_/c[448] ), .Z(
        \ADD_/FAINST[448].FA_/n2 ) );
  XOR \ADD_/FAINST[448].FA_/U1  ( .A(a[448]), .B(\ADD_/c[448] ), .Z(
        \ADD_/FAINST[448].FA_/n1 ) );
  XOR \ADD_/FAINST[447].FA_/U5  ( .A(\ADD_/FAINST[447].FA_/n3 ), .B(
        \ADD_/c[447] ), .Z(\ADD_/c[448] ) );
  XOR \ADD_/FAINST[447].FA_/U4  ( .A(\ADD_/FAINST[447].FA_/n1 ), .B(b[447]), 
        .Z(c[447]) );
  AND \ADD_/FAINST[447].FA_/U3  ( .A(\ADD_/FAINST[447].FA_/n1 ), .B(
        \ADD_/FAINST[447].FA_/n2 ), .Z(\ADD_/FAINST[447].FA_/n3 ) );
  XOR \ADD_/FAINST[447].FA_/U2  ( .A(b[447]), .B(\ADD_/c[447] ), .Z(
        \ADD_/FAINST[447].FA_/n2 ) );
  XOR \ADD_/FAINST[447].FA_/U1  ( .A(a[447]), .B(\ADD_/c[447] ), .Z(
        \ADD_/FAINST[447].FA_/n1 ) );
  XOR \ADD_/FAINST[446].FA_/U5  ( .A(\ADD_/FAINST[446].FA_/n3 ), .B(
        \ADD_/c[446] ), .Z(\ADD_/c[447] ) );
  XOR \ADD_/FAINST[446].FA_/U4  ( .A(\ADD_/FAINST[446].FA_/n1 ), .B(b[446]), 
        .Z(c[446]) );
  AND \ADD_/FAINST[446].FA_/U3  ( .A(\ADD_/FAINST[446].FA_/n1 ), .B(
        \ADD_/FAINST[446].FA_/n2 ), .Z(\ADD_/FAINST[446].FA_/n3 ) );
  XOR \ADD_/FAINST[446].FA_/U2  ( .A(b[446]), .B(\ADD_/c[446] ), .Z(
        \ADD_/FAINST[446].FA_/n2 ) );
  XOR \ADD_/FAINST[446].FA_/U1  ( .A(a[446]), .B(\ADD_/c[446] ), .Z(
        \ADD_/FAINST[446].FA_/n1 ) );
  XOR \ADD_/FAINST[445].FA_/U5  ( .A(\ADD_/FAINST[445].FA_/n3 ), .B(
        \ADD_/c[445] ), .Z(\ADD_/c[446] ) );
  XOR \ADD_/FAINST[445].FA_/U4  ( .A(\ADD_/FAINST[445].FA_/n1 ), .B(b[445]), 
        .Z(c[445]) );
  AND \ADD_/FAINST[445].FA_/U3  ( .A(\ADD_/FAINST[445].FA_/n1 ), .B(
        \ADD_/FAINST[445].FA_/n2 ), .Z(\ADD_/FAINST[445].FA_/n3 ) );
  XOR \ADD_/FAINST[445].FA_/U2  ( .A(b[445]), .B(\ADD_/c[445] ), .Z(
        \ADD_/FAINST[445].FA_/n2 ) );
  XOR \ADD_/FAINST[445].FA_/U1  ( .A(a[445]), .B(\ADD_/c[445] ), .Z(
        \ADD_/FAINST[445].FA_/n1 ) );
  XOR \ADD_/FAINST[444].FA_/U5  ( .A(\ADD_/FAINST[444].FA_/n3 ), .B(
        \ADD_/c[444] ), .Z(\ADD_/c[445] ) );
  XOR \ADD_/FAINST[444].FA_/U4  ( .A(\ADD_/FAINST[444].FA_/n1 ), .B(b[444]), 
        .Z(c[444]) );
  AND \ADD_/FAINST[444].FA_/U3  ( .A(\ADD_/FAINST[444].FA_/n1 ), .B(
        \ADD_/FAINST[444].FA_/n2 ), .Z(\ADD_/FAINST[444].FA_/n3 ) );
  XOR \ADD_/FAINST[444].FA_/U2  ( .A(b[444]), .B(\ADD_/c[444] ), .Z(
        \ADD_/FAINST[444].FA_/n2 ) );
  XOR \ADD_/FAINST[444].FA_/U1  ( .A(a[444]), .B(\ADD_/c[444] ), .Z(
        \ADD_/FAINST[444].FA_/n1 ) );
  XOR \ADD_/FAINST[443].FA_/U5  ( .A(\ADD_/FAINST[443].FA_/n3 ), .B(
        \ADD_/c[443] ), .Z(\ADD_/c[444] ) );
  XOR \ADD_/FAINST[443].FA_/U4  ( .A(\ADD_/FAINST[443].FA_/n1 ), .B(b[443]), 
        .Z(c[443]) );
  AND \ADD_/FAINST[443].FA_/U3  ( .A(\ADD_/FAINST[443].FA_/n1 ), .B(
        \ADD_/FAINST[443].FA_/n2 ), .Z(\ADD_/FAINST[443].FA_/n3 ) );
  XOR \ADD_/FAINST[443].FA_/U2  ( .A(b[443]), .B(\ADD_/c[443] ), .Z(
        \ADD_/FAINST[443].FA_/n2 ) );
  XOR \ADD_/FAINST[443].FA_/U1  ( .A(a[443]), .B(\ADD_/c[443] ), .Z(
        \ADD_/FAINST[443].FA_/n1 ) );
  XOR \ADD_/FAINST[442].FA_/U5  ( .A(\ADD_/FAINST[442].FA_/n3 ), .B(
        \ADD_/c[442] ), .Z(\ADD_/c[443] ) );
  XOR \ADD_/FAINST[442].FA_/U4  ( .A(\ADD_/FAINST[442].FA_/n1 ), .B(b[442]), 
        .Z(c[442]) );
  AND \ADD_/FAINST[442].FA_/U3  ( .A(\ADD_/FAINST[442].FA_/n1 ), .B(
        \ADD_/FAINST[442].FA_/n2 ), .Z(\ADD_/FAINST[442].FA_/n3 ) );
  XOR \ADD_/FAINST[442].FA_/U2  ( .A(b[442]), .B(\ADD_/c[442] ), .Z(
        \ADD_/FAINST[442].FA_/n2 ) );
  XOR \ADD_/FAINST[442].FA_/U1  ( .A(a[442]), .B(\ADD_/c[442] ), .Z(
        \ADD_/FAINST[442].FA_/n1 ) );
  XOR \ADD_/FAINST[441].FA_/U5  ( .A(\ADD_/FAINST[441].FA_/n3 ), .B(
        \ADD_/c[441] ), .Z(\ADD_/c[442] ) );
  XOR \ADD_/FAINST[441].FA_/U4  ( .A(\ADD_/FAINST[441].FA_/n1 ), .B(b[441]), 
        .Z(c[441]) );
  AND \ADD_/FAINST[441].FA_/U3  ( .A(\ADD_/FAINST[441].FA_/n1 ), .B(
        \ADD_/FAINST[441].FA_/n2 ), .Z(\ADD_/FAINST[441].FA_/n3 ) );
  XOR \ADD_/FAINST[441].FA_/U2  ( .A(b[441]), .B(\ADD_/c[441] ), .Z(
        \ADD_/FAINST[441].FA_/n2 ) );
  XOR \ADD_/FAINST[441].FA_/U1  ( .A(a[441]), .B(\ADD_/c[441] ), .Z(
        \ADD_/FAINST[441].FA_/n1 ) );
  XOR \ADD_/FAINST[440].FA_/U5  ( .A(\ADD_/FAINST[440].FA_/n3 ), .B(
        \ADD_/c[440] ), .Z(\ADD_/c[441] ) );
  XOR \ADD_/FAINST[440].FA_/U4  ( .A(\ADD_/FAINST[440].FA_/n1 ), .B(b[440]), 
        .Z(c[440]) );
  AND \ADD_/FAINST[440].FA_/U3  ( .A(\ADD_/FAINST[440].FA_/n1 ), .B(
        \ADD_/FAINST[440].FA_/n2 ), .Z(\ADD_/FAINST[440].FA_/n3 ) );
  XOR \ADD_/FAINST[440].FA_/U2  ( .A(b[440]), .B(\ADD_/c[440] ), .Z(
        \ADD_/FAINST[440].FA_/n2 ) );
  XOR \ADD_/FAINST[440].FA_/U1  ( .A(a[440]), .B(\ADD_/c[440] ), .Z(
        \ADD_/FAINST[440].FA_/n1 ) );
  XOR \ADD_/FAINST[439].FA_/U5  ( .A(\ADD_/FAINST[439].FA_/n3 ), .B(
        \ADD_/c[439] ), .Z(\ADD_/c[440] ) );
  XOR \ADD_/FAINST[439].FA_/U4  ( .A(\ADD_/FAINST[439].FA_/n1 ), .B(b[439]), 
        .Z(c[439]) );
  AND \ADD_/FAINST[439].FA_/U3  ( .A(\ADD_/FAINST[439].FA_/n1 ), .B(
        \ADD_/FAINST[439].FA_/n2 ), .Z(\ADD_/FAINST[439].FA_/n3 ) );
  XOR \ADD_/FAINST[439].FA_/U2  ( .A(b[439]), .B(\ADD_/c[439] ), .Z(
        \ADD_/FAINST[439].FA_/n2 ) );
  XOR \ADD_/FAINST[439].FA_/U1  ( .A(a[439]), .B(\ADD_/c[439] ), .Z(
        \ADD_/FAINST[439].FA_/n1 ) );
  XOR \ADD_/FAINST[438].FA_/U5  ( .A(\ADD_/FAINST[438].FA_/n3 ), .B(
        \ADD_/c[438] ), .Z(\ADD_/c[439] ) );
  XOR \ADD_/FAINST[438].FA_/U4  ( .A(\ADD_/FAINST[438].FA_/n1 ), .B(b[438]), 
        .Z(c[438]) );
  AND \ADD_/FAINST[438].FA_/U3  ( .A(\ADD_/FAINST[438].FA_/n1 ), .B(
        \ADD_/FAINST[438].FA_/n2 ), .Z(\ADD_/FAINST[438].FA_/n3 ) );
  XOR \ADD_/FAINST[438].FA_/U2  ( .A(b[438]), .B(\ADD_/c[438] ), .Z(
        \ADD_/FAINST[438].FA_/n2 ) );
  XOR \ADD_/FAINST[438].FA_/U1  ( .A(a[438]), .B(\ADD_/c[438] ), .Z(
        \ADD_/FAINST[438].FA_/n1 ) );
  XOR \ADD_/FAINST[437].FA_/U5  ( .A(\ADD_/FAINST[437].FA_/n3 ), .B(
        \ADD_/c[437] ), .Z(\ADD_/c[438] ) );
  XOR \ADD_/FAINST[437].FA_/U4  ( .A(\ADD_/FAINST[437].FA_/n1 ), .B(b[437]), 
        .Z(c[437]) );
  AND \ADD_/FAINST[437].FA_/U3  ( .A(\ADD_/FAINST[437].FA_/n1 ), .B(
        \ADD_/FAINST[437].FA_/n2 ), .Z(\ADD_/FAINST[437].FA_/n3 ) );
  XOR \ADD_/FAINST[437].FA_/U2  ( .A(b[437]), .B(\ADD_/c[437] ), .Z(
        \ADD_/FAINST[437].FA_/n2 ) );
  XOR \ADD_/FAINST[437].FA_/U1  ( .A(a[437]), .B(\ADD_/c[437] ), .Z(
        \ADD_/FAINST[437].FA_/n1 ) );
  XOR \ADD_/FAINST[436].FA_/U5  ( .A(\ADD_/FAINST[436].FA_/n3 ), .B(
        \ADD_/c[436] ), .Z(\ADD_/c[437] ) );
  XOR \ADD_/FAINST[436].FA_/U4  ( .A(\ADD_/FAINST[436].FA_/n1 ), .B(b[436]), 
        .Z(c[436]) );
  AND \ADD_/FAINST[436].FA_/U3  ( .A(\ADD_/FAINST[436].FA_/n1 ), .B(
        \ADD_/FAINST[436].FA_/n2 ), .Z(\ADD_/FAINST[436].FA_/n3 ) );
  XOR \ADD_/FAINST[436].FA_/U2  ( .A(b[436]), .B(\ADD_/c[436] ), .Z(
        \ADD_/FAINST[436].FA_/n2 ) );
  XOR \ADD_/FAINST[436].FA_/U1  ( .A(a[436]), .B(\ADD_/c[436] ), .Z(
        \ADD_/FAINST[436].FA_/n1 ) );
  XOR \ADD_/FAINST[435].FA_/U5  ( .A(\ADD_/FAINST[435].FA_/n3 ), .B(
        \ADD_/c[435] ), .Z(\ADD_/c[436] ) );
  XOR \ADD_/FAINST[435].FA_/U4  ( .A(\ADD_/FAINST[435].FA_/n1 ), .B(b[435]), 
        .Z(c[435]) );
  AND \ADD_/FAINST[435].FA_/U3  ( .A(\ADD_/FAINST[435].FA_/n1 ), .B(
        \ADD_/FAINST[435].FA_/n2 ), .Z(\ADD_/FAINST[435].FA_/n3 ) );
  XOR \ADD_/FAINST[435].FA_/U2  ( .A(b[435]), .B(\ADD_/c[435] ), .Z(
        \ADD_/FAINST[435].FA_/n2 ) );
  XOR \ADD_/FAINST[435].FA_/U1  ( .A(a[435]), .B(\ADD_/c[435] ), .Z(
        \ADD_/FAINST[435].FA_/n1 ) );
  XOR \ADD_/FAINST[434].FA_/U5  ( .A(\ADD_/FAINST[434].FA_/n3 ), .B(
        \ADD_/c[434] ), .Z(\ADD_/c[435] ) );
  XOR \ADD_/FAINST[434].FA_/U4  ( .A(\ADD_/FAINST[434].FA_/n1 ), .B(b[434]), 
        .Z(c[434]) );
  AND \ADD_/FAINST[434].FA_/U3  ( .A(\ADD_/FAINST[434].FA_/n1 ), .B(
        \ADD_/FAINST[434].FA_/n2 ), .Z(\ADD_/FAINST[434].FA_/n3 ) );
  XOR \ADD_/FAINST[434].FA_/U2  ( .A(b[434]), .B(\ADD_/c[434] ), .Z(
        \ADD_/FAINST[434].FA_/n2 ) );
  XOR \ADD_/FAINST[434].FA_/U1  ( .A(a[434]), .B(\ADD_/c[434] ), .Z(
        \ADD_/FAINST[434].FA_/n1 ) );
  XOR \ADD_/FAINST[433].FA_/U5  ( .A(\ADD_/FAINST[433].FA_/n3 ), .B(
        \ADD_/c[433] ), .Z(\ADD_/c[434] ) );
  XOR \ADD_/FAINST[433].FA_/U4  ( .A(\ADD_/FAINST[433].FA_/n1 ), .B(b[433]), 
        .Z(c[433]) );
  AND \ADD_/FAINST[433].FA_/U3  ( .A(\ADD_/FAINST[433].FA_/n1 ), .B(
        \ADD_/FAINST[433].FA_/n2 ), .Z(\ADD_/FAINST[433].FA_/n3 ) );
  XOR \ADD_/FAINST[433].FA_/U2  ( .A(b[433]), .B(\ADD_/c[433] ), .Z(
        \ADD_/FAINST[433].FA_/n2 ) );
  XOR \ADD_/FAINST[433].FA_/U1  ( .A(a[433]), .B(\ADD_/c[433] ), .Z(
        \ADD_/FAINST[433].FA_/n1 ) );
  XOR \ADD_/FAINST[432].FA_/U5  ( .A(\ADD_/FAINST[432].FA_/n3 ), .B(
        \ADD_/c[432] ), .Z(\ADD_/c[433] ) );
  XOR \ADD_/FAINST[432].FA_/U4  ( .A(\ADD_/FAINST[432].FA_/n1 ), .B(b[432]), 
        .Z(c[432]) );
  AND \ADD_/FAINST[432].FA_/U3  ( .A(\ADD_/FAINST[432].FA_/n1 ), .B(
        \ADD_/FAINST[432].FA_/n2 ), .Z(\ADD_/FAINST[432].FA_/n3 ) );
  XOR \ADD_/FAINST[432].FA_/U2  ( .A(b[432]), .B(\ADD_/c[432] ), .Z(
        \ADD_/FAINST[432].FA_/n2 ) );
  XOR \ADD_/FAINST[432].FA_/U1  ( .A(a[432]), .B(\ADD_/c[432] ), .Z(
        \ADD_/FAINST[432].FA_/n1 ) );
  XOR \ADD_/FAINST[431].FA_/U5  ( .A(\ADD_/FAINST[431].FA_/n3 ), .B(
        \ADD_/c[431] ), .Z(\ADD_/c[432] ) );
  XOR \ADD_/FAINST[431].FA_/U4  ( .A(\ADD_/FAINST[431].FA_/n1 ), .B(b[431]), 
        .Z(c[431]) );
  AND \ADD_/FAINST[431].FA_/U3  ( .A(\ADD_/FAINST[431].FA_/n1 ), .B(
        \ADD_/FAINST[431].FA_/n2 ), .Z(\ADD_/FAINST[431].FA_/n3 ) );
  XOR \ADD_/FAINST[431].FA_/U2  ( .A(b[431]), .B(\ADD_/c[431] ), .Z(
        \ADD_/FAINST[431].FA_/n2 ) );
  XOR \ADD_/FAINST[431].FA_/U1  ( .A(a[431]), .B(\ADD_/c[431] ), .Z(
        \ADD_/FAINST[431].FA_/n1 ) );
  XOR \ADD_/FAINST[430].FA_/U5  ( .A(\ADD_/FAINST[430].FA_/n3 ), .B(
        \ADD_/c[430] ), .Z(\ADD_/c[431] ) );
  XOR \ADD_/FAINST[430].FA_/U4  ( .A(\ADD_/FAINST[430].FA_/n1 ), .B(b[430]), 
        .Z(c[430]) );
  AND \ADD_/FAINST[430].FA_/U3  ( .A(\ADD_/FAINST[430].FA_/n1 ), .B(
        \ADD_/FAINST[430].FA_/n2 ), .Z(\ADD_/FAINST[430].FA_/n3 ) );
  XOR \ADD_/FAINST[430].FA_/U2  ( .A(b[430]), .B(\ADD_/c[430] ), .Z(
        \ADD_/FAINST[430].FA_/n2 ) );
  XOR \ADD_/FAINST[430].FA_/U1  ( .A(a[430]), .B(\ADD_/c[430] ), .Z(
        \ADD_/FAINST[430].FA_/n1 ) );
  XOR \ADD_/FAINST[429].FA_/U5  ( .A(\ADD_/FAINST[429].FA_/n3 ), .B(
        \ADD_/c[429] ), .Z(\ADD_/c[430] ) );
  XOR \ADD_/FAINST[429].FA_/U4  ( .A(\ADD_/FAINST[429].FA_/n1 ), .B(b[429]), 
        .Z(c[429]) );
  AND \ADD_/FAINST[429].FA_/U3  ( .A(\ADD_/FAINST[429].FA_/n1 ), .B(
        \ADD_/FAINST[429].FA_/n2 ), .Z(\ADD_/FAINST[429].FA_/n3 ) );
  XOR \ADD_/FAINST[429].FA_/U2  ( .A(b[429]), .B(\ADD_/c[429] ), .Z(
        \ADD_/FAINST[429].FA_/n2 ) );
  XOR \ADD_/FAINST[429].FA_/U1  ( .A(a[429]), .B(\ADD_/c[429] ), .Z(
        \ADD_/FAINST[429].FA_/n1 ) );
  XOR \ADD_/FAINST[428].FA_/U5  ( .A(\ADD_/FAINST[428].FA_/n3 ), .B(
        \ADD_/c[428] ), .Z(\ADD_/c[429] ) );
  XOR \ADD_/FAINST[428].FA_/U4  ( .A(\ADD_/FAINST[428].FA_/n1 ), .B(b[428]), 
        .Z(c[428]) );
  AND \ADD_/FAINST[428].FA_/U3  ( .A(\ADD_/FAINST[428].FA_/n1 ), .B(
        \ADD_/FAINST[428].FA_/n2 ), .Z(\ADD_/FAINST[428].FA_/n3 ) );
  XOR \ADD_/FAINST[428].FA_/U2  ( .A(b[428]), .B(\ADD_/c[428] ), .Z(
        \ADD_/FAINST[428].FA_/n2 ) );
  XOR \ADD_/FAINST[428].FA_/U1  ( .A(a[428]), .B(\ADD_/c[428] ), .Z(
        \ADD_/FAINST[428].FA_/n1 ) );
  XOR \ADD_/FAINST[427].FA_/U5  ( .A(\ADD_/FAINST[427].FA_/n3 ), .B(
        \ADD_/c[427] ), .Z(\ADD_/c[428] ) );
  XOR \ADD_/FAINST[427].FA_/U4  ( .A(\ADD_/FAINST[427].FA_/n1 ), .B(b[427]), 
        .Z(c[427]) );
  AND \ADD_/FAINST[427].FA_/U3  ( .A(\ADD_/FAINST[427].FA_/n1 ), .B(
        \ADD_/FAINST[427].FA_/n2 ), .Z(\ADD_/FAINST[427].FA_/n3 ) );
  XOR \ADD_/FAINST[427].FA_/U2  ( .A(b[427]), .B(\ADD_/c[427] ), .Z(
        \ADD_/FAINST[427].FA_/n2 ) );
  XOR \ADD_/FAINST[427].FA_/U1  ( .A(a[427]), .B(\ADD_/c[427] ), .Z(
        \ADD_/FAINST[427].FA_/n1 ) );
  XOR \ADD_/FAINST[426].FA_/U5  ( .A(\ADD_/FAINST[426].FA_/n3 ), .B(
        \ADD_/c[426] ), .Z(\ADD_/c[427] ) );
  XOR \ADD_/FAINST[426].FA_/U4  ( .A(\ADD_/FAINST[426].FA_/n1 ), .B(b[426]), 
        .Z(c[426]) );
  AND \ADD_/FAINST[426].FA_/U3  ( .A(\ADD_/FAINST[426].FA_/n1 ), .B(
        \ADD_/FAINST[426].FA_/n2 ), .Z(\ADD_/FAINST[426].FA_/n3 ) );
  XOR \ADD_/FAINST[426].FA_/U2  ( .A(b[426]), .B(\ADD_/c[426] ), .Z(
        \ADD_/FAINST[426].FA_/n2 ) );
  XOR \ADD_/FAINST[426].FA_/U1  ( .A(a[426]), .B(\ADD_/c[426] ), .Z(
        \ADD_/FAINST[426].FA_/n1 ) );
  XOR \ADD_/FAINST[425].FA_/U5  ( .A(\ADD_/FAINST[425].FA_/n3 ), .B(
        \ADD_/c[425] ), .Z(\ADD_/c[426] ) );
  XOR \ADD_/FAINST[425].FA_/U4  ( .A(\ADD_/FAINST[425].FA_/n1 ), .B(b[425]), 
        .Z(c[425]) );
  AND \ADD_/FAINST[425].FA_/U3  ( .A(\ADD_/FAINST[425].FA_/n1 ), .B(
        \ADD_/FAINST[425].FA_/n2 ), .Z(\ADD_/FAINST[425].FA_/n3 ) );
  XOR \ADD_/FAINST[425].FA_/U2  ( .A(b[425]), .B(\ADD_/c[425] ), .Z(
        \ADD_/FAINST[425].FA_/n2 ) );
  XOR \ADD_/FAINST[425].FA_/U1  ( .A(a[425]), .B(\ADD_/c[425] ), .Z(
        \ADD_/FAINST[425].FA_/n1 ) );
  XOR \ADD_/FAINST[424].FA_/U5  ( .A(\ADD_/FAINST[424].FA_/n3 ), .B(
        \ADD_/c[424] ), .Z(\ADD_/c[425] ) );
  XOR \ADD_/FAINST[424].FA_/U4  ( .A(\ADD_/FAINST[424].FA_/n1 ), .B(b[424]), 
        .Z(c[424]) );
  AND \ADD_/FAINST[424].FA_/U3  ( .A(\ADD_/FAINST[424].FA_/n1 ), .B(
        \ADD_/FAINST[424].FA_/n2 ), .Z(\ADD_/FAINST[424].FA_/n3 ) );
  XOR \ADD_/FAINST[424].FA_/U2  ( .A(b[424]), .B(\ADD_/c[424] ), .Z(
        \ADD_/FAINST[424].FA_/n2 ) );
  XOR \ADD_/FAINST[424].FA_/U1  ( .A(a[424]), .B(\ADD_/c[424] ), .Z(
        \ADD_/FAINST[424].FA_/n1 ) );
  XOR \ADD_/FAINST[423].FA_/U5  ( .A(\ADD_/FAINST[423].FA_/n3 ), .B(
        \ADD_/c[423] ), .Z(\ADD_/c[424] ) );
  XOR \ADD_/FAINST[423].FA_/U4  ( .A(\ADD_/FAINST[423].FA_/n1 ), .B(b[423]), 
        .Z(c[423]) );
  AND \ADD_/FAINST[423].FA_/U3  ( .A(\ADD_/FAINST[423].FA_/n1 ), .B(
        \ADD_/FAINST[423].FA_/n2 ), .Z(\ADD_/FAINST[423].FA_/n3 ) );
  XOR \ADD_/FAINST[423].FA_/U2  ( .A(b[423]), .B(\ADD_/c[423] ), .Z(
        \ADD_/FAINST[423].FA_/n2 ) );
  XOR \ADD_/FAINST[423].FA_/U1  ( .A(a[423]), .B(\ADD_/c[423] ), .Z(
        \ADD_/FAINST[423].FA_/n1 ) );
  XOR \ADD_/FAINST[422].FA_/U5  ( .A(\ADD_/FAINST[422].FA_/n3 ), .B(
        \ADD_/c[422] ), .Z(\ADD_/c[423] ) );
  XOR \ADD_/FAINST[422].FA_/U4  ( .A(\ADD_/FAINST[422].FA_/n1 ), .B(b[422]), 
        .Z(c[422]) );
  AND \ADD_/FAINST[422].FA_/U3  ( .A(\ADD_/FAINST[422].FA_/n1 ), .B(
        \ADD_/FAINST[422].FA_/n2 ), .Z(\ADD_/FAINST[422].FA_/n3 ) );
  XOR \ADD_/FAINST[422].FA_/U2  ( .A(b[422]), .B(\ADD_/c[422] ), .Z(
        \ADD_/FAINST[422].FA_/n2 ) );
  XOR \ADD_/FAINST[422].FA_/U1  ( .A(a[422]), .B(\ADD_/c[422] ), .Z(
        \ADD_/FAINST[422].FA_/n1 ) );
  XOR \ADD_/FAINST[421].FA_/U5  ( .A(\ADD_/FAINST[421].FA_/n3 ), .B(
        \ADD_/c[421] ), .Z(\ADD_/c[422] ) );
  XOR \ADD_/FAINST[421].FA_/U4  ( .A(\ADD_/FAINST[421].FA_/n1 ), .B(b[421]), 
        .Z(c[421]) );
  AND \ADD_/FAINST[421].FA_/U3  ( .A(\ADD_/FAINST[421].FA_/n1 ), .B(
        \ADD_/FAINST[421].FA_/n2 ), .Z(\ADD_/FAINST[421].FA_/n3 ) );
  XOR \ADD_/FAINST[421].FA_/U2  ( .A(b[421]), .B(\ADD_/c[421] ), .Z(
        \ADD_/FAINST[421].FA_/n2 ) );
  XOR \ADD_/FAINST[421].FA_/U1  ( .A(a[421]), .B(\ADD_/c[421] ), .Z(
        \ADD_/FAINST[421].FA_/n1 ) );
  XOR \ADD_/FAINST[420].FA_/U5  ( .A(\ADD_/FAINST[420].FA_/n3 ), .B(
        \ADD_/c[420] ), .Z(\ADD_/c[421] ) );
  XOR \ADD_/FAINST[420].FA_/U4  ( .A(\ADD_/FAINST[420].FA_/n1 ), .B(b[420]), 
        .Z(c[420]) );
  AND \ADD_/FAINST[420].FA_/U3  ( .A(\ADD_/FAINST[420].FA_/n1 ), .B(
        \ADD_/FAINST[420].FA_/n2 ), .Z(\ADD_/FAINST[420].FA_/n3 ) );
  XOR \ADD_/FAINST[420].FA_/U2  ( .A(b[420]), .B(\ADD_/c[420] ), .Z(
        \ADD_/FAINST[420].FA_/n2 ) );
  XOR \ADD_/FAINST[420].FA_/U1  ( .A(a[420]), .B(\ADD_/c[420] ), .Z(
        \ADD_/FAINST[420].FA_/n1 ) );
  XOR \ADD_/FAINST[419].FA_/U5  ( .A(\ADD_/FAINST[419].FA_/n3 ), .B(
        \ADD_/c[419] ), .Z(\ADD_/c[420] ) );
  XOR \ADD_/FAINST[419].FA_/U4  ( .A(\ADD_/FAINST[419].FA_/n1 ), .B(b[419]), 
        .Z(c[419]) );
  AND \ADD_/FAINST[419].FA_/U3  ( .A(\ADD_/FAINST[419].FA_/n1 ), .B(
        \ADD_/FAINST[419].FA_/n2 ), .Z(\ADD_/FAINST[419].FA_/n3 ) );
  XOR \ADD_/FAINST[419].FA_/U2  ( .A(b[419]), .B(\ADD_/c[419] ), .Z(
        \ADD_/FAINST[419].FA_/n2 ) );
  XOR \ADD_/FAINST[419].FA_/U1  ( .A(a[419]), .B(\ADD_/c[419] ), .Z(
        \ADD_/FAINST[419].FA_/n1 ) );
  XOR \ADD_/FAINST[418].FA_/U5  ( .A(\ADD_/FAINST[418].FA_/n3 ), .B(
        \ADD_/c[418] ), .Z(\ADD_/c[419] ) );
  XOR \ADD_/FAINST[418].FA_/U4  ( .A(\ADD_/FAINST[418].FA_/n1 ), .B(b[418]), 
        .Z(c[418]) );
  AND \ADD_/FAINST[418].FA_/U3  ( .A(\ADD_/FAINST[418].FA_/n1 ), .B(
        \ADD_/FAINST[418].FA_/n2 ), .Z(\ADD_/FAINST[418].FA_/n3 ) );
  XOR \ADD_/FAINST[418].FA_/U2  ( .A(b[418]), .B(\ADD_/c[418] ), .Z(
        \ADD_/FAINST[418].FA_/n2 ) );
  XOR \ADD_/FAINST[418].FA_/U1  ( .A(a[418]), .B(\ADD_/c[418] ), .Z(
        \ADD_/FAINST[418].FA_/n1 ) );
  XOR \ADD_/FAINST[417].FA_/U5  ( .A(\ADD_/FAINST[417].FA_/n3 ), .B(
        \ADD_/c[417] ), .Z(\ADD_/c[418] ) );
  XOR \ADD_/FAINST[417].FA_/U4  ( .A(\ADD_/FAINST[417].FA_/n1 ), .B(b[417]), 
        .Z(c[417]) );
  AND \ADD_/FAINST[417].FA_/U3  ( .A(\ADD_/FAINST[417].FA_/n1 ), .B(
        \ADD_/FAINST[417].FA_/n2 ), .Z(\ADD_/FAINST[417].FA_/n3 ) );
  XOR \ADD_/FAINST[417].FA_/U2  ( .A(b[417]), .B(\ADD_/c[417] ), .Z(
        \ADD_/FAINST[417].FA_/n2 ) );
  XOR \ADD_/FAINST[417].FA_/U1  ( .A(a[417]), .B(\ADD_/c[417] ), .Z(
        \ADD_/FAINST[417].FA_/n1 ) );
  XOR \ADD_/FAINST[416].FA_/U5  ( .A(\ADD_/FAINST[416].FA_/n3 ), .B(
        \ADD_/c[416] ), .Z(\ADD_/c[417] ) );
  XOR \ADD_/FAINST[416].FA_/U4  ( .A(\ADD_/FAINST[416].FA_/n1 ), .B(b[416]), 
        .Z(c[416]) );
  AND \ADD_/FAINST[416].FA_/U3  ( .A(\ADD_/FAINST[416].FA_/n1 ), .B(
        \ADD_/FAINST[416].FA_/n2 ), .Z(\ADD_/FAINST[416].FA_/n3 ) );
  XOR \ADD_/FAINST[416].FA_/U2  ( .A(b[416]), .B(\ADD_/c[416] ), .Z(
        \ADD_/FAINST[416].FA_/n2 ) );
  XOR \ADD_/FAINST[416].FA_/U1  ( .A(a[416]), .B(\ADD_/c[416] ), .Z(
        \ADD_/FAINST[416].FA_/n1 ) );
  XOR \ADD_/FAINST[415].FA_/U5  ( .A(\ADD_/FAINST[415].FA_/n3 ), .B(
        \ADD_/c[415] ), .Z(\ADD_/c[416] ) );
  XOR \ADD_/FAINST[415].FA_/U4  ( .A(\ADD_/FAINST[415].FA_/n1 ), .B(b[415]), 
        .Z(c[415]) );
  AND \ADD_/FAINST[415].FA_/U3  ( .A(\ADD_/FAINST[415].FA_/n1 ), .B(
        \ADD_/FAINST[415].FA_/n2 ), .Z(\ADD_/FAINST[415].FA_/n3 ) );
  XOR \ADD_/FAINST[415].FA_/U2  ( .A(b[415]), .B(\ADD_/c[415] ), .Z(
        \ADD_/FAINST[415].FA_/n2 ) );
  XOR \ADD_/FAINST[415].FA_/U1  ( .A(a[415]), .B(\ADD_/c[415] ), .Z(
        \ADD_/FAINST[415].FA_/n1 ) );
  XOR \ADD_/FAINST[414].FA_/U5  ( .A(\ADD_/FAINST[414].FA_/n3 ), .B(
        \ADD_/c[414] ), .Z(\ADD_/c[415] ) );
  XOR \ADD_/FAINST[414].FA_/U4  ( .A(\ADD_/FAINST[414].FA_/n1 ), .B(b[414]), 
        .Z(c[414]) );
  AND \ADD_/FAINST[414].FA_/U3  ( .A(\ADD_/FAINST[414].FA_/n1 ), .B(
        \ADD_/FAINST[414].FA_/n2 ), .Z(\ADD_/FAINST[414].FA_/n3 ) );
  XOR \ADD_/FAINST[414].FA_/U2  ( .A(b[414]), .B(\ADD_/c[414] ), .Z(
        \ADD_/FAINST[414].FA_/n2 ) );
  XOR \ADD_/FAINST[414].FA_/U1  ( .A(a[414]), .B(\ADD_/c[414] ), .Z(
        \ADD_/FAINST[414].FA_/n1 ) );
  XOR \ADD_/FAINST[413].FA_/U5  ( .A(\ADD_/FAINST[413].FA_/n3 ), .B(
        \ADD_/c[413] ), .Z(\ADD_/c[414] ) );
  XOR \ADD_/FAINST[413].FA_/U4  ( .A(\ADD_/FAINST[413].FA_/n1 ), .B(b[413]), 
        .Z(c[413]) );
  AND \ADD_/FAINST[413].FA_/U3  ( .A(\ADD_/FAINST[413].FA_/n1 ), .B(
        \ADD_/FAINST[413].FA_/n2 ), .Z(\ADD_/FAINST[413].FA_/n3 ) );
  XOR \ADD_/FAINST[413].FA_/U2  ( .A(b[413]), .B(\ADD_/c[413] ), .Z(
        \ADD_/FAINST[413].FA_/n2 ) );
  XOR \ADD_/FAINST[413].FA_/U1  ( .A(a[413]), .B(\ADD_/c[413] ), .Z(
        \ADD_/FAINST[413].FA_/n1 ) );
  XOR \ADD_/FAINST[412].FA_/U5  ( .A(\ADD_/FAINST[412].FA_/n3 ), .B(
        \ADD_/c[412] ), .Z(\ADD_/c[413] ) );
  XOR \ADD_/FAINST[412].FA_/U4  ( .A(\ADD_/FAINST[412].FA_/n1 ), .B(b[412]), 
        .Z(c[412]) );
  AND \ADD_/FAINST[412].FA_/U3  ( .A(\ADD_/FAINST[412].FA_/n1 ), .B(
        \ADD_/FAINST[412].FA_/n2 ), .Z(\ADD_/FAINST[412].FA_/n3 ) );
  XOR \ADD_/FAINST[412].FA_/U2  ( .A(b[412]), .B(\ADD_/c[412] ), .Z(
        \ADD_/FAINST[412].FA_/n2 ) );
  XOR \ADD_/FAINST[412].FA_/U1  ( .A(a[412]), .B(\ADD_/c[412] ), .Z(
        \ADD_/FAINST[412].FA_/n1 ) );
  XOR \ADD_/FAINST[411].FA_/U5  ( .A(\ADD_/FAINST[411].FA_/n3 ), .B(
        \ADD_/c[411] ), .Z(\ADD_/c[412] ) );
  XOR \ADD_/FAINST[411].FA_/U4  ( .A(\ADD_/FAINST[411].FA_/n1 ), .B(b[411]), 
        .Z(c[411]) );
  AND \ADD_/FAINST[411].FA_/U3  ( .A(\ADD_/FAINST[411].FA_/n1 ), .B(
        \ADD_/FAINST[411].FA_/n2 ), .Z(\ADD_/FAINST[411].FA_/n3 ) );
  XOR \ADD_/FAINST[411].FA_/U2  ( .A(b[411]), .B(\ADD_/c[411] ), .Z(
        \ADD_/FAINST[411].FA_/n2 ) );
  XOR \ADD_/FAINST[411].FA_/U1  ( .A(a[411]), .B(\ADD_/c[411] ), .Z(
        \ADD_/FAINST[411].FA_/n1 ) );
  XOR \ADD_/FAINST[410].FA_/U5  ( .A(\ADD_/FAINST[410].FA_/n3 ), .B(
        \ADD_/c[410] ), .Z(\ADD_/c[411] ) );
  XOR \ADD_/FAINST[410].FA_/U4  ( .A(\ADD_/FAINST[410].FA_/n1 ), .B(b[410]), 
        .Z(c[410]) );
  AND \ADD_/FAINST[410].FA_/U3  ( .A(\ADD_/FAINST[410].FA_/n1 ), .B(
        \ADD_/FAINST[410].FA_/n2 ), .Z(\ADD_/FAINST[410].FA_/n3 ) );
  XOR \ADD_/FAINST[410].FA_/U2  ( .A(b[410]), .B(\ADD_/c[410] ), .Z(
        \ADD_/FAINST[410].FA_/n2 ) );
  XOR \ADD_/FAINST[410].FA_/U1  ( .A(a[410]), .B(\ADD_/c[410] ), .Z(
        \ADD_/FAINST[410].FA_/n1 ) );
  XOR \ADD_/FAINST[409].FA_/U5  ( .A(\ADD_/FAINST[409].FA_/n3 ), .B(
        \ADD_/c[409] ), .Z(\ADD_/c[410] ) );
  XOR \ADD_/FAINST[409].FA_/U4  ( .A(\ADD_/FAINST[409].FA_/n1 ), .B(b[409]), 
        .Z(c[409]) );
  AND \ADD_/FAINST[409].FA_/U3  ( .A(\ADD_/FAINST[409].FA_/n1 ), .B(
        \ADD_/FAINST[409].FA_/n2 ), .Z(\ADD_/FAINST[409].FA_/n3 ) );
  XOR \ADD_/FAINST[409].FA_/U2  ( .A(b[409]), .B(\ADD_/c[409] ), .Z(
        \ADD_/FAINST[409].FA_/n2 ) );
  XOR \ADD_/FAINST[409].FA_/U1  ( .A(a[409]), .B(\ADD_/c[409] ), .Z(
        \ADD_/FAINST[409].FA_/n1 ) );
  XOR \ADD_/FAINST[408].FA_/U5  ( .A(\ADD_/FAINST[408].FA_/n3 ), .B(
        \ADD_/c[408] ), .Z(\ADD_/c[409] ) );
  XOR \ADD_/FAINST[408].FA_/U4  ( .A(\ADD_/FAINST[408].FA_/n1 ), .B(b[408]), 
        .Z(c[408]) );
  AND \ADD_/FAINST[408].FA_/U3  ( .A(\ADD_/FAINST[408].FA_/n1 ), .B(
        \ADD_/FAINST[408].FA_/n2 ), .Z(\ADD_/FAINST[408].FA_/n3 ) );
  XOR \ADD_/FAINST[408].FA_/U2  ( .A(b[408]), .B(\ADD_/c[408] ), .Z(
        \ADD_/FAINST[408].FA_/n2 ) );
  XOR \ADD_/FAINST[408].FA_/U1  ( .A(a[408]), .B(\ADD_/c[408] ), .Z(
        \ADD_/FAINST[408].FA_/n1 ) );
  XOR \ADD_/FAINST[407].FA_/U5  ( .A(\ADD_/FAINST[407].FA_/n3 ), .B(
        \ADD_/c[407] ), .Z(\ADD_/c[408] ) );
  XOR \ADD_/FAINST[407].FA_/U4  ( .A(\ADD_/FAINST[407].FA_/n1 ), .B(b[407]), 
        .Z(c[407]) );
  AND \ADD_/FAINST[407].FA_/U3  ( .A(\ADD_/FAINST[407].FA_/n1 ), .B(
        \ADD_/FAINST[407].FA_/n2 ), .Z(\ADD_/FAINST[407].FA_/n3 ) );
  XOR \ADD_/FAINST[407].FA_/U2  ( .A(b[407]), .B(\ADD_/c[407] ), .Z(
        \ADD_/FAINST[407].FA_/n2 ) );
  XOR \ADD_/FAINST[407].FA_/U1  ( .A(a[407]), .B(\ADD_/c[407] ), .Z(
        \ADD_/FAINST[407].FA_/n1 ) );
  XOR \ADD_/FAINST[406].FA_/U5  ( .A(\ADD_/FAINST[406].FA_/n3 ), .B(
        \ADD_/c[406] ), .Z(\ADD_/c[407] ) );
  XOR \ADD_/FAINST[406].FA_/U4  ( .A(\ADD_/FAINST[406].FA_/n1 ), .B(b[406]), 
        .Z(c[406]) );
  AND \ADD_/FAINST[406].FA_/U3  ( .A(\ADD_/FAINST[406].FA_/n1 ), .B(
        \ADD_/FAINST[406].FA_/n2 ), .Z(\ADD_/FAINST[406].FA_/n3 ) );
  XOR \ADD_/FAINST[406].FA_/U2  ( .A(b[406]), .B(\ADD_/c[406] ), .Z(
        \ADD_/FAINST[406].FA_/n2 ) );
  XOR \ADD_/FAINST[406].FA_/U1  ( .A(a[406]), .B(\ADD_/c[406] ), .Z(
        \ADD_/FAINST[406].FA_/n1 ) );
  XOR \ADD_/FAINST[405].FA_/U5  ( .A(\ADD_/FAINST[405].FA_/n3 ), .B(
        \ADD_/c[405] ), .Z(\ADD_/c[406] ) );
  XOR \ADD_/FAINST[405].FA_/U4  ( .A(\ADD_/FAINST[405].FA_/n1 ), .B(b[405]), 
        .Z(c[405]) );
  AND \ADD_/FAINST[405].FA_/U3  ( .A(\ADD_/FAINST[405].FA_/n1 ), .B(
        \ADD_/FAINST[405].FA_/n2 ), .Z(\ADD_/FAINST[405].FA_/n3 ) );
  XOR \ADD_/FAINST[405].FA_/U2  ( .A(b[405]), .B(\ADD_/c[405] ), .Z(
        \ADD_/FAINST[405].FA_/n2 ) );
  XOR \ADD_/FAINST[405].FA_/U1  ( .A(a[405]), .B(\ADD_/c[405] ), .Z(
        \ADD_/FAINST[405].FA_/n1 ) );
  XOR \ADD_/FAINST[404].FA_/U5  ( .A(\ADD_/FAINST[404].FA_/n3 ), .B(
        \ADD_/c[404] ), .Z(\ADD_/c[405] ) );
  XOR \ADD_/FAINST[404].FA_/U4  ( .A(\ADD_/FAINST[404].FA_/n1 ), .B(b[404]), 
        .Z(c[404]) );
  AND \ADD_/FAINST[404].FA_/U3  ( .A(\ADD_/FAINST[404].FA_/n1 ), .B(
        \ADD_/FAINST[404].FA_/n2 ), .Z(\ADD_/FAINST[404].FA_/n3 ) );
  XOR \ADD_/FAINST[404].FA_/U2  ( .A(b[404]), .B(\ADD_/c[404] ), .Z(
        \ADD_/FAINST[404].FA_/n2 ) );
  XOR \ADD_/FAINST[404].FA_/U1  ( .A(a[404]), .B(\ADD_/c[404] ), .Z(
        \ADD_/FAINST[404].FA_/n1 ) );
  XOR \ADD_/FAINST[403].FA_/U5  ( .A(\ADD_/FAINST[403].FA_/n3 ), .B(
        \ADD_/c[403] ), .Z(\ADD_/c[404] ) );
  XOR \ADD_/FAINST[403].FA_/U4  ( .A(\ADD_/FAINST[403].FA_/n1 ), .B(b[403]), 
        .Z(c[403]) );
  AND \ADD_/FAINST[403].FA_/U3  ( .A(\ADD_/FAINST[403].FA_/n1 ), .B(
        \ADD_/FAINST[403].FA_/n2 ), .Z(\ADD_/FAINST[403].FA_/n3 ) );
  XOR \ADD_/FAINST[403].FA_/U2  ( .A(b[403]), .B(\ADD_/c[403] ), .Z(
        \ADD_/FAINST[403].FA_/n2 ) );
  XOR \ADD_/FAINST[403].FA_/U1  ( .A(a[403]), .B(\ADD_/c[403] ), .Z(
        \ADD_/FAINST[403].FA_/n1 ) );
  XOR \ADD_/FAINST[402].FA_/U5  ( .A(\ADD_/FAINST[402].FA_/n3 ), .B(
        \ADD_/c[402] ), .Z(\ADD_/c[403] ) );
  XOR \ADD_/FAINST[402].FA_/U4  ( .A(\ADD_/FAINST[402].FA_/n1 ), .B(b[402]), 
        .Z(c[402]) );
  AND \ADD_/FAINST[402].FA_/U3  ( .A(\ADD_/FAINST[402].FA_/n1 ), .B(
        \ADD_/FAINST[402].FA_/n2 ), .Z(\ADD_/FAINST[402].FA_/n3 ) );
  XOR \ADD_/FAINST[402].FA_/U2  ( .A(b[402]), .B(\ADD_/c[402] ), .Z(
        \ADD_/FAINST[402].FA_/n2 ) );
  XOR \ADD_/FAINST[402].FA_/U1  ( .A(a[402]), .B(\ADD_/c[402] ), .Z(
        \ADD_/FAINST[402].FA_/n1 ) );
  XOR \ADD_/FAINST[401].FA_/U5  ( .A(\ADD_/FAINST[401].FA_/n3 ), .B(
        \ADD_/c[401] ), .Z(\ADD_/c[402] ) );
  XOR \ADD_/FAINST[401].FA_/U4  ( .A(\ADD_/FAINST[401].FA_/n1 ), .B(b[401]), 
        .Z(c[401]) );
  AND \ADD_/FAINST[401].FA_/U3  ( .A(\ADD_/FAINST[401].FA_/n1 ), .B(
        \ADD_/FAINST[401].FA_/n2 ), .Z(\ADD_/FAINST[401].FA_/n3 ) );
  XOR \ADD_/FAINST[401].FA_/U2  ( .A(b[401]), .B(\ADD_/c[401] ), .Z(
        \ADD_/FAINST[401].FA_/n2 ) );
  XOR \ADD_/FAINST[401].FA_/U1  ( .A(a[401]), .B(\ADD_/c[401] ), .Z(
        \ADD_/FAINST[401].FA_/n1 ) );
  XOR \ADD_/FAINST[400].FA_/U5  ( .A(\ADD_/FAINST[400].FA_/n3 ), .B(
        \ADD_/c[400] ), .Z(\ADD_/c[401] ) );
  XOR \ADD_/FAINST[400].FA_/U4  ( .A(\ADD_/FAINST[400].FA_/n1 ), .B(b[400]), 
        .Z(c[400]) );
  AND \ADD_/FAINST[400].FA_/U3  ( .A(\ADD_/FAINST[400].FA_/n1 ), .B(
        \ADD_/FAINST[400].FA_/n2 ), .Z(\ADD_/FAINST[400].FA_/n3 ) );
  XOR \ADD_/FAINST[400].FA_/U2  ( .A(b[400]), .B(\ADD_/c[400] ), .Z(
        \ADD_/FAINST[400].FA_/n2 ) );
  XOR \ADD_/FAINST[400].FA_/U1  ( .A(a[400]), .B(\ADD_/c[400] ), .Z(
        \ADD_/FAINST[400].FA_/n1 ) );
  XOR \ADD_/FAINST[399].FA_/U5  ( .A(\ADD_/FAINST[399].FA_/n3 ), .B(
        \ADD_/c[399] ), .Z(\ADD_/c[400] ) );
  XOR \ADD_/FAINST[399].FA_/U4  ( .A(\ADD_/FAINST[399].FA_/n1 ), .B(b[399]), 
        .Z(c[399]) );
  AND \ADD_/FAINST[399].FA_/U3  ( .A(\ADD_/FAINST[399].FA_/n1 ), .B(
        \ADD_/FAINST[399].FA_/n2 ), .Z(\ADD_/FAINST[399].FA_/n3 ) );
  XOR \ADD_/FAINST[399].FA_/U2  ( .A(b[399]), .B(\ADD_/c[399] ), .Z(
        \ADD_/FAINST[399].FA_/n2 ) );
  XOR \ADD_/FAINST[399].FA_/U1  ( .A(a[399]), .B(\ADD_/c[399] ), .Z(
        \ADD_/FAINST[399].FA_/n1 ) );
  XOR \ADD_/FAINST[398].FA_/U5  ( .A(\ADD_/FAINST[398].FA_/n3 ), .B(
        \ADD_/c[398] ), .Z(\ADD_/c[399] ) );
  XOR \ADD_/FAINST[398].FA_/U4  ( .A(\ADD_/FAINST[398].FA_/n1 ), .B(b[398]), 
        .Z(c[398]) );
  AND \ADD_/FAINST[398].FA_/U3  ( .A(\ADD_/FAINST[398].FA_/n1 ), .B(
        \ADD_/FAINST[398].FA_/n2 ), .Z(\ADD_/FAINST[398].FA_/n3 ) );
  XOR \ADD_/FAINST[398].FA_/U2  ( .A(b[398]), .B(\ADD_/c[398] ), .Z(
        \ADD_/FAINST[398].FA_/n2 ) );
  XOR \ADD_/FAINST[398].FA_/U1  ( .A(a[398]), .B(\ADD_/c[398] ), .Z(
        \ADD_/FAINST[398].FA_/n1 ) );
  XOR \ADD_/FAINST[397].FA_/U5  ( .A(\ADD_/FAINST[397].FA_/n3 ), .B(
        \ADD_/c[397] ), .Z(\ADD_/c[398] ) );
  XOR \ADD_/FAINST[397].FA_/U4  ( .A(\ADD_/FAINST[397].FA_/n1 ), .B(b[397]), 
        .Z(c[397]) );
  AND \ADD_/FAINST[397].FA_/U3  ( .A(\ADD_/FAINST[397].FA_/n1 ), .B(
        \ADD_/FAINST[397].FA_/n2 ), .Z(\ADD_/FAINST[397].FA_/n3 ) );
  XOR \ADD_/FAINST[397].FA_/U2  ( .A(b[397]), .B(\ADD_/c[397] ), .Z(
        \ADD_/FAINST[397].FA_/n2 ) );
  XOR \ADD_/FAINST[397].FA_/U1  ( .A(a[397]), .B(\ADD_/c[397] ), .Z(
        \ADD_/FAINST[397].FA_/n1 ) );
  XOR \ADD_/FAINST[396].FA_/U5  ( .A(\ADD_/FAINST[396].FA_/n3 ), .B(
        \ADD_/c[396] ), .Z(\ADD_/c[397] ) );
  XOR \ADD_/FAINST[396].FA_/U4  ( .A(\ADD_/FAINST[396].FA_/n1 ), .B(b[396]), 
        .Z(c[396]) );
  AND \ADD_/FAINST[396].FA_/U3  ( .A(\ADD_/FAINST[396].FA_/n1 ), .B(
        \ADD_/FAINST[396].FA_/n2 ), .Z(\ADD_/FAINST[396].FA_/n3 ) );
  XOR \ADD_/FAINST[396].FA_/U2  ( .A(b[396]), .B(\ADD_/c[396] ), .Z(
        \ADD_/FAINST[396].FA_/n2 ) );
  XOR \ADD_/FAINST[396].FA_/U1  ( .A(a[396]), .B(\ADD_/c[396] ), .Z(
        \ADD_/FAINST[396].FA_/n1 ) );
  XOR \ADD_/FAINST[395].FA_/U5  ( .A(\ADD_/FAINST[395].FA_/n3 ), .B(
        \ADD_/c[395] ), .Z(\ADD_/c[396] ) );
  XOR \ADD_/FAINST[395].FA_/U4  ( .A(\ADD_/FAINST[395].FA_/n1 ), .B(b[395]), 
        .Z(c[395]) );
  AND \ADD_/FAINST[395].FA_/U3  ( .A(\ADD_/FAINST[395].FA_/n1 ), .B(
        \ADD_/FAINST[395].FA_/n2 ), .Z(\ADD_/FAINST[395].FA_/n3 ) );
  XOR \ADD_/FAINST[395].FA_/U2  ( .A(b[395]), .B(\ADD_/c[395] ), .Z(
        \ADD_/FAINST[395].FA_/n2 ) );
  XOR \ADD_/FAINST[395].FA_/U1  ( .A(a[395]), .B(\ADD_/c[395] ), .Z(
        \ADD_/FAINST[395].FA_/n1 ) );
  XOR \ADD_/FAINST[394].FA_/U5  ( .A(\ADD_/FAINST[394].FA_/n3 ), .B(
        \ADD_/c[394] ), .Z(\ADD_/c[395] ) );
  XOR \ADD_/FAINST[394].FA_/U4  ( .A(\ADD_/FAINST[394].FA_/n1 ), .B(b[394]), 
        .Z(c[394]) );
  AND \ADD_/FAINST[394].FA_/U3  ( .A(\ADD_/FAINST[394].FA_/n1 ), .B(
        \ADD_/FAINST[394].FA_/n2 ), .Z(\ADD_/FAINST[394].FA_/n3 ) );
  XOR \ADD_/FAINST[394].FA_/U2  ( .A(b[394]), .B(\ADD_/c[394] ), .Z(
        \ADD_/FAINST[394].FA_/n2 ) );
  XOR \ADD_/FAINST[394].FA_/U1  ( .A(a[394]), .B(\ADD_/c[394] ), .Z(
        \ADD_/FAINST[394].FA_/n1 ) );
  XOR \ADD_/FAINST[393].FA_/U5  ( .A(\ADD_/FAINST[393].FA_/n3 ), .B(
        \ADD_/c[393] ), .Z(\ADD_/c[394] ) );
  XOR \ADD_/FAINST[393].FA_/U4  ( .A(\ADD_/FAINST[393].FA_/n1 ), .B(b[393]), 
        .Z(c[393]) );
  AND \ADD_/FAINST[393].FA_/U3  ( .A(\ADD_/FAINST[393].FA_/n1 ), .B(
        \ADD_/FAINST[393].FA_/n2 ), .Z(\ADD_/FAINST[393].FA_/n3 ) );
  XOR \ADD_/FAINST[393].FA_/U2  ( .A(b[393]), .B(\ADD_/c[393] ), .Z(
        \ADD_/FAINST[393].FA_/n2 ) );
  XOR \ADD_/FAINST[393].FA_/U1  ( .A(a[393]), .B(\ADD_/c[393] ), .Z(
        \ADD_/FAINST[393].FA_/n1 ) );
  XOR \ADD_/FAINST[392].FA_/U5  ( .A(\ADD_/FAINST[392].FA_/n3 ), .B(
        \ADD_/c[392] ), .Z(\ADD_/c[393] ) );
  XOR \ADD_/FAINST[392].FA_/U4  ( .A(\ADD_/FAINST[392].FA_/n1 ), .B(b[392]), 
        .Z(c[392]) );
  AND \ADD_/FAINST[392].FA_/U3  ( .A(\ADD_/FAINST[392].FA_/n1 ), .B(
        \ADD_/FAINST[392].FA_/n2 ), .Z(\ADD_/FAINST[392].FA_/n3 ) );
  XOR \ADD_/FAINST[392].FA_/U2  ( .A(b[392]), .B(\ADD_/c[392] ), .Z(
        \ADD_/FAINST[392].FA_/n2 ) );
  XOR \ADD_/FAINST[392].FA_/U1  ( .A(a[392]), .B(\ADD_/c[392] ), .Z(
        \ADD_/FAINST[392].FA_/n1 ) );
  XOR \ADD_/FAINST[391].FA_/U5  ( .A(\ADD_/FAINST[391].FA_/n3 ), .B(
        \ADD_/c[391] ), .Z(\ADD_/c[392] ) );
  XOR \ADD_/FAINST[391].FA_/U4  ( .A(\ADD_/FAINST[391].FA_/n1 ), .B(b[391]), 
        .Z(c[391]) );
  AND \ADD_/FAINST[391].FA_/U3  ( .A(\ADD_/FAINST[391].FA_/n1 ), .B(
        \ADD_/FAINST[391].FA_/n2 ), .Z(\ADD_/FAINST[391].FA_/n3 ) );
  XOR \ADD_/FAINST[391].FA_/U2  ( .A(b[391]), .B(\ADD_/c[391] ), .Z(
        \ADD_/FAINST[391].FA_/n2 ) );
  XOR \ADD_/FAINST[391].FA_/U1  ( .A(a[391]), .B(\ADD_/c[391] ), .Z(
        \ADD_/FAINST[391].FA_/n1 ) );
  XOR \ADD_/FAINST[390].FA_/U5  ( .A(\ADD_/FAINST[390].FA_/n3 ), .B(
        \ADD_/c[390] ), .Z(\ADD_/c[391] ) );
  XOR \ADD_/FAINST[390].FA_/U4  ( .A(\ADD_/FAINST[390].FA_/n1 ), .B(b[390]), 
        .Z(c[390]) );
  AND \ADD_/FAINST[390].FA_/U3  ( .A(\ADD_/FAINST[390].FA_/n1 ), .B(
        \ADD_/FAINST[390].FA_/n2 ), .Z(\ADD_/FAINST[390].FA_/n3 ) );
  XOR \ADD_/FAINST[390].FA_/U2  ( .A(b[390]), .B(\ADD_/c[390] ), .Z(
        \ADD_/FAINST[390].FA_/n2 ) );
  XOR \ADD_/FAINST[390].FA_/U1  ( .A(a[390]), .B(\ADD_/c[390] ), .Z(
        \ADD_/FAINST[390].FA_/n1 ) );
  XOR \ADD_/FAINST[389].FA_/U5  ( .A(\ADD_/FAINST[389].FA_/n3 ), .B(
        \ADD_/c[389] ), .Z(\ADD_/c[390] ) );
  XOR \ADD_/FAINST[389].FA_/U4  ( .A(\ADD_/FAINST[389].FA_/n1 ), .B(b[389]), 
        .Z(c[389]) );
  AND \ADD_/FAINST[389].FA_/U3  ( .A(\ADD_/FAINST[389].FA_/n1 ), .B(
        \ADD_/FAINST[389].FA_/n2 ), .Z(\ADD_/FAINST[389].FA_/n3 ) );
  XOR \ADD_/FAINST[389].FA_/U2  ( .A(b[389]), .B(\ADD_/c[389] ), .Z(
        \ADD_/FAINST[389].FA_/n2 ) );
  XOR \ADD_/FAINST[389].FA_/U1  ( .A(a[389]), .B(\ADD_/c[389] ), .Z(
        \ADD_/FAINST[389].FA_/n1 ) );
  XOR \ADD_/FAINST[388].FA_/U5  ( .A(\ADD_/FAINST[388].FA_/n3 ), .B(
        \ADD_/c[388] ), .Z(\ADD_/c[389] ) );
  XOR \ADD_/FAINST[388].FA_/U4  ( .A(\ADD_/FAINST[388].FA_/n1 ), .B(b[388]), 
        .Z(c[388]) );
  AND \ADD_/FAINST[388].FA_/U3  ( .A(\ADD_/FAINST[388].FA_/n1 ), .B(
        \ADD_/FAINST[388].FA_/n2 ), .Z(\ADD_/FAINST[388].FA_/n3 ) );
  XOR \ADD_/FAINST[388].FA_/U2  ( .A(b[388]), .B(\ADD_/c[388] ), .Z(
        \ADD_/FAINST[388].FA_/n2 ) );
  XOR \ADD_/FAINST[388].FA_/U1  ( .A(a[388]), .B(\ADD_/c[388] ), .Z(
        \ADD_/FAINST[388].FA_/n1 ) );
  XOR \ADD_/FAINST[387].FA_/U5  ( .A(\ADD_/FAINST[387].FA_/n3 ), .B(
        \ADD_/c[387] ), .Z(\ADD_/c[388] ) );
  XOR \ADD_/FAINST[387].FA_/U4  ( .A(\ADD_/FAINST[387].FA_/n1 ), .B(b[387]), 
        .Z(c[387]) );
  AND \ADD_/FAINST[387].FA_/U3  ( .A(\ADD_/FAINST[387].FA_/n1 ), .B(
        \ADD_/FAINST[387].FA_/n2 ), .Z(\ADD_/FAINST[387].FA_/n3 ) );
  XOR \ADD_/FAINST[387].FA_/U2  ( .A(b[387]), .B(\ADD_/c[387] ), .Z(
        \ADD_/FAINST[387].FA_/n2 ) );
  XOR \ADD_/FAINST[387].FA_/U1  ( .A(a[387]), .B(\ADD_/c[387] ), .Z(
        \ADD_/FAINST[387].FA_/n1 ) );
  XOR \ADD_/FAINST[386].FA_/U5  ( .A(\ADD_/FAINST[386].FA_/n3 ), .B(
        \ADD_/c[386] ), .Z(\ADD_/c[387] ) );
  XOR \ADD_/FAINST[386].FA_/U4  ( .A(\ADD_/FAINST[386].FA_/n1 ), .B(b[386]), 
        .Z(c[386]) );
  AND \ADD_/FAINST[386].FA_/U3  ( .A(\ADD_/FAINST[386].FA_/n1 ), .B(
        \ADD_/FAINST[386].FA_/n2 ), .Z(\ADD_/FAINST[386].FA_/n3 ) );
  XOR \ADD_/FAINST[386].FA_/U2  ( .A(b[386]), .B(\ADD_/c[386] ), .Z(
        \ADD_/FAINST[386].FA_/n2 ) );
  XOR \ADD_/FAINST[386].FA_/U1  ( .A(a[386]), .B(\ADD_/c[386] ), .Z(
        \ADD_/FAINST[386].FA_/n1 ) );
  XOR \ADD_/FAINST[385].FA_/U5  ( .A(\ADD_/FAINST[385].FA_/n3 ), .B(
        \ADD_/c[385] ), .Z(\ADD_/c[386] ) );
  XOR \ADD_/FAINST[385].FA_/U4  ( .A(\ADD_/FAINST[385].FA_/n1 ), .B(b[385]), 
        .Z(c[385]) );
  AND \ADD_/FAINST[385].FA_/U3  ( .A(\ADD_/FAINST[385].FA_/n1 ), .B(
        \ADD_/FAINST[385].FA_/n2 ), .Z(\ADD_/FAINST[385].FA_/n3 ) );
  XOR \ADD_/FAINST[385].FA_/U2  ( .A(b[385]), .B(\ADD_/c[385] ), .Z(
        \ADD_/FAINST[385].FA_/n2 ) );
  XOR \ADD_/FAINST[385].FA_/U1  ( .A(a[385]), .B(\ADD_/c[385] ), .Z(
        \ADD_/FAINST[385].FA_/n1 ) );
  XOR \ADD_/FAINST[384].FA_/U5  ( .A(\ADD_/FAINST[384].FA_/n3 ), .B(
        \ADD_/c[384] ), .Z(\ADD_/c[385] ) );
  XOR \ADD_/FAINST[384].FA_/U4  ( .A(\ADD_/FAINST[384].FA_/n1 ), .B(b[384]), 
        .Z(c[384]) );
  AND \ADD_/FAINST[384].FA_/U3  ( .A(\ADD_/FAINST[384].FA_/n1 ), .B(
        \ADD_/FAINST[384].FA_/n2 ), .Z(\ADD_/FAINST[384].FA_/n3 ) );
  XOR \ADD_/FAINST[384].FA_/U2  ( .A(b[384]), .B(\ADD_/c[384] ), .Z(
        \ADD_/FAINST[384].FA_/n2 ) );
  XOR \ADD_/FAINST[384].FA_/U1  ( .A(a[384]), .B(\ADD_/c[384] ), .Z(
        \ADD_/FAINST[384].FA_/n1 ) );
  XOR \ADD_/FAINST[383].FA_/U5  ( .A(\ADD_/FAINST[383].FA_/n3 ), .B(
        \ADD_/c[383] ), .Z(\ADD_/c[384] ) );
  XOR \ADD_/FAINST[383].FA_/U4  ( .A(\ADD_/FAINST[383].FA_/n1 ), .B(b[383]), 
        .Z(c[383]) );
  AND \ADD_/FAINST[383].FA_/U3  ( .A(\ADD_/FAINST[383].FA_/n1 ), .B(
        \ADD_/FAINST[383].FA_/n2 ), .Z(\ADD_/FAINST[383].FA_/n3 ) );
  XOR \ADD_/FAINST[383].FA_/U2  ( .A(b[383]), .B(\ADD_/c[383] ), .Z(
        \ADD_/FAINST[383].FA_/n2 ) );
  XOR \ADD_/FAINST[383].FA_/U1  ( .A(a[383]), .B(\ADD_/c[383] ), .Z(
        \ADD_/FAINST[383].FA_/n1 ) );
  XOR \ADD_/FAINST[382].FA_/U5  ( .A(\ADD_/FAINST[382].FA_/n3 ), .B(
        \ADD_/c[382] ), .Z(\ADD_/c[383] ) );
  XOR \ADD_/FAINST[382].FA_/U4  ( .A(\ADD_/FAINST[382].FA_/n1 ), .B(b[382]), 
        .Z(c[382]) );
  AND \ADD_/FAINST[382].FA_/U3  ( .A(\ADD_/FAINST[382].FA_/n1 ), .B(
        \ADD_/FAINST[382].FA_/n2 ), .Z(\ADD_/FAINST[382].FA_/n3 ) );
  XOR \ADD_/FAINST[382].FA_/U2  ( .A(b[382]), .B(\ADD_/c[382] ), .Z(
        \ADD_/FAINST[382].FA_/n2 ) );
  XOR \ADD_/FAINST[382].FA_/U1  ( .A(a[382]), .B(\ADD_/c[382] ), .Z(
        \ADD_/FAINST[382].FA_/n1 ) );
  XOR \ADD_/FAINST[381].FA_/U5  ( .A(\ADD_/FAINST[381].FA_/n3 ), .B(
        \ADD_/c[381] ), .Z(\ADD_/c[382] ) );
  XOR \ADD_/FAINST[381].FA_/U4  ( .A(\ADD_/FAINST[381].FA_/n1 ), .B(b[381]), 
        .Z(c[381]) );
  AND \ADD_/FAINST[381].FA_/U3  ( .A(\ADD_/FAINST[381].FA_/n1 ), .B(
        \ADD_/FAINST[381].FA_/n2 ), .Z(\ADD_/FAINST[381].FA_/n3 ) );
  XOR \ADD_/FAINST[381].FA_/U2  ( .A(b[381]), .B(\ADD_/c[381] ), .Z(
        \ADD_/FAINST[381].FA_/n2 ) );
  XOR \ADD_/FAINST[381].FA_/U1  ( .A(a[381]), .B(\ADD_/c[381] ), .Z(
        \ADD_/FAINST[381].FA_/n1 ) );
  XOR \ADD_/FAINST[380].FA_/U5  ( .A(\ADD_/FAINST[380].FA_/n3 ), .B(
        \ADD_/c[380] ), .Z(\ADD_/c[381] ) );
  XOR \ADD_/FAINST[380].FA_/U4  ( .A(\ADD_/FAINST[380].FA_/n1 ), .B(b[380]), 
        .Z(c[380]) );
  AND \ADD_/FAINST[380].FA_/U3  ( .A(\ADD_/FAINST[380].FA_/n1 ), .B(
        \ADD_/FAINST[380].FA_/n2 ), .Z(\ADD_/FAINST[380].FA_/n3 ) );
  XOR \ADD_/FAINST[380].FA_/U2  ( .A(b[380]), .B(\ADD_/c[380] ), .Z(
        \ADD_/FAINST[380].FA_/n2 ) );
  XOR \ADD_/FAINST[380].FA_/U1  ( .A(a[380]), .B(\ADD_/c[380] ), .Z(
        \ADD_/FAINST[380].FA_/n1 ) );
  XOR \ADD_/FAINST[379].FA_/U5  ( .A(\ADD_/FAINST[379].FA_/n3 ), .B(
        \ADD_/c[379] ), .Z(\ADD_/c[380] ) );
  XOR \ADD_/FAINST[379].FA_/U4  ( .A(\ADD_/FAINST[379].FA_/n1 ), .B(b[379]), 
        .Z(c[379]) );
  AND \ADD_/FAINST[379].FA_/U3  ( .A(\ADD_/FAINST[379].FA_/n1 ), .B(
        \ADD_/FAINST[379].FA_/n2 ), .Z(\ADD_/FAINST[379].FA_/n3 ) );
  XOR \ADD_/FAINST[379].FA_/U2  ( .A(b[379]), .B(\ADD_/c[379] ), .Z(
        \ADD_/FAINST[379].FA_/n2 ) );
  XOR \ADD_/FAINST[379].FA_/U1  ( .A(a[379]), .B(\ADD_/c[379] ), .Z(
        \ADD_/FAINST[379].FA_/n1 ) );
  XOR \ADD_/FAINST[378].FA_/U5  ( .A(\ADD_/FAINST[378].FA_/n3 ), .B(
        \ADD_/c[378] ), .Z(\ADD_/c[379] ) );
  XOR \ADD_/FAINST[378].FA_/U4  ( .A(\ADD_/FAINST[378].FA_/n1 ), .B(b[378]), 
        .Z(c[378]) );
  AND \ADD_/FAINST[378].FA_/U3  ( .A(\ADD_/FAINST[378].FA_/n1 ), .B(
        \ADD_/FAINST[378].FA_/n2 ), .Z(\ADD_/FAINST[378].FA_/n3 ) );
  XOR \ADD_/FAINST[378].FA_/U2  ( .A(b[378]), .B(\ADD_/c[378] ), .Z(
        \ADD_/FAINST[378].FA_/n2 ) );
  XOR \ADD_/FAINST[378].FA_/U1  ( .A(a[378]), .B(\ADD_/c[378] ), .Z(
        \ADD_/FAINST[378].FA_/n1 ) );
  XOR \ADD_/FAINST[377].FA_/U5  ( .A(\ADD_/FAINST[377].FA_/n3 ), .B(
        \ADD_/c[377] ), .Z(\ADD_/c[378] ) );
  XOR \ADD_/FAINST[377].FA_/U4  ( .A(\ADD_/FAINST[377].FA_/n1 ), .B(b[377]), 
        .Z(c[377]) );
  AND \ADD_/FAINST[377].FA_/U3  ( .A(\ADD_/FAINST[377].FA_/n1 ), .B(
        \ADD_/FAINST[377].FA_/n2 ), .Z(\ADD_/FAINST[377].FA_/n3 ) );
  XOR \ADD_/FAINST[377].FA_/U2  ( .A(b[377]), .B(\ADD_/c[377] ), .Z(
        \ADD_/FAINST[377].FA_/n2 ) );
  XOR \ADD_/FAINST[377].FA_/U1  ( .A(a[377]), .B(\ADD_/c[377] ), .Z(
        \ADD_/FAINST[377].FA_/n1 ) );
  XOR \ADD_/FAINST[376].FA_/U5  ( .A(\ADD_/FAINST[376].FA_/n3 ), .B(
        \ADD_/c[376] ), .Z(\ADD_/c[377] ) );
  XOR \ADD_/FAINST[376].FA_/U4  ( .A(\ADD_/FAINST[376].FA_/n1 ), .B(b[376]), 
        .Z(c[376]) );
  AND \ADD_/FAINST[376].FA_/U3  ( .A(\ADD_/FAINST[376].FA_/n1 ), .B(
        \ADD_/FAINST[376].FA_/n2 ), .Z(\ADD_/FAINST[376].FA_/n3 ) );
  XOR \ADD_/FAINST[376].FA_/U2  ( .A(b[376]), .B(\ADD_/c[376] ), .Z(
        \ADD_/FAINST[376].FA_/n2 ) );
  XOR \ADD_/FAINST[376].FA_/U1  ( .A(a[376]), .B(\ADD_/c[376] ), .Z(
        \ADD_/FAINST[376].FA_/n1 ) );
  XOR \ADD_/FAINST[375].FA_/U5  ( .A(\ADD_/FAINST[375].FA_/n3 ), .B(
        \ADD_/c[375] ), .Z(\ADD_/c[376] ) );
  XOR \ADD_/FAINST[375].FA_/U4  ( .A(\ADD_/FAINST[375].FA_/n1 ), .B(b[375]), 
        .Z(c[375]) );
  AND \ADD_/FAINST[375].FA_/U3  ( .A(\ADD_/FAINST[375].FA_/n1 ), .B(
        \ADD_/FAINST[375].FA_/n2 ), .Z(\ADD_/FAINST[375].FA_/n3 ) );
  XOR \ADD_/FAINST[375].FA_/U2  ( .A(b[375]), .B(\ADD_/c[375] ), .Z(
        \ADD_/FAINST[375].FA_/n2 ) );
  XOR \ADD_/FAINST[375].FA_/U1  ( .A(a[375]), .B(\ADD_/c[375] ), .Z(
        \ADD_/FAINST[375].FA_/n1 ) );
  XOR \ADD_/FAINST[374].FA_/U5  ( .A(\ADD_/FAINST[374].FA_/n3 ), .B(
        \ADD_/c[374] ), .Z(\ADD_/c[375] ) );
  XOR \ADD_/FAINST[374].FA_/U4  ( .A(\ADD_/FAINST[374].FA_/n1 ), .B(b[374]), 
        .Z(c[374]) );
  AND \ADD_/FAINST[374].FA_/U3  ( .A(\ADD_/FAINST[374].FA_/n1 ), .B(
        \ADD_/FAINST[374].FA_/n2 ), .Z(\ADD_/FAINST[374].FA_/n3 ) );
  XOR \ADD_/FAINST[374].FA_/U2  ( .A(b[374]), .B(\ADD_/c[374] ), .Z(
        \ADD_/FAINST[374].FA_/n2 ) );
  XOR \ADD_/FAINST[374].FA_/U1  ( .A(a[374]), .B(\ADD_/c[374] ), .Z(
        \ADD_/FAINST[374].FA_/n1 ) );
  XOR \ADD_/FAINST[373].FA_/U5  ( .A(\ADD_/FAINST[373].FA_/n3 ), .B(
        \ADD_/c[373] ), .Z(\ADD_/c[374] ) );
  XOR \ADD_/FAINST[373].FA_/U4  ( .A(\ADD_/FAINST[373].FA_/n1 ), .B(b[373]), 
        .Z(c[373]) );
  AND \ADD_/FAINST[373].FA_/U3  ( .A(\ADD_/FAINST[373].FA_/n1 ), .B(
        \ADD_/FAINST[373].FA_/n2 ), .Z(\ADD_/FAINST[373].FA_/n3 ) );
  XOR \ADD_/FAINST[373].FA_/U2  ( .A(b[373]), .B(\ADD_/c[373] ), .Z(
        \ADD_/FAINST[373].FA_/n2 ) );
  XOR \ADD_/FAINST[373].FA_/U1  ( .A(a[373]), .B(\ADD_/c[373] ), .Z(
        \ADD_/FAINST[373].FA_/n1 ) );
  XOR \ADD_/FAINST[372].FA_/U5  ( .A(\ADD_/FAINST[372].FA_/n3 ), .B(
        \ADD_/c[372] ), .Z(\ADD_/c[373] ) );
  XOR \ADD_/FAINST[372].FA_/U4  ( .A(\ADD_/FAINST[372].FA_/n1 ), .B(b[372]), 
        .Z(c[372]) );
  AND \ADD_/FAINST[372].FA_/U3  ( .A(\ADD_/FAINST[372].FA_/n1 ), .B(
        \ADD_/FAINST[372].FA_/n2 ), .Z(\ADD_/FAINST[372].FA_/n3 ) );
  XOR \ADD_/FAINST[372].FA_/U2  ( .A(b[372]), .B(\ADD_/c[372] ), .Z(
        \ADD_/FAINST[372].FA_/n2 ) );
  XOR \ADD_/FAINST[372].FA_/U1  ( .A(a[372]), .B(\ADD_/c[372] ), .Z(
        \ADD_/FAINST[372].FA_/n1 ) );
  XOR \ADD_/FAINST[371].FA_/U5  ( .A(\ADD_/FAINST[371].FA_/n3 ), .B(
        \ADD_/c[371] ), .Z(\ADD_/c[372] ) );
  XOR \ADD_/FAINST[371].FA_/U4  ( .A(\ADD_/FAINST[371].FA_/n1 ), .B(b[371]), 
        .Z(c[371]) );
  AND \ADD_/FAINST[371].FA_/U3  ( .A(\ADD_/FAINST[371].FA_/n1 ), .B(
        \ADD_/FAINST[371].FA_/n2 ), .Z(\ADD_/FAINST[371].FA_/n3 ) );
  XOR \ADD_/FAINST[371].FA_/U2  ( .A(b[371]), .B(\ADD_/c[371] ), .Z(
        \ADD_/FAINST[371].FA_/n2 ) );
  XOR \ADD_/FAINST[371].FA_/U1  ( .A(a[371]), .B(\ADD_/c[371] ), .Z(
        \ADD_/FAINST[371].FA_/n1 ) );
  XOR \ADD_/FAINST[370].FA_/U5  ( .A(\ADD_/FAINST[370].FA_/n3 ), .B(
        \ADD_/c[370] ), .Z(\ADD_/c[371] ) );
  XOR \ADD_/FAINST[370].FA_/U4  ( .A(\ADD_/FAINST[370].FA_/n1 ), .B(b[370]), 
        .Z(c[370]) );
  AND \ADD_/FAINST[370].FA_/U3  ( .A(\ADD_/FAINST[370].FA_/n1 ), .B(
        \ADD_/FAINST[370].FA_/n2 ), .Z(\ADD_/FAINST[370].FA_/n3 ) );
  XOR \ADD_/FAINST[370].FA_/U2  ( .A(b[370]), .B(\ADD_/c[370] ), .Z(
        \ADD_/FAINST[370].FA_/n2 ) );
  XOR \ADD_/FAINST[370].FA_/U1  ( .A(a[370]), .B(\ADD_/c[370] ), .Z(
        \ADD_/FAINST[370].FA_/n1 ) );
  XOR \ADD_/FAINST[369].FA_/U5  ( .A(\ADD_/FAINST[369].FA_/n3 ), .B(
        \ADD_/c[369] ), .Z(\ADD_/c[370] ) );
  XOR \ADD_/FAINST[369].FA_/U4  ( .A(\ADD_/FAINST[369].FA_/n1 ), .B(b[369]), 
        .Z(c[369]) );
  AND \ADD_/FAINST[369].FA_/U3  ( .A(\ADD_/FAINST[369].FA_/n1 ), .B(
        \ADD_/FAINST[369].FA_/n2 ), .Z(\ADD_/FAINST[369].FA_/n3 ) );
  XOR \ADD_/FAINST[369].FA_/U2  ( .A(b[369]), .B(\ADD_/c[369] ), .Z(
        \ADD_/FAINST[369].FA_/n2 ) );
  XOR \ADD_/FAINST[369].FA_/U1  ( .A(a[369]), .B(\ADD_/c[369] ), .Z(
        \ADD_/FAINST[369].FA_/n1 ) );
  XOR \ADD_/FAINST[368].FA_/U5  ( .A(\ADD_/FAINST[368].FA_/n3 ), .B(
        \ADD_/c[368] ), .Z(\ADD_/c[369] ) );
  XOR \ADD_/FAINST[368].FA_/U4  ( .A(\ADD_/FAINST[368].FA_/n1 ), .B(b[368]), 
        .Z(c[368]) );
  AND \ADD_/FAINST[368].FA_/U3  ( .A(\ADD_/FAINST[368].FA_/n1 ), .B(
        \ADD_/FAINST[368].FA_/n2 ), .Z(\ADD_/FAINST[368].FA_/n3 ) );
  XOR \ADD_/FAINST[368].FA_/U2  ( .A(b[368]), .B(\ADD_/c[368] ), .Z(
        \ADD_/FAINST[368].FA_/n2 ) );
  XOR \ADD_/FAINST[368].FA_/U1  ( .A(a[368]), .B(\ADD_/c[368] ), .Z(
        \ADD_/FAINST[368].FA_/n1 ) );
  XOR \ADD_/FAINST[367].FA_/U5  ( .A(\ADD_/FAINST[367].FA_/n3 ), .B(
        \ADD_/c[367] ), .Z(\ADD_/c[368] ) );
  XOR \ADD_/FAINST[367].FA_/U4  ( .A(\ADD_/FAINST[367].FA_/n1 ), .B(b[367]), 
        .Z(c[367]) );
  AND \ADD_/FAINST[367].FA_/U3  ( .A(\ADD_/FAINST[367].FA_/n1 ), .B(
        \ADD_/FAINST[367].FA_/n2 ), .Z(\ADD_/FAINST[367].FA_/n3 ) );
  XOR \ADD_/FAINST[367].FA_/U2  ( .A(b[367]), .B(\ADD_/c[367] ), .Z(
        \ADD_/FAINST[367].FA_/n2 ) );
  XOR \ADD_/FAINST[367].FA_/U1  ( .A(a[367]), .B(\ADD_/c[367] ), .Z(
        \ADD_/FAINST[367].FA_/n1 ) );
  XOR \ADD_/FAINST[366].FA_/U5  ( .A(\ADD_/FAINST[366].FA_/n3 ), .B(
        \ADD_/c[366] ), .Z(\ADD_/c[367] ) );
  XOR \ADD_/FAINST[366].FA_/U4  ( .A(\ADD_/FAINST[366].FA_/n1 ), .B(b[366]), 
        .Z(c[366]) );
  AND \ADD_/FAINST[366].FA_/U3  ( .A(\ADD_/FAINST[366].FA_/n1 ), .B(
        \ADD_/FAINST[366].FA_/n2 ), .Z(\ADD_/FAINST[366].FA_/n3 ) );
  XOR \ADD_/FAINST[366].FA_/U2  ( .A(b[366]), .B(\ADD_/c[366] ), .Z(
        \ADD_/FAINST[366].FA_/n2 ) );
  XOR \ADD_/FAINST[366].FA_/U1  ( .A(a[366]), .B(\ADD_/c[366] ), .Z(
        \ADD_/FAINST[366].FA_/n1 ) );
  XOR \ADD_/FAINST[365].FA_/U5  ( .A(\ADD_/FAINST[365].FA_/n3 ), .B(
        \ADD_/c[365] ), .Z(\ADD_/c[366] ) );
  XOR \ADD_/FAINST[365].FA_/U4  ( .A(\ADD_/FAINST[365].FA_/n1 ), .B(b[365]), 
        .Z(c[365]) );
  AND \ADD_/FAINST[365].FA_/U3  ( .A(\ADD_/FAINST[365].FA_/n1 ), .B(
        \ADD_/FAINST[365].FA_/n2 ), .Z(\ADD_/FAINST[365].FA_/n3 ) );
  XOR \ADD_/FAINST[365].FA_/U2  ( .A(b[365]), .B(\ADD_/c[365] ), .Z(
        \ADD_/FAINST[365].FA_/n2 ) );
  XOR \ADD_/FAINST[365].FA_/U1  ( .A(a[365]), .B(\ADD_/c[365] ), .Z(
        \ADD_/FAINST[365].FA_/n1 ) );
  XOR \ADD_/FAINST[364].FA_/U5  ( .A(\ADD_/FAINST[364].FA_/n3 ), .B(
        \ADD_/c[364] ), .Z(\ADD_/c[365] ) );
  XOR \ADD_/FAINST[364].FA_/U4  ( .A(\ADD_/FAINST[364].FA_/n1 ), .B(b[364]), 
        .Z(c[364]) );
  AND \ADD_/FAINST[364].FA_/U3  ( .A(\ADD_/FAINST[364].FA_/n1 ), .B(
        \ADD_/FAINST[364].FA_/n2 ), .Z(\ADD_/FAINST[364].FA_/n3 ) );
  XOR \ADD_/FAINST[364].FA_/U2  ( .A(b[364]), .B(\ADD_/c[364] ), .Z(
        \ADD_/FAINST[364].FA_/n2 ) );
  XOR \ADD_/FAINST[364].FA_/U1  ( .A(a[364]), .B(\ADD_/c[364] ), .Z(
        \ADD_/FAINST[364].FA_/n1 ) );
  XOR \ADD_/FAINST[363].FA_/U5  ( .A(\ADD_/FAINST[363].FA_/n3 ), .B(
        \ADD_/c[363] ), .Z(\ADD_/c[364] ) );
  XOR \ADD_/FAINST[363].FA_/U4  ( .A(\ADD_/FAINST[363].FA_/n1 ), .B(b[363]), 
        .Z(c[363]) );
  AND \ADD_/FAINST[363].FA_/U3  ( .A(\ADD_/FAINST[363].FA_/n1 ), .B(
        \ADD_/FAINST[363].FA_/n2 ), .Z(\ADD_/FAINST[363].FA_/n3 ) );
  XOR \ADD_/FAINST[363].FA_/U2  ( .A(b[363]), .B(\ADD_/c[363] ), .Z(
        \ADD_/FAINST[363].FA_/n2 ) );
  XOR \ADD_/FAINST[363].FA_/U1  ( .A(a[363]), .B(\ADD_/c[363] ), .Z(
        \ADD_/FAINST[363].FA_/n1 ) );
  XOR \ADD_/FAINST[362].FA_/U5  ( .A(\ADD_/FAINST[362].FA_/n3 ), .B(
        \ADD_/c[362] ), .Z(\ADD_/c[363] ) );
  XOR \ADD_/FAINST[362].FA_/U4  ( .A(\ADD_/FAINST[362].FA_/n1 ), .B(b[362]), 
        .Z(c[362]) );
  AND \ADD_/FAINST[362].FA_/U3  ( .A(\ADD_/FAINST[362].FA_/n1 ), .B(
        \ADD_/FAINST[362].FA_/n2 ), .Z(\ADD_/FAINST[362].FA_/n3 ) );
  XOR \ADD_/FAINST[362].FA_/U2  ( .A(b[362]), .B(\ADD_/c[362] ), .Z(
        \ADD_/FAINST[362].FA_/n2 ) );
  XOR \ADD_/FAINST[362].FA_/U1  ( .A(a[362]), .B(\ADD_/c[362] ), .Z(
        \ADD_/FAINST[362].FA_/n1 ) );
  XOR \ADD_/FAINST[361].FA_/U5  ( .A(\ADD_/FAINST[361].FA_/n3 ), .B(
        \ADD_/c[361] ), .Z(\ADD_/c[362] ) );
  XOR \ADD_/FAINST[361].FA_/U4  ( .A(\ADD_/FAINST[361].FA_/n1 ), .B(b[361]), 
        .Z(c[361]) );
  AND \ADD_/FAINST[361].FA_/U3  ( .A(\ADD_/FAINST[361].FA_/n1 ), .B(
        \ADD_/FAINST[361].FA_/n2 ), .Z(\ADD_/FAINST[361].FA_/n3 ) );
  XOR \ADD_/FAINST[361].FA_/U2  ( .A(b[361]), .B(\ADD_/c[361] ), .Z(
        \ADD_/FAINST[361].FA_/n2 ) );
  XOR \ADD_/FAINST[361].FA_/U1  ( .A(a[361]), .B(\ADD_/c[361] ), .Z(
        \ADD_/FAINST[361].FA_/n1 ) );
  XOR \ADD_/FAINST[360].FA_/U5  ( .A(\ADD_/FAINST[360].FA_/n3 ), .B(
        \ADD_/c[360] ), .Z(\ADD_/c[361] ) );
  XOR \ADD_/FAINST[360].FA_/U4  ( .A(\ADD_/FAINST[360].FA_/n1 ), .B(b[360]), 
        .Z(c[360]) );
  AND \ADD_/FAINST[360].FA_/U3  ( .A(\ADD_/FAINST[360].FA_/n1 ), .B(
        \ADD_/FAINST[360].FA_/n2 ), .Z(\ADD_/FAINST[360].FA_/n3 ) );
  XOR \ADD_/FAINST[360].FA_/U2  ( .A(b[360]), .B(\ADD_/c[360] ), .Z(
        \ADD_/FAINST[360].FA_/n2 ) );
  XOR \ADD_/FAINST[360].FA_/U1  ( .A(a[360]), .B(\ADD_/c[360] ), .Z(
        \ADD_/FAINST[360].FA_/n1 ) );
  XOR \ADD_/FAINST[359].FA_/U5  ( .A(\ADD_/FAINST[359].FA_/n3 ), .B(
        \ADD_/c[359] ), .Z(\ADD_/c[360] ) );
  XOR \ADD_/FAINST[359].FA_/U4  ( .A(\ADD_/FAINST[359].FA_/n1 ), .B(b[359]), 
        .Z(c[359]) );
  AND \ADD_/FAINST[359].FA_/U3  ( .A(\ADD_/FAINST[359].FA_/n1 ), .B(
        \ADD_/FAINST[359].FA_/n2 ), .Z(\ADD_/FAINST[359].FA_/n3 ) );
  XOR \ADD_/FAINST[359].FA_/U2  ( .A(b[359]), .B(\ADD_/c[359] ), .Z(
        \ADD_/FAINST[359].FA_/n2 ) );
  XOR \ADD_/FAINST[359].FA_/U1  ( .A(a[359]), .B(\ADD_/c[359] ), .Z(
        \ADD_/FAINST[359].FA_/n1 ) );
  XOR \ADD_/FAINST[358].FA_/U5  ( .A(\ADD_/FAINST[358].FA_/n3 ), .B(
        \ADD_/c[358] ), .Z(\ADD_/c[359] ) );
  XOR \ADD_/FAINST[358].FA_/U4  ( .A(\ADD_/FAINST[358].FA_/n1 ), .B(b[358]), 
        .Z(c[358]) );
  AND \ADD_/FAINST[358].FA_/U3  ( .A(\ADD_/FAINST[358].FA_/n1 ), .B(
        \ADD_/FAINST[358].FA_/n2 ), .Z(\ADD_/FAINST[358].FA_/n3 ) );
  XOR \ADD_/FAINST[358].FA_/U2  ( .A(b[358]), .B(\ADD_/c[358] ), .Z(
        \ADD_/FAINST[358].FA_/n2 ) );
  XOR \ADD_/FAINST[358].FA_/U1  ( .A(a[358]), .B(\ADD_/c[358] ), .Z(
        \ADD_/FAINST[358].FA_/n1 ) );
  XOR \ADD_/FAINST[357].FA_/U5  ( .A(\ADD_/FAINST[357].FA_/n3 ), .B(
        \ADD_/c[357] ), .Z(\ADD_/c[358] ) );
  XOR \ADD_/FAINST[357].FA_/U4  ( .A(\ADD_/FAINST[357].FA_/n1 ), .B(b[357]), 
        .Z(c[357]) );
  AND \ADD_/FAINST[357].FA_/U3  ( .A(\ADD_/FAINST[357].FA_/n1 ), .B(
        \ADD_/FAINST[357].FA_/n2 ), .Z(\ADD_/FAINST[357].FA_/n3 ) );
  XOR \ADD_/FAINST[357].FA_/U2  ( .A(b[357]), .B(\ADD_/c[357] ), .Z(
        \ADD_/FAINST[357].FA_/n2 ) );
  XOR \ADD_/FAINST[357].FA_/U1  ( .A(a[357]), .B(\ADD_/c[357] ), .Z(
        \ADD_/FAINST[357].FA_/n1 ) );
  XOR \ADD_/FAINST[356].FA_/U5  ( .A(\ADD_/FAINST[356].FA_/n3 ), .B(
        \ADD_/c[356] ), .Z(\ADD_/c[357] ) );
  XOR \ADD_/FAINST[356].FA_/U4  ( .A(\ADD_/FAINST[356].FA_/n1 ), .B(b[356]), 
        .Z(c[356]) );
  AND \ADD_/FAINST[356].FA_/U3  ( .A(\ADD_/FAINST[356].FA_/n1 ), .B(
        \ADD_/FAINST[356].FA_/n2 ), .Z(\ADD_/FAINST[356].FA_/n3 ) );
  XOR \ADD_/FAINST[356].FA_/U2  ( .A(b[356]), .B(\ADD_/c[356] ), .Z(
        \ADD_/FAINST[356].FA_/n2 ) );
  XOR \ADD_/FAINST[356].FA_/U1  ( .A(a[356]), .B(\ADD_/c[356] ), .Z(
        \ADD_/FAINST[356].FA_/n1 ) );
  XOR \ADD_/FAINST[355].FA_/U5  ( .A(\ADD_/FAINST[355].FA_/n3 ), .B(
        \ADD_/c[355] ), .Z(\ADD_/c[356] ) );
  XOR \ADD_/FAINST[355].FA_/U4  ( .A(\ADD_/FAINST[355].FA_/n1 ), .B(b[355]), 
        .Z(c[355]) );
  AND \ADD_/FAINST[355].FA_/U3  ( .A(\ADD_/FAINST[355].FA_/n1 ), .B(
        \ADD_/FAINST[355].FA_/n2 ), .Z(\ADD_/FAINST[355].FA_/n3 ) );
  XOR \ADD_/FAINST[355].FA_/U2  ( .A(b[355]), .B(\ADD_/c[355] ), .Z(
        \ADD_/FAINST[355].FA_/n2 ) );
  XOR \ADD_/FAINST[355].FA_/U1  ( .A(a[355]), .B(\ADD_/c[355] ), .Z(
        \ADD_/FAINST[355].FA_/n1 ) );
  XOR \ADD_/FAINST[354].FA_/U5  ( .A(\ADD_/FAINST[354].FA_/n3 ), .B(
        \ADD_/c[354] ), .Z(\ADD_/c[355] ) );
  XOR \ADD_/FAINST[354].FA_/U4  ( .A(\ADD_/FAINST[354].FA_/n1 ), .B(b[354]), 
        .Z(c[354]) );
  AND \ADD_/FAINST[354].FA_/U3  ( .A(\ADD_/FAINST[354].FA_/n1 ), .B(
        \ADD_/FAINST[354].FA_/n2 ), .Z(\ADD_/FAINST[354].FA_/n3 ) );
  XOR \ADD_/FAINST[354].FA_/U2  ( .A(b[354]), .B(\ADD_/c[354] ), .Z(
        \ADD_/FAINST[354].FA_/n2 ) );
  XOR \ADD_/FAINST[354].FA_/U1  ( .A(a[354]), .B(\ADD_/c[354] ), .Z(
        \ADD_/FAINST[354].FA_/n1 ) );
  XOR \ADD_/FAINST[353].FA_/U5  ( .A(\ADD_/FAINST[353].FA_/n3 ), .B(
        \ADD_/c[353] ), .Z(\ADD_/c[354] ) );
  XOR \ADD_/FAINST[353].FA_/U4  ( .A(\ADD_/FAINST[353].FA_/n1 ), .B(b[353]), 
        .Z(c[353]) );
  AND \ADD_/FAINST[353].FA_/U3  ( .A(\ADD_/FAINST[353].FA_/n1 ), .B(
        \ADD_/FAINST[353].FA_/n2 ), .Z(\ADD_/FAINST[353].FA_/n3 ) );
  XOR \ADD_/FAINST[353].FA_/U2  ( .A(b[353]), .B(\ADD_/c[353] ), .Z(
        \ADD_/FAINST[353].FA_/n2 ) );
  XOR \ADD_/FAINST[353].FA_/U1  ( .A(a[353]), .B(\ADD_/c[353] ), .Z(
        \ADD_/FAINST[353].FA_/n1 ) );
  XOR \ADD_/FAINST[352].FA_/U5  ( .A(\ADD_/FAINST[352].FA_/n3 ), .B(
        \ADD_/c[352] ), .Z(\ADD_/c[353] ) );
  XOR \ADD_/FAINST[352].FA_/U4  ( .A(\ADD_/FAINST[352].FA_/n1 ), .B(b[352]), 
        .Z(c[352]) );
  AND \ADD_/FAINST[352].FA_/U3  ( .A(\ADD_/FAINST[352].FA_/n1 ), .B(
        \ADD_/FAINST[352].FA_/n2 ), .Z(\ADD_/FAINST[352].FA_/n3 ) );
  XOR \ADD_/FAINST[352].FA_/U2  ( .A(b[352]), .B(\ADD_/c[352] ), .Z(
        \ADD_/FAINST[352].FA_/n2 ) );
  XOR \ADD_/FAINST[352].FA_/U1  ( .A(a[352]), .B(\ADD_/c[352] ), .Z(
        \ADD_/FAINST[352].FA_/n1 ) );
  XOR \ADD_/FAINST[351].FA_/U5  ( .A(\ADD_/FAINST[351].FA_/n3 ), .B(
        \ADD_/c[351] ), .Z(\ADD_/c[352] ) );
  XOR \ADD_/FAINST[351].FA_/U4  ( .A(\ADD_/FAINST[351].FA_/n1 ), .B(b[351]), 
        .Z(c[351]) );
  AND \ADD_/FAINST[351].FA_/U3  ( .A(\ADD_/FAINST[351].FA_/n1 ), .B(
        \ADD_/FAINST[351].FA_/n2 ), .Z(\ADD_/FAINST[351].FA_/n3 ) );
  XOR \ADD_/FAINST[351].FA_/U2  ( .A(b[351]), .B(\ADD_/c[351] ), .Z(
        \ADD_/FAINST[351].FA_/n2 ) );
  XOR \ADD_/FAINST[351].FA_/U1  ( .A(a[351]), .B(\ADD_/c[351] ), .Z(
        \ADD_/FAINST[351].FA_/n1 ) );
  XOR \ADD_/FAINST[350].FA_/U5  ( .A(\ADD_/FAINST[350].FA_/n3 ), .B(
        \ADD_/c[350] ), .Z(\ADD_/c[351] ) );
  XOR \ADD_/FAINST[350].FA_/U4  ( .A(\ADD_/FAINST[350].FA_/n1 ), .B(b[350]), 
        .Z(c[350]) );
  AND \ADD_/FAINST[350].FA_/U3  ( .A(\ADD_/FAINST[350].FA_/n1 ), .B(
        \ADD_/FAINST[350].FA_/n2 ), .Z(\ADD_/FAINST[350].FA_/n3 ) );
  XOR \ADD_/FAINST[350].FA_/U2  ( .A(b[350]), .B(\ADD_/c[350] ), .Z(
        \ADD_/FAINST[350].FA_/n2 ) );
  XOR \ADD_/FAINST[350].FA_/U1  ( .A(a[350]), .B(\ADD_/c[350] ), .Z(
        \ADD_/FAINST[350].FA_/n1 ) );
  XOR \ADD_/FAINST[349].FA_/U5  ( .A(\ADD_/FAINST[349].FA_/n3 ), .B(
        \ADD_/c[349] ), .Z(\ADD_/c[350] ) );
  XOR \ADD_/FAINST[349].FA_/U4  ( .A(\ADD_/FAINST[349].FA_/n1 ), .B(b[349]), 
        .Z(c[349]) );
  AND \ADD_/FAINST[349].FA_/U3  ( .A(\ADD_/FAINST[349].FA_/n1 ), .B(
        \ADD_/FAINST[349].FA_/n2 ), .Z(\ADD_/FAINST[349].FA_/n3 ) );
  XOR \ADD_/FAINST[349].FA_/U2  ( .A(b[349]), .B(\ADD_/c[349] ), .Z(
        \ADD_/FAINST[349].FA_/n2 ) );
  XOR \ADD_/FAINST[349].FA_/U1  ( .A(a[349]), .B(\ADD_/c[349] ), .Z(
        \ADD_/FAINST[349].FA_/n1 ) );
  XOR \ADD_/FAINST[348].FA_/U5  ( .A(\ADD_/FAINST[348].FA_/n3 ), .B(
        \ADD_/c[348] ), .Z(\ADD_/c[349] ) );
  XOR \ADD_/FAINST[348].FA_/U4  ( .A(\ADD_/FAINST[348].FA_/n1 ), .B(b[348]), 
        .Z(c[348]) );
  AND \ADD_/FAINST[348].FA_/U3  ( .A(\ADD_/FAINST[348].FA_/n1 ), .B(
        \ADD_/FAINST[348].FA_/n2 ), .Z(\ADD_/FAINST[348].FA_/n3 ) );
  XOR \ADD_/FAINST[348].FA_/U2  ( .A(b[348]), .B(\ADD_/c[348] ), .Z(
        \ADD_/FAINST[348].FA_/n2 ) );
  XOR \ADD_/FAINST[348].FA_/U1  ( .A(a[348]), .B(\ADD_/c[348] ), .Z(
        \ADD_/FAINST[348].FA_/n1 ) );
  XOR \ADD_/FAINST[347].FA_/U5  ( .A(\ADD_/FAINST[347].FA_/n3 ), .B(
        \ADD_/c[347] ), .Z(\ADD_/c[348] ) );
  XOR \ADD_/FAINST[347].FA_/U4  ( .A(\ADD_/FAINST[347].FA_/n1 ), .B(b[347]), 
        .Z(c[347]) );
  AND \ADD_/FAINST[347].FA_/U3  ( .A(\ADD_/FAINST[347].FA_/n1 ), .B(
        \ADD_/FAINST[347].FA_/n2 ), .Z(\ADD_/FAINST[347].FA_/n3 ) );
  XOR \ADD_/FAINST[347].FA_/U2  ( .A(b[347]), .B(\ADD_/c[347] ), .Z(
        \ADD_/FAINST[347].FA_/n2 ) );
  XOR \ADD_/FAINST[347].FA_/U1  ( .A(a[347]), .B(\ADD_/c[347] ), .Z(
        \ADD_/FAINST[347].FA_/n1 ) );
  XOR \ADD_/FAINST[346].FA_/U5  ( .A(\ADD_/FAINST[346].FA_/n3 ), .B(
        \ADD_/c[346] ), .Z(\ADD_/c[347] ) );
  XOR \ADD_/FAINST[346].FA_/U4  ( .A(\ADD_/FAINST[346].FA_/n1 ), .B(b[346]), 
        .Z(c[346]) );
  AND \ADD_/FAINST[346].FA_/U3  ( .A(\ADD_/FAINST[346].FA_/n1 ), .B(
        \ADD_/FAINST[346].FA_/n2 ), .Z(\ADD_/FAINST[346].FA_/n3 ) );
  XOR \ADD_/FAINST[346].FA_/U2  ( .A(b[346]), .B(\ADD_/c[346] ), .Z(
        \ADD_/FAINST[346].FA_/n2 ) );
  XOR \ADD_/FAINST[346].FA_/U1  ( .A(a[346]), .B(\ADD_/c[346] ), .Z(
        \ADD_/FAINST[346].FA_/n1 ) );
  XOR \ADD_/FAINST[345].FA_/U5  ( .A(\ADD_/FAINST[345].FA_/n3 ), .B(
        \ADD_/c[345] ), .Z(\ADD_/c[346] ) );
  XOR \ADD_/FAINST[345].FA_/U4  ( .A(\ADD_/FAINST[345].FA_/n1 ), .B(b[345]), 
        .Z(c[345]) );
  AND \ADD_/FAINST[345].FA_/U3  ( .A(\ADD_/FAINST[345].FA_/n1 ), .B(
        \ADD_/FAINST[345].FA_/n2 ), .Z(\ADD_/FAINST[345].FA_/n3 ) );
  XOR \ADD_/FAINST[345].FA_/U2  ( .A(b[345]), .B(\ADD_/c[345] ), .Z(
        \ADD_/FAINST[345].FA_/n2 ) );
  XOR \ADD_/FAINST[345].FA_/U1  ( .A(a[345]), .B(\ADD_/c[345] ), .Z(
        \ADD_/FAINST[345].FA_/n1 ) );
  XOR \ADD_/FAINST[344].FA_/U5  ( .A(\ADD_/FAINST[344].FA_/n3 ), .B(
        \ADD_/c[344] ), .Z(\ADD_/c[345] ) );
  XOR \ADD_/FAINST[344].FA_/U4  ( .A(\ADD_/FAINST[344].FA_/n1 ), .B(b[344]), 
        .Z(c[344]) );
  AND \ADD_/FAINST[344].FA_/U3  ( .A(\ADD_/FAINST[344].FA_/n1 ), .B(
        \ADD_/FAINST[344].FA_/n2 ), .Z(\ADD_/FAINST[344].FA_/n3 ) );
  XOR \ADD_/FAINST[344].FA_/U2  ( .A(b[344]), .B(\ADD_/c[344] ), .Z(
        \ADD_/FAINST[344].FA_/n2 ) );
  XOR \ADD_/FAINST[344].FA_/U1  ( .A(a[344]), .B(\ADD_/c[344] ), .Z(
        \ADD_/FAINST[344].FA_/n1 ) );
  XOR \ADD_/FAINST[343].FA_/U5  ( .A(\ADD_/FAINST[343].FA_/n3 ), .B(
        \ADD_/c[343] ), .Z(\ADD_/c[344] ) );
  XOR \ADD_/FAINST[343].FA_/U4  ( .A(\ADD_/FAINST[343].FA_/n1 ), .B(b[343]), 
        .Z(c[343]) );
  AND \ADD_/FAINST[343].FA_/U3  ( .A(\ADD_/FAINST[343].FA_/n1 ), .B(
        \ADD_/FAINST[343].FA_/n2 ), .Z(\ADD_/FAINST[343].FA_/n3 ) );
  XOR \ADD_/FAINST[343].FA_/U2  ( .A(b[343]), .B(\ADD_/c[343] ), .Z(
        \ADD_/FAINST[343].FA_/n2 ) );
  XOR \ADD_/FAINST[343].FA_/U1  ( .A(a[343]), .B(\ADD_/c[343] ), .Z(
        \ADD_/FAINST[343].FA_/n1 ) );
  XOR \ADD_/FAINST[342].FA_/U5  ( .A(\ADD_/FAINST[342].FA_/n3 ), .B(
        \ADD_/c[342] ), .Z(\ADD_/c[343] ) );
  XOR \ADD_/FAINST[342].FA_/U4  ( .A(\ADD_/FAINST[342].FA_/n1 ), .B(b[342]), 
        .Z(c[342]) );
  AND \ADD_/FAINST[342].FA_/U3  ( .A(\ADD_/FAINST[342].FA_/n1 ), .B(
        \ADD_/FAINST[342].FA_/n2 ), .Z(\ADD_/FAINST[342].FA_/n3 ) );
  XOR \ADD_/FAINST[342].FA_/U2  ( .A(b[342]), .B(\ADD_/c[342] ), .Z(
        \ADD_/FAINST[342].FA_/n2 ) );
  XOR \ADD_/FAINST[342].FA_/U1  ( .A(a[342]), .B(\ADD_/c[342] ), .Z(
        \ADD_/FAINST[342].FA_/n1 ) );
  XOR \ADD_/FAINST[341].FA_/U5  ( .A(\ADD_/FAINST[341].FA_/n3 ), .B(
        \ADD_/c[341] ), .Z(\ADD_/c[342] ) );
  XOR \ADD_/FAINST[341].FA_/U4  ( .A(\ADD_/FAINST[341].FA_/n1 ), .B(b[341]), 
        .Z(c[341]) );
  AND \ADD_/FAINST[341].FA_/U3  ( .A(\ADD_/FAINST[341].FA_/n1 ), .B(
        \ADD_/FAINST[341].FA_/n2 ), .Z(\ADD_/FAINST[341].FA_/n3 ) );
  XOR \ADD_/FAINST[341].FA_/U2  ( .A(b[341]), .B(\ADD_/c[341] ), .Z(
        \ADD_/FAINST[341].FA_/n2 ) );
  XOR \ADD_/FAINST[341].FA_/U1  ( .A(a[341]), .B(\ADD_/c[341] ), .Z(
        \ADD_/FAINST[341].FA_/n1 ) );
  XOR \ADD_/FAINST[340].FA_/U5  ( .A(\ADD_/FAINST[340].FA_/n3 ), .B(
        \ADD_/c[340] ), .Z(\ADD_/c[341] ) );
  XOR \ADD_/FAINST[340].FA_/U4  ( .A(\ADD_/FAINST[340].FA_/n1 ), .B(b[340]), 
        .Z(c[340]) );
  AND \ADD_/FAINST[340].FA_/U3  ( .A(\ADD_/FAINST[340].FA_/n1 ), .B(
        \ADD_/FAINST[340].FA_/n2 ), .Z(\ADD_/FAINST[340].FA_/n3 ) );
  XOR \ADD_/FAINST[340].FA_/U2  ( .A(b[340]), .B(\ADD_/c[340] ), .Z(
        \ADD_/FAINST[340].FA_/n2 ) );
  XOR \ADD_/FAINST[340].FA_/U1  ( .A(a[340]), .B(\ADD_/c[340] ), .Z(
        \ADD_/FAINST[340].FA_/n1 ) );
  XOR \ADD_/FAINST[339].FA_/U5  ( .A(\ADD_/FAINST[339].FA_/n3 ), .B(
        \ADD_/c[339] ), .Z(\ADD_/c[340] ) );
  XOR \ADD_/FAINST[339].FA_/U4  ( .A(\ADD_/FAINST[339].FA_/n1 ), .B(b[339]), 
        .Z(c[339]) );
  AND \ADD_/FAINST[339].FA_/U3  ( .A(\ADD_/FAINST[339].FA_/n1 ), .B(
        \ADD_/FAINST[339].FA_/n2 ), .Z(\ADD_/FAINST[339].FA_/n3 ) );
  XOR \ADD_/FAINST[339].FA_/U2  ( .A(b[339]), .B(\ADD_/c[339] ), .Z(
        \ADD_/FAINST[339].FA_/n2 ) );
  XOR \ADD_/FAINST[339].FA_/U1  ( .A(a[339]), .B(\ADD_/c[339] ), .Z(
        \ADD_/FAINST[339].FA_/n1 ) );
  XOR \ADD_/FAINST[338].FA_/U5  ( .A(\ADD_/FAINST[338].FA_/n3 ), .B(
        \ADD_/c[338] ), .Z(\ADD_/c[339] ) );
  XOR \ADD_/FAINST[338].FA_/U4  ( .A(\ADD_/FAINST[338].FA_/n1 ), .B(b[338]), 
        .Z(c[338]) );
  AND \ADD_/FAINST[338].FA_/U3  ( .A(\ADD_/FAINST[338].FA_/n1 ), .B(
        \ADD_/FAINST[338].FA_/n2 ), .Z(\ADD_/FAINST[338].FA_/n3 ) );
  XOR \ADD_/FAINST[338].FA_/U2  ( .A(b[338]), .B(\ADD_/c[338] ), .Z(
        \ADD_/FAINST[338].FA_/n2 ) );
  XOR \ADD_/FAINST[338].FA_/U1  ( .A(a[338]), .B(\ADD_/c[338] ), .Z(
        \ADD_/FAINST[338].FA_/n1 ) );
  XOR \ADD_/FAINST[337].FA_/U5  ( .A(\ADD_/FAINST[337].FA_/n3 ), .B(
        \ADD_/c[337] ), .Z(\ADD_/c[338] ) );
  XOR \ADD_/FAINST[337].FA_/U4  ( .A(\ADD_/FAINST[337].FA_/n1 ), .B(b[337]), 
        .Z(c[337]) );
  AND \ADD_/FAINST[337].FA_/U3  ( .A(\ADD_/FAINST[337].FA_/n1 ), .B(
        \ADD_/FAINST[337].FA_/n2 ), .Z(\ADD_/FAINST[337].FA_/n3 ) );
  XOR \ADD_/FAINST[337].FA_/U2  ( .A(b[337]), .B(\ADD_/c[337] ), .Z(
        \ADD_/FAINST[337].FA_/n2 ) );
  XOR \ADD_/FAINST[337].FA_/U1  ( .A(a[337]), .B(\ADD_/c[337] ), .Z(
        \ADD_/FAINST[337].FA_/n1 ) );
  XOR \ADD_/FAINST[336].FA_/U5  ( .A(\ADD_/FAINST[336].FA_/n3 ), .B(
        \ADD_/c[336] ), .Z(\ADD_/c[337] ) );
  XOR \ADD_/FAINST[336].FA_/U4  ( .A(\ADD_/FAINST[336].FA_/n1 ), .B(b[336]), 
        .Z(c[336]) );
  AND \ADD_/FAINST[336].FA_/U3  ( .A(\ADD_/FAINST[336].FA_/n1 ), .B(
        \ADD_/FAINST[336].FA_/n2 ), .Z(\ADD_/FAINST[336].FA_/n3 ) );
  XOR \ADD_/FAINST[336].FA_/U2  ( .A(b[336]), .B(\ADD_/c[336] ), .Z(
        \ADD_/FAINST[336].FA_/n2 ) );
  XOR \ADD_/FAINST[336].FA_/U1  ( .A(a[336]), .B(\ADD_/c[336] ), .Z(
        \ADD_/FAINST[336].FA_/n1 ) );
  XOR \ADD_/FAINST[335].FA_/U5  ( .A(\ADD_/FAINST[335].FA_/n3 ), .B(
        \ADD_/c[335] ), .Z(\ADD_/c[336] ) );
  XOR \ADD_/FAINST[335].FA_/U4  ( .A(\ADD_/FAINST[335].FA_/n1 ), .B(b[335]), 
        .Z(c[335]) );
  AND \ADD_/FAINST[335].FA_/U3  ( .A(\ADD_/FAINST[335].FA_/n1 ), .B(
        \ADD_/FAINST[335].FA_/n2 ), .Z(\ADD_/FAINST[335].FA_/n3 ) );
  XOR \ADD_/FAINST[335].FA_/U2  ( .A(b[335]), .B(\ADD_/c[335] ), .Z(
        \ADD_/FAINST[335].FA_/n2 ) );
  XOR \ADD_/FAINST[335].FA_/U1  ( .A(a[335]), .B(\ADD_/c[335] ), .Z(
        \ADD_/FAINST[335].FA_/n1 ) );
  XOR \ADD_/FAINST[334].FA_/U5  ( .A(\ADD_/FAINST[334].FA_/n3 ), .B(
        \ADD_/c[334] ), .Z(\ADD_/c[335] ) );
  XOR \ADD_/FAINST[334].FA_/U4  ( .A(\ADD_/FAINST[334].FA_/n1 ), .B(b[334]), 
        .Z(c[334]) );
  AND \ADD_/FAINST[334].FA_/U3  ( .A(\ADD_/FAINST[334].FA_/n1 ), .B(
        \ADD_/FAINST[334].FA_/n2 ), .Z(\ADD_/FAINST[334].FA_/n3 ) );
  XOR \ADD_/FAINST[334].FA_/U2  ( .A(b[334]), .B(\ADD_/c[334] ), .Z(
        \ADD_/FAINST[334].FA_/n2 ) );
  XOR \ADD_/FAINST[334].FA_/U1  ( .A(a[334]), .B(\ADD_/c[334] ), .Z(
        \ADD_/FAINST[334].FA_/n1 ) );
  XOR \ADD_/FAINST[333].FA_/U5  ( .A(\ADD_/FAINST[333].FA_/n3 ), .B(
        \ADD_/c[333] ), .Z(\ADD_/c[334] ) );
  XOR \ADD_/FAINST[333].FA_/U4  ( .A(\ADD_/FAINST[333].FA_/n1 ), .B(b[333]), 
        .Z(c[333]) );
  AND \ADD_/FAINST[333].FA_/U3  ( .A(\ADD_/FAINST[333].FA_/n1 ), .B(
        \ADD_/FAINST[333].FA_/n2 ), .Z(\ADD_/FAINST[333].FA_/n3 ) );
  XOR \ADD_/FAINST[333].FA_/U2  ( .A(b[333]), .B(\ADD_/c[333] ), .Z(
        \ADD_/FAINST[333].FA_/n2 ) );
  XOR \ADD_/FAINST[333].FA_/U1  ( .A(a[333]), .B(\ADD_/c[333] ), .Z(
        \ADD_/FAINST[333].FA_/n1 ) );
  XOR \ADD_/FAINST[332].FA_/U5  ( .A(\ADD_/FAINST[332].FA_/n3 ), .B(
        \ADD_/c[332] ), .Z(\ADD_/c[333] ) );
  XOR \ADD_/FAINST[332].FA_/U4  ( .A(\ADD_/FAINST[332].FA_/n1 ), .B(b[332]), 
        .Z(c[332]) );
  AND \ADD_/FAINST[332].FA_/U3  ( .A(\ADD_/FAINST[332].FA_/n1 ), .B(
        \ADD_/FAINST[332].FA_/n2 ), .Z(\ADD_/FAINST[332].FA_/n3 ) );
  XOR \ADD_/FAINST[332].FA_/U2  ( .A(b[332]), .B(\ADD_/c[332] ), .Z(
        \ADD_/FAINST[332].FA_/n2 ) );
  XOR \ADD_/FAINST[332].FA_/U1  ( .A(a[332]), .B(\ADD_/c[332] ), .Z(
        \ADD_/FAINST[332].FA_/n1 ) );
  XOR \ADD_/FAINST[331].FA_/U5  ( .A(\ADD_/FAINST[331].FA_/n3 ), .B(
        \ADD_/c[331] ), .Z(\ADD_/c[332] ) );
  XOR \ADD_/FAINST[331].FA_/U4  ( .A(\ADD_/FAINST[331].FA_/n1 ), .B(b[331]), 
        .Z(c[331]) );
  AND \ADD_/FAINST[331].FA_/U3  ( .A(\ADD_/FAINST[331].FA_/n1 ), .B(
        \ADD_/FAINST[331].FA_/n2 ), .Z(\ADD_/FAINST[331].FA_/n3 ) );
  XOR \ADD_/FAINST[331].FA_/U2  ( .A(b[331]), .B(\ADD_/c[331] ), .Z(
        \ADD_/FAINST[331].FA_/n2 ) );
  XOR \ADD_/FAINST[331].FA_/U1  ( .A(a[331]), .B(\ADD_/c[331] ), .Z(
        \ADD_/FAINST[331].FA_/n1 ) );
  XOR \ADD_/FAINST[330].FA_/U5  ( .A(\ADD_/FAINST[330].FA_/n3 ), .B(
        \ADD_/c[330] ), .Z(\ADD_/c[331] ) );
  XOR \ADD_/FAINST[330].FA_/U4  ( .A(\ADD_/FAINST[330].FA_/n1 ), .B(b[330]), 
        .Z(c[330]) );
  AND \ADD_/FAINST[330].FA_/U3  ( .A(\ADD_/FAINST[330].FA_/n1 ), .B(
        \ADD_/FAINST[330].FA_/n2 ), .Z(\ADD_/FAINST[330].FA_/n3 ) );
  XOR \ADD_/FAINST[330].FA_/U2  ( .A(b[330]), .B(\ADD_/c[330] ), .Z(
        \ADD_/FAINST[330].FA_/n2 ) );
  XOR \ADD_/FAINST[330].FA_/U1  ( .A(a[330]), .B(\ADD_/c[330] ), .Z(
        \ADD_/FAINST[330].FA_/n1 ) );
  XOR \ADD_/FAINST[329].FA_/U5  ( .A(\ADD_/FAINST[329].FA_/n3 ), .B(
        \ADD_/c[329] ), .Z(\ADD_/c[330] ) );
  XOR \ADD_/FAINST[329].FA_/U4  ( .A(\ADD_/FAINST[329].FA_/n1 ), .B(b[329]), 
        .Z(c[329]) );
  AND \ADD_/FAINST[329].FA_/U3  ( .A(\ADD_/FAINST[329].FA_/n1 ), .B(
        \ADD_/FAINST[329].FA_/n2 ), .Z(\ADD_/FAINST[329].FA_/n3 ) );
  XOR \ADD_/FAINST[329].FA_/U2  ( .A(b[329]), .B(\ADD_/c[329] ), .Z(
        \ADD_/FAINST[329].FA_/n2 ) );
  XOR \ADD_/FAINST[329].FA_/U1  ( .A(a[329]), .B(\ADD_/c[329] ), .Z(
        \ADD_/FAINST[329].FA_/n1 ) );
  XOR \ADD_/FAINST[328].FA_/U5  ( .A(\ADD_/FAINST[328].FA_/n3 ), .B(
        \ADD_/c[328] ), .Z(\ADD_/c[329] ) );
  XOR \ADD_/FAINST[328].FA_/U4  ( .A(\ADD_/FAINST[328].FA_/n1 ), .B(b[328]), 
        .Z(c[328]) );
  AND \ADD_/FAINST[328].FA_/U3  ( .A(\ADD_/FAINST[328].FA_/n1 ), .B(
        \ADD_/FAINST[328].FA_/n2 ), .Z(\ADD_/FAINST[328].FA_/n3 ) );
  XOR \ADD_/FAINST[328].FA_/U2  ( .A(b[328]), .B(\ADD_/c[328] ), .Z(
        \ADD_/FAINST[328].FA_/n2 ) );
  XOR \ADD_/FAINST[328].FA_/U1  ( .A(a[328]), .B(\ADD_/c[328] ), .Z(
        \ADD_/FAINST[328].FA_/n1 ) );
  XOR \ADD_/FAINST[327].FA_/U5  ( .A(\ADD_/FAINST[327].FA_/n3 ), .B(
        \ADD_/c[327] ), .Z(\ADD_/c[328] ) );
  XOR \ADD_/FAINST[327].FA_/U4  ( .A(\ADD_/FAINST[327].FA_/n1 ), .B(b[327]), 
        .Z(c[327]) );
  AND \ADD_/FAINST[327].FA_/U3  ( .A(\ADD_/FAINST[327].FA_/n1 ), .B(
        \ADD_/FAINST[327].FA_/n2 ), .Z(\ADD_/FAINST[327].FA_/n3 ) );
  XOR \ADD_/FAINST[327].FA_/U2  ( .A(b[327]), .B(\ADD_/c[327] ), .Z(
        \ADD_/FAINST[327].FA_/n2 ) );
  XOR \ADD_/FAINST[327].FA_/U1  ( .A(a[327]), .B(\ADD_/c[327] ), .Z(
        \ADD_/FAINST[327].FA_/n1 ) );
  XOR \ADD_/FAINST[326].FA_/U5  ( .A(\ADD_/FAINST[326].FA_/n3 ), .B(
        \ADD_/c[326] ), .Z(\ADD_/c[327] ) );
  XOR \ADD_/FAINST[326].FA_/U4  ( .A(\ADD_/FAINST[326].FA_/n1 ), .B(b[326]), 
        .Z(c[326]) );
  AND \ADD_/FAINST[326].FA_/U3  ( .A(\ADD_/FAINST[326].FA_/n1 ), .B(
        \ADD_/FAINST[326].FA_/n2 ), .Z(\ADD_/FAINST[326].FA_/n3 ) );
  XOR \ADD_/FAINST[326].FA_/U2  ( .A(b[326]), .B(\ADD_/c[326] ), .Z(
        \ADD_/FAINST[326].FA_/n2 ) );
  XOR \ADD_/FAINST[326].FA_/U1  ( .A(a[326]), .B(\ADD_/c[326] ), .Z(
        \ADD_/FAINST[326].FA_/n1 ) );
  XOR \ADD_/FAINST[325].FA_/U5  ( .A(\ADD_/FAINST[325].FA_/n3 ), .B(
        \ADD_/c[325] ), .Z(\ADD_/c[326] ) );
  XOR \ADD_/FAINST[325].FA_/U4  ( .A(\ADD_/FAINST[325].FA_/n1 ), .B(b[325]), 
        .Z(c[325]) );
  AND \ADD_/FAINST[325].FA_/U3  ( .A(\ADD_/FAINST[325].FA_/n1 ), .B(
        \ADD_/FAINST[325].FA_/n2 ), .Z(\ADD_/FAINST[325].FA_/n3 ) );
  XOR \ADD_/FAINST[325].FA_/U2  ( .A(b[325]), .B(\ADD_/c[325] ), .Z(
        \ADD_/FAINST[325].FA_/n2 ) );
  XOR \ADD_/FAINST[325].FA_/U1  ( .A(a[325]), .B(\ADD_/c[325] ), .Z(
        \ADD_/FAINST[325].FA_/n1 ) );
  XOR \ADD_/FAINST[324].FA_/U5  ( .A(\ADD_/FAINST[324].FA_/n3 ), .B(
        \ADD_/c[324] ), .Z(\ADD_/c[325] ) );
  XOR \ADD_/FAINST[324].FA_/U4  ( .A(\ADD_/FAINST[324].FA_/n1 ), .B(b[324]), 
        .Z(c[324]) );
  AND \ADD_/FAINST[324].FA_/U3  ( .A(\ADD_/FAINST[324].FA_/n1 ), .B(
        \ADD_/FAINST[324].FA_/n2 ), .Z(\ADD_/FAINST[324].FA_/n3 ) );
  XOR \ADD_/FAINST[324].FA_/U2  ( .A(b[324]), .B(\ADD_/c[324] ), .Z(
        \ADD_/FAINST[324].FA_/n2 ) );
  XOR \ADD_/FAINST[324].FA_/U1  ( .A(a[324]), .B(\ADD_/c[324] ), .Z(
        \ADD_/FAINST[324].FA_/n1 ) );
  XOR \ADD_/FAINST[323].FA_/U5  ( .A(\ADD_/FAINST[323].FA_/n3 ), .B(
        \ADD_/c[323] ), .Z(\ADD_/c[324] ) );
  XOR \ADD_/FAINST[323].FA_/U4  ( .A(\ADD_/FAINST[323].FA_/n1 ), .B(b[323]), 
        .Z(c[323]) );
  AND \ADD_/FAINST[323].FA_/U3  ( .A(\ADD_/FAINST[323].FA_/n1 ), .B(
        \ADD_/FAINST[323].FA_/n2 ), .Z(\ADD_/FAINST[323].FA_/n3 ) );
  XOR \ADD_/FAINST[323].FA_/U2  ( .A(b[323]), .B(\ADD_/c[323] ), .Z(
        \ADD_/FAINST[323].FA_/n2 ) );
  XOR \ADD_/FAINST[323].FA_/U1  ( .A(a[323]), .B(\ADD_/c[323] ), .Z(
        \ADD_/FAINST[323].FA_/n1 ) );
  XOR \ADD_/FAINST[322].FA_/U5  ( .A(\ADD_/FAINST[322].FA_/n3 ), .B(
        \ADD_/c[322] ), .Z(\ADD_/c[323] ) );
  XOR \ADD_/FAINST[322].FA_/U4  ( .A(\ADD_/FAINST[322].FA_/n1 ), .B(b[322]), 
        .Z(c[322]) );
  AND \ADD_/FAINST[322].FA_/U3  ( .A(\ADD_/FAINST[322].FA_/n1 ), .B(
        \ADD_/FAINST[322].FA_/n2 ), .Z(\ADD_/FAINST[322].FA_/n3 ) );
  XOR \ADD_/FAINST[322].FA_/U2  ( .A(b[322]), .B(\ADD_/c[322] ), .Z(
        \ADD_/FAINST[322].FA_/n2 ) );
  XOR \ADD_/FAINST[322].FA_/U1  ( .A(a[322]), .B(\ADD_/c[322] ), .Z(
        \ADD_/FAINST[322].FA_/n1 ) );
  XOR \ADD_/FAINST[321].FA_/U5  ( .A(\ADD_/FAINST[321].FA_/n3 ), .B(
        \ADD_/c[321] ), .Z(\ADD_/c[322] ) );
  XOR \ADD_/FAINST[321].FA_/U4  ( .A(\ADD_/FAINST[321].FA_/n1 ), .B(b[321]), 
        .Z(c[321]) );
  AND \ADD_/FAINST[321].FA_/U3  ( .A(\ADD_/FAINST[321].FA_/n1 ), .B(
        \ADD_/FAINST[321].FA_/n2 ), .Z(\ADD_/FAINST[321].FA_/n3 ) );
  XOR \ADD_/FAINST[321].FA_/U2  ( .A(b[321]), .B(\ADD_/c[321] ), .Z(
        \ADD_/FAINST[321].FA_/n2 ) );
  XOR \ADD_/FAINST[321].FA_/U1  ( .A(a[321]), .B(\ADD_/c[321] ), .Z(
        \ADD_/FAINST[321].FA_/n1 ) );
  XOR \ADD_/FAINST[320].FA_/U5  ( .A(\ADD_/FAINST[320].FA_/n3 ), .B(
        \ADD_/c[320] ), .Z(\ADD_/c[321] ) );
  XOR \ADD_/FAINST[320].FA_/U4  ( .A(\ADD_/FAINST[320].FA_/n1 ), .B(b[320]), 
        .Z(c[320]) );
  AND \ADD_/FAINST[320].FA_/U3  ( .A(\ADD_/FAINST[320].FA_/n1 ), .B(
        \ADD_/FAINST[320].FA_/n2 ), .Z(\ADD_/FAINST[320].FA_/n3 ) );
  XOR \ADD_/FAINST[320].FA_/U2  ( .A(b[320]), .B(\ADD_/c[320] ), .Z(
        \ADD_/FAINST[320].FA_/n2 ) );
  XOR \ADD_/FAINST[320].FA_/U1  ( .A(a[320]), .B(\ADD_/c[320] ), .Z(
        \ADD_/FAINST[320].FA_/n1 ) );
  XOR \ADD_/FAINST[319].FA_/U5  ( .A(\ADD_/FAINST[319].FA_/n3 ), .B(
        \ADD_/c[319] ), .Z(\ADD_/c[320] ) );
  XOR \ADD_/FAINST[319].FA_/U4  ( .A(\ADD_/FAINST[319].FA_/n1 ), .B(b[319]), 
        .Z(c[319]) );
  AND \ADD_/FAINST[319].FA_/U3  ( .A(\ADD_/FAINST[319].FA_/n1 ), .B(
        \ADD_/FAINST[319].FA_/n2 ), .Z(\ADD_/FAINST[319].FA_/n3 ) );
  XOR \ADD_/FAINST[319].FA_/U2  ( .A(b[319]), .B(\ADD_/c[319] ), .Z(
        \ADD_/FAINST[319].FA_/n2 ) );
  XOR \ADD_/FAINST[319].FA_/U1  ( .A(a[319]), .B(\ADD_/c[319] ), .Z(
        \ADD_/FAINST[319].FA_/n1 ) );
  XOR \ADD_/FAINST[318].FA_/U5  ( .A(\ADD_/FAINST[318].FA_/n3 ), .B(
        \ADD_/c[318] ), .Z(\ADD_/c[319] ) );
  XOR \ADD_/FAINST[318].FA_/U4  ( .A(\ADD_/FAINST[318].FA_/n1 ), .B(b[318]), 
        .Z(c[318]) );
  AND \ADD_/FAINST[318].FA_/U3  ( .A(\ADD_/FAINST[318].FA_/n1 ), .B(
        \ADD_/FAINST[318].FA_/n2 ), .Z(\ADD_/FAINST[318].FA_/n3 ) );
  XOR \ADD_/FAINST[318].FA_/U2  ( .A(b[318]), .B(\ADD_/c[318] ), .Z(
        \ADD_/FAINST[318].FA_/n2 ) );
  XOR \ADD_/FAINST[318].FA_/U1  ( .A(a[318]), .B(\ADD_/c[318] ), .Z(
        \ADD_/FAINST[318].FA_/n1 ) );
  XOR \ADD_/FAINST[317].FA_/U5  ( .A(\ADD_/FAINST[317].FA_/n3 ), .B(
        \ADD_/c[317] ), .Z(\ADD_/c[318] ) );
  XOR \ADD_/FAINST[317].FA_/U4  ( .A(\ADD_/FAINST[317].FA_/n1 ), .B(b[317]), 
        .Z(c[317]) );
  AND \ADD_/FAINST[317].FA_/U3  ( .A(\ADD_/FAINST[317].FA_/n1 ), .B(
        \ADD_/FAINST[317].FA_/n2 ), .Z(\ADD_/FAINST[317].FA_/n3 ) );
  XOR \ADD_/FAINST[317].FA_/U2  ( .A(b[317]), .B(\ADD_/c[317] ), .Z(
        \ADD_/FAINST[317].FA_/n2 ) );
  XOR \ADD_/FAINST[317].FA_/U1  ( .A(a[317]), .B(\ADD_/c[317] ), .Z(
        \ADD_/FAINST[317].FA_/n1 ) );
  XOR \ADD_/FAINST[316].FA_/U5  ( .A(\ADD_/FAINST[316].FA_/n3 ), .B(
        \ADD_/c[316] ), .Z(\ADD_/c[317] ) );
  XOR \ADD_/FAINST[316].FA_/U4  ( .A(\ADD_/FAINST[316].FA_/n1 ), .B(b[316]), 
        .Z(c[316]) );
  AND \ADD_/FAINST[316].FA_/U3  ( .A(\ADD_/FAINST[316].FA_/n1 ), .B(
        \ADD_/FAINST[316].FA_/n2 ), .Z(\ADD_/FAINST[316].FA_/n3 ) );
  XOR \ADD_/FAINST[316].FA_/U2  ( .A(b[316]), .B(\ADD_/c[316] ), .Z(
        \ADD_/FAINST[316].FA_/n2 ) );
  XOR \ADD_/FAINST[316].FA_/U1  ( .A(a[316]), .B(\ADD_/c[316] ), .Z(
        \ADD_/FAINST[316].FA_/n1 ) );
  XOR \ADD_/FAINST[315].FA_/U5  ( .A(\ADD_/FAINST[315].FA_/n3 ), .B(
        \ADD_/c[315] ), .Z(\ADD_/c[316] ) );
  XOR \ADD_/FAINST[315].FA_/U4  ( .A(\ADD_/FAINST[315].FA_/n1 ), .B(b[315]), 
        .Z(c[315]) );
  AND \ADD_/FAINST[315].FA_/U3  ( .A(\ADD_/FAINST[315].FA_/n1 ), .B(
        \ADD_/FAINST[315].FA_/n2 ), .Z(\ADD_/FAINST[315].FA_/n3 ) );
  XOR \ADD_/FAINST[315].FA_/U2  ( .A(b[315]), .B(\ADD_/c[315] ), .Z(
        \ADD_/FAINST[315].FA_/n2 ) );
  XOR \ADD_/FAINST[315].FA_/U1  ( .A(a[315]), .B(\ADD_/c[315] ), .Z(
        \ADD_/FAINST[315].FA_/n1 ) );
  XOR \ADD_/FAINST[314].FA_/U5  ( .A(\ADD_/FAINST[314].FA_/n3 ), .B(
        \ADD_/c[314] ), .Z(\ADD_/c[315] ) );
  XOR \ADD_/FAINST[314].FA_/U4  ( .A(\ADD_/FAINST[314].FA_/n1 ), .B(b[314]), 
        .Z(c[314]) );
  AND \ADD_/FAINST[314].FA_/U3  ( .A(\ADD_/FAINST[314].FA_/n1 ), .B(
        \ADD_/FAINST[314].FA_/n2 ), .Z(\ADD_/FAINST[314].FA_/n3 ) );
  XOR \ADD_/FAINST[314].FA_/U2  ( .A(b[314]), .B(\ADD_/c[314] ), .Z(
        \ADD_/FAINST[314].FA_/n2 ) );
  XOR \ADD_/FAINST[314].FA_/U1  ( .A(a[314]), .B(\ADD_/c[314] ), .Z(
        \ADD_/FAINST[314].FA_/n1 ) );
  XOR \ADD_/FAINST[313].FA_/U5  ( .A(\ADD_/FAINST[313].FA_/n3 ), .B(
        \ADD_/c[313] ), .Z(\ADD_/c[314] ) );
  XOR \ADD_/FAINST[313].FA_/U4  ( .A(\ADD_/FAINST[313].FA_/n1 ), .B(b[313]), 
        .Z(c[313]) );
  AND \ADD_/FAINST[313].FA_/U3  ( .A(\ADD_/FAINST[313].FA_/n1 ), .B(
        \ADD_/FAINST[313].FA_/n2 ), .Z(\ADD_/FAINST[313].FA_/n3 ) );
  XOR \ADD_/FAINST[313].FA_/U2  ( .A(b[313]), .B(\ADD_/c[313] ), .Z(
        \ADD_/FAINST[313].FA_/n2 ) );
  XOR \ADD_/FAINST[313].FA_/U1  ( .A(a[313]), .B(\ADD_/c[313] ), .Z(
        \ADD_/FAINST[313].FA_/n1 ) );
  XOR \ADD_/FAINST[312].FA_/U5  ( .A(\ADD_/FAINST[312].FA_/n3 ), .B(
        \ADD_/c[312] ), .Z(\ADD_/c[313] ) );
  XOR \ADD_/FAINST[312].FA_/U4  ( .A(\ADD_/FAINST[312].FA_/n1 ), .B(b[312]), 
        .Z(c[312]) );
  AND \ADD_/FAINST[312].FA_/U3  ( .A(\ADD_/FAINST[312].FA_/n1 ), .B(
        \ADD_/FAINST[312].FA_/n2 ), .Z(\ADD_/FAINST[312].FA_/n3 ) );
  XOR \ADD_/FAINST[312].FA_/U2  ( .A(b[312]), .B(\ADD_/c[312] ), .Z(
        \ADD_/FAINST[312].FA_/n2 ) );
  XOR \ADD_/FAINST[312].FA_/U1  ( .A(a[312]), .B(\ADD_/c[312] ), .Z(
        \ADD_/FAINST[312].FA_/n1 ) );
  XOR \ADD_/FAINST[311].FA_/U5  ( .A(\ADD_/FAINST[311].FA_/n3 ), .B(
        \ADD_/c[311] ), .Z(\ADD_/c[312] ) );
  XOR \ADD_/FAINST[311].FA_/U4  ( .A(\ADD_/FAINST[311].FA_/n1 ), .B(b[311]), 
        .Z(c[311]) );
  AND \ADD_/FAINST[311].FA_/U3  ( .A(\ADD_/FAINST[311].FA_/n1 ), .B(
        \ADD_/FAINST[311].FA_/n2 ), .Z(\ADD_/FAINST[311].FA_/n3 ) );
  XOR \ADD_/FAINST[311].FA_/U2  ( .A(b[311]), .B(\ADD_/c[311] ), .Z(
        \ADD_/FAINST[311].FA_/n2 ) );
  XOR \ADD_/FAINST[311].FA_/U1  ( .A(a[311]), .B(\ADD_/c[311] ), .Z(
        \ADD_/FAINST[311].FA_/n1 ) );
  XOR \ADD_/FAINST[310].FA_/U5  ( .A(\ADD_/FAINST[310].FA_/n3 ), .B(
        \ADD_/c[310] ), .Z(\ADD_/c[311] ) );
  XOR \ADD_/FAINST[310].FA_/U4  ( .A(\ADD_/FAINST[310].FA_/n1 ), .B(b[310]), 
        .Z(c[310]) );
  AND \ADD_/FAINST[310].FA_/U3  ( .A(\ADD_/FAINST[310].FA_/n1 ), .B(
        \ADD_/FAINST[310].FA_/n2 ), .Z(\ADD_/FAINST[310].FA_/n3 ) );
  XOR \ADD_/FAINST[310].FA_/U2  ( .A(b[310]), .B(\ADD_/c[310] ), .Z(
        \ADD_/FAINST[310].FA_/n2 ) );
  XOR \ADD_/FAINST[310].FA_/U1  ( .A(a[310]), .B(\ADD_/c[310] ), .Z(
        \ADD_/FAINST[310].FA_/n1 ) );
  XOR \ADD_/FAINST[309].FA_/U5  ( .A(\ADD_/FAINST[309].FA_/n3 ), .B(
        \ADD_/c[309] ), .Z(\ADD_/c[310] ) );
  XOR \ADD_/FAINST[309].FA_/U4  ( .A(\ADD_/FAINST[309].FA_/n1 ), .B(b[309]), 
        .Z(c[309]) );
  AND \ADD_/FAINST[309].FA_/U3  ( .A(\ADD_/FAINST[309].FA_/n1 ), .B(
        \ADD_/FAINST[309].FA_/n2 ), .Z(\ADD_/FAINST[309].FA_/n3 ) );
  XOR \ADD_/FAINST[309].FA_/U2  ( .A(b[309]), .B(\ADD_/c[309] ), .Z(
        \ADD_/FAINST[309].FA_/n2 ) );
  XOR \ADD_/FAINST[309].FA_/U1  ( .A(a[309]), .B(\ADD_/c[309] ), .Z(
        \ADD_/FAINST[309].FA_/n1 ) );
  XOR \ADD_/FAINST[308].FA_/U5  ( .A(\ADD_/FAINST[308].FA_/n3 ), .B(
        \ADD_/c[308] ), .Z(\ADD_/c[309] ) );
  XOR \ADD_/FAINST[308].FA_/U4  ( .A(\ADD_/FAINST[308].FA_/n1 ), .B(b[308]), 
        .Z(c[308]) );
  AND \ADD_/FAINST[308].FA_/U3  ( .A(\ADD_/FAINST[308].FA_/n1 ), .B(
        \ADD_/FAINST[308].FA_/n2 ), .Z(\ADD_/FAINST[308].FA_/n3 ) );
  XOR \ADD_/FAINST[308].FA_/U2  ( .A(b[308]), .B(\ADD_/c[308] ), .Z(
        \ADD_/FAINST[308].FA_/n2 ) );
  XOR \ADD_/FAINST[308].FA_/U1  ( .A(a[308]), .B(\ADD_/c[308] ), .Z(
        \ADD_/FAINST[308].FA_/n1 ) );
  XOR \ADD_/FAINST[307].FA_/U5  ( .A(\ADD_/FAINST[307].FA_/n3 ), .B(
        \ADD_/c[307] ), .Z(\ADD_/c[308] ) );
  XOR \ADD_/FAINST[307].FA_/U4  ( .A(\ADD_/FAINST[307].FA_/n1 ), .B(b[307]), 
        .Z(c[307]) );
  AND \ADD_/FAINST[307].FA_/U3  ( .A(\ADD_/FAINST[307].FA_/n1 ), .B(
        \ADD_/FAINST[307].FA_/n2 ), .Z(\ADD_/FAINST[307].FA_/n3 ) );
  XOR \ADD_/FAINST[307].FA_/U2  ( .A(b[307]), .B(\ADD_/c[307] ), .Z(
        \ADD_/FAINST[307].FA_/n2 ) );
  XOR \ADD_/FAINST[307].FA_/U1  ( .A(a[307]), .B(\ADD_/c[307] ), .Z(
        \ADD_/FAINST[307].FA_/n1 ) );
  XOR \ADD_/FAINST[306].FA_/U5  ( .A(\ADD_/FAINST[306].FA_/n3 ), .B(
        \ADD_/c[306] ), .Z(\ADD_/c[307] ) );
  XOR \ADD_/FAINST[306].FA_/U4  ( .A(\ADD_/FAINST[306].FA_/n1 ), .B(b[306]), 
        .Z(c[306]) );
  AND \ADD_/FAINST[306].FA_/U3  ( .A(\ADD_/FAINST[306].FA_/n1 ), .B(
        \ADD_/FAINST[306].FA_/n2 ), .Z(\ADD_/FAINST[306].FA_/n3 ) );
  XOR \ADD_/FAINST[306].FA_/U2  ( .A(b[306]), .B(\ADD_/c[306] ), .Z(
        \ADD_/FAINST[306].FA_/n2 ) );
  XOR \ADD_/FAINST[306].FA_/U1  ( .A(a[306]), .B(\ADD_/c[306] ), .Z(
        \ADD_/FAINST[306].FA_/n1 ) );
  XOR \ADD_/FAINST[305].FA_/U5  ( .A(\ADD_/FAINST[305].FA_/n3 ), .B(
        \ADD_/c[305] ), .Z(\ADD_/c[306] ) );
  XOR \ADD_/FAINST[305].FA_/U4  ( .A(\ADD_/FAINST[305].FA_/n1 ), .B(b[305]), 
        .Z(c[305]) );
  AND \ADD_/FAINST[305].FA_/U3  ( .A(\ADD_/FAINST[305].FA_/n1 ), .B(
        \ADD_/FAINST[305].FA_/n2 ), .Z(\ADD_/FAINST[305].FA_/n3 ) );
  XOR \ADD_/FAINST[305].FA_/U2  ( .A(b[305]), .B(\ADD_/c[305] ), .Z(
        \ADD_/FAINST[305].FA_/n2 ) );
  XOR \ADD_/FAINST[305].FA_/U1  ( .A(a[305]), .B(\ADD_/c[305] ), .Z(
        \ADD_/FAINST[305].FA_/n1 ) );
  XOR \ADD_/FAINST[304].FA_/U5  ( .A(\ADD_/FAINST[304].FA_/n3 ), .B(
        \ADD_/c[304] ), .Z(\ADD_/c[305] ) );
  XOR \ADD_/FAINST[304].FA_/U4  ( .A(\ADD_/FAINST[304].FA_/n1 ), .B(b[304]), 
        .Z(c[304]) );
  AND \ADD_/FAINST[304].FA_/U3  ( .A(\ADD_/FAINST[304].FA_/n1 ), .B(
        \ADD_/FAINST[304].FA_/n2 ), .Z(\ADD_/FAINST[304].FA_/n3 ) );
  XOR \ADD_/FAINST[304].FA_/U2  ( .A(b[304]), .B(\ADD_/c[304] ), .Z(
        \ADD_/FAINST[304].FA_/n2 ) );
  XOR \ADD_/FAINST[304].FA_/U1  ( .A(a[304]), .B(\ADD_/c[304] ), .Z(
        \ADD_/FAINST[304].FA_/n1 ) );
  XOR \ADD_/FAINST[303].FA_/U5  ( .A(\ADD_/FAINST[303].FA_/n3 ), .B(
        \ADD_/c[303] ), .Z(\ADD_/c[304] ) );
  XOR \ADD_/FAINST[303].FA_/U4  ( .A(\ADD_/FAINST[303].FA_/n1 ), .B(b[303]), 
        .Z(c[303]) );
  AND \ADD_/FAINST[303].FA_/U3  ( .A(\ADD_/FAINST[303].FA_/n1 ), .B(
        \ADD_/FAINST[303].FA_/n2 ), .Z(\ADD_/FAINST[303].FA_/n3 ) );
  XOR \ADD_/FAINST[303].FA_/U2  ( .A(b[303]), .B(\ADD_/c[303] ), .Z(
        \ADD_/FAINST[303].FA_/n2 ) );
  XOR \ADD_/FAINST[303].FA_/U1  ( .A(a[303]), .B(\ADD_/c[303] ), .Z(
        \ADD_/FAINST[303].FA_/n1 ) );
  XOR \ADD_/FAINST[302].FA_/U5  ( .A(\ADD_/FAINST[302].FA_/n3 ), .B(
        \ADD_/c[302] ), .Z(\ADD_/c[303] ) );
  XOR \ADD_/FAINST[302].FA_/U4  ( .A(\ADD_/FAINST[302].FA_/n1 ), .B(b[302]), 
        .Z(c[302]) );
  AND \ADD_/FAINST[302].FA_/U3  ( .A(\ADD_/FAINST[302].FA_/n1 ), .B(
        \ADD_/FAINST[302].FA_/n2 ), .Z(\ADD_/FAINST[302].FA_/n3 ) );
  XOR \ADD_/FAINST[302].FA_/U2  ( .A(b[302]), .B(\ADD_/c[302] ), .Z(
        \ADD_/FAINST[302].FA_/n2 ) );
  XOR \ADD_/FAINST[302].FA_/U1  ( .A(a[302]), .B(\ADD_/c[302] ), .Z(
        \ADD_/FAINST[302].FA_/n1 ) );
  XOR \ADD_/FAINST[301].FA_/U5  ( .A(\ADD_/FAINST[301].FA_/n3 ), .B(
        \ADD_/c[301] ), .Z(\ADD_/c[302] ) );
  XOR \ADD_/FAINST[301].FA_/U4  ( .A(\ADD_/FAINST[301].FA_/n1 ), .B(b[301]), 
        .Z(c[301]) );
  AND \ADD_/FAINST[301].FA_/U3  ( .A(\ADD_/FAINST[301].FA_/n1 ), .B(
        \ADD_/FAINST[301].FA_/n2 ), .Z(\ADD_/FAINST[301].FA_/n3 ) );
  XOR \ADD_/FAINST[301].FA_/U2  ( .A(b[301]), .B(\ADD_/c[301] ), .Z(
        \ADD_/FAINST[301].FA_/n2 ) );
  XOR \ADD_/FAINST[301].FA_/U1  ( .A(a[301]), .B(\ADD_/c[301] ), .Z(
        \ADD_/FAINST[301].FA_/n1 ) );
  XOR \ADD_/FAINST[300].FA_/U5  ( .A(\ADD_/FAINST[300].FA_/n3 ), .B(
        \ADD_/c[300] ), .Z(\ADD_/c[301] ) );
  XOR \ADD_/FAINST[300].FA_/U4  ( .A(\ADD_/FAINST[300].FA_/n1 ), .B(b[300]), 
        .Z(c[300]) );
  AND \ADD_/FAINST[300].FA_/U3  ( .A(\ADD_/FAINST[300].FA_/n1 ), .B(
        \ADD_/FAINST[300].FA_/n2 ), .Z(\ADD_/FAINST[300].FA_/n3 ) );
  XOR \ADD_/FAINST[300].FA_/U2  ( .A(b[300]), .B(\ADD_/c[300] ), .Z(
        \ADD_/FAINST[300].FA_/n2 ) );
  XOR \ADD_/FAINST[300].FA_/U1  ( .A(a[300]), .B(\ADD_/c[300] ), .Z(
        \ADD_/FAINST[300].FA_/n1 ) );
  XOR \ADD_/FAINST[299].FA_/U5  ( .A(\ADD_/FAINST[299].FA_/n3 ), .B(
        \ADD_/c[299] ), .Z(\ADD_/c[300] ) );
  XOR \ADD_/FAINST[299].FA_/U4  ( .A(\ADD_/FAINST[299].FA_/n1 ), .B(b[299]), 
        .Z(c[299]) );
  AND \ADD_/FAINST[299].FA_/U3  ( .A(\ADD_/FAINST[299].FA_/n1 ), .B(
        \ADD_/FAINST[299].FA_/n2 ), .Z(\ADD_/FAINST[299].FA_/n3 ) );
  XOR \ADD_/FAINST[299].FA_/U2  ( .A(b[299]), .B(\ADD_/c[299] ), .Z(
        \ADD_/FAINST[299].FA_/n2 ) );
  XOR \ADD_/FAINST[299].FA_/U1  ( .A(a[299]), .B(\ADD_/c[299] ), .Z(
        \ADD_/FAINST[299].FA_/n1 ) );
  XOR \ADD_/FAINST[298].FA_/U5  ( .A(\ADD_/FAINST[298].FA_/n3 ), .B(
        \ADD_/c[298] ), .Z(\ADD_/c[299] ) );
  XOR \ADD_/FAINST[298].FA_/U4  ( .A(\ADD_/FAINST[298].FA_/n1 ), .B(b[298]), 
        .Z(c[298]) );
  AND \ADD_/FAINST[298].FA_/U3  ( .A(\ADD_/FAINST[298].FA_/n1 ), .B(
        \ADD_/FAINST[298].FA_/n2 ), .Z(\ADD_/FAINST[298].FA_/n3 ) );
  XOR \ADD_/FAINST[298].FA_/U2  ( .A(b[298]), .B(\ADD_/c[298] ), .Z(
        \ADD_/FAINST[298].FA_/n2 ) );
  XOR \ADD_/FAINST[298].FA_/U1  ( .A(a[298]), .B(\ADD_/c[298] ), .Z(
        \ADD_/FAINST[298].FA_/n1 ) );
  XOR \ADD_/FAINST[297].FA_/U5  ( .A(\ADD_/FAINST[297].FA_/n3 ), .B(
        \ADD_/c[297] ), .Z(\ADD_/c[298] ) );
  XOR \ADD_/FAINST[297].FA_/U4  ( .A(\ADD_/FAINST[297].FA_/n1 ), .B(b[297]), 
        .Z(c[297]) );
  AND \ADD_/FAINST[297].FA_/U3  ( .A(\ADD_/FAINST[297].FA_/n1 ), .B(
        \ADD_/FAINST[297].FA_/n2 ), .Z(\ADD_/FAINST[297].FA_/n3 ) );
  XOR \ADD_/FAINST[297].FA_/U2  ( .A(b[297]), .B(\ADD_/c[297] ), .Z(
        \ADD_/FAINST[297].FA_/n2 ) );
  XOR \ADD_/FAINST[297].FA_/U1  ( .A(a[297]), .B(\ADD_/c[297] ), .Z(
        \ADD_/FAINST[297].FA_/n1 ) );
  XOR \ADD_/FAINST[296].FA_/U5  ( .A(\ADD_/FAINST[296].FA_/n3 ), .B(
        \ADD_/c[296] ), .Z(\ADD_/c[297] ) );
  XOR \ADD_/FAINST[296].FA_/U4  ( .A(\ADD_/FAINST[296].FA_/n1 ), .B(b[296]), 
        .Z(c[296]) );
  AND \ADD_/FAINST[296].FA_/U3  ( .A(\ADD_/FAINST[296].FA_/n1 ), .B(
        \ADD_/FAINST[296].FA_/n2 ), .Z(\ADD_/FAINST[296].FA_/n3 ) );
  XOR \ADD_/FAINST[296].FA_/U2  ( .A(b[296]), .B(\ADD_/c[296] ), .Z(
        \ADD_/FAINST[296].FA_/n2 ) );
  XOR \ADD_/FAINST[296].FA_/U1  ( .A(a[296]), .B(\ADD_/c[296] ), .Z(
        \ADD_/FAINST[296].FA_/n1 ) );
  XOR \ADD_/FAINST[295].FA_/U5  ( .A(\ADD_/FAINST[295].FA_/n3 ), .B(
        \ADD_/c[295] ), .Z(\ADD_/c[296] ) );
  XOR \ADD_/FAINST[295].FA_/U4  ( .A(\ADD_/FAINST[295].FA_/n1 ), .B(b[295]), 
        .Z(c[295]) );
  AND \ADD_/FAINST[295].FA_/U3  ( .A(\ADD_/FAINST[295].FA_/n1 ), .B(
        \ADD_/FAINST[295].FA_/n2 ), .Z(\ADD_/FAINST[295].FA_/n3 ) );
  XOR \ADD_/FAINST[295].FA_/U2  ( .A(b[295]), .B(\ADD_/c[295] ), .Z(
        \ADD_/FAINST[295].FA_/n2 ) );
  XOR \ADD_/FAINST[295].FA_/U1  ( .A(a[295]), .B(\ADD_/c[295] ), .Z(
        \ADD_/FAINST[295].FA_/n1 ) );
  XOR \ADD_/FAINST[294].FA_/U5  ( .A(\ADD_/FAINST[294].FA_/n3 ), .B(
        \ADD_/c[294] ), .Z(\ADD_/c[295] ) );
  XOR \ADD_/FAINST[294].FA_/U4  ( .A(\ADD_/FAINST[294].FA_/n1 ), .B(b[294]), 
        .Z(c[294]) );
  AND \ADD_/FAINST[294].FA_/U3  ( .A(\ADD_/FAINST[294].FA_/n1 ), .B(
        \ADD_/FAINST[294].FA_/n2 ), .Z(\ADD_/FAINST[294].FA_/n3 ) );
  XOR \ADD_/FAINST[294].FA_/U2  ( .A(b[294]), .B(\ADD_/c[294] ), .Z(
        \ADD_/FAINST[294].FA_/n2 ) );
  XOR \ADD_/FAINST[294].FA_/U1  ( .A(a[294]), .B(\ADD_/c[294] ), .Z(
        \ADD_/FAINST[294].FA_/n1 ) );
  XOR \ADD_/FAINST[293].FA_/U5  ( .A(\ADD_/FAINST[293].FA_/n3 ), .B(
        \ADD_/c[293] ), .Z(\ADD_/c[294] ) );
  XOR \ADD_/FAINST[293].FA_/U4  ( .A(\ADD_/FAINST[293].FA_/n1 ), .B(b[293]), 
        .Z(c[293]) );
  AND \ADD_/FAINST[293].FA_/U3  ( .A(\ADD_/FAINST[293].FA_/n1 ), .B(
        \ADD_/FAINST[293].FA_/n2 ), .Z(\ADD_/FAINST[293].FA_/n3 ) );
  XOR \ADD_/FAINST[293].FA_/U2  ( .A(b[293]), .B(\ADD_/c[293] ), .Z(
        \ADD_/FAINST[293].FA_/n2 ) );
  XOR \ADD_/FAINST[293].FA_/U1  ( .A(a[293]), .B(\ADD_/c[293] ), .Z(
        \ADD_/FAINST[293].FA_/n1 ) );
  XOR \ADD_/FAINST[292].FA_/U5  ( .A(\ADD_/FAINST[292].FA_/n3 ), .B(
        \ADD_/c[292] ), .Z(\ADD_/c[293] ) );
  XOR \ADD_/FAINST[292].FA_/U4  ( .A(\ADD_/FAINST[292].FA_/n1 ), .B(b[292]), 
        .Z(c[292]) );
  AND \ADD_/FAINST[292].FA_/U3  ( .A(\ADD_/FAINST[292].FA_/n1 ), .B(
        \ADD_/FAINST[292].FA_/n2 ), .Z(\ADD_/FAINST[292].FA_/n3 ) );
  XOR \ADD_/FAINST[292].FA_/U2  ( .A(b[292]), .B(\ADD_/c[292] ), .Z(
        \ADD_/FAINST[292].FA_/n2 ) );
  XOR \ADD_/FAINST[292].FA_/U1  ( .A(a[292]), .B(\ADD_/c[292] ), .Z(
        \ADD_/FAINST[292].FA_/n1 ) );
  XOR \ADD_/FAINST[291].FA_/U5  ( .A(\ADD_/FAINST[291].FA_/n3 ), .B(
        \ADD_/c[291] ), .Z(\ADD_/c[292] ) );
  XOR \ADD_/FAINST[291].FA_/U4  ( .A(\ADD_/FAINST[291].FA_/n1 ), .B(b[291]), 
        .Z(c[291]) );
  AND \ADD_/FAINST[291].FA_/U3  ( .A(\ADD_/FAINST[291].FA_/n1 ), .B(
        \ADD_/FAINST[291].FA_/n2 ), .Z(\ADD_/FAINST[291].FA_/n3 ) );
  XOR \ADD_/FAINST[291].FA_/U2  ( .A(b[291]), .B(\ADD_/c[291] ), .Z(
        \ADD_/FAINST[291].FA_/n2 ) );
  XOR \ADD_/FAINST[291].FA_/U1  ( .A(a[291]), .B(\ADD_/c[291] ), .Z(
        \ADD_/FAINST[291].FA_/n1 ) );
  XOR \ADD_/FAINST[290].FA_/U5  ( .A(\ADD_/FAINST[290].FA_/n3 ), .B(
        \ADD_/c[290] ), .Z(\ADD_/c[291] ) );
  XOR \ADD_/FAINST[290].FA_/U4  ( .A(\ADD_/FAINST[290].FA_/n1 ), .B(b[290]), 
        .Z(c[290]) );
  AND \ADD_/FAINST[290].FA_/U3  ( .A(\ADD_/FAINST[290].FA_/n1 ), .B(
        \ADD_/FAINST[290].FA_/n2 ), .Z(\ADD_/FAINST[290].FA_/n3 ) );
  XOR \ADD_/FAINST[290].FA_/U2  ( .A(b[290]), .B(\ADD_/c[290] ), .Z(
        \ADD_/FAINST[290].FA_/n2 ) );
  XOR \ADD_/FAINST[290].FA_/U1  ( .A(a[290]), .B(\ADD_/c[290] ), .Z(
        \ADD_/FAINST[290].FA_/n1 ) );
  XOR \ADD_/FAINST[289].FA_/U5  ( .A(\ADD_/FAINST[289].FA_/n3 ), .B(
        \ADD_/c[289] ), .Z(\ADD_/c[290] ) );
  XOR \ADD_/FAINST[289].FA_/U4  ( .A(\ADD_/FAINST[289].FA_/n1 ), .B(b[289]), 
        .Z(c[289]) );
  AND \ADD_/FAINST[289].FA_/U3  ( .A(\ADD_/FAINST[289].FA_/n1 ), .B(
        \ADD_/FAINST[289].FA_/n2 ), .Z(\ADD_/FAINST[289].FA_/n3 ) );
  XOR \ADD_/FAINST[289].FA_/U2  ( .A(b[289]), .B(\ADD_/c[289] ), .Z(
        \ADD_/FAINST[289].FA_/n2 ) );
  XOR \ADD_/FAINST[289].FA_/U1  ( .A(a[289]), .B(\ADD_/c[289] ), .Z(
        \ADD_/FAINST[289].FA_/n1 ) );
  XOR \ADD_/FAINST[288].FA_/U5  ( .A(\ADD_/FAINST[288].FA_/n3 ), .B(
        \ADD_/c[288] ), .Z(\ADD_/c[289] ) );
  XOR \ADD_/FAINST[288].FA_/U4  ( .A(\ADD_/FAINST[288].FA_/n1 ), .B(b[288]), 
        .Z(c[288]) );
  AND \ADD_/FAINST[288].FA_/U3  ( .A(\ADD_/FAINST[288].FA_/n1 ), .B(
        \ADD_/FAINST[288].FA_/n2 ), .Z(\ADD_/FAINST[288].FA_/n3 ) );
  XOR \ADD_/FAINST[288].FA_/U2  ( .A(b[288]), .B(\ADD_/c[288] ), .Z(
        \ADD_/FAINST[288].FA_/n2 ) );
  XOR \ADD_/FAINST[288].FA_/U1  ( .A(a[288]), .B(\ADD_/c[288] ), .Z(
        \ADD_/FAINST[288].FA_/n1 ) );
  XOR \ADD_/FAINST[287].FA_/U5  ( .A(\ADD_/FAINST[287].FA_/n3 ), .B(
        \ADD_/c[287] ), .Z(\ADD_/c[288] ) );
  XOR \ADD_/FAINST[287].FA_/U4  ( .A(\ADD_/FAINST[287].FA_/n1 ), .B(b[287]), 
        .Z(c[287]) );
  AND \ADD_/FAINST[287].FA_/U3  ( .A(\ADD_/FAINST[287].FA_/n1 ), .B(
        \ADD_/FAINST[287].FA_/n2 ), .Z(\ADD_/FAINST[287].FA_/n3 ) );
  XOR \ADD_/FAINST[287].FA_/U2  ( .A(b[287]), .B(\ADD_/c[287] ), .Z(
        \ADD_/FAINST[287].FA_/n2 ) );
  XOR \ADD_/FAINST[287].FA_/U1  ( .A(a[287]), .B(\ADD_/c[287] ), .Z(
        \ADD_/FAINST[287].FA_/n1 ) );
  XOR \ADD_/FAINST[286].FA_/U5  ( .A(\ADD_/FAINST[286].FA_/n3 ), .B(
        \ADD_/c[286] ), .Z(\ADD_/c[287] ) );
  XOR \ADD_/FAINST[286].FA_/U4  ( .A(\ADD_/FAINST[286].FA_/n1 ), .B(b[286]), 
        .Z(c[286]) );
  AND \ADD_/FAINST[286].FA_/U3  ( .A(\ADD_/FAINST[286].FA_/n1 ), .B(
        \ADD_/FAINST[286].FA_/n2 ), .Z(\ADD_/FAINST[286].FA_/n3 ) );
  XOR \ADD_/FAINST[286].FA_/U2  ( .A(b[286]), .B(\ADD_/c[286] ), .Z(
        \ADD_/FAINST[286].FA_/n2 ) );
  XOR \ADD_/FAINST[286].FA_/U1  ( .A(a[286]), .B(\ADD_/c[286] ), .Z(
        \ADD_/FAINST[286].FA_/n1 ) );
  XOR \ADD_/FAINST[285].FA_/U5  ( .A(\ADD_/FAINST[285].FA_/n3 ), .B(
        \ADD_/c[285] ), .Z(\ADD_/c[286] ) );
  XOR \ADD_/FAINST[285].FA_/U4  ( .A(\ADD_/FAINST[285].FA_/n1 ), .B(b[285]), 
        .Z(c[285]) );
  AND \ADD_/FAINST[285].FA_/U3  ( .A(\ADD_/FAINST[285].FA_/n1 ), .B(
        \ADD_/FAINST[285].FA_/n2 ), .Z(\ADD_/FAINST[285].FA_/n3 ) );
  XOR \ADD_/FAINST[285].FA_/U2  ( .A(b[285]), .B(\ADD_/c[285] ), .Z(
        \ADD_/FAINST[285].FA_/n2 ) );
  XOR \ADD_/FAINST[285].FA_/U1  ( .A(a[285]), .B(\ADD_/c[285] ), .Z(
        \ADD_/FAINST[285].FA_/n1 ) );
  XOR \ADD_/FAINST[284].FA_/U5  ( .A(\ADD_/FAINST[284].FA_/n3 ), .B(
        \ADD_/c[284] ), .Z(\ADD_/c[285] ) );
  XOR \ADD_/FAINST[284].FA_/U4  ( .A(\ADD_/FAINST[284].FA_/n1 ), .B(b[284]), 
        .Z(c[284]) );
  AND \ADD_/FAINST[284].FA_/U3  ( .A(\ADD_/FAINST[284].FA_/n1 ), .B(
        \ADD_/FAINST[284].FA_/n2 ), .Z(\ADD_/FAINST[284].FA_/n3 ) );
  XOR \ADD_/FAINST[284].FA_/U2  ( .A(b[284]), .B(\ADD_/c[284] ), .Z(
        \ADD_/FAINST[284].FA_/n2 ) );
  XOR \ADD_/FAINST[284].FA_/U1  ( .A(a[284]), .B(\ADD_/c[284] ), .Z(
        \ADD_/FAINST[284].FA_/n1 ) );
  XOR \ADD_/FAINST[283].FA_/U5  ( .A(\ADD_/FAINST[283].FA_/n3 ), .B(
        \ADD_/c[283] ), .Z(\ADD_/c[284] ) );
  XOR \ADD_/FAINST[283].FA_/U4  ( .A(\ADD_/FAINST[283].FA_/n1 ), .B(b[283]), 
        .Z(c[283]) );
  AND \ADD_/FAINST[283].FA_/U3  ( .A(\ADD_/FAINST[283].FA_/n1 ), .B(
        \ADD_/FAINST[283].FA_/n2 ), .Z(\ADD_/FAINST[283].FA_/n3 ) );
  XOR \ADD_/FAINST[283].FA_/U2  ( .A(b[283]), .B(\ADD_/c[283] ), .Z(
        \ADD_/FAINST[283].FA_/n2 ) );
  XOR \ADD_/FAINST[283].FA_/U1  ( .A(a[283]), .B(\ADD_/c[283] ), .Z(
        \ADD_/FAINST[283].FA_/n1 ) );
  XOR \ADD_/FAINST[282].FA_/U5  ( .A(\ADD_/FAINST[282].FA_/n3 ), .B(
        \ADD_/c[282] ), .Z(\ADD_/c[283] ) );
  XOR \ADD_/FAINST[282].FA_/U4  ( .A(\ADD_/FAINST[282].FA_/n1 ), .B(b[282]), 
        .Z(c[282]) );
  AND \ADD_/FAINST[282].FA_/U3  ( .A(\ADD_/FAINST[282].FA_/n1 ), .B(
        \ADD_/FAINST[282].FA_/n2 ), .Z(\ADD_/FAINST[282].FA_/n3 ) );
  XOR \ADD_/FAINST[282].FA_/U2  ( .A(b[282]), .B(\ADD_/c[282] ), .Z(
        \ADD_/FAINST[282].FA_/n2 ) );
  XOR \ADD_/FAINST[282].FA_/U1  ( .A(a[282]), .B(\ADD_/c[282] ), .Z(
        \ADD_/FAINST[282].FA_/n1 ) );
  XOR \ADD_/FAINST[281].FA_/U5  ( .A(\ADD_/FAINST[281].FA_/n3 ), .B(
        \ADD_/c[281] ), .Z(\ADD_/c[282] ) );
  XOR \ADD_/FAINST[281].FA_/U4  ( .A(\ADD_/FAINST[281].FA_/n1 ), .B(b[281]), 
        .Z(c[281]) );
  AND \ADD_/FAINST[281].FA_/U3  ( .A(\ADD_/FAINST[281].FA_/n1 ), .B(
        \ADD_/FAINST[281].FA_/n2 ), .Z(\ADD_/FAINST[281].FA_/n3 ) );
  XOR \ADD_/FAINST[281].FA_/U2  ( .A(b[281]), .B(\ADD_/c[281] ), .Z(
        \ADD_/FAINST[281].FA_/n2 ) );
  XOR \ADD_/FAINST[281].FA_/U1  ( .A(a[281]), .B(\ADD_/c[281] ), .Z(
        \ADD_/FAINST[281].FA_/n1 ) );
  XOR \ADD_/FAINST[280].FA_/U5  ( .A(\ADD_/FAINST[280].FA_/n3 ), .B(
        \ADD_/c[280] ), .Z(\ADD_/c[281] ) );
  XOR \ADD_/FAINST[280].FA_/U4  ( .A(\ADD_/FAINST[280].FA_/n1 ), .B(b[280]), 
        .Z(c[280]) );
  AND \ADD_/FAINST[280].FA_/U3  ( .A(\ADD_/FAINST[280].FA_/n1 ), .B(
        \ADD_/FAINST[280].FA_/n2 ), .Z(\ADD_/FAINST[280].FA_/n3 ) );
  XOR \ADD_/FAINST[280].FA_/U2  ( .A(b[280]), .B(\ADD_/c[280] ), .Z(
        \ADD_/FAINST[280].FA_/n2 ) );
  XOR \ADD_/FAINST[280].FA_/U1  ( .A(a[280]), .B(\ADD_/c[280] ), .Z(
        \ADD_/FAINST[280].FA_/n1 ) );
  XOR \ADD_/FAINST[279].FA_/U5  ( .A(\ADD_/FAINST[279].FA_/n3 ), .B(
        \ADD_/c[279] ), .Z(\ADD_/c[280] ) );
  XOR \ADD_/FAINST[279].FA_/U4  ( .A(\ADD_/FAINST[279].FA_/n1 ), .B(b[279]), 
        .Z(c[279]) );
  AND \ADD_/FAINST[279].FA_/U3  ( .A(\ADD_/FAINST[279].FA_/n1 ), .B(
        \ADD_/FAINST[279].FA_/n2 ), .Z(\ADD_/FAINST[279].FA_/n3 ) );
  XOR \ADD_/FAINST[279].FA_/U2  ( .A(b[279]), .B(\ADD_/c[279] ), .Z(
        \ADD_/FAINST[279].FA_/n2 ) );
  XOR \ADD_/FAINST[279].FA_/U1  ( .A(a[279]), .B(\ADD_/c[279] ), .Z(
        \ADD_/FAINST[279].FA_/n1 ) );
  XOR \ADD_/FAINST[278].FA_/U5  ( .A(\ADD_/FAINST[278].FA_/n3 ), .B(
        \ADD_/c[278] ), .Z(\ADD_/c[279] ) );
  XOR \ADD_/FAINST[278].FA_/U4  ( .A(\ADD_/FAINST[278].FA_/n1 ), .B(b[278]), 
        .Z(c[278]) );
  AND \ADD_/FAINST[278].FA_/U3  ( .A(\ADD_/FAINST[278].FA_/n1 ), .B(
        \ADD_/FAINST[278].FA_/n2 ), .Z(\ADD_/FAINST[278].FA_/n3 ) );
  XOR \ADD_/FAINST[278].FA_/U2  ( .A(b[278]), .B(\ADD_/c[278] ), .Z(
        \ADD_/FAINST[278].FA_/n2 ) );
  XOR \ADD_/FAINST[278].FA_/U1  ( .A(a[278]), .B(\ADD_/c[278] ), .Z(
        \ADD_/FAINST[278].FA_/n1 ) );
  XOR \ADD_/FAINST[277].FA_/U5  ( .A(\ADD_/FAINST[277].FA_/n3 ), .B(
        \ADD_/c[277] ), .Z(\ADD_/c[278] ) );
  XOR \ADD_/FAINST[277].FA_/U4  ( .A(\ADD_/FAINST[277].FA_/n1 ), .B(b[277]), 
        .Z(c[277]) );
  AND \ADD_/FAINST[277].FA_/U3  ( .A(\ADD_/FAINST[277].FA_/n1 ), .B(
        \ADD_/FAINST[277].FA_/n2 ), .Z(\ADD_/FAINST[277].FA_/n3 ) );
  XOR \ADD_/FAINST[277].FA_/U2  ( .A(b[277]), .B(\ADD_/c[277] ), .Z(
        \ADD_/FAINST[277].FA_/n2 ) );
  XOR \ADD_/FAINST[277].FA_/U1  ( .A(a[277]), .B(\ADD_/c[277] ), .Z(
        \ADD_/FAINST[277].FA_/n1 ) );
  XOR \ADD_/FAINST[276].FA_/U5  ( .A(\ADD_/FAINST[276].FA_/n3 ), .B(
        \ADD_/c[276] ), .Z(\ADD_/c[277] ) );
  XOR \ADD_/FAINST[276].FA_/U4  ( .A(\ADD_/FAINST[276].FA_/n1 ), .B(b[276]), 
        .Z(c[276]) );
  AND \ADD_/FAINST[276].FA_/U3  ( .A(\ADD_/FAINST[276].FA_/n1 ), .B(
        \ADD_/FAINST[276].FA_/n2 ), .Z(\ADD_/FAINST[276].FA_/n3 ) );
  XOR \ADD_/FAINST[276].FA_/U2  ( .A(b[276]), .B(\ADD_/c[276] ), .Z(
        \ADD_/FAINST[276].FA_/n2 ) );
  XOR \ADD_/FAINST[276].FA_/U1  ( .A(a[276]), .B(\ADD_/c[276] ), .Z(
        \ADD_/FAINST[276].FA_/n1 ) );
  XOR \ADD_/FAINST[275].FA_/U5  ( .A(\ADD_/FAINST[275].FA_/n3 ), .B(
        \ADD_/c[275] ), .Z(\ADD_/c[276] ) );
  XOR \ADD_/FAINST[275].FA_/U4  ( .A(\ADD_/FAINST[275].FA_/n1 ), .B(b[275]), 
        .Z(c[275]) );
  AND \ADD_/FAINST[275].FA_/U3  ( .A(\ADD_/FAINST[275].FA_/n1 ), .B(
        \ADD_/FAINST[275].FA_/n2 ), .Z(\ADD_/FAINST[275].FA_/n3 ) );
  XOR \ADD_/FAINST[275].FA_/U2  ( .A(b[275]), .B(\ADD_/c[275] ), .Z(
        \ADD_/FAINST[275].FA_/n2 ) );
  XOR \ADD_/FAINST[275].FA_/U1  ( .A(a[275]), .B(\ADD_/c[275] ), .Z(
        \ADD_/FAINST[275].FA_/n1 ) );
  XOR \ADD_/FAINST[274].FA_/U5  ( .A(\ADD_/FAINST[274].FA_/n3 ), .B(
        \ADD_/c[274] ), .Z(\ADD_/c[275] ) );
  XOR \ADD_/FAINST[274].FA_/U4  ( .A(\ADD_/FAINST[274].FA_/n1 ), .B(b[274]), 
        .Z(c[274]) );
  AND \ADD_/FAINST[274].FA_/U3  ( .A(\ADD_/FAINST[274].FA_/n1 ), .B(
        \ADD_/FAINST[274].FA_/n2 ), .Z(\ADD_/FAINST[274].FA_/n3 ) );
  XOR \ADD_/FAINST[274].FA_/U2  ( .A(b[274]), .B(\ADD_/c[274] ), .Z(
        \ADD_/FAINST[274].FA_/n2 ) );
  XOR \ADD_/FAINST[274].FA_/U1  ( .A(a[274]), .B(\ADD_/c[274] ), .Z(
        \ADD_/FAINST[274].FA_/n1 ) );
  XOR \ADD_/FAINST[273].FA_/U5  ( .A(\ADD_/FAINST[273].FA_/n3 ), .B(
        \ADD_/c[273] ), .Z(\ADD_/c[274] ) );
  XOR \ADD_/FAINST[273].FA_/U4  ( .A(\ADD_/FAINST[273].FA_/n1 ), .B(b[273]), 
        .Z(c[273]) );
  AND \ADD_/FAINST[273].FA_/U3  ( .A(\ADD_/FAINST[273].FA_/n1 ), .B(
        \ADD_/FAINST[273].FA_/n2 ), .Z(\ADD_/FAINST[273].FA_/n3 ) );
  XOR \ADD_/FAINST[273].FA_/U2  ( .A(b[273]), .B(\ADD_/c[273] ), .Z(
        \ADD_/FAINST[273].FA_/n2 ) );
  XOR \ADD_/FAINST[273].FA_/U1  ( .A(a[273]), .B(\ADD_/c[273] ), .Z(
        \ADD_/FAINST[273].FA_/n1 ) );
  XOR \ADD_/FAINST[272].FA_/U5  ( .A(\ADD_/FAINST[272].FA_/n3 ), .B(
        \ADD_/c[272] ), .Z(\ADD_/c[273] ) );
  XOR \ADD_/FAINST[272].FA_/U4  ( .A(\ADD_/FAINST[272].FA_/n1 ), .B(b[272]), 
        .Z(c[272]) );
  AND \ADD_/FAINST[272].FA_/U3  ( .A(\ADD_/FAINST[272].FA_/n1 ), .B(
        \ADD_/FAINST[272].FA_/n2 ), .Z(\ADD_/FAINST[272].FA_/n3 ) );
  XOR \ADD_/FAINST[272].FA_/U2  ( .A(b[272]), .B(\ADD_/c[272] ), .Z(
        \ADD_/FAINST[272].FA_/n2 ) );
  XOR \ADD_/FAINST[272].FA_/U1  ( .A(a[272]), .B(\ADD_/c[272] ), .Z(
        \ADD_/FAINST[272].FA_/n1 ) );
  XOR \ADD_/FAINST[271].FA_/U5  ( .A(\ADD_/FAINST[271].FA_/n3 ), .B(
        \ADD_/c[271] ), .Z(\ADD_/c[272] ) );
  XOR \ADD_/FAINST[271].FA_/U4  ( .A(\ADD_/FAINST[271].FA_/n1 ), .B(b[271]), 
        .Z(c[271]) );
  AND \ADD_/FAINST[271].FA_/U3  ( .A(\ADD_/FAINST[271].FA_/n1 ), .B(
        \ADD_/FAINST[271].FA_/n2 ), .Z(\ADD_/FAINST[271].FA_/n3 ) );
  XOR \ADD_/FAINST[271].FA_/U2  ( .A(b[271]), .B(\ADD_/c[271] ), .Z(
        \ADD_/FAINST[271].FA_/n2 ) );
  XOR \ADD_/FAINST[271].FA_/U1  ( .A(a[271]), .B(\ADD_/c[271] ), .Z(
        \ADD_/FAINST[271].FA_/n1 ) );
  XOR \ADD_/FAINST[270].FA_/U5  ( .A(\ADD_/FAINST[270].FA_/n3 ), .B(
        \ADD_/c[270] ), .Z(\ADD_/c[271] ) );
  XOR \ADD_/FAINST[270].FA_/U4  ( .A(\ADD_/FAINST[270].FA_/n1 ), .B(b[270]), 
        .Z(c[270]) );
  AND \ADD_/FAINST[270].FA_/U3  ( .A(\ADD_/FAINST[270].FA_/n1 ), .B(
        \ADD_/FAINST[270].FA_/n2 ), .Z(\ADD_/FAINST[270].FA_/n3 ) );
  XOR \ADD_/FAINST[270].FA_/U2  ( .A(b[270]), .B(\ADD_/c[270] ), .Z(
        \ADD_/FAINST[270].FA_/n2 ) );
  XOR \ADD_/FAINST[270].FA_/U1  ( .A(a[270]), .B(\ADD_/c[270] ), .Z(
        \ADD_/FAINST[270].FA_/n1 ) );
  XOR \ADD_/FAINST[269].FA_/U5  ( .A(\ADD_/FAINST[269].FA_/n3 ), .B(
        \ADD_/c[269] ), .Z(\ADD_/c[270] ) );
  XOR \ADD_/FAINST[269].FA_/U4  ( .A(\ADD_/FAINST[269].FA_/n1 ), .B(b[269]), 
        .Z(c[269]) );
  AND \ADD_/FAINST[269].FA_/U3  ( .A(\ADD_/FAINST[269].FA_/n1 ), .B(
        \ADD_/FAINST[269].FA_/n2 ), .Z(\ADD_/FAINST[269].FA_/n3 ) );
  XOR \ADD_/FAINST[269].FA_/U2  ( .A(b[269]), .B(\ADD_/c[269] ), .Z(
        \ADD_/FAINST[269].FA_/n2 ) );
  XOR \ADD_/FAINST[269].FA_/U1  ( .A(a[269]), .B(\ADD_/c[269] ), .Z(
        \ADD_/FAINST[269].FA_/n1 ) );
  XOR \ADD_/FAINST[268].FA_/U5  ( .A(\ADD_/FAINST[268].FA_/n3 ), .B(
        \ADD_/c[268] ), .Z(\ADD_/c[269] ) );
  XOR \ADD_/FAINST[268].FA_/U4  ( .A(\ADD_/FAINST[268].FA_/n1 ), .B(b[268]), 
        .Z(c[268]) );
  AND \ADD_/FAINST[268].FA_/U3  ( .A(\ADD_/FAINST[268].FA_/n1 ), .B(
        \ADD_/FAINST[268].FA_/n2 ), .Z(\ADD_/FAINST[268].FA_/n3 ) );
  XOR \ADD_/FAINST[268].FA_/U2  ( .A(b[268]), .B(\ADD_/c[268] ), .Z(
        \ADD_/FAINST[268].FA_/n2 ) );
  XOR \ADD_/FAINST[268].FA_/U1  ( .A(a[268]), .B(\ADD_/c[268] ), .Z(
        \ADD_/FAINST[268].FA_/n1 ) );
  XOR \ADD_/FAINST[267].FA_/U5  ( .A(\ADD_/FAINST[267].FA_/n3 ), .B(
        \ADD_/c[267] ), .Z(\ADD_/c[268] ) );
  XOR \ADD_/FAINST[267].FA_/U4  ( .A(\ADD_/FAINST[267].FA_/n1 ), .B(b[267]), 
        .Z(c[267]) );
  AND \ADD_/FAINST[267].FA_/U3  ( .A(\ADD_/FAINST[267].FA_/n1 ), .B(
        \ADD_/FAINST[267].FA_/n2 ), .Z(\ADD_/FAINST[267].FA_/n3 ) );
  XOR \ADD_/FAINST[267].FA_/U2  ( .A(b[267]), .B(\ADD_/c[267] ), .Z(
        \ADD_/FAINST[267].FA_/n2 ) );
  XOR \ADD_/FAINST[267].FA_/U1  ( .A(a[267]), .B(\ADD_/c[267] ), .Z(
        \ADD_/FAINST[267].FA_/n1 ) );
  XOR \ADD_/FAINST[266].FA_/U5  ( .A(\ADD_/FAINST[266].FA_/n3 ), .B(
        \ADD_/c[266] ), .Z(\ADD_/c[267] ) );
  XOR \ADD_/FAINST[266].FA_/U4  ( .A(\ADD_/FAINST[266].FA_/n1 ), .B(b[266]), 
        .Z(c[266]) );
  AND \ADD_/FAINST[266].FA_/U3  ( .A(\ADD_/FAINST[266].FA_/n1 ), .B(
        \ADD_/FAINST[266].FA_/n2 ), .Z(\ADD_/FAINST[266].FA_/n3 ) );
  XOR \ADD_/FAINST[266].FA_/U2  ( .A(b[266]), .B(\ADD_/c[266] ), .Z(
        \ADD_/FAINST[266].FA_/n2 ) );
  XOR \ADD_/FAINST[266].FA_/U1  ( .A(a[266]), .B(\ADD_/c[266] ), .Z(
        \ADD_/FAINST[266].FA_/n1 ) );
  XOR \ADD_/FAINST[265].FA_/U5  ( .A(\ADD_/FAINST[265].FA_/n3 ), .B(
        \ADD_/c[265] ), .Z(\ADD_/c[266] ) );
  XOR \ADD_/FAINST[265].FA_/U4  ( .A(\ADD_/FAINST[265].FA_/n1 ), .B(b[265]), 
        .Z(c[265]) );
  AND \ADD_/FAINST[265].FA_/U3  ( .A(\ADD_/FAINST[265].FA_/n1 ), .B(
        \ADD_/FAINST[265].FA_/n2 ), .Z(\ADD_/FAINST[265].FA_/n3 ) );
  XOR \ADD_/FAINST[265].FA_/U2  ( .A(b[265]), .B(\ADD_/c[265] ), .Z(
        \ADD_/FAINST[265].FA_/n2 ) );
  XOR \ADD_/FAINST[265].FA_/U1  ( .A(a[265]), .B(\ADD_/c[265] ), .Z(
        \ADD_/FAINST[265].FA_/n1 ) );
  XOR \ADD_/FAINST[264].FA_/U5  ( .A(\ADD_/FAINST[264].FA_/n3 ), .B(
        \ADD_/c[264] ), .Z(\ADD_/c[265] ) );
  XOR \ADD_/FAINST[264].FA_/U4  ( .A(\ADD_/FAINST[264].FA_/n1 ), .B(b[264]), 
        .Z(c[264]) );
  AND \ADD_/FAINST[264].FA_/U3  ( .A(\ADD_/FAINST[264].FA_/n1 ), .B(
        \ADD_/FAINST[264].FA_/n2 ), .Z(\ADD_/FAINST[264].FA_/n3 ) );
  XOR \ADD_/FAINST[264].FA_/U2  ( .A(b[264]), .B(\ADD_/c[264] ), .Z(
        \ADD_/FAINST[264].FA_/n2 ) );
  XOR \ADD_/FAINST[264].FA_/U1  ( .A(a[264]), .B(\ADD_/c[264] ), .Z(
        \ADD_/FAINST[264].FA_/n1 ) );
  XOR \ADD_/FAINST[263].FA_/U5  ( .A(\ADD_/FAINST[263].FA_/n3 ), .B(
        \ADD_/c[263] ), .Z(\ADD_/c[264] ) );
  XOR \ADD_/FAINST[263].FA_/U4  ( .A(\ADD_/FAINST[263].FA_/n1 ), .B(b[263]), 
        .Z(c[263]) );
  AND \ADD_/FAINST[263].FA_/U3  ( .A(\ADD_/FAINST[263].FA_/n1 ), .B(
        \ADD_/FAINST[263].FA_/n2 ), .Z(\ADD_/FAINST[263].FA_/n3 ) );
  XOR \ADD_/FAINST[263].FA_/U2  ( .A(b[263]), .B(\ADD_/c[263] ), .Z(
        \ADD_/FAINST[263].FA_/n2 ) );
  XOR \ADD_/FAINST[263].FA_/U1  ( .A(a[263]), .B(\ADD_/c[263] ), .Z(
        \ADD_/FAINST[263].FA_/n1 ) );
  XOR \ADD_/FAINST[262].FA_/U5  ( .A(\ADD_/FAINST[262].FA_/n3 ), .B(
        \ADD_/c[262] ), .Z(\ADD_/c[263] ) );
  XOR \ADD_/FAINST[262].FA_/U4  ( .A(\ADD_/FAINST[262].FA_/n1 ), .B(b[262]), 
        .Z(c[262]) );
  AND \ADD_/FAINST[262].FA_/U3  ( .A(\ADD_/FAINST[262].FA_/n1 ), .B(
        \ADD_/FAINST[262].FA_/n2 ), .Z(\ADD_/FAINST[262].FA_/n3 ) );
  XOR \ADD_/FAINST[262].FA_/U2  ( .A(b[262]), .B(\ADD_/c[262] ), .Z(
        \ADD_/FAINST[262].FA_/n2 ) );
  XOR \ADD_/FAINST[262].FA_/U1  ( .A(a[262]), .B(\ADD_/c[262] ), .Z(
        \ADD_/FAINST[262].FA_/n1 ) );
  XOR \ADD_/FAINST[261].FA_/U5  ( .A(\ADD_/FAINST[261].FA_/n3 ), .B(
        \ADD_/c[261] ), .Z(\ADD_/c[262] ) );
  XOR \ADD_/FAINST[261].FA_/U4  ( .A(\ADD_/FAINST[261].FA_/n1 ), .B(b[261]), 
        .Z(c[261]) );
  AND \ADD_/FAINST[261].FA_/U3  ( .A(\ADD_/FAINST[261].FA_/n1 ), .B(
        \ADD_/FAINST[261].FA_/n2 ), .Z(\ADD_/FAINST[261].FA_/n3 ) );
  XOR \ADD_/FAINST[261].FA_/U2  ( .A(b[261]), .B(\ADD_/c[261] ), .Z(
        \ADD_/FAINST[261].FA_/n2 ) );
  XOR \ADD_/FAINST[261].FA_/U1  ( .A(a[261]), .B(\ADD_/c[261] ), .Z(
        \ADD_/FAINST[261].FA_/n1 ) );
  XOR \ADD_/FAINST[260].FA_/U5  ( .A(\ADD_/FAINST[260].FA_/n3 ), .B(
        \ADD_/c[260] ), .Z(\ADD_/c[261] ) );
  XOR \ADD_/FAINST[260].FA_/U4  ( .A(\ADD_/FAINST[260].FA_/n1 ), .B(b[260]), 
        .Z(c[260]) );
  AND \ADD_/FAINST[260].FA_/U3  ( .A(\ADD_/FAINST[260].FA_/n1 ), .B(
        \ADD_/FAINST[260].FA_/n2 ), .Z(\ADD_/FAINST[260].FA_/n3 ) );
  XOR \ADD_/FAINST[260].FA_/U2  ( .A(b[260]), .B(\ADD_/c[260] ), .Z(
        \ADD_/FAINST[260].FA_/n2 ) );
  XOR \ADD_/FAINST[260].FA_/U1  ( .A(a[260]), .B(\ADD_/c[260] ), .Z(
        \ADD_/FAINST[260].FA_/n1 ) );
  XOR \ADD_/FAINST[259].FA_/U5  ( .A(\ADD_/FAINST[259].FA_/n3 ), .B(
        \ADD_/c[259] ), .Z(\ADD_/c[260] ) );
  XOR \ADD_/FAINST[259].FA_/U4  ( .A(\ADD_/FAINST[259].FA_/n1 ), .B(b[259]), 
        .Z(c[259]) );
  AND \ADD_/FAINST[259].FA_/U3  ( .A(\ADD_/FAINST[259].FA_/n1 ), .B(
        \ADD_/FAINST[259].FA_/n2 ), .Z(\ADD_/FAINST[259].FA_/n3 ) );
  XOR \ADD_/FAINST[259].FA_/U2  ( .A(b[259]), .B(\ADD_/c[259] ), .Z(
        \ADD_/FAINST[259].FA_/n2 ) );
  XOR \ADD_/FAINST[259].FA_/U1  ( .A(a[259]), .B(\ADD_/c[259] ), .Z(
        \ADD_/FAINST[259].FA_/n1 ) );
  XOR \ADD_/FAINST[258].FA_/U5  ( .A(\ADD_/FAINST[258].FA_/n3 ), .B(
        \ADD_/c[258] ), .Z(\ADD_/c[259] ) );
  XOR \ADD_/FAINST[258].FA_/U4  ( .A(\ADD_/FAINST[258].FA_/n1 ), .B(b[258]), 
        .Z(c[258]) );
  AND \ADD_/FAINST[258].FA_/U3  ( .A(\ADD_/FAINST[258].FA_/n1 ), .B(
        \ADD_/FAINST[258].FA_/n2 ), .Z(\ADD_/FAINST[258].FA_/n3 ) );
  XOR \ADD_/FAINST[258].FA_/U2  ( .A(b[258]), .B(\ADD_/c[258] ), .Z(
        \ADD_/FAINST[258].FA_/n2 ) );
  XOR \ADD_/FAINST[258].FA_/U1  ( .A(a[258]), .B(\ADD_/c[258] ), .Z(
        \ADD_/FAINST[258].FA_/n1 ) );
  XOR \ADD_/FAINST[257].FA_/U5  ( .A(\ADD_/FAINST[257].FA_/n3 ), .B(
        \ADD_/c[257] ), .Z(\ADD_/c[258] ) );
  XOR \ADD_/FAINST[257].FA_/U4  ( .A(\ADD_/FAINST[257].FA_/n1 ), .B(b[257]), 
        .Z(c[257]) );
  AND \ADD_/FAINST[257].FA_/U3  ( .A(\ADD_/FAINST[257].FA_/n1 ), .B(
        \ADD_/FAINST[257].FA_/n2 ), .Z(\ADD_/FAINST[257].FA_/n3 ) );
  XOR \ADD_/FAINST[257].FA_/U2  ( .A(b[257]), .B(\ADD_/c[257] ), .Z(
        \ADD_/FAINST[257].FA_/n2 ) );
  XOR \ADD_/FAINST[257].FA_/U1  ( .A(a[257]), .B(\ADD_/c[257] ), .Z(
        \ADD_/FAINST[257].FA_/n1 ) );
  XOR \ADD_/FAINST[256].FA_/U5  ( .A(\ADD_/FAINST[256].FA_/n3 ), .B(
        \ADD_/c[256] ), .Z(\ADD_/c[257] ) );
  XOR \ADD_/FAINST[256].FA_/U4  ( .A(\ADD_/FAINST[256].FA_/n1 ), .B(b[256]), 
        .Z(c[256]) );
  AND \ADD_/FAINST[256].FA_/U3  ( .A(\ADD_/FAINST[256].FA_/n1 ), .B(
        \ADD_/FAINST[256].FA_/n2 ), .Z(\ADD_/FAINST[256].FA_/n3 ) );
  XOR \ADD_/FAINST[256].FA_/U2  ( .A(b[256]), .B(\ADD_/c[256] ), .Z(
        \ADD_/FAINST[256].FA_/n2 ) );
  XOR \ADD_/FAINST[256].FA_/U1  ( .A(a[256]), .B(\ADD_/c[256] ), .Z(
        \ADD_/FAINST[256].FA_/n1 ) );
  XOR \ADD_/FAINST[255].FA_/U5  ( .A(\ADD_/FAINST[255].FA_/n3 ), .B(
        \ADD_/c[255] ), .Z(\ADD_/c[256] ) );
  XOR \ADD_/FAINST[255].FA_/U4  ( .A(\ADD_/FAINST[255].FA_/n1 ), .B(b[255]), 
        .Z(c[255]) );
  AND \ADD_/FAINST[255].FA_/U3  ( .A(\ADD_/FAINST[255].FA_/n1 ), .B(
        \ADD_/FAINST[255].FA_/n2 ), .Z(\ADD_/FAINST[255].FA_/n3 ) );
  XOR \ADD_/FAINST[255].FA_/U2  ( .A(b[255]), .B(\ADD_/c[255] ), .Z(
        \ADD_/FAINST[255].FA_/n2 ) );
  XOR \ADD_/FAINST[255].FA_/U1  ( .A(a[255]), .B(\ADD_/c[255] ), .Z(
        \ADD_/FAINST[255].FA_/n1 ) );
  XOR \ADD_/FAINST[254].FA_/U5  ( .A(\ADD_/FAINST[254].FA_/n3 ), .B(
        \ADD_/c[254] ), .Z(\ADD_/c[255] ) );
  XOR \ADD_/FAINST[254].FA_/U4  ( .A(\ADD_/FAINST[254].FA_/n1 ), .B(b[254]), 
        .Z(c[254]) );
  AND \ADD_/FAINST[254].FA_/U3  ( .A(\ADD_/FAINST[254].FA_/n1 ), .B(
        \ADD_/FAINST[254].FA_/n2 ), .Z(\ADD_/FAINST[254].FA_/n3 ) );
  XOR \ADD_/FAINST[254].FA_/U2  ( .A(b[254]), .B(\ADD_/c[254] ), .Z(
        \ADD_/FAINST[254].FA_/n2 ) );
  XOR \ADD_/FAINST[254].FA_/U1  ( .A(a[254]), .B(\ADD_/c[254] ), .Z(
        \ADD_/FAINST[254].FA_/n1 ) );
  XOR \ADD_/FAINST[253].FA_/U5  ( .A(\ADD_/FAINST[253].FA_/n3 ), .B(
        \ADD_/c[253] ), .Z(\ADD_/c[254] ) );
  XOR \ADD_/FAINST[253].FA_/U4  ( .A(\ADD_/FAINST[253].FA_/n1 ), .B(b[253]), 
        .Z(c[253]) );
  AND \ADD_/FAINST[253].FA_/U3  ( .A(\ADD_/FAINST[253].FA_/n1 ), .B(
        \ADD_/FAINST[253].FA_/n2 ), .Z(\ADD_/FAINST[253].FA_/n3 ) );
  XOR \ADD_/FAINST[253].FA_/U2  ( .A(b[253]), .B(\ADD_/c[253] ), .Z(
        \ADD_/FAINST[253].FA_/n2 ) );
  XOR \ADD_/FAINST[253].FA_/U1  ( .A(a[253]), .B(\ADD_/c[253] ), .Z(
        \ADD_/FAINST[253].FA_/n1 ) );
  XOR \ADD_/FAINST[252].FA_/U5  ( .A(\ADD_/FAINST[252].FA_/n3 ), .B(
        \ADD_/c[252] ), .Z(\ADD_/c[253] ) );
  XOR \ADD_/FAINST[252].FA_/U4  ( .A(\ADD_/FAINST[252].FA_/n1 ), .B(b[252]), 
        .Z(c[252]) );
  AND \ADD_/FAINST[252].FA_/U3  ( .A(\ADD_/FAINST[252].FA_/n1 ), .B(
        \ADD_/FAINST[252].FA_/n2 ), .Z(\ADD_/FAINST[252].FA_/n3 ) );
  XOR \ADD_/FAINST[252].FA_/U2  ( .A(b[252]), .B(\ADD_/c[252] ), .Z(
        \ADD_/FAINST[252].FA_/n2 ) );
  XOR \ADD_/FAINST[252].FA_/U1  ( .A(a[252]), .B(\ADD_/c[252] ), .Z(
        \ADD_/FAINST[252].FA_/n1 ) );
  XOR \ADD_/FAINST[251].FA_/U5  ( .A(\ADD_/FAINST[251].FA_/n3 ), .B(
        \ADD_/c[251] ), .Z(\ADD_/c[252] ) );
  XOR \ADD_/FAINST[251].FA_/U4  ( .A(\ADD_/FAINST[251].FA_/n1 ), .B(b[251]), 
        .Z(c[251]) );
  AND \ADD_/FAINST[251].FA_/U3  ( .A(\ADD_/FAINST[251].FA_/n1 ), .B(
        \ADD_/FAINST[251].FA_/n2 ), .Z(\ADD_/FAINST[251].FA_/n3 ) );
  XOR \ADD_/FAINST[251].FA_/U2  ( .A(b[251]), .B(\ADD_/c[251] ), .Z(
        \ADD_/FAINST[251].FA_/n2 ) );
  XOR \ADD_/FAINST[251].FA_/U1  ( .A(a[251]), .B(\ADD_/c[251] ), .Z(
        \ADD_/FAINST[251].FA_/n1 ) );
  XOR \ADD_/FAINST[250].FA_/U5  ( .A(\ADD_/FAINST[250].FA_/n3 ), .B(
        \ADD_/c[250] ), .Z(\ADD_/c[251] ) );
  XOR \ADD_/FAINST[250].FA_/U4  ( .A(\ADD_/FAINST[250].FA_/n1 ), .B(b[250]), 
        .Z(c[250]) );
  AND \ADD_/FAINST[250].FA_/U3  ( .A(\ADD_/FAINST[250].FA_/n1 ), .B(
        \ADD_/FAINST[250].FA_/n2 ), .Z(\ADD_/FAINST[250].FA_/n3 ) );
  XOR \ADD_/FAINST[250].FA_/U2  ( .A(b[250]), .B(\ADD_/c[250] ), .Z(
        \ADD_/FAINST[250].FA_/n2 ) );
  XOR \ADD_/FAINST[250].FA_/U1  ( .A(a[250]), .B(\ADD_/c[250] ), .Z(
        \ADD_/FAINST[250].FA_/n1 ) );
  XOR \ADD_/FAINST[249].FA_/U5  ( .A(\ADD_/FAINST[249].FA_/n3 ), .B(
        \ADD_/c[249] ), .Z(\ADD_/c[250] ) );
  XOR \ADD_/FAINST[249].FA_/U4  ( .A(\ADD_/FAINST[249].FA_/n1 ), .B(b[249]), 
        .Z(c[249]) );
  AND \ADD_/FAINST[249].FA_/U3  ( .A(\ADD_/FAINST[249].FA_/n1 ), .B(
        \ADD_/FAINST[249].FA_/n2 ), .Z(\ADD_/FAINST[249].FA_/n3 ) );
  XOR \ADD_/FAINST[249].FA_/U2  ( .A(b[249]), .B(\ADD_/c[249] ), .Z(
        \ADD_/FAINST[249].FA_/n2 ) );
  XOR \ADD_/FAINST[249].FA_/U1  ( .A(a[249]), .B(\ADD_/c[249] ), .Z(
        \ADD_/FAINST[249].FA_/n1 ) );
  XOR \ADD_/FAINST[248].FA_/U5  ( .A(\ADD_/FAINST[248].FA_/n3 ), .B(
        \ADD_/c[248] ), .Z(\ADD_/c[249] ) );
  XOR \ADD_/FAINST[248].FA_/U4  ( .A(\ADD_/FAINST[248].FA_/n1 ), .B(b[248]), 
        .Z(c[248]) );
  AND \ADD_/FAINST[248].FA_/U3  ( .A(\ADD_/FAINST[248].FA_/n1 ), .B(
        \ADD_/FAINST[248].FA_/n2 ), .Z(\ADD_/FAINST[248].FA_/n3 ) );
  XOR \ADD_/FAINST[248].FA_/U2  ( .A(b[248]), .B(\ADD_/c[248] ), .Z(
        \ADD_/FAINST[248].FA_/n2 ) );
  XOR \ADD_/FAINST[248].FA_/U1  ( .A(a[248]), .B(\ADD_/c[248] ), .Z(
        \ADD_/FAINST[248].FA_/n1 ) );
  XOR \ADD_/FAINST[247].FA_/U5  ( .A(\ADD_/FAINST[247].FA_/n3 ), .B(
        \ADD_/c[247] ), .Z(\ADD_/c[248] ) );
  XOR \ADD_/FAINST[247].FA_/U4  ( .A(\ADD_/FAINST[247].FA_/n1 ), .B(b[247]), 
        .Z(c[247]) );
  AND \ADD_/FAINST[247].FA_/U3  ( .A(\ADD_/FAINST[247].FA_/n1 ), .B(
        \ADD_/FAINST[247].FA_/n2 ), .Z(\ADD_/FAINST[247].FA_/n3 ) );
  XOR \ADD_/FAINST[247].FA_/U2  ( .A(b[247]), .B(\ADD_/c[247] ), .Z(
        \ADD_/FAINST[247].FA_/n2 ) );
  XOR \ADD_/FAINST[247].FA_/U1  ( .A(a[247]), .B(\ADD_/c[247] ), .Z(
        \ADD_/FAINST[247].FA_/n1 ) );
  XOR \ADD_/FAINST[246].FA_/U5  ( .A(\ADD_/FAINST[246].FA_/n3 ), .B(
        \ADD_/c[246] ), .Z(\ADD_/c[247] ) );
  XOR \ADD_/FAINST[246].FA_/U4  ( .A(\ADD_/FAINST[246].FA_/n1 ), .B(b[246]), 
        .Z(c[246]) );
  AND \ADD_/FAINST[246].FA_/U3  ( .A(\ADD_/FAINST[246].FA_/n1 ), .B(
        \ADD_/FAINST[246].FA_/n2 ), .Z(\ADD_/FAINST[246].FA_/n3 ) );
  XOR \ADD_/FAINST[246].FA_/U2  ( .A(b[246]), .B(\ADD_/c[246] ), .Z(
        \ADD_/FAINST[246].FA_/n2 ) );
  XOR \ADD_/FAINST[246].FA_/U1  ( .A(a[246]), .B(\ADD_/c[246] ), .Z(
        \ADD_/FAINST[246].FA_/n1 ) );
  XOR \ADD_/FAINST[245].FA_/U5  ( .A(\ADD_/FAINST[245].FA_/n3 ), .B(
        \ADD_/c[245] ), .Z(\ADD_/c[246] ) );
  XOR \ADD_/FAINST[245].FA_/U4  ( .A(\ADD_/FAINST[245].FA_/n1 ), .B(b[245]), 
        .Z(c[245]) );
  AND \ADD_/FAINST[245].FA_/U3  ( .A(\ADD_/FAINST[245].FA_/n1 ), .B(
        \ADD_/FAINST[245].FA_/n2 ), .Z(\ADD_/FAINST[245].FA_/n3 ) );
  XOR \ADD_/FAINST[245].FA_/U2  ( .A(b[245]), .B(\ADD_/c[245] ), .Z(
        \ADD_/FAINST[245].FA_/n2 ) );
  XOR \ADD_/FAINST[245].FA_/U1  ( .A(a[245]), .B(\ADD_/c[245] ), .Z(
        \ADD_/FAINST[245].FA_/n1 ) );
  XOR \ADD_/FAINST[244].FA_/U5  ( .A(\ADD_/FAINST[244].FA_/n3 ), .B(
        \ADD_/c[244] ), .Z(\ADD_/c[245] ) );
  XOR \ADD_/FAINST[244].FA_/U4  ( .A(\ADD_/FAINST[244].FA_/n1 ), .B(b[244]), 
        .Z(c[244]) );
  AND \ADD_/FAINST[244].FA_/U3  ( .A(\ADD_/FAINST[244].FA_/n1 ), .B(
        \ADD_/FAINST[244].FA_/n2 ), .Z(\ADD_/FAINST[244].FA_/n3 ) );
  XOR \ADD_/FAINST[244].FA_/U2  ( .A(b[244]), .B(\ADD_/c[244] ), .Z(
        \ADD_/FAINST[244].FA_/n2 ) );
  XOR \ADD_/FAINST[244].FA_/U1  ( .A(a[244]), .B(\ADD_/c[244] ), .Z(
        \ADD_/FAINST[244].FA_/n1 ) );
  XOR \ADD_/FAINST[243].FA_/U5  ( .A(\ADD_/FAINST[243].FA_/n3 ), .B(
        \ADD_/c[243] ), .Z(\ADD_/c[244] ) );
  XOR \ADD_/FAINST[243].FA_/U4  ( .A(\ADD_/FAINST[243].FA_/n1 ), .B(b[243]), 
        .Z(c[243]) );
  AND \ADD_/FAINST[243].FA_/U3  ( .A(\ADD_/FAINST[243].FA_/n1 ), .B(
        \ADD_/FAINST[243].FA_/n2 ), .Z(\ADD_/FAINST[243].FA_/n3 ) );
  XOR \ADD_/FAINST[243].FA_/U2  ( .A(b[243]), .B(\ADD_/c[243] ), .Z(
        \ADD_/FAINST[243].FA_/n2 ) );
  XOR \ADD_/FAINST[243].FA_/U1  ( .A(a[243]), .B(\ADD_/c[243] ), .Z(
        \ADD_/FAINST[243].FA_/n1 ) );
  XOR \ADD_/FAINST[242].FA_/U5  ( .A(\ADD_/FAINST[242].FA_/n3 ), .B(
        \ADD_/c[242] ), .Z(\ADD_/c[243] ) );
  XOR \ADD_/FAINST[242].FA_/U4  ( .A(\ADD_/FAINST[242].FA_/n1 ), .B(b[242]), 
        .Z(c[242]) );
  AND \ADD_/FAINST[242].FA_/U3  ( .A(\ADD_/FAINST[242].FA_/n1 ), .B(
        \ADD_/FAINST[242].FA_/n2 ), .Z(\ADD_/FAINST[242].FA_/n3 ) );
  XOR \ADD_/FAINST[242].FA_/U2  ( .A(b[242]), .B(\ADD_/c[242] ), .Z(
        \ADD_/FAINST[242].FA_/n2 ) );
  XOR \ADD_/FAINST[242].FA_/U1  ( .A(a[242]), .B(\ADD_/c[242] ), .Z(
        \ADD_/FAINST[242].FA_/n1 ) );
  XOR \ADD_/FAINST[241].FA_/U5  ( .A(\ADD_/FAINST[241].FA_/n3 ), .B(
        \ADD_/c[241] ), .Z(\ADD_/c[242] ) );
  XOR \ADD_/FAINST[241].FA_/U4  ( .A(\ADD_/FAINST[241].FA_/n1 ), .B(b[241]), 
        .Z(c[241]) );
  AND \ADD_/FAINST[241].FA_/U3  ( .A(\ADD_/FAINST[241].FA_/n1 ), .B(
        \ADD_/FAINST[241].FA_/n2 ), .Z(\ADD_/FAINST[241].FA_/n3 ) );
  XOR \ADD_/FAINST[241].FA_/U2  ( .A(b[241]), .B(\ADD_/c[241] ), .Z(
        \ADD_/FAINST[241].FA_/n2 ) );
  XOR \ADD_/FAINST[241].FA_/U1  ( .A(a[241]), .B(\ADD_/c[241] ), .Z(
        \ADD_/FAINST[241].FA_/n1 ) );
  XOR \ADD_/FAINST[240].FA_/U5  ( .A(\ADD_/FAINST[240].FA_/n3 ), .B(
        \ADD_/c[240] ), .Z(\ADD_/c[241] ) );
  XOR \ADD_/FAINST[240].FA_/U4  ( .A(\ADD_/FAINST[240].FA_/n1 ), .B(b[240]), 
        .Z(c[240]) );
  AND \ADD_/FAINST[240].FA_/U3  ( .A(\ADD_/FAINST[240].FA_/n1 ), .B(
        \ADD_/FAINST[240].FA_/n2 ), .Z(\ADD_/FAINST[240].FA_/n3 ) );
  XOR \ADD_/FAINST[240].FA_/U2  ( .A(b[240]), .B(\ADD_/c[240] ), .Z(
        \ADD_/FAINST[240].FA_/n2 ) );
  XOR \ADD_/FAINST[240].FA_/U1  ( .A(a[240]), .B(\ADD_/c[240] ), .Z(
        \ADD_/FAINST[240].FA_/n1 ) );
  XOR \ADD_/FAINST[239].FA_/U5  ( .A(\ADD_/FAINST[239].FA_/n3 ), .B(
        \ADD_/c[239] ), .Z(\ADD_/c[240] ) );
  XOR \ADD_/FAINST[239].FA_/U4  ( .A(\ADD_/FAINST[239].FA_/n1 ), .B(b[239]), 
        .Z(c[239]) );
  AND \ADD_/FAINST[239].FA_/U3  ( .A(\ADD_/FAINST[239].FA_/n1 ), .B(
        \ADD_/FAINST[239].FA_/n2 ), .Z(\ADD_/FAINST[239].FA_/n3 ) );
  XOR \ADD_/FAINST[239].FA_/U2  ( .A(b[239]), .B(\ADD_/c[239] ), .Z(
        \ADD_/FAINST[239].FA_/n2 ) );
  XOR \ADD_/FAINST[239].FA_/U1  ( .A(a[239]), .B(\ADD_/c[239] ), .Z(
        \ADD_/FAINST[239].FA_/n1 ) );
  XOR \ADD_/FAINST[238].FA_/U5  ( .A(\ADD_/FAINST[238].FA_/n3 ), .B(
        \ADD_/c[238] ), .Z(\ADD_/c[239] ) );
  XOR \ADD_/FAINST[238].FA_/U4  ( .A(\ADD_/FAINST[238].FA_/n1 ), .B(b[238]), 
        .Z(c[238]) );
  AND \ADD_/FAINST[238].FA_/U3  ( .A(\ADD_/FAINST[238].FA_/n1 ), .B(
        \ADD_/FAINST[238].FA_/n2 ), .Z(\ADD_/FAINST[238].FA_/n3 ) );
  XOR \ADD_/FAINST[238].FA_/U2  ( .A(b[238]), .B(\ADD_/c[238] ), .Z(
        \ADD_/FAINST[238].FA_/n2 ) );
  XOR \ADD_/FAINST[238].FA_/U1  ( .A(a[238]), .B(\ADD_/c[238] ), .Z(
        \ADD_/FAINST[238].FA_/n1 ) );
  XOR \ADD_/FAINST[237].FA_/U5  ( .A(\ADD_/FAINST[237].FA_/n3 ), .B(
        \ADD_/c[237] ), .Z(\ADD_/c[238] ) );
  XOR \ADD_/FAINST[237].FA_/U4  ( .A(\ADD_/FAINST[237].FA_/n1 ), .B(b[237]), 
        .Z(c[237]) );
  AND \ADD_/FAINST[237].FA_/U3  ( .A(\ADD_/FAINST[237].FA_/n1 ), .B(
        \ADD_/FAINST[237].FA_/n2 ), .Z(\ADD_/FAINST[237].FA_/n3 ) );
  XOR \ADD_/FAINST[237].FA_/U2  ( .A(b[237]), .B(\ADD_/c[237] ), .Z(
        \ADD_/FAINST[237].FA_/n2 ) );
  XOR \ADD_/FAINST[237].FA_/U1  ( .A(a[237]), .B(\ADD_/c[237] ), .Z(
        \ADD_/FAINST[237].FA_/n1 ) );
  XOR \ADD_/FAINST[236].FA_/U5  ( .A(\ADD_/FAINST[236].FA_/n3 ), .B(
        \ADD_/c[236] ), .Z(\ADD_/c[237] ) );
  XOR \ADD_/FAINST[236].FA_/U4  ( .A(\ADD_/FAINST[236].FA_/n1 ), .B(b[236]), 
        .Z(c[236]) );
  AND \ADD_/FAINST[236].FA_/U3  ( .A(\ADD_/FAINST[236].FA_/n1 ), .B(
        \ADD_/FAINST[236].FA_/n2 ), .Z(\ADD_/FAINST[236].FA_/n3 ) );
  XOR \ADD_/FAINST[236].FA_/U2  ( .A(b[236]), .B(\ADD_/c[236] ), .Z(
        \ADD_/FAINST[236].FA_/n2 ) );
  XOR \ADD_/FAINST[236].FA_/U1  ( .A(a[236]), .B(\ADD_/c[236] ), .Z(
        \ADD_/FAINST[236].FA_/n1 ) );
  XOR \ADD_/FAINST[235].FA_/U5  ( .A(\ADD_/FAINST[235].FA_/n3 ), .B(
        \ADD_/c[235] ), .Z(\ADD_/c[236] ) );
  XOR \ADD_/FAINST[235].FA_/U4  ( .A(\ADD_/FAINST[235].FA_/n1 ), .B(b[235]), 
        .Z(c[235]) );
  AND \ADD_/FAINST[235].FA_/U3  ( .A(\ADD_/FAINST[235].FA_/n1 ), .B(
        \ADD_/FAINST[235].FA_/n2 ), .Z(\ADD_/FAINST[235].FA_/n3 ) );
  XOR \ADD_/FAINST[235].FA_/U2  ( .A(b[235]), .B(\ADD_/c[235] ), .Z(
        \ADD_/FAINST[235].FA_/n2 ) );
  XOR \ADD_/FAINST[235].FA_/U1  ( .A(a[235]), .B(\ADD_/c[235] ), .Z(
        \ADD_/FAINST[235].FA_/n1 ) );
  XOR \ADD_/FAINST[234].FA_/U5  ( .A(\ADD_/FAINST[234].FA_/n3 ), .B(
        \ADD_/c[234] ), .Z(\ADD_/c[235] ) );
  XOR \ADD_/FAINST[234].FA_/U4  ( .A(\ADD_/FAINST[234].FA_/n1 ), .B(b[234]), 
        .Z(c[234]) );
  AND \ADD_/FAINST[234].FA_/U3  ( .A(\ADD_/FAINST[234].FA_/n1 ), .B(
        \ADD_/FAINST[234].FA_/n2 ), .Z(\ADD_/FAINST[234].FA_/n3 ) );
  XOR \ADD_/FAINST[234].FA_/U2  ( .A(b[234]), .B(\ADD_/c[234] ), .Z(
        \ADD_/FAINST[234].FA_/n2 ) );
  XOR \ADD_/FAINST[234].FA_/U1  ( .A(a[234]), .B(\ADD_/c[234] ), .Z(
        \ADD_/FAINST[234].FA_/n1 ) );
  XOR \ADD_/FAINST[233].FA_/U5  ( .A(\ADD_/FAINST[233].FA_/n3 ), .B(
        \ADD_/c[233] ), .Z(\ADD_/c[234] ) );
  XOR \ADD_/FAINST[233].FA_/U4  ( .A(\ADD_/FAINST[233].FA_/n1 ), .B(b[233]), 
        .Z(c[233]) );
  AND \ADD_/FAINST[233].FA_/U3  ( .A(\ADD_/FAINST[233].FA_/n1 ), .B(
        \ADD_/FAINST[233].FA_/n2 ), .Z(\ADD_/FAINST[233].FA_/n3 ) );
  XOR \ADD_/FAINST[233].FA_/U2  ( .A(b[233]), .B(\ADD_/c[233] ), .Z(
        \ADD_/FAINST[233].FA_/n2 ) );
  XOR \ADD_/FAINST[233].FA_/U1  ( .A(a[233]), .B(\ADD_/c[233] ), .Z(
        \ADD_/FAINST[233].FA_/n1 ) );
  XOR \ADD_/FAINST[232].FA_/U5  ( .A(\ADD_/FAINST[232].FA_/n3 ), .B(
        \ADD_/c[232] ), .Z(\ADD_/c[233] ) );
  XOR \ADD_/FAINST[232].FA_/U4  ( .A(\ADD_/FAINST[232].FA_/n1 ), .B(b[232]), 
        .Z(c[232]) );
  AND \ADD_/FAINST[232].FA_/U3  ( .A(\ADD_/FAINST[232].FA_/n1 ), .B(
        \ADD_/FAINST[232].FA_/n2 ), .Z(\ADD_/FAINST[232].FA_/n3 ) );
  XOR \ADD_/FAINST[232].FA_/U2  ( .A(b[232]), .B(\ADD_/c[232] ), .Z(
        \ADD_/FAINST[232].FA_/n2 ) );
  XOR \ADD_/FAINST[232].FA_/U1  ( .A(a[232]), .B(\ADD_/c[232] ), .Z(
        \ADD_/FAINST[232].FA_/n1 ) );
  XOR \ADD_/FAINST[231].FA_/U5  ( .A(\ADD_/FAINST[231].FA_/n3 ), .B(
        \ADD_/c[231] ), .Z(\ADD_/c[232] ) );
  XOR \ADD_/FAINST[231].FA_/U4  ( .A(\ADD_/FAINST[231].FA_/n1 ), .B(b[231]), 
        .Z(c[231]) );
  AND \ADD_/FAINST[231].FA_/U3  ( .A(\ADD_/FAINST[231].FA_/n1 ), .B(
        \ADD_/FAINST[231].FA_/n2 ), .Z(\ADD_/FAINST[231].FA_/n3 ) );
  XOR \ADD_/FAINST[231].FA_/U2  ( .A(b[231]), .B(\ADD_/c[231] ), .Z(
        \ADD_/FAINST[231].FA_/n2 ) );
  XOR \ADD_/FAINST[231].FA_/U1  ( .A(a[231]), .B(\ADD_/c[231] ), .Z(
        \ADD_/FAINST[231].FA_/n1 ) );
  XOR \ADD_/FAINST[230].FA_/U5  ( .A(\ADD_/FAINST[230].FA_/n3 ), .B(
        \ADD_/c[230] ), .Z(\ADD_/c[231] ) );
  XOR \ADD_/FAINST[230].FA_/U4  ( .A(\ADD_/FAINST[230].FA_/n1 ), .B(b[230]), 
        .Z(c[230]) );
  AND \ADD_/FAINST[230].FA_/U3  ( .A(\ADD_/FAINST[230].FA_/n1 ), .B(
        \ADD_/FAINST[230].FA_/n2 ), .Z(\ADD_/FAINST[230].FA_/n3 ) );
  XOR \ADD_/FAINST[230].FA_/U2  ( .A(b[230]), .B(\ADD_/c[230] ), .Z(
        \ADD_/FAINST[230].FA_/n2 ) );
  XOR \ADD_/FAINST[230].FA_/U1  ( .A(a[230]), .B(\ADD_/c[230] ), .Z(
        \ADD_/FAINST[230].FA_/n1 ) );
  XOR \ADD_/FAINST[229].FA_/U5  ( .A(\ADD_/FAINST[229].FA_/n3 ), .B(
        \ADD_/c[229] ), .Z(\ADD_/c[230] ) );
  XOR \ADD_/FAINST[229].FA_/U4  ( .A(\ADD_/FAINST[229].FA_/n1 ), .B(b[229]), 
        .Z(c[229]) );
  AND \ADD_/FAINST[229].FA_/U3  ( .A(\ADD_/FAINST[229].FA_/n1 ), .B(
        \ADD_/FAINST[229].FA_/n2 ), .Z(\ADD_/FAINST[229].FA_/n3 ) );
  XOR \ADD_/FAINST[229].FA_/U2  ( .A(b[229]), .B(\ADD_/c[229] ), .Z(
        \ADD_/FAINST[229].FA_/n2 ) );
  XOR \ADD_/FAINST[229].FA_/U1  ( .A(a[229]), .B(\ADD_/c[229] ), .Z(
        \ADD_/FAINST[229].FA_/n1 ) );
  XOR \ADD_/FAINST[228].FA_/U5  ( .A(\ADD_/FAINST[228].FA_/n3 ), .B(
        \ADD_/c[228] ), .Z(\ADD_/c[229] ) );
  XOR \ADD_/FAINST[228].FA_/U4  ( .A(\ADD_/FAINST[228].FA_/n1 ), .B(b[228]), 
        .Z(c[228]) );
  AND \ADD_/FAINST[228].FA_/U3  ( .A(\ADD_/FAINST[228].FA_/n1 ), .B(
        \ADD_/FAINST[228].FA_/n2 ), .Z(\ADD_/FAINST[228].FA_/n3 ) );
  XOR \ADD_/FAINST[228].FA_/U2  ( .A(b[228]), .B(\ADD_/c[228] ), .Z(
        \ADD_/FAINST[228].FA_/n2 ) );
  XOR \ADD_/FAINST[228].FA_/U1  ( .A(a[228]), .B(\ADD_/c[228] ), .Z(
        \ADD_/FAINST[228].FA_/n1 ) );
  XOR \ADD_/FAINST[227].FA_/U5  ( .A(\ADD_/FAINST[227].FA_/n3 ), .B(
        \ADD_/c[227] ), .Z(\ADD_/c[228] ) );
  XOR \ADD_/FAINST[227].FA_/U4  ( .A(\ADD_/FAINST[227].FA_/n1 ), .B(b[227]), 
        .Z(c[227]) );
  AND \ADD_/FAINST[227].FA_/U3  ( .A(\ADD_/FAINST[227].FA_/n1 ), .B(
        \ADD_/FAINST[227].FA_/n2 ), .Z(\ADD_/FAINST[227].FA_/n3 ) );
  XOR \ADD_/FAINST[227].FA_/U2  ( .A(b[227]), .B(\ADD_/c[227] ), .Z(
        \ADD_/FAINST[227].FA_/n2 ) );
  XOR \ADD_/FAINST[227].FA_/U1  ( .A(a[227]), .B(\ADD_/c[227] ), .Z(
        \ADD_/FAINST[227].FA_/n1 ) );
  XOR \ADD_/FAINST[226].FA_/U5  ( .A(\ADD_/FAINST[226].FA_/n3 ), .B(
        \ADD_/c[226] ), .Z(\ADD_/c[227] ) );
  XOR \ADD_/FAINST[226].FA_/U4  ( .A(\ADD_/FAINST[226].FA_/n1 ), .B(b[226]), 
        .Z(c[226]) );
  AND \ADD_/FAINST[226].FA_/U3  ( .A(\ADD_/FAINST[226].FA_/n1 ), .B(
        \ADD_/FAINST[226].FA_/n2 ), .Z(\ADD_/FAINST[226].FA_/n3 ) );
  XOR \ADD_/FAINST[226].FA_/U2  ( .A(b[226]), .B(\ADD_/c[226] ), .Z(
        \ADD_/FAINST[226].FA_/n2 ) );
  XOR \ADD_/FAINST[226].FA_/U1  ( .A(a[226]), .B(\ADD_/c[226] ), .Z(
        \ADD_/FAINST[226].FA_/n1 ) );
  XOR \ADD_/FAINST[225].FA_/U5  ( .A(\ADD_/FAINST[225].FA_/n3 ), .B(
        \ADD_/c[225] ), .Z(\ADD_/c[226] ) );
  XOR \ADD_/FAINST[225].FA_/U4  ( .A(\ADD_/FAINST[225].FA_/n1 ), .B(b[225]), 
        .Z(c[225]) );
  AND \ADD_/FAINST[225].FA_/U3  ( .A(\ADD_/FAINST[225].FA_/n1 ), .B(
        \ADD_/FAINST[225].FA_/n2 ), .Z(\ADD_/FAINST[225].FA_/n3 ) );
  XOR \ADD_/FAINST[225].FA_/U2  ( .A(b[225]), .B(\ADD_/c[225] ), .Z(
        \ADD_/FAINST[225].FA_/n2 ) );
  XOR \ADD_/FAINST[225].FA_/U1  ( .A(a[225]), .B(\ADD_/c[225] ), .Z(
        \ADD_/FAINST[225].FA_/n1 ) );
  XOR \ADD_/FAINST[224].FA_/U5  ( .A(\ADD_/FAINST[224].FA_/n3 ), .B(
        \ADD_/c[224] ), .Z(\ADD_/c[225] ) );
  XOR \ADD_/FAINST[224].FA_/U4  ( .A(\ADD_/FAINST[224].FA_/n1 ), .B(b[224]), 
        .Z(c[224]) );
  AND \ADD_/FAINST[224].FA_/U3  ( .A(\ADD_/FAINST[224].FA_/n1 ), .B(
        \ADD_/FAINST[224].FA_/n2 ), .Z(\ADD_/FAINST[224].FA_/n3 ) );
  XOR \ADD_/FAINST[224].FA_/U2  ( .A(b[224]), .B(\ADD_/c[224] ), .Z(
        \ADD_/FAINST[224].FA_/n2 ) );
  XOR \ADD_/FAINST[224].FA_/U1  ( .A(a[224]), .B(\ADD_/c[224] ), .Z(
        \ADD_/FAINST[224].FA_/n1 ) );
  XOR \ADD_/FAINST[223].FA_/U5  ( .A(\ADD_/FAINST[223].FA_/n3 ), .B(
        \ADD_/c[223] ), .Z(\ADD_/c[224] ) );
  XOR \ADD_/FAINST[223].FA_/U4  ( .A(\ADD_/FAINST[223].FA_/n1 ), .B(b[223]), 
        .Z(c[223]) );
  AND \ADD_/FAINST[223].FA_/U3  ( .A(\ADD_/FAINST[223].FA_/n1 ), .B(
        \ADD_/FAINST[223].FA_/n2 ), .Z(\ADD_/FAINST[223].FA_/n3 ) );
  XOR \ADD_/FAINST[223].FA_/U2  ( .A(b[223]), .B(\ADD_/c[223] ), .Z(
        \ADD_/FAINST[223].FA_/n2 ) );
  XOR \ADD_/FAINST[223].FA_/U1  ( .A(a[223]), .B(\ADD_/c[223] ), .Z(
        \ADD_/FAINST[223].FA_/n1 ) );
  XOR \ADD_/FAINST[222].FA_/U5  ( .A(\ADD_/FAINST[222].FA_/n3 ), .B(
        \ADD_/c[222] ), .Z(\ADD_/c[223] ) );
  XOR \ADD_/FAINST[222].FA_/U4  ( .A(\ADD_/FAINST[222].FA_/n1 ), .B(b[222]), 
        .Z(c[222]) );
  AND \ADD_/FAINST[222].FA_/U3  ( .A(\ADD_/FAINST[222].FA_/n1 ), .B(
        \ADD_/FAINST[222].FA_/n2 ), .Z(\ADD_/FAINST[222].FA_/n3 ) );
  XOR \ADD_/FAINST[222].FA_/U2  ( .A(b[222]), .B(\ADD_/c[222] ), .Z(
        \ADD_/FAINST[222].FA_/n2 ) );
  XOR \ADD_/FAINST[222].FA_/U1  ( .A(a[222]), .B(\ADD_/c[222] ), .Z(
        \ADD_/FAINST[222].FA_/n1 ) );
  XOR \ADD_/FAINST[221].FA_/U5  ( .A(\ADD_/FAINST[221].FA_/n3 ), .B(
        \ADD_/c[221] ), .Z(\ADD_/c[222] ) );
  XOR \ADD_/FAINST[221].FA_/U4  ( .A(\ADD_/FAINST[221].FA_/n1 ), .B(b[221]), 
        .Z(c[221]) );
  AND \ADD_/FAINST[221].FA_/U3  ( .A(\ADD_/FAINST[221].FA_/n1 ), .B(
        \ADD_/FAINST[221].FA_/n2 ), .Z(\ADD_/FAINST[221].FA_/n3 ) );
  XOR \ADD_/FAINST[221].FA_/U2  ( .A(b[221]), .B(\ADD_/c[221] ), .Z(
        \ADD_/FAINST[221].FA_/n2 ) );
  XOR \ADD_/FAINST[221].FA_/U1  ( .A(a[221]), .B(\ADD_/c[221] ), .Z(
        \ADD_/FAINST[221].FA_/n1 ) );
  XOR \ADD_/FAINST[220].FA_/U5  ( .A(\ADD_/FAINST[220].FA_/n3 ), .B(
        \ADD_/c[220] ), .Z(\ADD_/c[221] ) );
  XOR \ADD_/FAINST[220].FA_/U4  ( .A(\ADD_/FAINST[220].FA_/n1 ), .B(b[220]), 
        .Z(c[220]) );
  AND \ADD_/FAINST[220].FA_/U3  ( .A(\ADD_/FAINST[220].FA_/n1 ), .B(
        \ADD_/FAINST[220].FA_/n2 ), .Z(\ADD_/FAINST[220].FA_/n3 ) );
  XOR \ADD_/FAINST[220].FA_/U2  ( .A(b[220]), .B(\ADD_/c[220] ), .Z(
        \ADD_/FAINST[220].FA_/n2 ) );
  XOR \ADD_/FAINST[220].FA_/U1  ( .A(a[220]), .B(\ADD_/c[220] ), .Z(
        \ADD_/FAINST[220].FA_/n1 ) );
  XOR \ADD_/FAINST[219].FA_/U5  ( .A(\ADD_/FAINST[219].FA_/n3 ), .B(
        \ADD_/c[219] ), .Z(\ADD_/c[220] ) );
  XOR \ADD_/FAINST[219].FA_/U4  ( .A(\ADD_/FAINST[219].FA_/n1 ), .B(b[219]), 
        .Z(c[219]) );
  AND \ADD_/FAINST[219].FA_/U3  ( .A(\ADD_/FAINST[219].FA_/n1 ), .B(
        \ADD_/FAINST[219].FA_/n2 ), .Z(\ADD_/FAINST[219].FA_/n3 ) );
  XOR \ADD_/FAINST[219].FA_/U2  ( .A(b[219]), .B(\ADD_/c[219] ), .Z(
        \ADD_/FAINST[219].FA_/n2 ) );
  XOR \ADD_/FAINST[219].FA_/U1  ( .A(a[219]), .B(\ADD_/c[219] ), .Z(
        \ADD_/FAINST[219].FA_/n1 ) );
  XOR \ADD_/FAINST[218].FA_/U5  ( .A(\ADD_/FAINST[218].FA_/n3 ), .B(
        \ADD_/c[218] ), .Z(\ADD_/c[219] ) );
  XOR \ADD_/FAINST[218].FA_/U4  ( .A(\ADD_/FAINST[218].FA_/n1 ), .B(b[218]), 
        .Z(c[218]) );
  AND \ADD_/FAINST[218].FA_/U3  ( .A(\ADD_/FAINST[218].FA_/n1 ), .B(
        \ADD_/FAINST[218].FA_/n2 ), .Z(\ADD_/FAINST[218].FA_/n3 ) );
  XOR \ADD_/FAINST[218].FA_/U2  ( .A(b[218]), .B(\ADD_/c[218] ), .Z(
        \ADD_/FAINST[218].FA_/n2 ) );
  XOR \ADD_/FAINST[218].FA_/U1  ( .A(a[218]), .B(\ADD_/c[218] ), .Z(
        \ADD_/FAINST[218].FA_/n1 ) );
  XOR \ADD_/FAINST[217].FA_/U5  ( .A(\ADD_/FAINST[217].FA_/n3 ), .B(
        \ADD_/c[217] ), .Z(\ADD_/c[218] ) );
  XOR \ADD_/FAINST[217].FA_/U4  ( .A(\ADD_/FAINST[217].FA_/n1 ), .B(b[217]), 
        .Z(c[217]) );
  AND \ADD_/FAINST[217].FA_/U3  ( .A(\ADD_/FAINST[217].FA_/n1 ), .B(
        \ADD_/FAINST[217].FA_/n2 ), .Z(\ADD_/FAINST[217].FA_/n3 ) );
  XOR \ADD_/FAINST[217].FA_/U2  ( .A(b[217]), .B(\ADD_/c[217] ), .Z(
        \ADD_/FAINST[217].FA_/n2 ) );
  XOR \ADD_/FAINST[217].FA_/U1  ( .A(a[217]), .B(\ADD_/c[217] ), .Z(
        \ADD_/FAINST[217].FA_/n1 ) );
  XOR \ADD_/FAINST[216].FA_/U5  ( .A(\ADD_/FAINST[216].FA_/n3 ), .B(
        \ADD_/c[216] ), .Z(\ADD_/c[217] ) );
  XOR \ADD_/FAINST[216].FA_/U4  ( .A(\ADD_/FAINST[216].FA_/n1 ), .B(b[216]), 
        .Z(c[216]) );
  AND \ADD_/FAINST[216].FA_/U3  ( .A(\ADD_/FAINST[216].FA_/n1 ), .B(
        \ADD_/FAINST[216].FA_/n2 ), .Z(\ADD_/FAINST[216].FA_/n3 ) );
  XOR \ADD_/FAINST[216].FA_/U2  ( .A(b[216]), .B(\ADD_/c[216] ), .Z(
        \ADD_/FAINST[216].FA_/n2 ) );
  XOR \ADD_/FAINST[216].FA_/U1  ( .A(a[216]), .B(\ADD_/c[216] ), .Z(
        \ADD_/FAINST[216].FA_/n1 ) );
  XOR \ADD_/FAINST[215].FA_/U5  ( .A(\ADD_/FAINST[215].FA_/n3 ), .B(
        \ADD_/c[215] ), .Z(\ADD_/c[216] ) );
  XOR \ADD_/FAINST[215].FA_/U4  ( .A(\ADD_/FAINST[215].FA_/n1 ), .B(b[215]), 
        .Z(c[215]) );
  AND \ADD_/FAINST[215].FA_/U3  ( .A(\ADD_/FAINST[215].FA_/n1 ), .B(
        \ADD_/FAINST[215].FA_/n2 ), .Z(\ADD_/FAINST[215].FA_/n3 ) );
  XOR \ADD_/FAINST[215].FA_/U2  ( .A(b[215]), .B(\ADD_/c[215] ), .Z(
        \ADD_/FAINST[215].FA_/n2 ) );
  XOR \ADD_/FAINST[215].FA_/U1  ( .A(a[215]), .B(\ADD_/c[215] ), .Z(
        \ADD_/FAINST[215].FA_/n1 ) );
  XOR \ADD_/FAINST[214].FA_/U5  ( .A(\ADD_/FAINST[214].FA_/n3 ), .B(
        \ADD_/c[214] ), .Z(\ADD_/c[215] ) );
  XOR \ADD_/FAINST[214].FA_/U4  ( .A(\ADD_/FAINST[214].FA_/n1 ), .B(b[214]), 
        .Z(c[214]) );
  AND \ADD_/FAINST[214].FA_/U3  ( .A(\ADD_/FAINST[214].FA_/n1 ), .B(
        \ADD_/FAINST[214].FA_/n2 ), .Z(\ADD_/FAINST[214].FA_/n3 ) );
  XOR \ADD_/FAINST[214].FA_/U2  ( .A(b[214]), .B(\ADD_/c[214] ), .Z(
        \ADD_/FAINST[214].FA_/n2 ) );
  XOR \ADD_/FAINST[214].FA_/U1  ( .A(a[214]), .B(\ADD_/c[214] ), .Z(
        \ADD_/FAINST[214].FA_/n1 ) );
  XOR \ADD_/FAINST[213].FA_/U5  ( .A(\ADD_/FAINST[213].FA_/n3 ), .B(
        \ADD_/c[213] ), .Z(\ADD_/c[214] ) );
  XOR \ADD_/FAINST[213].FA_/U4  ( .A(\ADD_/FAINST[213].FA_/n1 ), .B(b[213]), 
        .Z(c[213]) );
  AND \ADD_/FAINST[213].FA_/U3  ( .A(\ADD_/FAINST[213].FA_/n1 ), .B(
        \ADD_/FAINST[213].FA_/n2 ), .Z(\ADD_/FAINST[213].FA_/n3 ) );
  XOR \ADD_/FAINST[213].FA_/U2  ( .A(b[213]), .B(\ADD_/c[213] ), .Z(
        \ADD_/FAINST[213].FA_/n2 ) );
  XOR \ADD_/FAINST[213].FA_/U1  ( .A(a[213]), .B(\ADD_/c[213] ), .Z(
        \ADD_/FAINST[213].FA_/n1 ) );
  XOR \ADD_/FAINST[212].FA_/U5  ( .A(\ADD_/FAINST[212].FA_/n3 ), .B(
        \ADD_/c[212] ), .Z(\ADD_/c[213] ) );
  XOR \ADD_/FAINST[212].FA_/U4  ( .A(\ADD_/FAINST[212].FA_/n1 ), .B(b[212]), 
        .Z(c[212]) );
  AND \ADD_/FAINST[212].FA_/U3  ( .A(\ADD_/FAINST[212].FA_/n1 ), .B(
        \ADD_/FAINST[212].FA_/n2 ), .Z(\ADD_/FAINST[212].FA_/n3 ) );
  XOR \ADD_/FAINST[212].FA_/U2  ( .A(b[212]), .B(\ADD_/c[212] ), .Z(
        \ADD_/FAINST[212].FA_/n2 ) );
  XOR \ADD_/FAINST[212].FA_/U1  ( .A(a[212]), .B(\ADD_/c[212] ), .Z(
        \ADD_/FAINST[212].FA_/n1 ) );
  XOR \ADD_/FAINST[211].FA_/U5  ( .A(\ADD_/FAINST[211].FA_/n3 ), .B(
        \ADD_/c[211] ), .Z(\ADD_/c[212] ) );
  XOR \ADD_/FAINST[211].FA_/U4  ( .A(\ADD_/FAINST[211].FA_/n1 ), .B(b[211]), 
        .Z(c[211]) );
  AND \ADD_/FAINST[211].FA_/U3  ( .A(\ADD_/FAINST[211].FA_/n1 ), .B(
        \ADD_/FAINST[211].FA_/n2 ), .Z(\ADD_/FAINST[211].FA_/n3 ) );
  XOR \ADD_/FAINST[211].FA_/U2  ( .A(b[211]), .B(\ADD_/c[211] ), .Z(
        \ADD_/FAINST[211].FA_/n2 ) );
  XOR \ADD_/FAINST[211].FA_/U1  ( .A(a[211]), .B(\ADD_/c[211] ), .Z(
        \ADD_/FAINST[211].FA_/n1 ) );
  XOR \ADD_/FAINST[210].FA_/U5  ( .A(\ADD_/FAINST[210].FA_/n3 ), .B(
        \ADD_/c[210] ), .Z(\ADD_/c[211] ) );
  XOR \ADD_/FAINST[210].FA_/U4  ( .A(\ADD_/FAINST[210].FA_/n1 ), .B(b[210]), 
        .Z(c[210]) );
  AND \ADD_/FAINST[210].FA_/U3  ( .A(\ADD_/FAINST[210].FA_/n1 ), .B(
        \ADD_/FAINST[210].FA_/n2 ), .Z(\ADD_/FAINST[210].FA_/n3 ) );
  XOR \ADD_/FAINST[210].FA_/U2  ( .A(b[210]), .B(\ADD_/c[210] ), .Z(
        \ADD_/FAINST[210].FA_/n2 ) );
  XOR \ADD_/FAINST[210].FA_/U1  ( .A(a[210]), .B(\ADD_/c[210] ), .Z(
        \ADD_/FAINST[210].FA_/n1 ) );
  XOR \ADD_/FAINST[209].FA_/U5  ( .A(\ADD_/FAINST[209].FA_/n3 ), .B(
        \ADD_/c[209] ), .Z(\ADD_/c[210] ) );
  XOR \ADD_/FAINST[209].FA_/U4  ( .A(\ADD_/FAINST[209].FA_/n1 ), .B(b[209]), 
        .Z(c[209]) );
  AND \ADD_/FAINST[209].FA_/U3  ( .A(\ADD_/FAINST[209].FA_/n1 ), .B(
        \ADD_/FAINST[209].FA_/n2 ), .Z(\ADD_/FAINST[209].FA_/n3 ) );
  XOR \ADD_/FAINST[209].FA_/U2  ( .A(b[209]), .B(\ADD_/c[209] ), .Z(
        \ADD_/FAINST[209].FA_/n2 ) );
  XOR \ADD_/FAINST[209].FA_/U1  ( .A(a[209]), .B(\ADD_/c[209] ), .Z(
        \ADD_/FAINST[209].FA_/n1 ) );
  XOR \ADD_/FAINST[208].FA_/U5  ( .A(\ADD_/FAINST[208].FA_/n3 ), .B(
        \ADD_/c[208] ), .Z(\ADD_/c[209] ) );
  XOR \ADD_/FAINST[208].FA_/U4  ( .A(\ADD_/FAINST[208].FA_/n1 ), .B(b[208]), 
        .Z(c[208]) );
  AND \ADD_/FAINST[208].FA_/U3  ( .A(\ADD_/FAINST[208].FA_/n1 ), .B(
        \ADD_/FAINST[208].FA_/n2 ), .Z(\ADD_/FAINST[208].FA_/n3 ) );
  XOR \ADD_/FAINST[208].FA_/U2  ( .A(b[208]), .B(\ADD_/c[208] ), .Z(
        \ADD_/FAINST[208].FA_/n2 ) );
  XOR \ADD_/FAINST[208].FA_/U1  ( .A(a[208]), .B(\ADD_/c[208] ), .Z(
        \ADD_/FAINST[208].FA_/n1 ) );
  XOR \ADD_/FAINST[207].FA_/U5  ( .A(\ADD_/FAINST[207].FA_/n3 ), .B(
        \ADD_/c[207] ), .Z(\ADD_/c[208] ) );
  XOR \ADD_/FAINST[207].FA_/U4  ( .A(\ADD_/FAINST[207].FA_/n1 ), .B(b[207]), 
        .Z(c[207]) );
  AND \ADD_/FAINST[207].FA_/U3  ( .A(\ADD_/FAINST[207].FA_/n1 ), .B(
        \ADD_/FAINST[207].FA_/n2 ), .Z(\ADD_/FAINST[207].FA_/n3 ) );
  XOR \ADD_/FAINST[207].FA_/U2  ( .A(b[207]), .B(\ADD_/c[207] ), .Z(
        \ADD_/FAINST[207].FA_/n2 ) );
  XOR \ADD_/FAINST[207].FA_/U1  ( .A(a[207]), .B(\ADD_/c[207] ), .Z(
        \ADD_/FAINST[207].FA_/n1 ) );
  XOR \ADD_/FAINST[206].FA_/U5  ( .A(\ADD_/FAINST[206].FA_/n3 ), .B(
        \ADD_/c[206] ), .Z(\ADD_/c[207] ) );
  XOR \ADD_/FAINST[206].FA_/U4  ( .A(\ADD_/FAINST[206].FA_/n1 ), .B(b[206]), 
        .Z(c[206]) );
  AND \ADD_/FAINST[206].FA_/U3  ( .A(\ADD_/FAINST[206].FA_/n1 ), .B(
        \ADD_/FAINST[206].FA_/n2 ), .Z(\ADD_/FAINST[206].FA_/n3 ) );
  XOR \ADD_/FAINST[206].FA_/U2  ( .A(b[206]), .B(\ADD_/c[206] ), .Z(
        \ADD_/FAINST[206].FA_/n2 ) );
  XOR \ADD_/FAINST[206].FA_/U1  ( .A(a[206]), .B(\ADD_/c[206] ), .Z(
        \ADD_/FAINST[206].FA_/n1 ) );
  XOR \ADD_/FAINST[205].FA_/U5  ( .A(\ADD_/FAINST[205].FA_/n3 ), .B(
        \ADD_/c[205] ), .Z(\ADD_/c[206] ) );
  XOR \ADD_/FAINST[205].FA_/U4  ( .A(\ADD_/FAINST[205].FA_/n1 ), .B(b[205]), 
        .Z(c[205]) );
  AND \ADD_/FAINST[205].FA_/U3  ( .A(\ADD_/FAINST[205].FA_/n1 ), .B(
        \ADD_/FAINST[205].FA_/n2 ), .Z(\ADD_/FAINST[205].FA_/n3 ) );
  XOR \ADD_/FAINST[205].FA_/U2  ( .A(b[205]), .B(\ADD_/c[205] ), .Z(
        \ADD_/FAINST[205].FA_/n2 ) );
  XOR \ADD_/FAINST[205].FA_/U1  ( .A(a[205]), .B(\ADD_/c[205] ), .Z(
        \ADD_/FAINST[205].FA_/n1 ) );
  XOR \ADD_/FAINST[204].FA_/U5  ( .A(\ADD_/FAINST[204].FA_/n3 ), .B(
        \ADD_/c[204] ), .Z(\ADD_/c[205] ) );
  XOR \ADD_/FAINST[204].FA_/U4  ( .A(\ADD_/FAINST[204].FA_/n1 ), .B(b[204]), 
        .Z(c[204]) );
  AND \ADD_/FAINST[204].FA_/U3  ( .A(\ADD_/FAINST[204].FA_/n1 ), .B(
        \ADD_/FAINST[204].FA_/n2 ), .Z(\ADD_/FAINST[204].FA_/n3 ) );
  XOR \ADD_/FAINST[204].FA_/U2  ( .A(b[204]), .B(\ADD_/c[204] ), .Z(
        \ADD_/FAINST[204].FA_/n2 ) );
  XOR \ADD_/FAINST[204].FA_/U1  ( .A(a[204]), .B(\ADD_/c[204] ), .Z(
        \ADD_/FAINST[204].FA_/n1 ) );
  XOR \ADD_/FAINST[203].FA_/U5  ( .A(\ADD_/FAINST[203].FA_/n3 ), .B(
        \ADD_/c[203] ), .Z(\ADD_/c[204] ) );
  XOR \ADD_/FAINST[203].FA_/U4  ( .A(\ADD_/FAINST[203].FA_/n1 ), .B(b[203]), 
        .Z(c[203]) );
  AND \ADD_/FAINST[203].FA_/U3  ( .A(\ADD_/FAINST[203].FA_/n1 ), .B(
        \ADD_/FAINST[203].FA_/n2 ), .Z(\ADD_/FAINST[203].FA_/n3 ) );
  XOR \ADD_/FAINST[203].FA_/U2  ( .A(b[203]), .B(\ADD_/c[203] ), .Z(
        \ADD_/FAINST[203].FA_/n2 ) );
  XOR \ADD_/FAINST[203].FA_/U1  ( .A(a[203]), .B(\ADD_/c[203] ), .Z(
        \ADD_/FAINST[203].FA_/n1 ) );
  XOR \ADD_/FAINST[202].FA_/U5  ( .A(\ADD_/FAINST[202].FA_/n3 ), .B(
        \ADD_/c[202] ), .Z(\ADD_/c[203] ) );
  XOR \ADD_/FAINST[202].FA_/U4  ( .A(\ADD_/FAINST[202].FA_/n1 ), .B(b[202]), 
        .Z(c[202]) );
  AND \ADD_/FAINST[202].FA_/U3  ( .A(\ADD_/FAINST[202].FA_/n1 ), .B(
        \ADD_/FAINST[202].FA_/n2 ), .Z(\ADD_/FAINST[202].FA_/n3 ) );
  XOR \ADD_/FAINST[202].FA_/U2  ( .A(b[202]), .B(\ADD_/c[202] ), .Z(
        \ADD_/FAINST[202].FA_/n2 ) );
  XOR \ADD_/FAINST[202].FA_/U1  ( .A(a[202]), .B(\ADD_/c[202] ), .Z(
        \ADD_/FAINST[202].FA_/n1 ) );
  XOR \ADD_/FAINST[201].FA_/U5  ( .A(\ADD_/FAINST[201].FA_/n3 ), .B(
        \ADD_/c[201] ), .Z(\ADD_/c[202] ) );
  XOR \ADD_/FAINST[201].FA_/U4  ( .A(\ADD_/FAINST[201].FA_/n1 ), .B(b[201]), 
        .Z(c[201]) );
  AND \ADD_/FAINST[201].FA_/U3  ( .A(\ADD_/FAINST[201].FA_/n1 ), .B(
        \ADD_/FAINST[201].FA_/n2 ), .Z(\ADD_/FAINST[201].FA_/n3 ) );
  XOR \ADD_/FAINST[201].FA_/U2  ( .A(b[201]), .B(\ADD_/c[201] ), .Z(
        \ADD_/FAINST[201].FA_/n2 ) );
  XOR \ADD_/FAINST[201].FA_/U1  ( .A(a[201]), .B(\ADD_/c[201] ), .Z(
        \ADD_/FAINST[201].FA_/n1 ) );
  XOR \ADD_/FAINST[200].FA_/U5  ( .A(\ADD_/FAINST[200].FA_/n3 ), .B(
        \ADD_/c[200] ), .Z(\ADD_/c[201] ) );
  XOR \ADD_/FAINST[200].FA_/U4  ( .A(\ADD_/FAINST[200].FA_/n1 ), .B(b[200]), 
        .Z(c[200]) );
  AND \ADD_/FAINST[200].FA_/U3  ( .A(\ADD_/FAINST[200].FA_/n1 ), .B(
        \ADD_/FAINST[200].FA_/n2 ), .Z(\ADD_/FAINST[200].FA_/n3 ) );
  XOR \ADD_/FAINST[200].FA_/U2  ( .A(b[200]), .B(\ADD_/c[200] ), .Z(
        \ADD_/FAINST[200].FA_/n2 ) );
  XOR \ADD_/FAINST[200].FA_/U1  ( .A(a[200]), .B(\ADD_/c[200] ), .Z(
        \ADD_/FAINST[200].FA_/n1 ) );
  XOR \ADD_/FAINST[199].FA_/U5  ( .A(\ADD_/FAINST[199].FA_/n3 ), .B(
        \ADD_/c[199] ), .Z(\ADD_/c[200] ) );
  XOR \ADD_/FAINST[199].FA_/U4  ( .A(\ADD_/FAINST[199].FA_/n1 ), .B(b[199]), 
        .Z(c[199]) );
  AND \ADD_/FAINST[199].FA_/U3  ( .A(\ADD_/FAINST[199].FA_/n1 ), .B(
        \ADD_/FAINST[199].FA_/n2 ), .Z(\ADD_/FAINST[199].FA_/n3 ) );
  XOR \ADD_/FAINST[199].FA_/U2  ( .A(b[199]), .B(\ADD_/c[199] ), .Z(
        \ADD_/FAINST[199].FA_/n2 ) );
  XOR \ADD_/FAINST[199].FA_/U1  ( .A(a[199]), .B(\ADD_/c[199] ), .Z(
        \ADD_/FAINST[199].FA_/n1 ) );
  XOR \ADD_/FAINST[198].FA_/U5  ( .A(\ADD_/FAINST[198].FA_/n3 ), .B(
        \ADD_/c[198] ), .Z(\ADD_/c[199] ) );
  XOR \ADD_/FAINST[198].FA_/U4  ( .A(\ADD_/FAINST[198].FA_/n1 ), .B(b[198]), 
        .Z(c[198]) );
  AND \ADD_/FAINST[198].FA_/U3  ( .A(\ADD_/FAINST[198].FA_/n1 ), .B(
        \ADD_/FAINST[198].FA_/n2 ), .Z(\ADD_/FAINST[198].FA_/n3 ) );
  XOR \ADD_/FAINST[198].FA_/U2  ( .A(b[198]), .B(\ADD_/c[198] ), .Z(
        \ADD_/FAINST[198].FA_/n2 ) );
  XOR \ADD_/FAINST[198].FA_/U1  ( .A(a[198]), .B(\ADD_/c[198] ), .Z(
        \ADD_/FAINST[198].FA_/n1 ) );
  XOR \ADD_/FAINST[197].FA_/U5  ( .A(\ADD_/FAINST[197].FA_/n3 ), .B(
        \ADD_/c[197] ), .Z(\ADD_/c[198] ) );
  XOR \ADD_/FAINST[197].FA_/U4  ( .A(\ADD_/FAINST[197].FA_/n1 ), .B(b[197]), 
        .Z(c[197]) );
  AND \ADD_/FAINST[197].FA_/U3  ( .A(\ADD_/FAINST[197].FA_/n1 ), .B(
        \ADD_/FAINST[197].FA_/n2 ), .Z(\ADD_/FAINST[197].FA_/n3 ) );
  XOR \ADD_/FAINST[197].FA_/U2  ( .A(b[197]), .B(\ADD_/c[197] ), .Z(
        \ADD_/FAINST[197].FA_/n2 ) );
  XOR \ADD_/FAINST[197].FA_/U1  ( .A(a[197]), .B(\ADD_/c[197] ), .Z(
        \ADD_/FAINST[197].FA_/n1 ) );
  XOR \ADD_/FAINST[196].FA_/U5  ( .A(\ADD_/FAINST[196].FA_/n3 ), .B(
        \ADD_/c[196] ), .Z(\ADD_/c[197] ) );
  XOR \ADD_/FAINST[196].FA_/U4  ( .A(\ADD_/FAINST[196].FA_/n1 ), .B(b[196]), 
        .Z(c[196]) );
  AND \ADD_/FAINST[196].FA_/U3  ( .A(\ADD_/FAINST[196].FA_/n1 ), .B(
        \ADD_/FAINST[196].FA_/n2 ), .Z(\ADD_/FAINST[196].FA_/n3 ) );
  XOR \ADD_/FAINST[196].FA_/U2  ( .A(b[196]), .B(\ADD_/c[196] ), .Z(
        \ADD_/FAINST[196].FA_/n2 ) );
  XOR \ADD_/FAINST[196].FA_/U1  ( .A(a[196]), .B(\ADD_/c[196] ), .Z(
        \ADD_/FAINST[196].FA_/n1 ) );
  XOR \ADD_/FAINST[195].FA_/U5  ( .A(\ADD_/FAINST[195].FA_/n3 ), .B(
        \ADD_/c[195] ), .Z(\ADD_/c[196] ) );
  XOR \ADD_/FAINST[195].FA_/U4  ( .A(\ADD_/FAINST[195].FA_/n1 ), .B(b[195]), 
        .Z(c[195]) );
  AND \ADD_/FAINST[195].FA_/U3  ( .A(\ADD_/FAINST[195].FA_/n1 ), .B(
        \ADD_/FAINST[195].FA_/n2 ), .Z(\ADD_/FAINST[195].FA_/n3 ) );
  XOR \ADD_/FAINST[195].FA_/U2  ( .A(b[195]), .B(\ADD_/c[195] ), .Z(
        \ADD_/FAINST[195].FA_/n2 ) );
  XOR \ADD_/FAINST[195].FA_/U1  ( .A(a[195]), .B(\ADD_/c[195] ), .Z(
        \ADD_/FAINST[195].FA_/n1 ) );
  XOR \ADD_/FAINST[194].FA_/U5  ( .A(\ADD_/FAINST[194].FA_/n3 ), .B(
        \ADD_/c[194] ), .Z(\ADD_/c[195] ) );
  XOR \ADD_/FAINST[194].FA_/U4  ( .A(\ADD_/FAINST[194].FA_/n1 ), .B(b[194]), 
        .Z(c[194]) );
  AND \ADD_/FAINST[194].FA_/U3  ( .A(\ADD_/FAINST[194].FA_/n1 ), .B(
        \ADD_/FAINST[194].FA_/n2 ), .Z(\ADD_/FAINST[194].FA_/n3 ) );
  XOR \ADD_/FAINST[194].FA_/U2  ( .A(b[194]), .B(\ADD_/c[194] ), .Z(
        \ADD_/FAINST[194].FA_/n2 ) );
  XOR \ADD_/FAINST[194].FA_/U1  ( .A(a[194]), .B(\ADD_/c[194] ), .Z(
        \ADD_/FAINST[194].FA_/n1 ) );
  XOR \ADD_/FAINST[193].FA_/U5  ( .A(\ADD_/FAINST[193].FA_/n3 ), .B(
        \ADD_/c[193] ), .Z(\ADD_/c[194] ) );
  XOR \ADD_/FAINST[193].FA_/U4  ( .A(\ADD_/FAINST[193].FA_/n1 ), .B(b[193]), 
        .Z(c[193]) );
  AND \ADD_/FAINST[193].FA_/U3  ( .A(\ADD_/FAINST[193].FA_/n1 ), .B(
        \ADD_/FAINST[193].FA_/n2 ), .Z(\ADD_/FAINST[193].FA_/n3 ) );
  XOR \ADD_/FAINST[193].FA_/U2  ( .A(b[193]), .B(\ADD_/c[193] ), .Z(
        \ADD_/FAINST[193].FA_/n2 ) );
  XOR \ADD_/FAINST[193].FA_/U1  ( .A(a[193]), .B(\ADD_/c[193] ), .Z(
        \ADD_/FAINST[193].FA_/n1 ) );
  XOR \ADD_/FAINST[192].FA_/U5  ( .A(\ADD_/FAINST[192].FA_/n3 ), .B(
        \ADD_/c[192] ), .Z(\ADD_/c[193] ) );
  XOR \ADD_/FAINST[192].FA_/U4  ( .A(\ADD_/FAINST[192].FA_/n1 ), .B(b[192]), 
        .Z(c[192]) );
  AND \ADD_/FAINST[192].FA_/U3  ( .A(\ADD_/FAINST[192].FA_/n1 ), .B(
        \ADD_/FAINST[192].FA_/n2 ), .Z(\ADD_/FAINST[192].FA_/n3 ) );
  XOR \ADD_/FAINST[192].FA_/U2  ( .A(b[192]), .B(\ADD_/c[192] ), .Z(
        \ADD_/FAINST[192].FA_/n2 ) );
  XOR \ADD_/FAINST[192].FA_/U1  ( .A(a[192]), .B(\ADD_/c[192] ), .Z(
        \ADD_/FAINST[192].FA_/n1 ) );
  XOR \ADD_/FAINST[191].FA_/U5  ( .A(\ADD_/FAINST[191].FA_/n3 ), .B(
        \ADD_/c[191] ), .Z(\ADD_/c[192] ) );
  XOR \ADD_/FAINST[191].FA_/U4  ( .A(\ADD_/FAINST[191].FA_/n1 ), .B(b[191]), 
        .Z(c[191]) );
  AND \ADD_/FAINST[191].FA_/U3  ( .A(\ADD_/FAINST[191].FA_/n1 ), .B(
        \ADD_/FAINST[191].FA_/n2 ), .Z(\ADD_/FAINST[191].FA_/n3 ) );
  XOR \ADD_/FAINST[191].FA_/U2  ( .A(b[191]), .B(\ADD_/c[191] ), .Z(
        \ADD_/FAINST[191].FA_/n2 ) );
  XOR \ADD_/FAINST[191].FA_/U1  ( .A(a[191]), .B(\ADD_/c[191] ), .Z(
        \ADD_/FAINST[191].FA_/n1 ) );
  XOR \ADD_/FAINST[190].FA_/U5  ( .A(\ADD_/FAINST[190].FA_/n3 ), .B(
        \ADD_/c[190] ), .Z(\ADD_/c[191] ) );
  XOR \ADD_/FAINST[190].FA_/U4  ( .A(\ADD_/FAINST[190].FA_/n1 ), .B(b[190]), 
        .Z(c[190]) );
  AND \ADD_/FAINST[190].FA_/U3  ( .A(\ADD_/FAINST[190].FA_/n1 ), .B(
        \ADD_/FAINST[190].FA_/n2 ), .Z(\ADD_/FAINST[190].FA_/n3 ) );
  XOR \ADD_/FAINST[190].FA_/U2  ( .A(b[190]), .B(\ADD_/c[190] ), .Z(
        \ADD_/FAINST[190].FA_/n2 ) );
  XOR \ADD_/FAINST[190].FA_/U1  ( .A(a[190]), .B(\ADD_/c[190] ), .Z(
        \ADD_/FAINST[190].FA_/n1 ) );
  XOR \ADD_/FAINST[189].FA_/U5  ( .A(\ADD_/FAINST[189].FA_/n3 ), .B(
        \ADD_/c[189] ), .Z(\ADD_/c[190] ) );
  XOR \ADD_/FAINST[189].FA_/U4  ( .A(\ADD_/FAINST[189].FA_/n1 ), .B(b[189]), 
        .Z(c[189]) );
  AND \ADD_/FAINST[189].FA_/U3  ( .A(\ADD_/FAINST[189].FA_/n1 ), .B(
        \ADD_/FAINST[189].FA_/n2 ), .Z(\ADD_/FAINST[189].FA_/n3 ) );
  XOR \ADD_/FAINST[189].FA_/U2  ( .A(b[189]), .B(\ADD_/c[189] ), .Z(
        \ADD_/FAINST[189].FA_/n2 ) );
  XOR \ADD_/FAINST[189].FA_/U1  ( .A(a[189]), .B(\ADD_/c[189] ), .Z(
        \ADD_/FAINST[189].FA_/n1 ) );
  XOR \ADD_/FAINST[188].FA_/U5  ( .A(\ADD_/FAINST[188].FA_/n3 ), .B(
        \ADD_/c[188] ), .Z(\ADD_/c[189] ) );
  XOR \ADD_/FAINST[188].FA_/U4  ( .A(\ADD_/FAINST[188].FA_/n1 ), .B(b[188]), 
        .Z(c[188]) );
  AND \ADD_/FAINST[188].FA_/U3  ( .A(\ADD_/FAINST[188].FA_/n1 ), .B(
        \ADD_/FAINST[188].FA_/n2 ), .Z(\ADD_/FAINST[188].FA_/n3 ) );
  XOR \ADD_/FAINST[188].FA_/U2  ( .A(b[188]), .B(\ADD_/c[188] ), .Z(
        \ADD_/FAINST[188].FA_/n2 ) );
  XOR \ADD_/FAINST[188].FA_/U1  ( .A(a[188]), .B(\ADD_/c[188] ), .Z(
        \ADD_/FAINST[188].FA_/n1 ) );
  XOR \ADD_/FAINST[187].FA_/U5  ( .A(\ADD_/FAINST[187].FA_/n3 ), .B(
        \ADD_/c[187] ), .Z(\ADD_/c[188] ) );
  XOR \ADD_/FAINST[187].FA_/U4  ( .A(\ADD_/FAINST[187].FA_/n1 ), .B(b[187]), 
        .Z(c[187]) );
  AND \ADD_/FAINST[187].FA_/U3  ( .A(\ADD_/FAINST[187].FA_/n1 ), .B(
        \ADD_/FAINST[187].FA_/n2 ), .Z(\ADD_/FAINST[187].FA_/n3 ) );
  XOR \ADD_/FAINST[187].FA_/U2  ( .A(b[187]), .B(\ADD_/c[187] ), .Z(
        \ADD_/FAINST[187].FA_/n2 ) );
  XOR \ADD_/FAINST[187].FA_/U1  ( .A(a[187]), .B(\ADD_/c[187] ), .Z(
        \ADD_/FAINST[187].FA_/n1 ) );
  XOR \ADD_/FAINST[186].FA_/U5  ( .A(\ADD_/FAINST[186].FA_/n3 ), .B(
        \ADD_/c[186] ), .Z(\ADD_/c[187] ) );
  XOR \ADD_/FAINST[186].FA_/U4  ( .A(\ADD_/FAINST[186].FA_/n1 ), .B(b[186]), 
        .Z(c[186]) );
  AND \ADD_/FAINST[186].FA_/U3  ( .A(\ADD_/FAINST[186].FA_/n1 ), .B(
        \ADD_/FAINST[186].FA_/n2 ), .Z(\ADD_/FAINST[186].FA_/n3 ) );
  XOR \ADD_/FAINST[186].FA_/U2  ( .A(b[186]), .B(\ADD_/c[186] ), .Z(
        \ADD_/FAINST[186].FA_/n2 ) );
  XOR \ADD_/FAINST[186].FA_/U1  ( .A(a[186]), .B(\ADD_/c[186] ), .Z(
        \ADD_/FAINST[186].FA_/n1 ) );
  XOR \ADD_/FAINST[185].FA_/U5  ( .A(\ADD_/FAINST[185].FA_/n3 ), .B(
        \ADD_/c[185] ), .Z(\ADD_/c[186] ) );
  XOR \ADD_/FAINST[185].FA_/U4  ( .A(\ADD_/FAINST[185].FA_/n1 ), .B(b[185]), 
        .Z(c[185]) );
  AND \ADD_/FAINST[185].FA_/U3  ( .A(\ADD_/FAINST[185].FA_/n1 ), .B(
        \ADD_/FAINST[185].FA_/n2 ), .Z(\ADD_/FAINST[185].FA_/n3 ) );
  XOR \ADD_/FAINST[185].FA_/U2  ( .A(b[185]), .B(\ADD_/c[185] ), .Z(
        \ADD_/FAINST[185].FA_/n2 ) );
  XOR \ADD_/FAINST[185].FA_/U1  ( .A(a[185]), .B(\ADD_/c[185] ), .Z(
        \ADD_/FAINST[185].FA_/n1 ) );
  XOR \ADD_/FAINST[184].FA_/U5  ( .A(\ADD_/FAINST[184].FA_/n3 ), .B(
        \ADD_/c[184] ), .Z(\ADD_/c[185] ) );
  XOR \ADD_/FAINST[184].FA_/U4  ( .A(\ADD_/FAINST[184].FA_/n1 ), .B(b[184]), 
        .Z(c[184]) );
  AND \ADD_/FAINST[184].FA_/U3  ( .A(\ADD_/FAINST[184].FA_/n1 ), .B(
        \ADD_/FAINST[184].FA_/n2 ), .Z(\ADD_/FAINST[184].FA_/n3 ) );
  XOR \ADD_/FAINST[184].FA_/U2  ( .A(b[184]), .B(\ADD_/c[184] ), .Z(
        \ADD_/FAINST[184].FA_/n2 ) );
  XOR \ADD_/FAINST[184].FA_/U1  ( .A(a[184]), .B(\ADD_/c[184] ), .Z(
        \ADD_/FAINST[184].FA_/n1 ) );
  XOR \ADD_/FAINST[183].FA_/U5  ( .A(\ADD_/FAINST[183].FA_/n3 ), .B(
        \ADD_/c[183] ), .Z(\ADD_/c[184] ) );
  XOR \ADD_/FAINST[183].FA_/U4  ( .A(\ADD_/FAINST[183].FA_/n1 ), .B(b[183]), 
        .Z(c[183]) );
  AND \ADD_/FAINST[183].FA_/U3  ( .A(\ADD_/FAINST[183].FA_/n1 ), .B(
        \ADD_/FAINST[183].FA_/n2 ), .Z(\ADD_/FAINST[183].FA_/n3 ) );
  XOR \ADD_/FAINST[183].FA_/U2  ( .A(b[183]), .B(\ADD_/c[183] ), .Z(
        \ADD_/FAINST[183].FA_/n2 ) );
  XOR \ADD_/FAINST[183].FA_/U1  ( .A(a[183]), .B(\ADD_/c[183] ), .Z(
        \ADD_/FAINST[183].FA_/n1 ) );
  XOR \ADD_/FAINST[182].FA_/U5  ( .A(\ADD_/FAINST[182].FA_/n3 ), .B(
        \ADD_/c[182] ), .Z(\ADD_/c[183] ) );
  XOR \ADD_/FAINST[182].FA_/U4  ( .A(\ADD_/FAINST[182].FA_/n1 ), .B(b[182]), 
        .Z(c[182]) );
  AND \ADD_/FAINST[182].FA_/U3  ( .A(\ADD_/FAINST[182].FA_/n1 ), .B(
        \ADD_/FAINST[182].FA_/n2 ), .Z(\ADD_/FAINST[182].FA_/n3 ) );
  XOR \ADD_/FAINST[182].FA_/U2  ( .A(b[182]), .B(\ADD_/c[182] ), .Z(
        \ADD_/FAINST[182].FA_/n2 ) );
  XOR \ADD_/FAINST[182].FA_/U1  ( .A(a[182]), .B(\ADD_/c[182] ), .Z(
        \ADD_/FAINST[182].FA_/n1 ) );
  XOR \ADD_/FAINST[181].FA_/U5  ( .A(\ADD_/FAINST[181].FA_/n3 ), .B(
        \ADD_/c[181] ), .Z(\ADD_/c[182] ) );
  XOR \ADD_/FAINST[181].FA_/U4  ( .A(\ADD_/FAINST[181].FA_/n1 ), .B(b[181]), 
        .Z(c[181]) );
  AND \ADD_/FAINST[181].FA_/U3  ( .A(\ADD_/FAINST[181].FA_/n1 ), .B(
        \ADD_/FAINST[181].FA_/n2 ), .Z(\ADD_/FAINST[181].FA_/n3 ) );
  XOR \ADD_/FAINST[181].FA_/U2  ( .A(b[181]), .B(\ADD_/c[181] ), .Z(
        \ADD_/FAINST[181].FA_/n2 ) );
  XOR \ADD_/FAINST[181].FA_/U1  ( .A(a[181]), .B(\ADD_/c[181] ), .Z(
        \ADD_/FAINST[181].FA_/n1 ) );
  XOR \ADD_/FAINST[180].FA_/U5  ( .A(\ADD_/FAINST[180].FA_/n3 ), .B(
        \ADD_/c[180] ), .Z(\ADD_/c[181] ) );
  XOR \ADD_/FAINST[180].FA_/U4  ( .A(\ADD_/FAINST[180].FA_/n1 ), .B(b[180]), 
        .Z(c[180]) );
  AND \ADD_/FAINST[180].FA_/U3  ( .A(\ADD_/FAINST[180].FA_/n1 ), .B(
        \ADD_/FAINST[180].FA_/n2 ), .Z(\ADD_/FAINST[180].FA_/n3 ) );
  XOR \ADD_/FAINST[180].FA_/U2  ( .A(b[180]), .B(\ADD_/c[180] ), .Z(
        \ADD_/FAINST[180].FA_/n2 ) );
  XOR \ADD_/FAINST[180].FA_/U1  ( .A(a[180]), .B(\ADD_/c[180] ), .Z(
        \ADD_/FAINST[180].FA_/n1 ) );
  XOR \ADD_/FAINST[179].FA_/U5  ( .A(\ADD_/FAINST[179].FA_/n3 ), .B(
        \ADD_/c[179] ), .Z(\ADD_/c[180] ) );
  XOR \ADD_/FAINST[179].FA_/U4  ( .A(\ADD_/FAINST[179].FA_/n1 ), .B(b[179]), 
        .Z(c[179]) );
  AND \ADD_/FAINST[179].FA_/U3  ( .A(\ADD_/FAINST[179].FA_/n1 ), .B(
        \ADD_/FAINST[179].FA_/n2 ), .Z(\ADD_/FAINST[179].FA_/n3 ) );
  XOR \ADD_/FAINST[179].FA_/U2  ( .A(b[179]), .B(\ADD_/c[179] ), .Z(
        \ADD_/FAINST[179].FA_/n2 ) );
  XOR \ADD_/FAINST[179].FA_/U1  ( .A(a[179]), .B(\ADD_/c[179] ), .Z(
        \ADD_/FAINST[179].FA_/n1 ) );
  XOR \ADD_/FAINST[178].FA_/U5  ( .A(\ADD_/FAINST[178].FA_/n3 ), .B(
        \ADD_/c[178] ), .Z(\ADD_/c[179] ) );
  XOR \ADD_/FAINST[178].FA_/U4  ( .A(\ADD_/FAINST[178].FA_/n1 ), .B(b[178]), 
        .Z(c[178]) );
  AND \ADD_/FAINST[178].FA_/U3  ( .A(\ADD_/FAINST[178].FA_/n1 ), .B(
        \ADD_/FAINST[178].FA_/n2 ), .Z(\ADD_/FAINST[178].FA_/n3 ) );
  XOR \ADD_/FAINST[178].FA_/U2  ( .A(b[178]), .B(\ADD_/c[178] ), .Z(
        \ADD_/FAINST[178].FA_/n2 ) );
  XOR \ADD_/FAINST[178].FA_/U1  ( .A(a[178]), .B(\ADD_/c[178] ), .Z(
        \ADD_/FAINST[178].FA_/n1 ) );
  XOR \ADD_/FAINST[177].FA_/U5  ( .A(\ADD_/FAINST[177].FA_/n3 ), .B(
        \ADD_/c[177] ), .Z(\ADD_/c[178] ) );
  XOR \ADD_/FAINST[177].FA_/U4  ( .A(\ADD_/FAINST[177].FA_/n1 ), .B(b[177]), 
        .Z(c[177]) );
  AND \ADD_/FAINST[177].FA_/U3  ( .A(\ADD_/FAINST[177].FA_/n1 ), .B(
        \ADD_/FAINST[177].FA_/n2 ), .Z(\ADD_/FAINST[177].FA_/n3 ) );
  XOR \ADD_/FAINST[177].FA_/U2  ( .A(b[177]), .B(\ADD_/c[177] ), .Z(
        \ADD_/FAINST[177].FA_/n2 ) );
  XOR \ADD_/FAINST[177].FA_/U1  ( .A(a[177]), .B(\ADD_/c[177] ), .Z(
        \ADD_/FAINST[177].FA_/n1 ) );
  XOR \ADD_/FAINST[176].FA_/U5  ( .A(\ADD_/FAINST[176].FA_/n3 ), .B(
        \ADD_/c[176] ), .Z(\ADD_/c[177] ) );
  XOR \ADD_/FAINST[176].FA_/U4  ( .A(\ADD_/FAINST[176].FA_/n1 ), .B(b[176]), 
        .Z(c[176]) );
  AND \ADD_/FAINST[176].FA_/U3  ( .A(\ADD_/FAINST[176].FA_/n1 ), .B(
        \ADD_/FAINST[176].FA_/n2 ), .Z(\ADD_/FAINST[176].FA_/n3 ) );
  XOR \ADD_/FAINST[176].FA_/U2  ( .A(b[176]), .B(\ADD_/c[176] ), .Z(
        \ADD_/FAINST[176].FA_/n2 ) );
  XOR \ADD_/FAINST[176].FA_/U1  ( .A(a[176]), .B(\ADD_/c[176] ), .Z(
        \ADD_/FAINST[176].FA_/n1 ) );
  XOR \ADD_/FAINST[175].FA_/U5  ( .A(\ADD_/FAINST[175].FA_/n3 ), .B(
        \ADD_/c[175] ), .Z(\ADD_/c[176] ) );
  XOR \ADD_/FAINST[175].FA_/U4  ( .A(\ADD_/FAINST[175].FA_/n1 ), .B(b[175]), 
        .Z(c[175]) );
  AND \ADD_/FAINST[175].FA_/U3  ( .A(\ADD_/FAINST[175].FA_/n1 ), .B(
        \ADD_/FAINST[175].FA_/n2 ), .Z(\ADD_/FAINST[175].FA_/n3 ) );
  XOR \ADD_/FAINST[175].FA_/U2  ( .A(b[175]), .B(\ADD_/c[175] ), .Z(
        \ADD_/FAINST[175].FA_/n2 ) );
  XOR \ADD_/FAINST[175].FA_/U1  ( .A(a[175]), .B(\ADD_/c[175] ), .Z(
        \ADD_/FAINST[175].FA_/n1 ) );
  XOR \ADD_/FAINST[174].FA_/U5  ( .A(\ADD_/FAINST[174].FA_/n3 ), .B(
        \ADD_/c[174] ), .Z(\ADD_/c[175] ) );
  XOR \ADD_/FAINST[174].FA_/U4  ( .A(\ADD_/FAINST[174].FA_/n1 ), .B(b[174]), 
        .Z(c[174]) );
  AND \ADD_/FAINST[174].FA_/U3  ( .A(\ADD_/FAINST[174].FA_/n1 ), .B(
        \ADD_/FAINST[174].FA_/n2 ), .Z(\ADD_/FAINST[174].FA_/n3 ) );
  XOR \ADD_/FAINST[174].FA_/U2  ( .A(b[174]), .B(\ADD_/c[174] ), .Z(
        \ADD_/FAINST[174].FA_/n2 ) );
  XOR \ADD_/FAINST[174].FA_/U1  ( .A(a[174]), .B(\ADD_/c[174] ), .Z(
        \ADD_/FAINST[174].FA_/n1 ) );
  XOR \ADD_/FAINST[173].FA_/U5  ( .A(\ADD_/FAINST[173].FA_/n3 ), .B(
        \ADD_/c[173] ), .Z(\ADD_/c[174] ) );
  XOR \ADD_/FAINST[173].FA_/U4  ( .A(\ADD_/FAINST[173].FA_/n1 ), .B(b[173]), 
        .Z(c[173]) );
  AND \ADD_/FAINST[173].FA_/U3  ( .A(\ADD_/FAINST[173].FA_/n1 ), .B(
        \ADD_/FAINST[173].FA_/n2 ), .Z(\ADD_/FAINST[173].FA_/n3 ) );
  XOR \ADD_/FAINST[173].FA_/U2  ( .A(b[173]), .B(\ADD_/c[173] ), .Z(
        \ADD_/FAINST[173].FA_/n2 ) );
  XOR \ADD_/FAINST[173].FA_/U1  ( .A(a[173]), .B(\ADD_/c[173] ), .Z(
        \ADD_/FAINST[173].FA_/n1 ) );
  XOR \ADD_/FAINST[172].FA_/U5  ( .A(\ADD_/FAINST[172].FA_/n3 ), .B(
        \ADD_/c[172] ), .Z(\ADD_/c[173] ) );
  XOR \ADD_/FAINST[172].FA_/U4  ( .A(\ADD_/FAINST[172].FA_/n1 ), .B(b[172]), 
        .Z(c[172]) );
  AND \ADD_/FAINST[172].FA_/U3  ( .A(\ADD_/FAINST[172].FA_/n1 ), .B(
        \ADD_/FAINST[172].FA_/n2 ), .Z(\ADD_/FAINST[172].FA_/n3 ) );
  XOR \ADD_/FAINST[172].FA_/U2  ( .A(b[172]), .B(\ADD_/c[172] ), .Z(
        \ADD_/FAINST[172].FA_/n2 ) );
  XOR \ADD_/FAINST[172].FA_/U1  ( .A(a[172]), .B(\ADD_/c[172] ), .Z(
        \ADD_/FAINST[172].FA_/n1 ) );
  XOR \ADD_/FAINST[171].FA_/U5  ( .A(\ADD_/FAINST[171].FA_/n3 ), .B(
        \ADD_/c[171] ), .Z(\ADD_/c[172] ) );
  XOR \ADD_/FAINST[171].FA_/U4  ( .A(\ADD_/FAINST[171].FA_/n1 ), .B(b[171]), 
        .Z(c[171]) );
  AND \ADD_/FAINST[171].FA_/U3  ( .A(\ADD_/FAINST[171].FA_/n1 ), .B(
        \ADD_/FAINST[171].FA_/n2 ), .Z(\ADD_/FAINST[171].FA_/n3 ) );
  XOR \ADD_/FAINST[171].FA_/U2  ( .A(b[171]), .B(\ADD_/c[171] ), .Z(
        \ADD_/FAINST[171].FA_/n2 ) );
  XOR \ADD_/FAINST[171].FA_/U1  ( .A(a[171]), .B(\ADD_/c[171] ), .Z(
        \ADD_/FAINST[171].FA_/n1 ) );
  XOR \ADD_/FAINST[170].FA_/U5  ( .A(\ADD_/FAINST[170].FA_/n3 ), .B(
        \ADD_/c[170] ), .Z(\ADD_/c[171] ) );
  XOR \ADD_/FAINST[170].FA_/U4  ( .A(\ADD_/FAINST[170].FA_/n1 ), .B(b[170]), 
        .Z(c[170]) );
  AND \ADD_/FAINST[170].FA_/U3  ( .A(\ADD_/FAINST[170].FA_/n1 ), .B(
        \ADD_/FAINST[170].FA_/n2 ), .Z(\ADD_/FAINST[170].FA_/n3 ) );
  XOR \ADD_/FAINST[170].FA_/U2  ( .A(b[170]), .B(\ADD_/c[170] ), .Z(
        \ADD_/FAINST[170].FA_/n2 ) );
  XOR \ADD_/FAINST[170].FA_/U1  ( .A(a[170]), .B(\ADD_/c[170] ), .Z(
        \ADD_/FAINST[170].FA_/n1 ) );
  XOR \ADD_/FAINST[169].FA_/U5  ( .A(\ADD_/FAINST[169].FA_/n3 ), .B(
        \ADD_/c[169] ), .Z(\ADD_/c[170] ) );
  XOR \ADD_/FAINST[169].FA_/U4  ( .A(\ADD_/FAINST[169].FA_/n1 ), .B(b[169]), 
        .Z(c[169]) );
  AND \ADD_/FAINST[169].FA_/U3  ( .A(\ADD_/FAINST[169].FA_/n1 ), .B(
        \ADD_/FAINST[169].FA_/n2 ), .Z(\ADD_/FAINST[169].FA_/n3 ) );
  XOR \ADD_/FAINST[169].FA_/U2  ( .A(b[169]), .B(\ADD_/c[169] ), .Z(
        \ADD_/FAINST[169].FA_/n2 ) );
  XOR \ADD_/FAINST[169].FA_/U1  ( .A(a[169]), .B(\ADD_/c[169] ), .Z(
        \ADD_/FAINST[169].FA_/n1 ) );
  XOR \ADD_/FAINST[168].FA_/U5  ( .A(\ADD_/FAINST[168].FA_/n3 ), .B(
        \ADD_/c[168] ), .Z(\ADD_/c[169] ) );
  XOR \ADD_/FAINST[168].FA_/U4  ( .A(\ADD_/FAINST[168].FA_/n1 ), .B(b[168]), 
        .Z(c[168]) );
  AND \ADD_/FAINST[168].FA_/U3  ( .A(\ADD_/FAINST[168].FA_/n1 ), .B(
        \ADD_/FAINST[168].FA_/n2 ), .Z(\ADD_/FAINST[168].FA_/n3 ) );
  XOR \ADD_/FAINST[168].FA_/U2  ( .A(b[168]), .B(\ADD_/c[168] ), .Z(
        \ADD_/FAINST[168].FA_/n2 ) );
  XOR \ADD_/FAINST[168].FA_/U1  ( .A(a[168]), .B(\ADD_/c[168] ), .Z(
        \ADD_/FAINST[168].FA_/n1 ) );
  XOR \ADD_/FAINST[167].FA_/U5  ( .A(\ADD_/FAINST[167].FA_/n3 ), .B(
        \ADD_/c[167] ), .Z(\ADD_/c[168] ) );
  XOR \ADD_/FAINST[167].FA_/U4  ( .A(\ADD_/FAINST[167].FA_/n1 ), .B(b[167]), 
        .Z(c[167]) );
  AND \ADD_/FAINST[167].FA_/U3  ( .A(\ADD_/FAINST[167].FA_/n1 ), .B(
        \ADD_/FAINST[167].FA_/n2 ), .Z(\ADD_/FAINST[167].FA_/n3 ) );
  XOR \ADD_/FAINST[167].FA_/U2  ( .A(b[167]), .B(\ADD_/c[167] ), .Z(
        \ADD_/FAINST[167].FA_/n2 ) );
  XOR \ADD_/FAINST[167].FA_/U1  ( .A(a[167]), .B(\ADD_/c[167] ), .Z(
        \ADD_/FAINST[167].FA_/n1 ) );
  XOR \ADD_/FAINST[166].FA_/U5  ( .A(\ADD_/FAINST[166].FA_/n3 ), .B(
        \ADD_/c[166] ), .Z(\ADD_/c[167] ) );
  XOR \ADD_/FAINST[166].FA_/U4  ( .A(\ADD_/FAINST[166].FA_/n1 ), .B(b[166]), 
        .Z(c[166]) );
  AND \ADD_/FAINST[166].FA_/U3  ( .A(\ADD_/FAINST[166].FA_/n1 ), .B(
        \ADD_/FAINST[166].FA_/n2 ), .Z(\ADD_/FAINST[166].FA_/n3 ) );
  XOR \ADD_/FAINST[166].FA_/U2  ( .A(b[166]), .B(\ADD_/c[166] ), .Z(
        \ADD_/FAINST[166].FA_/n2 ) );
  XOR \ADD_/FAINST[166].FA_/U1  ( .A(a[166]), .B(\ADD_/c[166] ), .Z(
        \ADD_/FAINST[166].FA_/n1 ) );
  XOR \ADD_/FAINST[165].FA_/U5  ( .A(\ADD_/FAINST[165].FA_/n3 ), .B(
        \ADD_/c[165] ), .Z(\ADD_/c[166] ) );
  XOR \ADD_/FAINST[165].FA_/U4  ( .A(\ADD_/FAINST[165].FA_/n1 ), .B(b[165]), 
        .Z(c[165]) );
  AND \ADD_/FAINST[165].FA_/U3  ( .A(\ADD_/FAINST[165].FA_/n1 ), .B(
        \ADD_/FAINST[165].FA_/n2 ), .Z(\ADD_/FAINST[165].FA_/n3 ) );
  XOR \ADD_/FAINST[165].FA_/U2  ( .A(b[165]), .B(\ADD_/c[165] ), .Z(
        \ADD_/FAINST[165].FA_/n2 ) );
  XOR \ADD_/FAINST[165].FA_/U1  ( .A(a[165]), .B(\ADD_/c[165] ), .Z(
        \ADD_/FAINST[165].FA_/n1 ) );
  XOR \ADD_/FAINST[164].FA_/U5  ( .A(\ADD_/FAINST[164].FA_/n3 ), .B(
        \ADD_/c[164] ), .Z(\ADD_/c[165] ) );
  XOR \ADD_/FAINST[164].FA_/U4  ( .A(\ADD_/FAINST[164].FA_/n1 ), .B(b[164]), 
        .Z(c[164]) );
  AND \ADD_/FAINST[164].FA_/U3  ( .A(\ADD_/FAINST[164].FA_/n1 ), .B(
        \ADD_/FAINST[164].FA_/n2 ), .Z(\ADD_/FAINST[164].FA_/n3 ) );
  XOR \ADD_/FAINST[164].FA_/U2  ( .A(b[164]), .B(\ADD_/c[164] ), .Z(
        \ADD_/FAINST[164].FA_/n2 ) );
  XOR \ADD_/FAINST[164].FA_/U1  ( .A(a[164]), .B(\ADD_/c[164] ), .Z(
        \ADD_/FAINST[164].FA_/n1 ) );
  XOR \ADD_/FAINST[163].FA_/U5  ( .A(\ADD_/FAINST[163].FA_/n3 ), .B(
        \ADD_/c[163] ), .Z(\ADD_/c[164] ) );
  XOR \ADD_/FAINST[163].FA_/U4  ( .A(\ADD_/FAINST[163].FA_/n1 ), .B(b[163]), 
        .Z(c[163]) );
  AND \ADD_/FAINST[163].FA_/U3  ( .A(\ADD_/FAINST[163].FA_/n1 ), .B(
        \ADD_/FAINST[163].FA_/n2 ), .Z(\ADD_/FAINST[163].FA_/n3 ) );
  XOR \ADD_/FAINST[163].FA_/U2  ( .A(b[163]), .B(\ADD_/c[163] ), .Z(
        \ADD_/FAINST[163].FA_/n2 ) );
  XOR \ADD_/FAINST[163].FA_/U1  ( .A(a[163]), .B(\ADD_/c[163] ), .Z(
        \ADD_/FAINST[163].FA_/n1 ) );
  XOR \ADD_/FAINST[162].FA_/U5  ( .A(\ADD_/FAINST[162].FA_/n3 ), .B(
        \ADD_/c[162] ), .Z(\ADD_/c[163] ) );
  XOR \ADD_/FAINST[162].FA_/U4  ( .A(\ADD_/FAINST[162].FA_/n1 ), .B(b[162]), 
        .Z(c[162]) );
  AND \ADD_/FAINST[162].FA_/U3  ( .A(\ADD_/FAINST[162].FA_/n1 ), .B(
        \ADD_/FAINST[162].FA_/n2 ), .Z(\ADD_/FAINST[162].FA_/n3 ) );
  XOR \ADD_/FAINST[162].FA_/U2  ( .A(b[162]), .B(\ADD_/c[162] ), .Z(
        \ADD_/FAINST[162].FA_/n2 ) );
  XOR \ADD_/FAINST[162].FA_/U1  ( .A(a[162]), .B(\ADD_/c[162] ), .Z(
        \ADD_/FAINST[162].FA_/n1 ) );
  XOR \ADD_/FAINST[161].FA_/U5  ( .A(\ADD_/FAINST[161].FA_/n3 ), .B(
        \ADD_/c[161] ), .Z(\ADD_/c[162] ) );
  XOR \ADD_/FAINST[161].FA_/U4  ( .A(\ADD_/FAINST[161].FA_/n1 ), .B(b[161]), 
        .Z(c[161]) );
  AND \ADD_/FAINST[161].FA_/U3  ( .A(\ADD_/FAINST[161].FA_/n1 ), .B(
        \ADD_/FAINST[161].FA_/n2 ), .Z(\ADD_/FAINST[161].FA_/n3 ) );
  XOR \ADD_/FAINST[161].FA_/U2  ( .A(b[161]), .B(\ADD_/c[161] ), .Z(
        \ADD_/FAINST[161].FA_/n2 ) );
  XOR \ADD_/FAINST[161].FA_/U1  ( .A(a[161]), .B(\ADD_/c[161] ), .Z(
        \ADD_/FAINST[161].FA_/n1 ) );
  XOR \ADD_/FAINST[160].FA_/U5  ( .A(\ADD_/FAINST[160].FA_/n3 ), .B(
        \ADD_/c[160] ), .Z(\ADD_/c[161] ) );
  XOR \ADD_/FAINST[160].FA_/U4  ( .A(\ADD_/FAINST[160].FA_/n1 ), .B(b[160]), 
        .Z(c[160]) );
  AND \ADD_/FAINST[160].FA_/U3  ( .A(\ADD_/FAINST[160].FA_/n1 ), .B(
        \ADD_/FAINST[160].FA_/n2 ), .Z(\ADD_/FAINST[160].FA_/n3 ) );
  XOR \ADD_/FAINST[160].FA_/U2  ( .A(b[160]), .B(\ADD_/c[160] ), .Z(
        \ADD_/FAINST[160].FA_/n2 ) );
  XOR \ADD_/FAINST[160].FA_/U1  ( .A(a[160]), .B(\ADD_/c[160] ), .Z(
        \ADD_/FAINST[160].FA_/n1 ) );
  XOR \ADD_/FAINST[159].FA_/U5  ( .A(\ADD_/FAINST[159].FA_/n3 ), .B(
        \ADD_/c[159] ), .Z(\ADD_/c[160] ) );
  XOR \ADD_/FAINST[159].FA_/U4  ( .A(\ADD_/FAINST[159].FA_/n1 ), .B(b[159]), 
        .Z(c[159]) );
  AND \ADD_/FAINST[159].FA_/U3  ( .A(\ADD_/FAINST[159].FA_/n1 ), .B(
        \ADD_/FAINST[159].FA_/n2 ), .Z(\ADD_/FAINST[159].FA_/n3 ) );
  XOR \ADD_/FAINST[159].FA_/U2  ( .A(b[159]), .B(\ADD_/c[159] ), .Z(
        \ADD_/FAINST[159].FA_/n2 ) );
  XOR \ADD_/FAINST[159].FA_/U1  ( .A(a[159]), .B(\ADD_/c[159] ), .Z(
        \ADD_/FAINST[159].FA_/n1 ) );
  XOR \ADD_/FAINST[158].FA_/U5  ( .A(\ADD_/FAINST[158].FA_/n3 ), .B(
        \ADD_/c[158] ), .Z(\ADD_/c[159] ) );
  XOR \ADD_/FAINST[158].FA_/U4  ( .A(\ADD_/FAINST[158].FA_/n1 ), .B(b[158]), 
        .Z(c[158]) );
  AND \ADD_/FAINST[158].FA_/U3  ( .A(\ADD_/FAINST[158].FA_/n1 ), .B(
        \ADD_/FAINST[158].FA_/n2 ), .Z(\ADD_/FAINST[158].FA_/n3 ) );
  XOR \ADD_/FAINST[158].FA_/U2  ( .A(b[158]), .B(\ADD_/c[158] ), .Z(
        \ADD_/FAINST[158].FA_/n2 ) );
  XOR \ADD_/FAINST[158].FA_/U1  ( .A(a[158]), .B(\ADD_/c[158] ), .Z(
        \ADD_/FAINST[158].FA_/n1 ) );
  XOR \ADD_/FAINST[157].FA_/U5  ( .A(\ADD_/FAINST[157].FA_/n3 ), .B(
        \ADD_/c[157] ), .Z(\ADD_/c[158] ) );
  XOR \ADD_/FAINST[157].FA_/U4  ( .A(\ADD_/FAINST[157].FA_/n1 ), .B(b[157]), 
        .Z(c[157]) );
  AND \ADD_/FAINST[157].FA_/U3  ( .A(\ADD_/FAINST[157].FA_/n1 ), .B(
        \ADD_/FAINST[157].FA_/n2 ), .Z(\ADD_/FAINST[157].FA_/n3 ) );
  XOR \ADD_/FAINST[157].FA_/U2  ( .A(b[157]), .B(\ADD_/c[157] ), .Z(
        \ADD_/FAINST[157].FA_/n2 ) );
  XOR \ADD_/FAINST[157].FA_/U1  ( .A(a[157]), .B(\ADD_/c[157] ), .Z(
        \ADD_/FAINST[157].FA_/n1 ) );
  XOR \ADD_/FAINST[156].FA_/U5  ( .A(\ADD_/FAINST[156].FA_/n3 ), .B(
        \ADD_/c[156] ), .Z(\ADD_/c[157] ) );
  XOR \ADD_/FAINST[156].FA_/U4  ( .A(\ADD_/FAINST[156].FA_/n1 ), .B(b[156]), 
        .Z(c[156]) );
  AND \ADD_/FAINST[156].FA_/U3  ( .A(\ADD_/FAINST[156].FA_/n1 ), .B(
        \ADD_/FAINST[156].FA_/n2 ), .Z(\ADD_/FAINST[156].FA_/n3 ) );
  XOR \ADD_/FAINST[156].FA_/U2  ( .A(b[156]), .B(\ADD_/c[156] ), .Z(
        \ADD_/FAINST[156].FA_/n2 ) );
  XOR \ADD_/FAINST[156].FA_/U1  ( .A(a[156]), .B(\ADD_/c[156] ), .Z(
        \ADD_/FAINST[156].FA_/n1 ) );
  XOR \ADD_/FAINST[155].FA_/U5  ( .A(\ADD_/FAINST[155].FA_/n3 ), .B(
        \ADD_/c[155] ), .Z(\ADD_/c[156] ) );
  XOR \ADD_/FAINST[155].FA_/U4  ( .A(\ADD_/FAINST[155].FA_/n1 ), .B(b[155]), 
        .Z(c[155]) );
  AND \ADD_/FAINST[155].FA_/U3  ( .A(\ADD_/FAINST[155].FA_/n1 ), .B(
        \ADD_/FAINST[155].FA_/n2 ), .Z(\ADD_/FAINST[155].FA_/n3 ) );
  XOR \ADD_/FAINST[155].FA_/U2  ( .A(b[155]), .B(\ADD_/c[155] ), .Z(
        \ADD_/FAINST[155].FA_/n2 ) );
  XOR \ADD_/FAINST[155].FA_/U1  ( .A(a[155]), .B(\ADD_/c[155] ), .Z(
        \ADD_/FAINST[155].FA_/n1 ) );
  XOR \ADD_/FAINST[154].FA_/U5  ( .A(\ADD_/FAINST[154].FA_/n3 ), .B(
        \ADD_/c[154] ), .Z(\ADD_/c[155] ) );
  XOR \ADD_/FAINST[154].FA_/U4  ( .A(\ADD_/FAINST[154].FA_/n1 ), .B(b[154]), 
        .Z(c[154]) );
  AND \ADD_/FAINST[154].FA_/U3  ( .A(\ADD_/FAINST[154].FA_/n1 ), .B(
        \ADD_/FAINST[154].FA_/n2 ), .Z(\ADD_/FAINST[154].FA_/n3 ) );
  XOR \ADD_/FAINST[154].FA_/U2  ( .A(b[154]), .B(\ADD_/c[154] ), .Z(
        \ADD_/FAINST[154].FA_/n2 ) );
  XOR \ADD_/FAINST[154].FA_/U1  ( .A(a[154]), .B(\ADD_/c[154] ), .Z(
        \ADD_/FAINST[154].FA_/n1 ) );
  XOR \ADD_/FAINST[153].FA_/U5  ( .A(\ADD_/FAINST[153].FA_/n3 ), .B(
        \ADD_/c[153] ), .Z(\ADD_/c[154] ) );
  XOR \ADD_/FAINST[153].FA_/U4  ( .A(\ADD_/FAINST[153].FA_/n1 ), .B(b[153]), 
        .Z(c[153]) );
  AND \ADD_/FAINST[153].FA_/U3  ( .A(\ADD_/FAINST[153].FA_/n1 ), .B(
        \ADD_/FAINST[153].FA_/n2 ), .Z(\ADD_/FAINST[153].FA_/n3 ) );
  XOR \ADD_/FAINST[153].FA_/U2  ( .A(b[153]), .B(\ADD_/c[153] ), .Z(
        \ADD_/FAINST[153].FA_/n2 ) );
  XOR \ADD_/FAINST[153].FA_/U1  ( .A(a[153]), .B(\ADD_/c[153] ), .Z(
        \ADD_/FAINST[153].FA_/n1 ) );
  XOR \ADD_/FAINST[152].FA_/U5  ( .A(\ADD_/FAINST[152].FA_/n3 ), .B(
        \ADD_/c[152] ), .Z(\ADD_/c[153] ) );
  XOR \ADD_/FAINST[152].FA_/U4  ( .A(\ADD_/FAINST[152].FA_/n1 ), .B(b[152]), 
        .Z(c[152]) );
  AND \ADD_/FAINST[152].FA_/U3  ( .A(\ADD_/FAINST[152].FA_/n1 ), .B(
        \ADD_/FAINST[152].FA_/n2 ), .Z(\ADD_/FAINST[152].FA_/n3 ) );
  XOR \ADD_/FAINST[152].FA_/U2  ( .A(b[152]), .B(\ADD_/c[152] ), .Z(
        \ADD_/FAINST[152].FA_/n2 ) );
  XOR \ADD_/FAINST[152].FA_/U1  ( .A(a[152]), .B(\ADD_/c[152] ), .Z(
        \ADD_/FAINST[152].FA_/n1 ) );
  XOR \ADD_/FAINST[151].FA_/U5  ( .A(\ADD_/FAINST[151].FA_/n3 ), .B(
        \ADD_/c[151] ), .Z(\ADD_/c[152] ) );
  XOR \ADD_/FAINST[151].FA_/U4  ( .A(\ADD_/FAINST[151].FA_/n1 ), .B(b[151]), 
        .Z(c[151]) );
  AND \ADD_/FAINST[151].FA_/U3  ( .A(\ADD_/FAINST[151].FA_/n1 ), .B(
        \ADD_/FAINST[151].FA_/n2 ), .Z(\ADD_/FAINST[151].FA_/n3 ) );
  XOR \ADD_/FAINST[151].FA_/U2  ( .A(b[151]), .B(\ADD_/c[151] ), .Z(
        \ADD_/FAINST[151].FA_/n2 ) );
  XOR \ADD_/FAINST[151].FA_/U1  ( .A(a[151]), .B(\ADD_/c[151] ), .Z(
        \ADD_/FAINST[151].FA_/n1 ) );
  XOR \ADD_/FAINST[150].FA_/U5  ( .A(\ADD_/FAINST[150].FA_/n3 ), .B(
        \ADD_/c[150] ), .Z(\ADD_/c[151] ) );
  XOR \ADD_/FAINST[150].FA_/U4  ( .A(\ADD_/FAINST[150].FA_/n1 ), .B(b[150]), 
        .Z(c[150]) );
  AND \ADD_/FAINST[150].FA_/U3  ( .A(\ADD_/FAINST[150].FA_/n1 ), .B(
        \ADD_/FAINST[150].FA_/n2 ), .Z(\ADD_/FAINST[150].FA_/n3 ) );
  XOR \ADD_/FAINST[150].FA_/U2  ( .A(b[150]), .B(\ADD_/c[150] ), .Z(
        \ADD_/FAINST[150].FA_/n2 ) );
  XOR \ADD_/FAINST[150].FA_/U1  ( .A(a[150]), .B(\ADD_/c[150] ), .Z(
        \ADD_/FAINST[150].FA_/n1 ) );
  XOR \ADD_/FAINST[149].FA_/U5  ( .A(\ADD_/FAINST[149].FA_/n3 ), .B(
        \ADD_/c[149] ), .Z(\ADD_/c[150] ) );
  XOR \ADD_/FAINST[149].FA_/U4  ( .A(\ADD_/FAINST[149].FA_/n1 ), .B(b[149]), 
        .Z(c[149]) );
  AND \ADD_/FAINST[149].FA_/U3  ( .A(\ADD_/FAINST[149].FA_/n1 ), .B(
        \ADD_/FAINST[149].FA_/n2 ), .Z(\ADD_/FAINST[149].FA_/n3 ) );
  XOR \ADD_/FAINST[149].FA_/U2  ( .A(b[149]), .B(\ADD_/c[149] ), .Z(
        \ADD_/FAINST[149].FA_/n2 ) );
  XOR \ADD_/FAINST[149].FA_/U1  ( .A(a[149]), .B(\ADD_/c[149] ), .Z(
        \ADD_/FAINST[149].FA_/n1 ) );
  XOR \ADD_/FAINST[148].FA_/U5  ( .A(\ADD_/FAINST[148].FA_/n3 ), .B(
        \ADD_/c[148] ), .Z(\ADD_/c[149] ) );
  XOR \ADD_/FAINST[148].FA_/U4  ( .A(\ADD_/FAINST[148].FA_/n1 ), .B(b[148]), 
        .Z(c[148]) );
  AND \ADD_/FAINST[148].FA_/U3  ( .A(\ADD_/FAINST[148].FA_/n1 ), .B(
        \ADD_/FAINST[148].FA_/n2 ), .Z(\ADD_/FAINST[148].FA_/n3 ) );
  XOR \ADD_/FAINST[148].FA_/U2  ( .A(b[148]), .B(\ADD_/c[148] ), .Z(
        \ADD_/FAINST[148].FA_/n2 ) );
  XOR \ADD_/FAINST[148].FA_/U1  ( .A(a[148]), .B(\ADD_/c[148] ), .Z(
        \ADD_/FAINST[148].FA_/n1 ) );
  XOR \ADD_/FAINST[147].FA_/U5  ( .A(\ADD_/FAINST[147].FA_/n3 ), .B(
        \ADD_/c[147] ), .Z(\ADD_/c[148] ) );
  XOR \ADD_/FAINST[147].FA_/U4  ( .A(\ADD_/FAINST[147].FA_/n1 ), .B(b[147]), 
        .Z(c[147]) );
  AND \ADD_/FAINST[147].FA_/U3  ( .A(\ADD_/FAINST[147].FA_/n1 ), .B(
        \ADD_/FAINST[147].FA_/n2 ), .Z(\ADD_/FAINST[147].FA_/n3 ) );
  XOR \ADD_/FAINST[147].FA_/U2  ( .A(b[147]), .B(\ADD_/c[147] ), .Z(
        \ADD_/FAINST[147].FA_/n2 ) );
  XOR \ADD_/FAINST[147].FA_/U1  ( .A(a[147]), .B(\ADD_/c[147] ), .Z(
        \ADD_/FAINST[147].FA_/n1 ) );
  XOR \ADD_/FAINST[146].FA_/U5  ( .A(\ADD_/FAINST[146].FA_/n3 ), .B(
        \ADD_/c[146] ), .Z(\ADD_/c[147] ) );
  XOR \ADD_/FAINST[146].FA_/U4  ( .A(\ADD_/FAINST[146].FA_/n1 ), .B(b[146]), 
        .Z(c[146]) );
  AND \ADD_/FAINST[146].FA_/U3  ( .A(\ADD_/FAINST[146].FA_/n1 ), .B(
        \ADD_/FAINST[146].FA_/n2 ), .Z(\ADD_/FAINST[146].FA_/n3 ) );
  XOR \ADD_/FAINST[146].FA_/U2  ( .A(b[146]), .B(\ADD_/c[146] ), .Z(
        \ADD_/FAINST[146].FA_/n2 ) );
  XOR \ADD_/FAINST[146].FA_/U1  ( .A(a[146]), .B(\ADD_/c[146] ), .Z(
        \ADD_/FAINST[146].FA_/n1 ) );
  XOR \ADD_/FAINST[145].FA_/U5  ( .A(\ADD_/FAINST[145].FA_/n3 ), .B(
        \ADD_/c[145] ), .Z(\ADD_/c[146] ) );
  XOR \ADD_/FAINST[145].FA_/U4  ( .A(\ADD_/FAINST[145].FA_/n1 ), .B(b[145]), 
        .Z(c[145]) );
  AND \ADD_/FAINST[145].FA_/U3  ( .A(\ADD_/FAINST[145].FA_/n1 ), .B(
        \ADD_/FAINST[145].FA_/n2 ), .Z(\ADD_/FAINST[145].FA_/n3 ) );
  XOR \ADD_/FAINST[145].FA_/U2  ( .A(b[145]), .B(\ADD_/c[145] ), .Z(
        \ADD_/FAINST[145].FA_/n2 ) );
  XOR \ADD_/FAINST[145].FA_/U1  ( .A(a[145]), .B(\ADD_/c[145] ), .Z(
        \ADD_/FAINST[145].FA_/n1 ) );
  XOR \ADD_/FAINST[144].FA_/U5  ( .A(\ADD_/FAINST[144].FA_/n3 ), .B(
        \ADD_/c[144] ), .Z(\ADD_/c[145] ) );
  XOR \ADD_/FAINST[144].FA_/U4  ( .A(\ADD_/FAINST[144].FA_/n1 ), .B(b[144]), 
        .Z(c[144]) );
  AND \ADD_/FAINST[144].FA_/U3  ( .A(\ADD_/FAINST[144].FA_/n1 ), .B(
        \ADD_/FAINST[144].FA_/n2 ), .Z(\ADD_/FAINST[144].FA_/n3 ) );
  XOR \ADD_/FAINST[144].FA_/U2  ( .A(b[144]), .B(\ADD_/c[144] ), .Z(
        \ADD_/FAINST[144].FA_/n2 ) );
  XOR \ADD_/FAINST[144].FA_/U1  ( .A(a[144]), .B(\ADD_/c[144] ), .Z(
        \ADD_/FAINST[144].FA_/n1 ) );
  XOR \ADD_/FAINST[143].FA_/U5  ( .A(\ADD_/FAINST[143].FA_/n3 ), .B(
        \ADD_/c[143] ), .Z(\ADD_/c[144] ) );
  XOR \ADD_/FAINST[143].FA_/U4  ( .A(\ADD_/FAINST[143].FA_/n1 ), .B(b[143]), 
        .Z(c[143]) );
  AND \ADD_/FAINST[143].FA_/U3  ( .A(\ADD_/FAINST[143].FA_/n1 ), .B(
        \ADD_/FAINST[143].FA_/n2 ), .Z(\ADD_/FAINST[143].FA_/n3 ) );
  XOR \ADD_/FAINST[143].FA_/U2  ( .A(b[143]), .B(\ADD_/c[143] ), .Z(
        \ADD_/FAINST[143].FA_/n2 ) );
  XOR \ADD_/FAINST[143].FA_/U1  ( .A(a[143]), .B(\ADD_/c[143] ), .Z(
        \ADD_/FAINST[143].FA_/n1 ) );
  XOR \ADD_/FAINST[142].FA_/U5  ( .A(\ADD_/FAINST[142].FA_/n3 ), .B(
        \ADD_/c[142] ), .Z(\ADD_/c[143] ) );
  XOR \ADD_/FAINST[142].FA_/U4  ( .A(\ADD_/FAINST[142].FA_/n1 ), .B(b[142]), 
        .Z(c[142]) );
  AND \ADD_/FAINST[142].FA_/U3  ( .A(\ADD_/FAINST[142].FA_/n1 ), .B(
        \ADD_/FAINST[142].FA_/n2 ), .Z(\ADD_/FAINST[142].FA_/n3 ) );
  XOR \ADD_/FAINST[142].FA_/U2  ( .A(b[142]), .B(\ADD_/c[142] ), .Z(
        \ADD_/FAINST[142].FA_/n2 ) );
  XOR \ADD_/FAINST[142].FA_/U1  ( .A(a[142]), .B(\ADD_/c[142] ), .Z(
        \ADD_/FAINST[142].FA_/n1 ) );
  XOR \ADD_/FAINST[141].FA_/U5  ( .A(\ADD_/FAINST[141].FA_/n3 ), .B(
        \ADD_/c[141] ), .Z(\ADD_/c[142] ) );
  XOR \ADD_/FAINST[141].FA_/U4  ( .A(\ADD_/FAINST[141].FA_/n1 ), .B(b[141]), 
        .Z(c[141]) );
  AND \ADD_/FAINST[141].FA_/U3  ( .A(\ADD_/FAINST[141].FA_/n1 ), .B(
        \ADD_/FAINST[141].FA_/n2 ), .Z(\ADD_/FAINST[141].FA_/n3 ) );
  XOR \ADD_/FAINST[141].FA_/U2  ( .A(b[141]), .B(\ADD_/c[141] ), .Z(
        \ADD_/FAINST[141].FA_/n2 ) );
  XOR \ADD_/FAINST[141].FA_/U1  ( .A(a[141]), .B(\ADD_/c[141] ), .Z(
        \ADD_/FAINST[141].FA_/n1 ) );
  XOR \ADD_/FAINST[140].FA_/U5  ( .A(\ADD_/FAINST[140].FA_/n3 ), .B(
        \ADD_/c[140] ), .Z(\ADD_/c[141] ) );
  XOR \ADD_/FAINST[140].FA_/U4  ( .A(\ADD_/FAINST[140].FA_/n1 ), .B(b[140]), 
        .Z(c[140]) );
  AND \ADD_/FAINST[140].FA_/U3  ( .A(\ADD_/FAINST[140].FA_/n1 ), .B(
        \ADD_/FAINST[140].FA_/n2 ), .Z(\ADD_/FAINST[140].FA_/n3 ) );
  XOR \ADD_/FAINST[140].FA_/U2  ( .A(b[140]), .B(\ADD_/c[140] ), .Z(
        \ADD_/FAINST[140].FA_/n2 ) );
  XOR \ADD_/FAINST[140].FA_/U1  ( .A(a[140]), .B(\ADD_/c[140] ), .Z(
        \ADD_/FAINST[140].FA_/n1 ) );
  XOR \ADD_/FAINST[139].FA_/U5  ( .A(\ADD_/FAINST[139].FA_/n3 ), .B(
        \ADD_/c[139] ), .Z(\ADD_/c[140] ) );
  XOR \ADD_/FAINST[139].FA_/U4  ( .A(\ADD_/FAINST[139].FA_/n1 ), .B(b[139]), 
        .Z(c[139]) );
  AND \ADD_/FAINST[139].FA_/U3  ( .A(\ADD_/FAINST[139].FA_/n1 ), .B(
        \ADD_/FAINST[139].FA_/n2 ), .Z(\ADD_/FAINST[139].FA_/n3 ) );
  XOR \ADD_/FAINST[139].FA_/U2  ( .A(b[139]), .B(\ADD_/c[139] ), .Z(
        \ADD_/FAINST[139].FA_/n2 ) );
  XOR \ADD_/FAINST[139].FA_/U1  ( .A(a[139]), .B(\ADD_/c[139] ), .Z(
        \ADD_/FAINST[139].FA_/n1 ) );
  XOR \ADD_/FAINST[138].FA_/U5  ( .A(\ADD_/FAINST[138].FA_/n3 ), .B(
        \ADD_/c[138] ), .Z(\ADD_/c[139] ) );
  XOR \ADD_/FAINST[138].FA_/U4  ( .A(\ADD_/FAINST[138].FA_/n1 ), .B(b[138]), 
        .Z(c[138]) );
  AND \ADD_/FAINST[138].FA_/U3  ( .A(\ADD_/FAINST[138].FA_/n1 ), .B(
        \ADD_/FAINST[138].FA_/n2 ), .Z(\ADD_/FAINST[138].FA_/n3 ) );
  XOR \ADD_/FAINST[138].FA_/U2  ( .A(b[138]), .B(\ADD_/c[138] ), .Z(
        \ADD_/FAINST[138].FA_/n2 ) );
  XOR \ADD_/FAINST[138].FA_/U1  ( .A(a[138]), .B(\ADD_/c[138] ), .Z(
        \ADD_/FAINST[138].FA_/n1 ) );
  XOR \ADD_/FAINST[137].FA_/U5  ( .A(\ADD_/FAINST[137].FA_/n3 ), .B(
        \ADD_/c[137] ), .Z(\ADD_/c[138] ) );
  XOR \ADD_/FAINST[137].FA_/U4  ( .A(\ADD_/FAINST[137].FA_/n1 ), .B(b[137]), 
        .Z(c[137]) );
  AND \ADD_/FAINST[137].FA_/U3  ( .A(\ADD_/FAINST[137].FA_/n1 ), .B(
        \ADD_/FAINST[137].FA_/n2 ), .Z(\ADD_/FAINST[137].FA_/n3 ) );
  XOR \ADD_/FAINST[137].FA_/U2  ( .A(b[137]), .B(\ADD_/c[137] ), .Z(
        \ADD_/FAINST[137].FA_/n2 ) );
  XOR \ADD_/FAINST[137].FA_/U1  ( .A(a[137]), .B(\ADD_/c[137] ), .Z(
        \ADD_/FAINST[137].FA_/n1 ) );
  XOR \ADD_/FAINST[136].FA_/U5  ( .A(\ADD_/FAINST[136].FA_/n3 ), .B(
        \ADD_/c[136] ), .Z(\ADD_/c[137] ) );
  XOR \ADD_/FAINST[136].FA_/U4  ( .A(\ADD_/FAINST[136].FA_/n1 ), .B(b[136]), 
        .Z(c[136]) );
  AND \ADD_/FAINST[136].FA_/U3  ( .A(\ADD_/FAINST[136].FA_/n1 ), .B(
        \ADD_/FAINST[136].FA_/n2 ), .Z(\ADD_/FAINST[136].FA_/n3 ) );
  XOR \ADD_/FAINST[136].FA_/U2  ( .A(b[136]), .B(\ADD_/c[136] ), .Z(
        \ADD_/FAINST[136].FA_/n2 ) );
  XOR \ADD_/FAINST[136].FA_/U1  ( .A(a[136]), .B(\ADD_/c[136] ), .Z(
        \ADD_/FAINST[136].FA_/n1 ) );
  XOR \ADD_/FAINST[135].FA_/U5  ( .A(\ADD_/FAINST[135].FA_/n3 ), .B(
        \ADD_/c[135] ), .Z(\ADD_/c[136] ) );
  XOR \ADD_/FAINST[135].FA_/U4  ( .A(\ADD_/FAINST[135].FA_/n1 ), .B(b[135]), 
        .Z(c[135]) );
  AND \ADD_/FAINST[135].FA_/U3  ( .A(\ADD_/FAINST[135].FA_/n1 ), .B(
        \ADD_/FAINST[135].FA_/n2 ), .Z(\ADD_/FAINST[135].FA_/n3 ) );
  XOR \ADD_/FAINST[135].FA_/U2  ( .A(b[135]), .B(\ADD_/c[135] ), .Z(
        \ADD_/FAINST[135].FA_/n2 ) );
  XOR \ADD_/FAINST[135].FA_/U1  ( .A(a[135]), .B(\ADD_/c[135] ), .Z(
        \ADD_/FAINST[135].FA_/n1 ) );
  XOR \ADD_/FAINST[134].FA_/U5  ( .A(\ADD_/FAINST[134].FA_/n3 ), .B(
        \ADD_/c[134] ), .Z(\ADD_/c[135] ) );
  XOR \ADD_/FAINST[134].FA_/U4  ( .A(\ADD_/FAINST[134].FA_/n1 ), .B(b[134]), 
        .Z(c[134]) );
  AND \ADD_/FAINST[134].FA_/U3  ( .A(\ADD_/FAINST[134].FA_/n1 ), .B(
        \ADD_/FAINST[134].FA_/n2 ), .Z(\ADD_/FAINST[134].FA_/n3 ) );
  XOR \ADD_/FAINST[134].FA_/U2  ( .A(b[134]), .B(\ADD_/c[134] ), .Z(
        \ADD_/FAINST[134].FA_/n2 ) );
  XOR \ADD_/FAINST[134].FA_/U1  ( .A(a[134]), .B(\ADD_/c[134] ), .Z(
        \ADD_/FAINST[134].FA_/n1 ) );
  XOR \ADD_/FAINST[133].FA_/U5  ( .A(\ADD_/FAINST[133].FA_/n3 ), .B(
        \ADD_/c[133] ), .Z(\ADD_/c[134] ) );
  XOR \ADD_/FAINST[133].FA_/U4  ( .A(\ADD_/FAINST[133].FA_/n1 ), .B(b[133]), 
        .Z(c[133]) );
  AND \ADD_/FAINST[133].FA_/U3  ( .A(\ADD_/FAINST[133].FA_/n1 ), .B(
        \ADD_/FAINST[133].FA_/n2 ), .Z(\ADD_/FAINST[133].FA_/n3 ) );
  XOR \ADD_/FAINST[133].FA_/U2  ( .A(b[133]), .B(\ADD_/c[133] ), .Z(
        \ADD_/FAINST[133].FA_/n2 ) );
  XOR \ADD_/FAINST[133].FA_/U1  ( .A(a[133]), .B(\ADD_/c[133] ), .Z(
        \ADD_/FAINST[133].FA_/n1 ) );
  XOR \ADD_/FAINST[132].FA_/U5  ( .A(\ADD_/FAINST[132].FA_/n3 ), .B(
        \ADD_/c[132] ), .Z(\ADD_/c[133] ) );
  XOR \ADD_/FAINST[132].FA_/U4  ( .A(\ADD_/FAINST[132].FA_/n1 ), .B(b[132]), 
        .Z(c[132]) );
  AND \ADD_/FAINST[132].FA_/U3  ( .A(\ADD_/FAINST[132].FA_/n1 ), .B(
        \ADD_/FAINST[132].FA_/n2 ), .Z(\ADD_/FAINST[132].FA_/n3 ) );
  XOR \ADD_/FAINST[132].FA_/U2  ( .A(b[132]), .B(\ADD_/c[132] ), .Z(
        \ADD_/FAINST[132].FA_/n2 ) );
  XOR \ADD_/FAINST[132].FA_/U1  ( .A(a[132]), .B(\ADD_/c[132] ), .Z(
        \ADD_/FAINST[132].FA_/n1 ) );
  XOR \ADD_/FAINST[131].FA_/U5  ( .A(\ADD_/FAINST[131].FA_/n3 ), .B(
        \ADD_/c[131] ), .Z(\ADD_/c[132] ) );
  XOR \ADD_/FAINST[131].FA_/U4  ( .A(\ADD_/FAINST[131].FA_/n1 ), .B(b[131]), 
        .Z(c[131]) );
  AND \ADD_/FAINST[131].FA_/U3  ( .A(\ADD_/FAINST[131].FA_/n1 ), .B(
        \ADD_/FAINST[131].FA_/n2 ), .Z(\ADD_/FAINST[131].FA_/n3 ) );
  XOR \ADD_/FAINST[131].FA_/U2  ( .A(b[131]), .B(\ADD_/c[131] ), .Z(
        \ADD_/FAINST[131].FA_/n2 ) );
  XOR \ADD_/FAINST[131].FA_/U1  ( .A(a[131]), .B(\ADD_/c[131] ), .Z(
        \ADD_/FAINST[131].FA_/n1 ) );
  XOR \ADD_/FAINST[130].FA_/U5  ( .A(\ADD_/FAINST[130].FA_/n3 ), .B(
        \ADD_/c[130] ), .Z(\ADD_/c[131] ) );
  XOR \ADD_/FAINST[130].FA_/U4  ( .A(\ADD_/FAINST[130].FA_/n1 ), .B(b[130]), 
        .Z(c[130]) );
  AND \ADD_/FAINST[130].FA_/U3  ( .A(\ADD_/FAINST[130].FA_/n1 ), .B(
        \ADD_/FAINST[130].FA_/n2 ), .Z(\ADD_/FAINST[130].FA_/n3 ) );
  XOR \ADD_/FAINST[130].FA_/U2  ( .A(b[130]), .B(\ADD_/c[130] ), .Z(
        \ADD_/FAINST[130].FA_/n2 ) );
  XOR \ADD_/FAINST[130].FA_/U1  ( .A(a[130]), .B(\ADD_/c[130] ), .Z(
        \ADD_/FAINST[130].FA_/n1 ) );
  XOR \ADD_/FAINST[129].FA_/U5  ( .A(\ADD_/FAINST[129].FA_/n3 ), .B(
        \ADD_/c[129] ), .Z(\ADD_/c[130] ) );
  XOR \ADD_/FAINST[129].FA_/U4  ( .A(\ADD_/FAINST[129].FA_/n1 ), .B(b[129]), 
        .Z(c[129]) );
  AND \ADD_/FAINST[129].FA_/U3  ( .A(\ADD_/FAINST[129].FA_/n1 ), .B(
        \ADD_/FAINST[129].FA_/n2 ), .Z(\ADD_/FAINST[129].FA_/n3 ) );
  XOR \ADD_/FAINST[129].FA_/U2  ( .A(b[129]), .B(\ADD_/c[129] ), .Z(
        \ADD_/FAINST[129].FA_/n2 ) );
  XOR \ADD_/FAINST[129].FA_/U1  ( .A(a[129]), .B(\ADD_/c[129] ), .Z(
        \ADD_/FAINST[129].FA_/n1 ) );
  XOR \ADD_/FAINST[128].FA_/U5  ( .A(\ADD_/FAINST[128].FA_/n3 ), .B(
        \ADD_/c[128] ), .Z(\ADD_/c[129] ) );
  XOR \ADD_/FAINST[128].FA_/U4  ( .A(\ADD_/FAINST[128].FA_/n1 ), .B(b[128]), 
        .Z(c[128]) );
  AND \ADD_/FAINST[128].FA_/U3  ( .A(\ADD_/FAINST[128].FA_/n1 ), .B(
        \ADD_/FAINST[128].FA_/n2 ), .Z(\ADD_/FAINST[128].FA_/n3 ) );
  XOR \ADD_/FAINST[128].FA_/U2  ( .A(b[128]), .B(\ADD_/c[128] ), .Z(
        \ADD_/FAINST[128].FA_/n2 ) );
  XOR \ADD_/FAINST[128].FA_/U1  ( .A(a[128]), .B(\ADD_/c[128] ), .Z(
        \ADD_/FAINST[128].FA_/n1 ) );
  XOR \ADD_/FAINST[127].FA_/U5  ( .A(\ADD_/FAINST[127].FA_/n3 ), .B(
        \ADD_/c[127] ), .Z(\ADD_/c[128] ) );
  XOR \ADD_/FAINST[127].FA_/U4  ( .A(\ADD_/FAINST[127].FA_/n1 ), .B(b[127]), 
        .Z(c[127]) );
  AND \ADD_/FAINST[127].FA_/U3  ( .A(\ADD_/FAINST[127].FA_/n1 ), .B(
        \ADD_/FAINST[127].FA_/n2 ), .Z(\ADD_/FAINST[127].FA_/n3 ) );
  XOR \ADD_/FAINST[127].FA_/U2  ( .A(b[127]), .B(\ADD_/c[127] ), .Z(
        \ADD_/FAINST[127].FA_/n2 ) );
  XOR \ADD_/FAINST[127].FA_/U1  ( .A(a[127]), .B(\ADD_/c[127] ), .Z(
        \ADD_/FAINST[127].FA_/n1 ) );
  XOR \ADD_/FAINST[126].FA_/U5  ( .A(\ADD_/FAINST[126].FA_/n3 ), .B(
        \ADD_/c[126] ), .Z(\ADD_/c[127] ) );
  XOR \ADD_/FAINST[126].FA_/U4  ( .A(\ADD_/FAINST[126].FA_/n1 ), .B(b[126]), 
        .Z(c[126]) );
  AND \ADD_/FAINST[126].FA_/U3  ( .A(\ADD_/FAINST[126].FA_/n1 ), .B(
        \ADD_/FAINST[126].FA_/n2 ), .Z(\ADD_/FAINST[126].FA_/n3 ) );
  XOR \ADD_/FAINST[126].FA_/U2  ( .A(b[126]), .B(\ADD_/c[126] ), .Z(
        \ADD_/FAINST[126].FA_/n2 ) );
  XOR \ADD_/FAINST[126].FA_/U1  ( .A(a[126]), .B(\ADD_/c[126] ), .Z(
        \ADD_/FAINST[126].FA_/n1 ) );
  XOR \ADD_/FAINST[125].FA_/U5  ( .A(\ADD_/FAINST[125].FA_/n3 ), .B(
        \ADD_/c[125] ), .Z(\ADD_/c[126] ) );
  XOR \ADD_/FAINST[125].FA_/U4  ( .A(\ADD_/FAINST[125].FA_/n1 ), .B(b[125]), 
        .Z(c[125]) );
  AND \ADD_/FAINST[125].FA_/U3  ( .A(\ADD_/FAINST[125].FA_/n1 ), .B(
        \ADD_/FAINST[125].FA_/n2 ), .Z(\ADD_/FAINST[125].FA_/n3 ) );
  XOR \ADD_/FAINST[125].FA_/U2  ( .A(b[125]), .B(\ADD_/c[125] ), .Z(
        \ADD_/FAINST[125].FA_/n2 ) );
  XOR \ADD_/FAINST[125].FA_/U1  ( .A(a[125]), .B(\ADD_/c[125] ), .Z(
        \ADD_/FAINST[125].FA_/n1 ) );
  XOR \ADD_/FAINST[124].FA_/U5  ( .A(\ADD_/FAINST[124].FA_/n3 ), .B(
        \ADD_/c[124] ), .Z(\ADD_/c[125] ) );
  XOR \ADD_/FAINST[124].FA_/U4  ( .A(\ADD_/FAINST[124].FA_/n1 ), .B(b[124]), 
        .Z(c[124]) );
  AND \ADD_/FAINST[124].FA_/U3  ( .A(\ADD_/FAINST[124].FA_/n1 ), .B(
        \ADD_/FAINST[124].FA_/n2 ), .Z(\ADD_/FAINST[124].FA_/n3 ) );
  XOR \ADD_/FAINST[124].FA_/U2  ( .A(b[124]), .B(\ADD_/c[124] ), .Z(
        \ADD_/FAINST[124].FA_/n2 ) );
  XOR \ADD_/FAINST[124].FA_/U1  ( .A(a[124]), .B(\ADD_/c[124] ), .Z(
        \ADD_/FAINST[124].FA_/n1 ) );
  XOR \ADD_/FAINST[123].FA_/U5  ( .A(\ADD_/FAINST[123].FA_/n3 ), .B(
        \ADD_/c[123] ), .Z(\ADD_/c[124] ) );
  XOR \ADD_/FAINST[123].FA_/U4  ( .A(\ADD_/FAINST[123].FA_/n1 ), .B(b[123]), 
        .Z(c[123]) );
  AND \ADD_/FAINST[123].FA_/U3  ( .A(\ADD_/FAINST[123].FA_/n1 ), .B(
        \ADD_/FAINST[123].FA_/n2 ), .Z(\ADD_/FAINST[123].FA_/n3 ) );
  XOR \ADD_/FAINST[123].FA_/U2  ( .A(b[123]), .B(\ADD_/c[123] ), .Z(
        \ADD_/FAINST[123].FA_/n2 ) );
  XOR \ADD_/FAINST[123].FA_/U1  ( .A(a[123]), .B(\ADD_/c[123] ), .Z(
        \ADD_/FAINST[123].FA_/n1 ) );
  XOR \ADD_/FAINST[122].FA_/U5  ( .A(\ADD_/FAINST[122].FA_/n3 ), .B(
        \ADD_/c[122] ), .Z(\ADD_/c[123] ) );
  XOR \ADD_/FAINST[122].FA_/U4  ( .A(\ADD_/FAINST[122].FA_/n1 ), .B(b[122]), 
        .Z(c[122]) );
  AND \ADD_/FAINST[122].FA_/U3  ( .A(\ADD_/FAINST[122].FA_/n1 ), .B(
        \ADD_/FAINST[122].FA_/n2 ), .Z(\ADD_/FAINST[122].FA_/n3 ) );
  XOR \ADD_/FAINST[122].FA_/U2  ( .A(b[122]), .B(\ADD_/c[122] ), .Z(
        \ADD_/FAINST[122].FA_/n2 ) );
  XOR \ADD_/FAINST[122].FA_/U1  ( .A(a[122]), .B(\ADD_/c[122] ), .Z(
        \ADD_/FAINST[122].FA_/n1 ) );
  XOR \ADD_/FAINST[121].FA_/U5  ( .A(\ADD_/FAINST[121].FA_/n3 ), .B(
        \ADD_/c[121] ), .Z(\ADD_/c[122] ) );
  XOR \ADD_/FAINST[121].FA_/U4  ( .A(\ADD_/FAINST[121].FA_/n1 ), .B(b[121]), 
        .Z(c[121]) );
  AND \ADD_/FAINST[121].FA_/U3  ( .A(\ADD_/FAINST[121].FA_/n1 ), .B(
        \ADD_/FAINST[121].FA_/n2 ), .Z(\ADD_/FAINST[121].FA_/n3 ) );
  XOR \ADD_/FAINST[121].FA_/U2  ( .A(b[121]), .B(\ADD_/c[121] ), .Z(
        \ADD_/FAINST[121].FA_/n2 ) );
  XOR \ADD_/FAINST[121].FA_/U1  ( .A(a[121]), .B(\ADD_/c[121] ), .Z(
        \ADD_/FAINST[121].FA_/n1 ) );
  XOR \ADD_/FAINST[120].FA_/U5  ( .A(\ADD_/FAINST[120].FA_/n3 ), .B(
        \ADD_/c[120] ), .Z(\ADD_/c[121] ) );
  XOR \ADD_/FAINST[120].FA_/U4  ( .A(\ADD_/FAINST[120].FA_/n1 ), .B(b[120]), 
        .Z(c[120]) );
  AND \ADD_/FAINST[120].FA_/U3  ( .A(\ADD_/FAINST[120].FA_/n1 ), .B(
        \ADD_/FAINST[120].FA_/n2 ), .Z(\ADD_/FAINST[120].FA_/n3 ) );
  XOR \ADD_/FAINST[120].FA_/U2  ( .A(b[120]), .B(\ADD_/c[120] ), .Z(
        \ADD_/FAINST[120].FA_/n2 ) );
  XOR \ADD_/FAINST[120].FA_/U1  ( .A(a[120]), .B(\ADD_/c[120] ), .Z(
        \ADD_/FAINST[120].FA_/n1 ) );
  XOR \ADD_/FAINST[119].FA_/U5  ( .A(\ADD_/FAINST[119].FA_/n3 ), .B(
        \ADD_/c[119] ), .Z(\ADD_/c[120] ) );
  XOR \ADD_/FAINST[119].FA_/U4  ( .A(\ADD_/FAINST[119].FA_/n1 ), .B(b[119]), 
        .Z(c[119]) );
  AND \ADD_/FAINST[119].FA_/U3  ( .A(\ADD_/FAINST[119].FA_/n1 ), .B(
        \ADD_/FAINST[119].FA_/n2 ), .Z(\ADD_/FAINST[119].FA_/n3 ) );
  XOR \ADD_/FAINST[119].FA_/U2  ( .A(b[119]), .B(\ADD_/c[119] ), .Z(
        \ADD_/FAINST[119].FA_/n2 ) );
  XOR \ADD_/FAINST[119].FA_/U1  ( .A(a[119]), .B(\ADD_/c[119] ), .Z(
        \ADD_/FAINST[119].FA_/n1 ) );
  XOR \ADD_/FAINST[118].FA_/U5  ( .A(\ADD_/FAINST[118].FA_/n3 ), .B(
        \ADD_/c[118] ), .Z(\ADD_/c[119] ) );
  XOR \ADD_/FAINST[118].FA_/U4  ( .A(\ADD_/FAINST[118].FA_/n1 ), .B(b[118]), 
        .Z(c[118]) );
  AND \ADD_/FAINST[118].FA_/U3  ( .A(\ADD_/FAINST[118].FA_/n1 ), .B(
        \ADD_/FAINST[118].FA_/n2 ), .Z(\ADD_/FAINST[118].FA_/n3 ) );
  XOR \ADD_/FAINST[118].FA_/U2  ( .A(b[118]), .B(\ADD_/c[118] ), .Z(
        \ADD_/FAINST[118].FA_/n2 ) );
  XOR \ADD_/FAINST[118].FA_/U1  ( .A(a[118]), .B(\ADD_/c[118] ), .Z(
        \ADD_/FAINST[118].FA_/n1 ) );
  XOR \ADD_/FAINST[117].FA_/U5  ( .A(\ADD_/FAINST[117].FA_/n3 ), .B(
        \ADD_/c[117] ), .Z(\ADD_/c[118] ) );
  XOR \ADD_/FAINST[117].FA_/U4  ( .A(\ADD_/FAINST[117].FA_/n1 ), .B(b[117]), 
        .Z(c[117]) );
  AND \ADD_/FAINST[117].FA_/U3  ( .A(\ADD_/FAINST[117].FA_/n1 ), .B(
        \ADD_/FAINST[117].FA_/n2 ), .Z(\ADD_/FAINST[117].FA_/n3 ) );
  XOR \ADD_/FAINST[117].FA_/U2  ( .A(b[117]), .B(\ADD_/c[117] ), .Z(
        \ADD_/FAINST[117].FA_/n2 ) );
  XOR \ADD_/FAINST[117].FA_/U1  ( .A(a[117]), .B(\ADD_/c[117] ), .Z(
        \ADD_/FAINST[117].FA_/n1 ) );
  XOR \ADD_/FAINST[116].FA_/U5  ( .A(\ADD_/FAINST[116].FA_/n3 ), .B(
        \ADD_/c[116] ), .Z(\ADD_/c[117] ) );
  XOR \ADD_/FAINST[116].FA_/U4  ( .A(\ADD_/FAINST[116].FA_/n1 ), .B(b[116]), 
        .Z(c[116]) );
  AND \ADD_/FAINST[116].FA_/U3  ( .A(\ADD_/FAINST[116].FA_/n1 ), .B(
        \ADD_/FAINST[116].FA_/n2 ), .Z(\ADD_/FAINST[116].FA_/n3 ) );
  XOR \ADD_/FAINST[116].FA_/U2  ( .A(b[116]), .B(\ADD_/c[116] ), .Z(
        \ADD_/FAINST[116].FA_/n2 ) );
  XOR \ADD_/FAINST[116].FA_/U1  ( .A(a[116]), .B(\ADD_/c[116] ), .Z(
        \ADD_/FAINST[116].FA_/n1 ) );
  XOR \ADD_/FAINST[115].FA_/U5  ( .A(\ADD_/FAINST[115].FA_/n3 ), .B(
        \ADD_/c[115] ), .Z(\ADD_/c[116] ) );
  XOR \ADD_/FAINST[115].FA_/U4  ( .A(\ADD_/FAINST[115].FA_/n1 ), .B(b[115]), 
        .Z(c[115]) );
  AND \ADD_/FAINST[115].FA_/U3  ( .A(\ADD_/FAINST[115].FA_/n1 ), .B(
        \ADD_/FAINST[115].FA_/n2 ), .Z(\ADD_/FAINST[115].FA_/n3 ) );
  XOR \ADD_/FAINST[115].FA_/U2  ( .A(b[115]), .B(\ADD_/c[115] ), .Z(
        \ADD_/FAINST[115].FA_/n2 ) );
  XOR \ADD_/FAINST[115].FA_/U1  ( .A(a[115]), .B(\ADD_/c[115] ), .Z(
        \ADD_/FAINST[115].FA_/n1 ) );
  XOR \ADD_/FAINST[114].FA_/U5  ( .A(\ADD_/FAINST[114].FA_/n3 ), .B(
        \ADD_/c[114] ), .Z(\ADD_/c[115] ) );
  XOR \ADD_/FAINST[114].FA_/U4  ( .A(\ADD_/FAINST[114].FA_/n1 ), .B(b[114]), 
        .Z(c[114]) );
  AND \ADD_/FAINST[114].FA_/U3  ( .A(\ADD_/FAINST[114].FA_/n1 ), .B(
        \ADD_/FAINST[114].FA_/n2 ), .Z(\ADD_/FAINST[114].FA_/n3 ) );
  XOR \ADD_/FAINST[114].FA_/U2  ( .A(b[114]), .B(\ADD_/c[114] ), .Z(
        \ADD_/FAINST[114].FA_/n2 ) );
  XOR \ADD_/FAINST[114].FA_/U1  ( .A(a[114]), .B(\ADD_/c[114] ), .Z(
        \ADD_/FAINST[114].FA_/n1 ) );
  XOR \ADD_/FAINST[113].FA_/U5  ( .A(\ADD_/FAINST[113].FA_/n3 ), .B(
        \ADD_/c[113] ), .Z(\ADD_/c[114] ) );
  XOR \ADD_/FAINST[113].FA_/U4  ( .A(\ADD_/FAINST[113].FA_/n1 ), .B(b[113]), 
        .Z(c[113]) );
  AND \ADD_/FAINST[113].FA_/U3  ( .A(\ADD_/FAINST[113].FA_/n1 ), .B(
        \ADD_/FAINST[113].FA_/n2 ), .Z(\ADD_/FAINST[113].FA_/n3 ) );
  XOR \ADD_/FAINST[113].FA_/U2  ( .A(b[113]), .B(\ADD_/c[113] ), .Z(
        \ADD_/FAINST[113].FA_/n2 ) );
  XOR \ADD_/FAINST[113].FA_/U1  ( .A(a[113]), .B(\ADD_/c[113] ), .Z(
        \ADD_/FAINST[113].FA_/n1 ) );
  XOR \ADD_/FAINST[112].FA_/U5  ( .A(\ADD_/FAINST[112].FA_/n3 ), .B(
        \ADD_/c[112] ), .Z(\ADD_/c[113] ) );
  XOR \ADD_/FAINST[112].FA_/U4  ( .A(\ADD_/FAINST[112].FA_/n1 ), .B(b[112]), 
        .Z(c[112]) );
  AND \ADD_/FAINST[112].FA_/U3  ( .A(\ADD_/FAINST[112].FA_/n1 ), .B(
        \ADD_/FAINST[112].FA_/n2 ), .Z(\ADD_/FAINST[112].FA_/n3 ) );
  XOR \ADD_/FAINST[112].FA_/U2  ( .A(b[112]), .B(\ADD_/c[112] ), .Z(
        \ADD_/FAINST[112].FA_/n2 ) );
  XOR \ADD_/FAINST[112].FA_/U1  ( .A(a[112]), .B(\ADD_/c[112] ), .Z(
        \ADD_/FAINST[112].FA_/n1 ) );
  XOR \ADD_/FAINST[111].FA_/U5  ( .A(\ADD_/FAINST[111].FA_/n3 ), .B(
        \ADD_/c[111] ), .Z(\ADD_/c[112] ) );
  XOR \ADD_/FAINST[111].FA_/U4  ( .A(\ADD_/FAINST[111].FA_/n1 ), .B(b[111]), 
        .Z(c[111]) );
  AND \ADD_/FAINST[111].FA_/U3  ( .A(\ADD_/FAINST[111].FA_/n1 ), .B(
        \ADD_/FAINST[111].FA_/n2 ), .Z(\ADD_/FAINST[111].FA_/n3 ) );
  XOR \ADD_/FAINST[111].FA_/U2  ( .A(b[111]), .B(\ADD_/c[111] ), .Z(
        \ADD_/FAINST[111].FA_/n2 ) );
  XOR \ADD_/FAINST[111].FA_/U1  ( .A(a[111]), .B(\ADD_/c[111] ), .Z(
        \ADD_/FAINST[111].FA_/n1 ) );
  XOR \ADD_/FAINST[110].FA_/U5  ( .A(\ADD_/FAINST[110].FA_/n3 ), .B(
        \ADD_/c[110] ), .Z(\ADD_/c[111] ) );
  XOR \ADD_/FAINST[110].FA_/U4  ( .A(\ADD_/FAINST[110].FA_/n1 ), .B(b[110]), 
        .Z(c[110]) );
  AND \ADD_/FAINST[110].FA_/U3  ( .A(\ADD_/FAINST[110].FA_/n1 ), .B(
        \ADD_/FAINST[110].FA_/n2 ), .Z(\ADD_/FAINST[110].FA_/n3 ) );
  XOR \ADD_/FAINST[110].FA_/U2  ( .A(b[110]), .B(\ADD_/c[110] ), .Z(
        \ADD_/FAINST[110].FA_/n2 ) );
  XOR \ADD_/FAINST[110].FA_/U1  ( .A(a[110]), .B(\ADD_/c[110] ), .Z(
        \ADD_/FAINST[110].FA_/n1 ) );
  XOR \ADD_/FAINST[109].FA_/U5  ( .A(\ADD_/FAINST[109].FA_/n3 ), .B(
        \ADD_/c[109] ), .Z(\ADD_/c[110] ) );
  XOR \ADD_/FAINST[109].FA_/U4  ( .A(\ADD_/FAINST[109].FA_/n1 ), .B(b[109]), 
        .Z(c[109]) );
  AND \ADD_/FAINST[109].FA_/U3  ( .A(\ADD_/FAINST[109].FA_/n1 ), .B(
        \ADD_/FAINST[109].FA_/n2 ), .Z(\ADD_/FAINST[109].FA_/n3 ) );
  XOR \ADD_/FAINST[109].FA_/U2  ( .A(b[109]), .B(\ADD_/c[109] ), .Z(
        \ADD_/FAINST[109].FA_/n2 ) );
  XOR \ADD_/FAINST[109].FA_/U1  ( .A(a[109]), .B(\ADD_/c[109] ), .Z(
        \ADD_/FAINST[109].FA_/n1 ) );
  XOR \ADD_/FAINST[108].FA_/U5  ( .A(\ADD_/FAINST[108].FA_/n3 ), .B(
        \ADD_/c[108] ), .Z(\ADD_/c[109] ) );
  XOR \ADD_/FAINST[108].FA_/U4  ( .A(\ADD_/FAINST[108].FA_/n1 ), .B(b[108]), 
        .Z(c[108]) );
  AND \ADD_/FAINST[108].FA_/U3  ( .A(\ADD_/FAINST[108].FA_/n1 ), .B(
        \ADD_/FAINST[108].FA_/n2 ), .Z(\ADD_/FAINST[108].FA_/n3 ) );
  XOR \ADD_/FAINST[108].FA_/U2  ( .A(b[108]), .B(\ADD_/c[108] ), .Z(
        \ADD_/FAINST[108].FA_/n2 ) );
  XOR \ADD_/FAINST[108].FA_/U1  ( .A(a[108]), .B(\ADD_/c[108] ), .Z(
        \ADD_/FAINST[108].FA_/n1 ) );
  XOR \ADD_/FAINST[107].FA_/U5  ( .A(\ADD_/FAINST[107].FA_/n3 ), .B(
        \ADD_/c[107] ), .Z(\ADD_/c[108] ) );
  XOR \ADD_/FAINST[107].FA_/U4  ( .A(\ADD_/FAINST[107].FA_/n1 ), .B(b[107]), 
        .Z(c[107]) );
  AND \ADD_/FAINST[107].FA_/U3  ( .A(\ADD_/FAINST[107].FA_/n1 ), .B(
        \ADD_/FAINST[107].FA_/n2 ), .Z(\ADD_/FAINST[107].FA_/n3 ) );
  XOR \ADD_/FAINST[107].FA_/U2  ( .A(b[107]), .B(\ADD_/c[107] ), .Z(
        \ADD_/FAINST[107].FA_/n2 ) );
  XOR \ADD_/FAINST[107].FA_/U1  ( .A(a[107]), .B(\ADD_/c[107] ), .Z(
        \ADD_/FAINST[107].FA_/n1 ) );
  XOR \ADD_/FAINST[106].FA_/U5  ( .A(\ADD_/FAINST[106].FA_/n3 ), .B(
        \ADD_/c[106] ), .Z(\ADD_/c[107] ) );
  XOR \ADD_/FAINST[106].FA_/U4  ( .A(\ADD_/FAINST[106].FA_/n1 ), .B(b[106]), 
        .Z(c[106]) );
  AND \ADD_/FAINST[106].FA_/U3  ( .A(\ADD_/FAINST[106].FA_/n1 ), .B(
        \ADD_/FAINST[106].FA_/n2 ), .Z(\ADD_/FAINST[106].FA_/n3 ) );
  XOR \ADD_/FAINST[106].FA_/U2  ( .A(b[106]), .B(\ADD_/c[106] ), .Z(
        \ADD_/FAINST[106].FA_/n2 ) );
  XOR \ADD_/FAINST[106].FA_/U1  ( .A(a[106]), .B(\ADD_/c[106] ), .Z(
        \ADD_/FAINST[106].FA_/n1 ) );
  XOR \ADD_/FAINST[105].FA_/U5  ( .A(\ADD_/FAINST[105].FA_/n3 ), .B(
        \ADD_/c[105] ), .Z(\ADD_/c[106] ) );
  XOR \ADD_/FAINST[105].FA_/U4  ( .A(\ADD_/FAINST[105].FA_/n1 ), .B(b[105]), 
        .Z(c[105]) );
  AND \ADD_/FAINST[105].FA_/U3  ( .A(\ADD_/FAINST[105].FA_/n1 ), .B(
        \ADD_/FAINST[105].FA_/n2 ), .Z(\ADD_/FAINST[105].FA_/n3 ) );
  XOR \ADD_/FAINST[105].FA_/U2  ( .A(b[105]), .B(\ADD_/c[105] ), .Z(
        \ADD_/FAINST[105].FA_/n2 ) );
  XOR \ADD_/FAINST[105].FA_/U1  ( .A(a[105]), .B(\ADD_/c[105] ), .Z(
        \ADD_/FAINST[105].FA_/n1 ) );
  XOR \ADD_/FAINST[104].FA_/U5  ( .A(\ADD_/FAINST[104].FA_/n3 ), .B(
        \ADD_/c[104] ), .Z(\ADD_/c[105] ) );
  XOR \ADD_/FAINST[104].FA_/U4  ( .A(\ADD_/FAINST[104].FA_/n1 ), .B(b[104]), 
        .Z(c[104]) );
  AND \ADD_/FAINST[104].FA_/U3  ( .A(\ADD_/FAINST[104].FA_/n1 ), .B(
        \ADD_/FAINST[104].FA_/n2 ), .Z(\ADD_/FAINST[104].FA_/n3 ) );
  XOR \ADD_/FAINST[104].FA_/U2  ( .A(b[104]), .B(\ADD_/c[104] ), .Z(
        \ADD_/FAINST[104].FA_/n2 ) );
  XOR \ADD_/FAINST[104].FA_/U1  ( .A(a[104]), .B(\ADD_/c[104] ), .Z(
        \ADD_/FAINST[104].FA_/n1 ) );
  XOR \ADD_/FAINST[103].FA_/U5  ( .A(\ADD_/FAINST[103].FA_/n3 ), .B(
        \ADD_/c[103] ), .Z(\ADD_/c[104] ) );
  XOR \ADD_/FAINST[103].FA_/U4  ( .A(\ADD_/FAINST[103].FA_/n1 ), .B(b[103]), 
        .Z(c[103]) );
  AND \ADD_/FAINST[103].FA_/U3  ( .A(\ADD_/FAINST[103].FA_/n1 ), .B(
        \ADD_/FAINST[103].FA_/n2 ), .Z(\ADD_/FAINST[103].FA_/n3 ) );
  XOR \ADD_/FAINST[103].FA_/U2  ( .A(b[103]), .B(\ADD_/c[103] ), .Z(
        \ADD_/FAINST[103].FA_/n2 ) );
  XOR \ADD_/FAINST[103].FA_/U1  ( .A(a[103]), .B(\ADD_/c[103] ), .Z(
        \ADD_/FAINST[103].FA_/n1 ) );
  XOR \ADD_/FAINST[102].FA_/U5  ( .A(\ADD_/FAINST[102].FA_/n3 ), .B(
        \ADD_/c[102] ), .Z(\ADD_/c[103] ) );
  XOR \ADD_/FAINST[102].FA_/U4  ( .A(\ADD_/FAINST[102].FA_/n1 ), .B(b[102]), 
        .Z(c[102]) );
  AND \ADD_/FAINST[102].FA_/U3  ( .A(\ADD_/FAINST[102].FA_/n1 ), .B(
        \ADD_/FAINST[102].FA_/n2 ), .Z(\ADD_/FAINST[102].FA_/n3 ) );
  XOR \ADD_/FAINST[102].FA_/U2  ( .A(b[102]), .B(\ADD_/c[102] ), .Z(
        \ADD_/FAINST[102].FA_/n2 ) );
  XOR \ADD_/FAINST[102].FA_/U1  ( .A(a[102]), .B(\ADD_/c[102] ), .Z(
        \ADD_/FAINST[102].FA_/n1 ) );
  XOR \ADD_/FAINST[101].FA_/U5  ( .A(\ADD_/FAINST[101].FA_/n3 ), .B(
        \ADD_/c[101] ), .Z(\ADD_/c[102] ) );
  XOR \ADD_/FAINST[101].FA_/U4  ( .A(\ADD_/FAINST[101].FA_/n1 ), .B(b[101]), 
        .Z(c[101]) );
  AND \ADD_/FAINST[101].FA_/U3  ( .A(\ADD_/FAINST[101].FA_/n1 ), .B(
        \ADD_/FAINST[101].FA_/n2 ), .Z(\ADD_/FAINST[101].FA_/n3 ) );
  XOR \ADD_/FAINST[101].FA_/U2  ( .A(b[101]), .B(\ADD_/c[101] ), .Z(
        \ADD_/FAINST[101].FA_/n2 ) );
  XOR \ADD_/FAINST[101].FA_/U1  ( .A(a[101]), .B(\ADD_/c[101] ), .Z(
        \ADD_/FAINST[101].FA_/n1 ) );
  XOR \ADD_/FAINST[100].FA_/U5  ( .A(\ADD_/FAINST[100].FA_/n3 ), .B(
        \ADD_/c[100] ), .Z(\ADD_/c[101] ) );
  XOR \ADD_/FAINST[100].FA_/U4  ( .A(\ADD_/FAINST[100].FA_/n1 ), .B(b[100]), 
        .Z(c[100]) );
  AND \ADD_/FAINST[100].FA_/U3  ( .A(\ADD_/FAINST[100].FA_/n1 ), .B(
        \ADD_/FAINST[100].FA_/n2 ), .Z(\ADD_/FAINST[100].FA_/n3 ) );
  XOR \ADD_/FAINST[100].FA_/U2  ( .A(b[100]), .B(\ADD_/c[100] ), .Z(
        \ADD_/FAINST[100].FA_/n2 ) );
  XOR \ADD_/FAINST[100].FA_/U1  ( .A(a[100]), .B(\ADD_/c[100] ), .Z(
        \ADD_/FAINST[100].FA_/n1 ) );
  XOR \ADD_/FAINST[99].FA_/U5  ( .A(\ADD_/FAINST[99].FA_/n3 ), .B(\ADD_/c[99] ), .Z(\ADD_/c[100] ) );
  XOR \ADD_/FAINST[99].FA_/U4  ( .A(\ADD_/FAINST[99].FA_/n1 ), .B(b[99]), .Z(
        c[99]) );
  AND \ADD_/FAINST[99].FA_/U3  ( .A(\ADD_/FAINST[99].FA_/n1 ), .B(
        \ADD_/FAINST[99].FA_/n2 ), .Z(\ADD_/FAINST[99].FA_/n3 ) );
  XOR \ADD_/FAINST[99].FA_/U2  ( .A(b[99]), .B(\ADD_/c[99] ), .Z(
        \ADD_/FAINST[99].FA_/n2 ) );
  XOR \ADD_/FAINST[99].FA_/U1  ( .A(a[99]), .B(\ADD_/c[99] ), .Z(
        \ADD_/FAINST[99].FA_/n1 ) );
  XOR \ADD_/FAINST[98].FA_/U5  ( .A(\ADD_/FAINST[98].FA_/n3 ), .B(\ADD_/c[98] ), .Z(\ADD_/c[99] ) );
  XOR \ADD_/FAINST[98].FA_/U4  ( .A(\ADD_/FAINST[98].FA_/n1 ), .B(b[98]), .Z(
        c[98]) );
  AND \ADD_/FAINST[98].FA_/U3  ( .A(\ADD_/FAINST[98].FA_/n1 ), .B(
        \ADD_/FAINST[98].FA_/n2 ), .Z(\ADD_/FAINST[98].FA_/n3 ) );
  XOR \ADD_/FAINST[98].FA_/U2  ( .A(b[98]), .B(\ADD_/c[98] ), .Z(
        \ADD_/FAINST[98].FA_/n2 ) );
  XOR \ADD_/FAINST[98].FA_/U1  ( .A(a[98]), .B(\ADD_/c[98] ), .Z(
        \ADD_/FAINST[98].FA_/n1 ) );
  XOR \ADD_/FAINST[97].FA_/U5  ( .A(\ADD_/FAINST[97].FA_/n3 ), .B(\ADD_/c[97] ), .Z(\ADD_/c[98] ) );
  XOR \ADD_/FAINST[97].FA_/U4  ( .A(\ADD_/FAINST[97].FA_/n1 ), .B(b[97]), .Z(
        c[97]) );
  AND \ADD_/FAINST[97].FA_/U3  ( .A(\ADD_/FAINST[97].FA_/n1 ), .B(
        \ADD_/FAINST[97].FA_/n2 ), .Z(\ADD_/FAINST[97].FA_/n3 ) );
  XOR \ADD_/FAINST[97].FA_/U2  ( .A(b[97]), .B(\ADD_/c[97] ), .Z(
        \ADD_/FAINST[97].FA_/n2 ) );
  XOR \ADD_/FAINST[97].FA_/U1  ( .A(a[97]), .B(\ADD_/c[97] ), .Z(
        \ADD_/FAINST[97].FA_/n1 ) );
  XOR \ADD_/FAINST[96].FA_/U5  ( .A(\ADD_/FAINST[96].FA_/n3 ), .B(\ADD_/c[96] ), .Z(\ADD_/c[97] ) );
  XOR \ADD_/FAINST[96].FA_/U4  ( .A(\ADD_/FAINST[96].FA_/n1 ), .B(b[96]), .Z(
        c[96]) );
  AND \ADD_/FAINST[96].FA_/U3  ( .A(\ADD_/FAINST[96].FA_/n1 ), .B(
        \ADD_/FAINST[96].FA_/n2 ), .Z(\ADD_/FAINST[96].FA_/n3 ) );
  XOR \ADD_/FAINST[96].FA_/U2  ( .A(b[96]), .B(\ADD_/c[96] ), .Z(
        \ADD_/FAINST[96].FA_/n2 ) );
  XOR \ADD_/FAINST[96].FA_/U1  ( .A(a[96]), .B(\ADD_/c[96] ), .Z(
        \ADD_/FAINST[96].FA_/n1 ) );
  XOR \ADD_/FAINST[95].FA_/U5  ( .A(\ADD_/FAINST[95].FA_/n3 ), .B(\ADD_/c[95] ), .Z(\ADD_/c[96] ) );
  XOR \ADD_/FAINST[95].FA_/U4  ( .A(\ADD_/FAINST[95].FA_/n1 ), .B(b[95]), .Z(
        c[95]) );
  AND \ADD_/FAINST[95].FA_/U3  ( .A(\ADD_/FAINST[95].FA_/n1 ), .B(
        \ADD_/FAINST[95].FA_/n2 ), .Z(\ADD_/FAINST[95].FA_/n3 ) );
  XOR \ADD_/FAINST[95].FA_/U2  ( .A(b[95]), .B(\ADD_/c[95] ), .Z(
        \ADD_/FAINST[95].FA_/n2 ) );
  XOR \ADD_/FAINST[95].FA_/U1  ( .A(a[95]), .B(\ADD_/c[95] ), .Z(
        \ADD_/FAINST[95].FA_/n1 ) );
  XOR \ADD_/FAINST[94].FA_/U5  ( .A(\ADD_/FAINST[94].FA_/n3 ), .B(\ADD_/c[94] ), .Z(\ADD_/c[95] ) );
  XOR \ADD_/FAINST[94].FA_/U4  ( .A(\ADD_/FAINST[94].FA_/n1 ), .B(b[94]), .Z(
        c[94]) );
  AND \ADD_/FAINST[94].FA_/U3  ( .A(\ADD_/FAINST[94].FA_/n1 ), .B(
        \ADD_/FAINST[94].FA_/n2 ), .Z(\ADD_/FAINST[94].FA_/n3 ) );
  XOR \ADD_/FAINST[94].FA_/U2  ( .A(b[94]), .B(\ADD_/c[94] ), .Z(
        \ADD_/FAINST[94].FA_/n2 ) );
  XOR \ADD_/FAINST[94].FA_/U1  ( .A(a[94]), .B(\ADD_/c[94] ), .Z(
        \ADD_/FAINST[94].FA_/n1 ) );
  XOR \ADD_/FAINST[93].FA_/U5  ( .A(\ADD_/FAINST[93].FA_/n3 ), .B(\ADD_/c[93] ), .Z(\ADD_/c[94] ) );
  XOR \ADD_/FAINST[93].FA_/U4  ( .A(\ADD_/FAINST[93].FA_/n1 ), .B(b[93]), .Z(
        c[93]) );
  AND \ADD_/FAINST[93].FA_/U3  ( .A(\ADD_/FAINST[93].FA_/n1 ), .B(
        \ADD_/FAINST[93].FA_/n2 ), .Z(\ADD_/FAINST[93].FA_/n3 ) );
  XOR \ADD_/FAINST[93].FA_/U2  ( .A(b[93]), .B(\ADD_/c[93] ), .Z(
        \ADD_/FAINST[93].FA_/n2 ) );
  XOR \ADD_/FAINST[93].FA_/U1  ( .A(a[93]), .B(\ADD_/c[93] ), .Z(
        \ADD_/FAINST[93].FA_/n1 ) );
  XOR \ADD_/FAINST[92].FA_/U5  ( .A(\ADD_/FAINST[92].FA_/n3 ), .B(\ADD_/c[92] ), .Z(\ADD_/c[93] ) );
  XOR \ADD_/FAINST[92].FA_/U4  ( .A(\ADD_/FAINST[92].FA_/n1 ), .B(b[92]), .Z(
        c[92]) );
  AND \ADD_/FAINST[92].FA_/U3  ( .A(\ADD_/FAINST[92].FA_/n1 ), .B(
        \ADD_/FAINST[92].FA_/n2 ), .Z(\ADD_/FAINST[92].FA_/n3 ) );
  XOR \ADD_/FAINST[92].FA_/U2  ( .A(b[92]), .B(\ADD_/c[92] ), .Z(
        \ADD_/FAINST[92].FA_/n2 ) );
  XOR \ADD_/FAINST[92].FA_/U1  ( .A(a[92]), .B(\ADD_/c[92] ), .Z(
        \ADD_/FAINST[92].FA_/n1 ) );
  XOR \ADD_/FAINST[91].FA_/U5  ( .A(\ADD_/FAINST[91].FA_/n3 ), .B(\ADD_/c[91] ), .Z(\ADD_/c[92] ) );
  XOR \ADD_/FAINST[91].FA_/U4  ( .A(\ADD_/FAINST[91].FA_/n1 ), .B(b[91]), .Z(
        c[91]) );
  AND \ADD_/FAINST[91].FA_/U3  ( .A(\ADD_/FAINST[91].FA_/n1 ), .B(
        \ADD_/FAINST[91].FA_/n2 ), .Z(\ADD_/FAINST[91].FA_/n3 ) );
  XOR \ADD_/FAINST[91].FA_/U2  ( .A(b[91]), .B(\ADD_/c[91] ), .Z(
        \ADD_/FAINST[91].FA_/n2 ) );
  XOR \ADD_/FAINST[91].FA_/U1  ( .A(a[91]), .B(\ADD_/c[91] ), .Z(
        \ADD_/FAINST[91].FA_/n1 ) );
  XOR \ADD_/FAINST[90].FA_/U5  ( .A(\ADD_/FAINST[90].FA_/n3 ), .B(\ADD_/c[90] ), .Z(\ADD_/c[91] ) );
  XOR \ADD_/FAINST[90].FA_/U4  ( .A(\ADD_/FAINST[90].FA_/n1 ), .B(b[90]), .Z(
        c[90]) );
  AND \ADD_/FAINST[90].FA_/U3  ( .A(\ADD_/FAINST[90].FA_/n1 ), .B(
        \ADD_/FAINST[90].FA_/n2 ), .Z(\ADD_/FAINST[90].FA_/n3 ) );
  XOR \ADD_/FAINST[90].FA_/U2  ( .A(b[90]), .B(\ADD_/c[90] ), .Z(
        \ADD_/FAINST[90].FA_/n2 ) );
  XOR \ADD_/FAINST[90].FA_/U1  ( .A(a[90]), .B(\ADD_/c[90] ), .Z(
        \ADD_/FAINST[90].FA_/n1 ) );
  XOR \ADD_/FAINST[89].FA_/U5  ( .A(\ADD_/FAINST[89].FA_/n3 ), .B(\ADD_/c[89] ), .Z(\ADD_/c[90] ) );
  XOR \ADD_/FAINST[89].FA_/U4  ( .A(\ADD_/FAINST[89].FA_/n1 ), .B(b[89]), .Z(
        c[89]) );
  AND \ADD_/FAINST[89].FA_/U3  ( .A(\ADD_/FAINST[89].FA_/n1 ), .B(
        \ADD_/FAINST[89].FA_/n2 ), .Z(\ADD_/FAINST[89].FA_/n3 ) );
  XOR \ADD_/FAINST[89].FA_/U2  ( .A(b[89]), .B(\ADD_/c[89] ), .Z(
        \ADD_/FAINST[89].FA_/n2 ) );
  XOR \ADD_/FAINST[89].FA_/U1  ( .A(a[89]), .B(\ADD_/c[89] ), .Z(
        \ADD_/FAINST[89].FA_/n1 ) );
  XOR \ADD_/FAINST[88].FA_/U5  ( .A(\ADD_/FAINST[88].FA_/n3 ), .B(\ADD_/c[88] ), .Z(\ADD_/c[89] ) );
  XOR \ADD_/FAINST[88].FA_/U4  ( .A(\ADD_/FAINST[88].FA_/n1 ), .B(b[88]), .Z(
        c[88]) );
  AND \ADD_/FAINST[88].FA_/U3  ( .A(\ADD_/FAINST[88].FA_/n1 ), .B(
        \ADD_/FAINST[88].FA_/n2 ), .Z(\ADD_/FAINST[88].FA_/n3 ) );
  XOR \ADD_/FAINST[88].FA_/U2  ( .A(b[88]), .B(\ADD_/c[88] ), .Z(
        \ADD_/FAINST[88].FA_/n2 ) );
  XOR \ADD_/FAINST[88].FA_/U1  ( .A(a[88]), .B(\ADD_/c[88] ), .Z(
        \ADD_/FAINST[88].FA_/n1 ) );
  XOR \ADD_/FAINST[87].FA_/U5  ( .A(\ADD_/FAINST[87].FA_/n3 ), .B(\ADD_/c[87] ), .Z(\ADD_/c[88] ) );
  XOR \ADD_/FAINST[87].FA_/U4  ( .A(\ADD_/FAINST[87].FA_/n1 ), .B(b[87]), .Z(
        c[87]) );
  AND \ADD_/FAINST[87].FA_/U3  ( .A(\ADD_/FAINST[87].FA_/n1 ), .B(
        \ADD_/FAINST[87].FA_/n2 ), .Z(\ADD_/FAINST[87].FA_/n3 ) );
  XOR \ADD_/FAINST[87].FA_/U2  ( .A(b[87]), .B(\ADD_/c[87] ), .Z(
        \ADD_/FAINST[87].FA_/n2 ) );
  XOR \ADD_/FAINST[87].FA_/U1  ( .A(a[87]), .B(\ADD_/c[87] ), .Z(
        \ADD_/FAINST[87].FA_/n1 ) );
  XOR \ADD_/FAINST[86].FA_/U5  ( .A(\ADD_/FAINST[86].FA_/n3 ), .B(\ADD_/c[86] ), .Z(\ADD_/c[87] ) );
  XOR \ADD_/FAINST[86].FA_/U4  ( .A(\ADD_/FAINST[86].FA_/n1 ), .B(b[86]), .Z(
        c[86]) );
  AND \ADD_/FAINST[86].FA_/U3  ( .A(\ADD_/FAINST[86].FA_/n1 ), .B(
        \ADD_/FAINST[86].FA_/n2 ), .Z(\ADD_/FAINST[86].FA_/n3 ) );
  XOR \ADD_/FAINST[86].FA_/U2  ( .A(b[86]), .B(\ADD_/c[86] ), .Z(
        \ADD_/FAINST[86].FA_/n2 ) );
  XOR \ADD_/FAINST[86].FA_/U1  ( .A(a[86]), .B(\ADD_/c[86] ), .Z(
        \ADD_/FAINST[86].FA_/n1 ) );
  XOR \ADD_/FAINST[85].FA_/U5  ( .A(\ADD_/FAINST[85].FA_/n3 ), .B(\ADD_/c[85] ), .Z(\ADD_/c[86] ) );
  XOR \ADD_/FAINST[85].FA_/U4  ( .A(\ADD_/FAINST[85].FA_/n1 ), .B(b[85]), .Z(
        c[85]) );
  AND \ADD_/FAINST[85].FA_/U3  ( .A(\ADD_/FAINST[85].FA_/n1 ), .B(
        \ADD_/FAINST[85].FA_/n2 ), .Z(\ADD_/FAINST[85].FA_/n3 ) );
  XOR \ADD_/FAINST[85].FA_/U2  ( .A(b[85]), .B(\ADD_/c[85] ), .Z(
        \ADD_/FAINST[85].FA_/n2 ) );
  XOR \ADD_/FAINST[85].FA_/U1  ( .A(a[85]), .B(\ADD_/c[85] ), .Z(
        \ADD_/FAINST[85].FA_/n1 ) );
  XOR \ADD_/FAINST[84].FA_/U5  ( .A(\ADD_/FAINST[84].FA_/n3 ), .B(\ADD_/c[84] ), .Z(\ADD_/c[85] ) );
  XOR \ADD_/FAINST[84].FA_/U4  ( .A(\ADD_/FAINST[84].FA_/n1 ), .B(b[84]), .Z(
        c[84]) );
  AND \ADD_/FAINST[84].FA_/U3  ( .A(\ADD_/FAINST[84].FA_/n1 ), .B(
        \ADD_/FAINST[84].FA_/n2 ), .Z(\ADD_/FAINST[84].FA_/n3 ) );
  XOR \ADD_/FAINST[84].FA_/U2  ( .A(b[84]), .B(\ADD_/c[84] ), .Z(
        \ADD_/FAINST[84].FA_/n2 ) );
  XOR \ADD_/FAINST[84].FA_/U1  ( .A(a[84]), .B(\ADD_/c[84] ), .Z(
        \ADD_/FAINST[84].FA_/n1 ) );
  XOR \ADD_/FAINST[83].FA_/U5  ( .A(\ADD_/FAINST[83].FA_/n3 ), .B(\ADD_/c[83] ), .Z(\ADD_/c[84] ) );
  XOR \ADD_/FAINST[83].FA_/U4  ( .A(\ADD_/FAINST[83].FA_/n1 ), .B(b[83]), .Z(
        c[83]) );
  AND \ADD_/FAINST[83].FA_/U3  ( .A(\ADD_/FAINST[83].FA_/n1 ), .B(
        \ADD_/FAINST[83].FA_/n2 ), .Z(\ADD_/FAINST[83].FA_/n3 ) );
  XOR \ADD_/FAINST[83].FA_/U2  ( .A(b[83]), .B(\ADD_/c[83] ), .Z(
        \ADD_/FAINST[83].FA_/n2 ) );
  XOR \ADD_/FAINST[83].FA_/U1  ( .A(a[83]), .B(\ADD_/c[83] ), .Z(
        \ADD_/FAINST[83].FA_/n1 ) );
  XOR \ADD_/FAINST[82].FA_/U5  ( .A(\ADD_/FAINST[82].FA_/n3 ), .B(\ADD_/c[82] ), .Z(\ADD_/c[83] ) );
  XOR \ADD_/FAINST[82].FA_/U4  ( .A(\ADD_/FAINST[82].FA_/n1 ), .B(b[82]), .Z(
        c[82]) );
  AND \ADD_/FAINST[82].FA_/U3  ( .A(\ADD_/FAINST[82].FA_/n1 ), .B(
        \ADD_/FAINST[82].FA_/n2 ), .Z(\ADD_/FAINST[82].FA_/n3 ) );
  XOR \ADD_/FAINST[82].FA_/U2  ( .A(b[82]), .B(\ADD_/c[82] ), .Z(
        \ADD_/FAINST[82].FA_/n2 ) );
  XOR \ADD_/FAINST[82].FA_/U1  ( .A(a[82]), .B(\ADD_/c[82] ), .Z(
        \ADD_/FAINST[82].FA_/n1 ) );
  XOR \ADD_/FAINST[81].FA_/U5  ( .A(\ADD_/FAINST[81].FA_/n3 ), .B(\ADD_/c[81] ), .Z(\ADD_/c[82] ) );
  XOR \ADD_/FAINST[81].FA_/U4  ( .A(\ADD_/FAINST[81].FA_/n1 ), .B(b[81]), .Z(
        c[81]) );
  AND \ADD_/FAINST[81].FA_/U3  ( .A(\ADD_/FAINST[81].FA_/n1 ), .B(
        \ADD_/FAINST[81].FA_/n2 ), .Z(\ADD_/FAINST[81].FA_/n3 ) );
  XOR \ADD_/FAINST[81].FA_/U2  ( .A(b[81]), .B(\ADD_/c[81] ), .Z(
        \ADD_/FAINST[81].FA_/n2 ) );
  XOR \ADD_/FAINST[81].FA_/U1  ( .A(a[81]), .B(\ADD_/c[81] ), .Z(
        \ADD_/FAINST[81].FA_/n1 ) );
  XOR \ADD_/FAINST[80].FA_/U5  ( .A(\ADD_/FAINST[80].FA_/n3 ), .B(\ADD_/c[80] ), .Z(\ADD_/c[81] ) );
  XOR \ADD_/FAINST[80].FA_/U4  ( .A(\ADD_/FAINST[80].FA_/n1 ), .B(b[80]), .Z(
        c[80]) );
  AND \ADD_/FAINST[80].FA_/U3  ( .A(\ADD_/FAINST[80].FA_/n1 ), .B(
        \ADD_/FAINST[80].FA_/n2 ), .Z(\ADD_/FAINST[80].FA_/n3 ) );
  XOR \ADD_/FAINST[80].FA_/U2  ( .A(b[80]), .B(\ADD_/c[80] ), .Z(
        \ADD_/FAINST[80].FA_/n2 ) );
  XOR \ADD_/FAINST[80].FA_/U1  ( .A(a[80]), .B(\ADD_/c[80] ), .Z(
        \ADD_/FAINST[80].FA_/n1 ) );
  XOR \ADD_/FAINST[79].FA_/U5  ( .A(\ADD_/FAINST[79].FA_/n3 ), .B(\ADD_/c[79] ), .Z(\ADD_/c[80] ) );
  XOR \ADD_/FAINST[79].FA_/U4  ( .A(\ADD_/FAINST[79].FA_/n1 ), .B(b[79]), .Z(
        c[79]) );
  AND \ADD_/FAINST[79].FA_/U3  ( .A(\ADD_/FAINST[79].FA_/n1 ), .B(
        \ADD_/FAINST[79].FA_/n2 ), .Z(\ADD_/FAINST[79].FA_/n3 ) );
  XOR \ADD_/FAINST[79].FA_/U2  ( .A(b[79]), .B(\ADD_/c[79] ), .Z(
        \ADD_/FAINST[79].FA_/n2 ) );
  XOR \ADD_/FAINST[79].FA_/U1  ( .A(a[79]), .B(\ADD_/c[79] ), .Z(
        \ADD_/FAINST[79].FA_/n1 ) );
  XOR \ADD_/FAINST[78].FA_/U5  ( .A(\ADD_/FAINST[78].FA_/n3 ), .B(\ADD_/c[78] ), .Z(\ADD_/c[79] ) );
  XOR \ADD_/FAINST[78].FA_/U4  ( .A(\ADD_/FAINST[78].FA_/n1 ), .B(b[78]), .Z(
        c[78]) );
  AND \ADD_/FAINST[78].FA_/U3  ( .A(\ADD_/FAINST[78].FA_/n1 ), .B(
        \ADD_/FAINST[78].FA_/n2 ), .Z(\ADD_/FAINST[78].FA_/n3 ) );
  XOR \ADD_/FAINST[78].FA_/U2  ( .A(b[78]), .B(\ADD_/c[78] ), .Z(
        \ADD_/FAINST[78].FA_/n2 ) );
  XOR \ADD_/FAINST[78].FA_/U1  ( .A(a[78]), .B(\ADD_/c[78] ), .Z(
        \ADD_/FAINST[78].FA_/n1 ) );
  XOR \ADD_/FAINST[77].FA_/U5  ( .A(\ADD_/FAINST[77].FA_/n3 ), .B(\ADD_/c[77] ), .Z(\ADD_/c[78] ) );
  XOR \ADD_/FAINST[77].FA_/U4  ( .A(\ADD_/FAINST[77].FA_/n1 ), .B(b[77]), .Z(
        c[77]) );
  AND \ADD_/FAINST[77].FA_/U3  ( .A(\ADD_/FAINST[77].FA_/n1 ), .B(
        \ADD_/FAINST[77].FA_/n2 ), .Z(\ADD_/FAINST[77].FA_/n3 ) );
  XOR \ADD_/FAINST[77].FA_/U2  ( .A(b[77]), .B(\ADD_/c[77] ), .Z(
        \ADD_/FAINST[77].FA_/n2 ) );
  XOR \ADD_/FAINST[77].FA_/U1  ( .A(a[77]), .B(\ADD_/c[77] ), .Z(
        \ADD_/FAINST[77].FA_/n1 ) );
  XOR \ADD_/FAINST[76].FA_/U5  ( .A(\ADD_/FAINST[76].FA_/n3 ), .B(\ADD_/c[76] ), .Z(\ADD_/c[77] ) );
  XOR \ADD_/FAINST[76].FA_/U4  ( .A(\ADD_/FAINST[76].FA_/n1 ), .B(b[76]), .Z(
        c[76]) );
  AND \ADD_/FAINST[76].FA_/U3  ( .A(\ADD_/FAINST[76].FA_/n1 ), .B(
        \ADD_/FAINST[76].FA_/n2 ), .Z(\ADD_/FAINST[76].FA_/n3 ) );
  XOR \ADD_/FAINST[76].FA_/U2  ( .A(b[76]), .B(\ADD_/c[76] ), .Z(
        \ADD_/FAINST[76].FA_/n2 ) );
  XOR \ADD_/FAINST[76].FA_/U1  ( .A(a[76]), .B(\ADD_/c[76] ), .Z(
        \ADD_/FAINST[76].FA_/n1 ) );
  XOR \ADD_/FAINST[75].FA_/U5  ( .A(\ADD_/FAINST[75].FA_/n3 ), .B(\ADD_/c[75] ), .Z(\ADD_/c[76] ) );
  XOR \ADD_/FAINST[75].FA_/U4  ( .A(\ADD_/FAINST[75].FA_/n1 ), .B(b[75]), .Z(
        c[75]) );
  AND \ADD_/FAINST[75].FA_/U3  ( .A(\ADD_/FAINST[75].FA_/n1 ), .B(
        \ADD_/FAINST[75].FA_/n2 ), .Z(\ADD_/FAINST[75].FA_/n3 ) );
  XOR \ADD_/FAINST[75].FA_/U2  ( .A(b[75]), .B(\ADD_/c[75] ), .Z(
        \ADD_/FAINST[75].FA_/n2 ) );
  XOR \ADD_/FAINST[75].FA_/U1  ( .A(a[75]), .B(\ADD_/c[75] ), .Z(
        \ADD_/FAINST[75].FA_/n1 ) );
  XOR \ADD_/FAINST[74].FA_/U5  ( .A(\ADD_/FAINST[74].FA_/n3 ), .B(\ADD_/c[74] ), .Z(\ADD_/c[75] ) );
  XOR \ADD_/FAINST[74].FA_/U4  ( .A(\ADD_/FAINST[74].FA_/n1 ), .B(b[74]), .Z(
        c[74]) );
  AND \ADD_/FAINST[74].FA_/U3  ( .A(\ADD_/FAINST[74].FA_/n1 ), .B(
        \ADD_/FAINST[74].FA_/n2 ), .Z(\ADD_/FAINST[74].FA_/n3 ) );
  XOR \ADD_/FAINST[74].FA_/U2  ( .A(b[74]), .B(\ADD_/c[74] ), .Z(
        \ADD_/FAINST[74].FA_/n2 ) );
  XOR \ADD_/FAINST[74].FA_/U1  ( .A(a[74]), .B(\ADD_/c[74] ), .Z(
        \ADD_/FAINST[74].FA_/n1 ) );
  XOR \ADD_/FAINST[73].FA_/U5  ( .A(\ADD_/FAINST[73].FA_/n3 ), .B(\ADD_/c[73] ), .Z(\ADD_/c[74] ) );
  XOR \ADD_/FAINST[73].FA_/U4  ( .A(\ADD_/FAINST[73].FA_/n1 ), .B(b[73]), .Z(
        c[73]) );
  AND \ADD_/FAINST[73].FA_/U3  ( .A(\ADD_/FAINST[73].FA_/n1 ), .B(
        \ADD_/FAINST[73].FA_/n2 ), .Z(\ADD_/FAINST[73].FA_/n3 ) );
  XOR \ADD_/FAINST[73].FA_/U2  ( .A(b[73]), .B(\ADD_/c[73] ), .Z(
        \ADD_/FAINST[73].FA_/n2 ) );
  XOR \ADD_/FAINST[73].FA_/U1  ( .A(a[73]), .B(\ADD_/c[73] ), .Z(
        \ADD_/FAINST[73].FA_/n1 ) );
  XOR \ADD_/FAINST[72].FA_/U5  ( .A(\ADD_/FAINST[72].FA_/n3 ), .B(\ADD_/c[72] ), .Z(\ADD_/c[73] ) );
  XOR \ADD_/FAINST[72].FA_/U4  ( .A(\ADD_/FAINST[72].FA_/n1 ), .B(b[72]), .Z(
        c[72]) );
  AND \ADD_/FAINST[72].FA_/U3  ( .A(\ADD_/FAINST[72].FA_/n1 ), .B(
        \ADD_/FAINST[72].FA_/n2 ), .Z(\ADD_/FAINST[72].FA_/n3 ) );
  XOR \ADD_/FAINST[72].FA_/U2  ( .A(b[72]), .B(\ADD_/c[72] ), .Z(
        \ADD_/FAINST[72].FA_/n2 ) );
  XOR \ADD_/FAINST[72].FA_/U1  ( .A(a[72]), .B(\ADD_/c[72] ), .Z(
        \ADD_/FAINST[72].FA_/n1 ) );
  XOR \ADD_/FAINST[71].FA_/U5  ( .A(\ADD_/FAINST[71].FA_/n3 ), .B(\ADD_/c[71] ), .Z(\ADD_/c[72] ) );
  XOR \ADD_/FAINST[71].FA_/U4  ( .A(\ADD_/FAINST[71].FA_/n1 ), .B(b[71]), .Z(
        c[71]) );
  AND \ADD_/FAINST[71].FA_/U3  ( .A(\ADD_/FAINST[71].FA_/n1 ), .B(
        \ADD_/FAINST[71].FA_/n2 ), .Z(\ADD_/FAINST[71].FA_/n3 ) );
  XOR \ADD_/FAINST[71].FA_/U2  ( .A(b[71]), .B(\ADD_/c[71] ), .Z(
        \ADD_/FAINST[71].FA_/n2 ) );
  XOR \ADD_/FAINST[71].FA_/U1  ( .A(a[71]), .B(\ADD_/c[71] ), .Z(
        \ADD_/FAINST[71].FA_/n1 ) );
  XOR \ADD_/FAINST[70].FA_/U5  ( .A(\ADD_/FAINST[70].FA_/n3 ), .B(\ADD_/c[70] ), .Z(\ADD_/c[71] ) );
  XOR \ADD_/FAINST[70].FA_/U4  ( .A(\ADD_/FAINST[70].FA_/n1 ), .B(b[70]), .Z(
        c[70]) );
  AND \ADD_/FAINST[70].FA_/U3  ( .A(\ADD_/FAINST[70].FA_/n1 ), .B(
        \ADD_/FAINST[70].FA_/n2 ), .Z(\ADD_/FAINST[70].FA_/n3 ) );
  XOR \ADD_/FAINST[70].FA_/U2  ( .A(b[70]), .B(\ADD_/c[70] ), .Z(
        \ADD_/FAINST[70].FA_/n2 ) );
  XOR \ADD_/FAINST[70].FA_/U1  ( .A(a[70]), .B(\ADD_/c[70] ), .Z(
        \ADD_/FAINST[70].FA_/n1 ) );
  XOR \ADD_/FAINST[69].FA_/U5  ( .A(\ADD_/FAINST[69].FA_/n3 ), .B(\ADD_/c[69] ), .Z(\ADD_/c[70] ) );
  XOR \ADD_/FAINST[69].FA_/U4  ( .A(\ADD_/FAINST[69].FA_/n1 ), .B(b[69]), .Z(
        c[69]) );
  AND \ADD_/FAINST[69].FA_/U3  ( .A(\ADD_/FAINST[69].FA_/n1 ), .B(
        \ADD_/FAINST[69].FA_/n2 ), .Z(\ADD_/FAINST[69].FA_/n3 ) );
  XOR \ADD_/FAINST[69].FA_/U2  ( .A(b[69]), .B(\ADD_/c[69] ), .Z(
        \ADD_/FAINST[69].FA_/n2 ) );
  XOR \ADD_/FAINST[69].FA_/U1  ( .A(a[69]), .B(\ADD_/c[69] ), .Z(
        \ADD_/FAINST[69].FA_/n1 ) );
  XOR \ADD_/FAINST[68].FA_/U5  ( .A(\ADD_/FAINST[68].FA_/n3 ), .B(\ADD_/c[68] ), .Z(\ADD_/c[69] ) );
  XOR \ADD_/FAINST[68].FA_/U4  ( .A(\ADD_/FAINST[68].FA_/n1 ), .B(b[68]), .Z(
        c[68]) );
  AND \ADD_/FAINST[68].FA_/U3  ( .A(\ADD_/FAINST[68].FA_/n1 ), .B(
        \ADD_/FAINST[68].FA_/n2 ), .Z(\ADD_/FAINST[68].FA_/n3 ) );
  XOR \ADD_/FAINST[68].FA_/U2  ( .A(b[68]), .B(\ADD_/c[68] ), .Z(
        \ADD_/FAINST[68].FA_/n2 ) );
  XOR \ADD_/FAINST[68].FA_/U1  ( .A(a[68]), .B(\ADD_/c[68] ), .Z(
        \ADD_/FAINST[68].FA_/n1 ) );
  XOR \ADD_/FAINST[67].FA_/U5  ( .A(\ADD_/FAINST[67].FA_/n3 ), .B(\ADD_/c[67] ), .Z(\ADD_/c[68] ) );
  XOR \ADD_/FAINST[67].FA_/U4  ( .A(\ADD_/FAINST[67].FA_/n1 ), .B(b[67]), .Z(
        c[67]) );
  AND \ADD_/FAINST[67].FA_/U3  ( .A(\ADD_/FAINST[67].FA_/n1 ), .B(
        \ADD_/FAINST[67].FA_/n2 ), .Z(\ADD_/FAINST[67].FA_/n3 ) );
  XOR \ADD_/FAINST[67].FA_/U2  ( .A(b[67]), .B(\ADD_/c[67] ), .Z(
        \ADD_/FAINST[67].FA_/n2 ) );
  XOR \ADD_/FAINST[67].FA_/U1  ( .A(a[67]), .B(\ADD_/c[67] ), .Z(
        \ADD_/FAINST[67].FA_/n1 ) );
  XOR \ADD_/FAINST[66].FA_/U5  ( .A(\ADD_/FAINST[66].FA_/n3 ), .B(\ADD_/c[66] ), .Z(\ADD_/c[67] ) );
  XOR \ADD_/FAINST[66].FA_/U4  ( .A(\ADD_/FAINST[66].FA_/n1 ), .B(b[66]), .Z(
        c[66]) );
  AND \ADD_/FAINST[66].FA_/U3  ( .A(\ADD_/FAINST[66].FA_/n1 ), .B(
        \ADD_/FAINST[66].FA_/n2 ), .Z(\ADD_/FAINST[66].FA_/n3 ) );
  XOR \ADD_/FAINST[66].FA_/U2  ( .A(b[66]), .B(\ADD_/c[66] ), .Z(
        \ADD_/FAINST[66].FA_/n2 ) );
  XOR \ADD_/FAINST[66].FA_/U1  ( .A(a[66]), .B(\ADD_/c[66] ), .Z(
        \ADD_/FAINST[66].FA_/n1 ) );
  XOR \ADD_/FAINST[65].FA_/U5  ( .A(\ADD_/FAINST[65].FA_/n3 ), .B(\ADD_/c[65] ), .Z(\ADD_/c[66] ) );
  XOR \ADD_/FAINST[65].FA_/U4  ( .A(\ADD_/FAINST[65].FA_/n1 ), .B(b[65]), .Z(
        c[65]) );
  AND \ADD_/FAINST[65].FA_/U3  ( .A(\ADD_/FAINST[65].FA_/n1 ), .B(
        \ADD_/FAINST[65].FA_/n2 ), .Z(\ADD_/FAINST[65].FA_/n3 ) );
  XOR \ADD_/FAINST[65].FA_/U2  ( .A(b[65]), .B(\ADD_/c[65] ), .Z(
        \ADD_/FAINST[65].FA_/n2 ) );
  XOR \ADD_/FAINST[65].FA_/U1  ( .A(a[65]), .B(\ADD_/c[65] ), .Z(
        \ADD_/FAINST[65].FA_/n1 ) );
  XOR \ADD_/FAINST[64].FA_/U5  ( .A(\ADD_/FAINST[64].FA_/n3 ), .B(\ADD_/c[64] ), .Z(\ADD_/c[65] ) );
  XOR \ADD_/FAINST[64].FA_/U4  ( .A(\ADD_/FAINST[64].FA_/n1 ), .B(b[64]), .Z(
        c[64]) );
  AND \ADD_/FAINST[64].FA_/U3  ( .A(\ADD_/FAINST[64].FA_/n1 ), .B(
        \ADD_/FAINST[64].FA_/n2 ), .Z(\ADD_/FAINST[64].FA_/n3 ) );
  XOR \ADD_/FAINST[64].FA_/U2  ( .A(b[64]), .B(\ADD_/c[64] ), .Z(
        \ADD_/FAINST[64].FA_/n2 ) );
  XOR \ADD_/FAINST[64].FA_/U1  ( .A(a[64]), .B(\ADD_/c[64] ), .Z(
        \ADD_/FAINST[64].FA_/n1 ) );
  XOR \ADD_/FAINST[63].FA_/U5  ( .A(\ADD_/FAINST[63].FA_/n3 ), .B(\ADD_/c[63] ), .Z(\ADD_/c[64] ) );
  XOR \ADD_/FAINST[63].FA_/U4  ( .A(\ADD_/FAINST[63].FA_/n1 ), .B(b[63]), .Z(
        c[63]) );
  AND \ADD_/FAINST[63].FA_/U3  ( .A(\ADD_/FAINST[63].FA_/n1 ), .B(
        \ADD_/FAINST[63].FA_/n2 ), .Z(\ADD_/FAINST[63].FA_/n3 ) );
  XOR \ADD_/FAINST[63].FA_/U2  ( .A(b[63]), .B(\ADD_/c[63] ), .Z(
        \ADD_/FAINST[63].FA_/n2 ) );
  XOR \ADD_/FAINST[63].FA_/U1  ( .A(a[63]), .B(\ADD_/c[63] ), .Z(
        \ADD_/FAINST[63].FA_/n1 ) );
  XOR \ADD_/FAINST[62].FA_/U5  ( .A(\ADD_/FAINST[62].FA_/n3 ), .B(\ADD_/c[62] ), .Z(\ADD_/c[63] ) );
  XOR \ADD_/FAINST[62].FA_/U4  ( .A(\ADD_/FAINST[62].FA_/n1 ), .B(b[62]), .Z(
        c[62]) );
  AND \ADD_/FAINST[62].FA_/U3  ( .A(\ADD_/FAINST[62].FA_/n1 ), .B(
        \ADD_/FAINST[62].FA_/n2 ), .Z(\ADD_/FAINST[62].FA_/n3 ) );
  XOR \ADD_/FAINST[62].FA_/U2  ( .A(b[62]), .B(\ADD_/c[62] ), .Z(
        \ADD_/FAINST[62].FA_/n2 ) );
  XOR \ADD_/FAINST[62].FA_/U1  ( .A(a[62]), .B(\ADD_/c[62] ), .Z(
        \ADD_/FAINST[62].FA_/n1 ) );
  XOR \ADD_/FAINST[61].FA_/U5  ( .A(\ADD_/FAINST[61].FA_/n3 ), .B(\ADD_/c[61] ), .Z(\ADD_/c[62] ) );
  XOR \ADD_/FAINST[61].FA_/U4  ( .A(\ADD_/FAINST[61].FA_/n1 ), .B(b[61]), .Z(
        c[61]) );
  AND \ADD_/FAINST[61].FA_/U3  ( .A(\ADD_/FAINST[61].FA_/n1 ), .B(
        \ADD_/FAINST[61].FA_/n2 ), .Z(\ADD_/FAINST[61].FA_/n3 ) );
  XOR \ADD_/FAINST[61].FA_/U2  ( .A(b[61]), .B(\ADD_/c[61] ), .Z(
        \ADD_/FAINST[61].FA_/n2 ) );
  XOR \ADD_/FAINST[61].FA_/U1  ( .A(a[61]), .B(\ADD_/c[61] ), .Z(
        \ADD_/FAINST[61].FA_/n1 ) );
  XOR \ADD_/FAINST[60].FA_/U5  ( .A(\ADD_/FAINST[60].FA_/n3 ), .B(\ADD_/c[60] ), .Z(\ADD_/c[61] ) );
  XOR \ADD_/FAINST[60].FA_/U4  ( .A(\ADD_/FAINST[60].FA_/n1 ), .B(b[60]), .Z(
        c[60]) );
  AND \ADD_/FAINST[60].FA_/U3  ( .A(\ADD_/FAINST[60].FA_/n1 ), .B(
        \ADD_/FAINST[60].FA_/n2 ), .Z(\ADD_/FAINST[60].FA_/n3 ) );
  XOR \ADD_/FAINST[60].FA_/U2  ( .A(b[60]), .B(\ADD_/c[60] ), .Z(
        \ADD_/FAINST[60].FA_/n2 ) );
  XOR \ADD_/FAINST[60].FA_/U1  ( .A(a[60]), .B(\ADD_/c[60] ), .Z(
        \ADD_/FAINST[60].FA_/n1 ) );
  XOR \ADD_/FAINST[59].FA_/U5  ( .A(\ADD_/FAINST[59].FA_/n3 ), .B(\ADD_/c[59] ), .Z(\ADD_/c[60] ) );
  XOR \ADD_/FAINST[59].FA_/U4  ( .A(\ADD_/FAINST[59].FA_/n1 ), .B(b[59]), .Z(
        c[59]) );
  AND \ADD_/FAINST[59].FA_/U3  ( .A(\ADD_/FAINST[59].FA_/n1 ), .B(
        \ADD_/FAINST[59].FA_/n2 ), .Z(\ADD_/FAINST[59].FA_/n3 ) );
  XOR \ADD_/FAINST[59].FA_/U2  ( .A(b[59]), .B(\ADD_/c[59] ), .Z(
        \ADD_/FAINST[59].FA_/n2 ) );
  XOR \ADD_/FAINST[59].FA_/U1  ( .A(a[59]), .B(\ADD_/c[59] ), .Z(
        \ADD_/FAINST[59].FA_/n1 ) );
  XOR \ADD_/FAINST[58].FA_/U5  ( .A(\ADD_/FAINST[58].FA_/n3 ), .B(\ADD_/c[58] ), .Z(\ADD_/c[59] ) );
  XOR \ADD_/FAINST[58].FA_/U4  ( .A(\ADD_/FAINST[58].FA_/n1 ), .B(b[58]), .Z(
        c[58]) );
  AND \ADD_/FAINST[58].FA_/U3  ( .A(\ADD_/FAINST[58].FA_/n1 ), .B(
        \ADD_/FAINST[58].FA_/n2 ), .Z(\ADD_/FAINST[58].FA_/n3 ) );
  XOR \ADD_/FAINST[58].FA_/U2  ( .A(b[58]), .B(\ADD_/c[58] ), .Z(
        \ADD_/FAINST[58].FA_/n2 ) );
  XOR \ADD_/FAINST[58].FA_/U1  ( .A(a[58]), .B(\ADD_/c[58] ), .Z(
        \ADD_/FAINST[58].FA_/n1 ) );
  XOR \ADD_/FAINST[57].FA_/U5  ( .A(\ADD_/FAINST[57].FA_/n3 ), .B(\ADD_/c[57] ), .Z(\ADD_/c[58] ) );
  XOR \ADD_/FAINST[57].FA_/U4  ( .A(\ADD_/FAINST[57].FA_/n1 ), .B(b[57]), .Z(
        c[57]) );
  AND \ADD_/FAINST[57].FA_/U3  ( .A(\ADD_/FAINST[57].FA_/n1 ), .B(
        \ADD_/FAINST[57].FA_/n2 ), .Z(\ADD_/FAINST[57].FA_/n3 ) );
  XOR \ADD_/FAINST[57].FA_/U2  ( .A(b[57]), .B(\ADD_/c[57] ), .Z(
        \ADD_/FAINST[57].FA_/n2 ) );
  XOR \ADD_/FAINST[57].FA_/U1  ( .A(a[57]), .B(\ADD_/c[57] ), .Z(
        \ADD_/FAINST[57].FA_/n1 ) );
  XOR \ADD_/FAINST[56].FA_/U5  ( .A(\ADD_/FAINST[56].FA_/n3 ), .B(\ADD_/c[56] ), .Z(\ADD_/c[57] ) );
  XOR \ADD_/FAINST[56].FA_/U4  ( .A(\ADD_/FAINST[56].FA_/n1 ), .B(b[56]), .Z(
        c[56]) );
  AND \ADD_/FAINST[56].FA_/U3  ( .A(\ADD_/FAINST[56].FA_/n1 ), .B(
        \ADD_/FAINST[56].FA_/n2 ), .Z(\ADD_/FAINST[56].FA_/n3 ) );
  XOR \ADD_/FAINST[56].FA_/U2  ( .A(b[56]), .B(\ADD_/c[56] ), .Z(
        \ADD_/FAINST[56].FA_/n2 ) );
  XOR \ADD_/FAINST[56].FA_/U1  ( .A(a[56]), .B(\ADD_/c[56] ), .Z(
        \ADD_/FAINST[56].FA_/n1 ) );
  XOR \ADD_/FAINST[55].FA_/U5  ( .A(\ADD_/FAINST[55].FA_/n3 ), .B(\ADD_/c[55] ), .Z(\ADD_/c[56] ) );
  XOR \ADD_/FAINST[55].FA_/U4  ( .A(\ADD_/FAINST[55].FA_/n1 ), .B(b[55]), .Z(
        c[55]) );
  AND \ADD_/FAINST[55].FA_/U3  ( .A(\ADD_/FAINST[55].FA_/n1 ), .B(
        \ADD_/FAINST[55].FA_/n2 ), .Z(\ADD_/FAINST[55].FA_/n3 ) );
  XOR \ADD_/FAINST[55].FA_/U2  ( .A(b[55]), .B(\ADD_/c[55] ), .Z(
        \ADD_/FAINST[55].FA_/n2 ) );
  XOR \ADD_/FAINST[55].FA_/U1  ( .A(a[55]), .B(\ADD_/c[55] ), .Z(
        \ADD_/FAINST[55].FA_/n1 ) );
  XOR \ADD_/FAINST[54].FA_/U5  ( .A(\ADD_/FAINST[54].FA_/n3 ), .B(\ADD_/c[54] ), .Z(\ADD_/c[55] ) );
  XOR \ADD_/FAINST[54].FA_/U4  ( .A(\ADD_/FAINST[54].FA_/n1 ), .B(b[54]), .Z(
        c[54]) );
  AND \ADD_/FAINST[54].FA_/U3  ( .A(\ADD_/FAINST[54].FA_/n1 ), .B(
        \ADD_/FAINST[54].FA_/n2 ), .Z(\ADD_/FAINST[54].FA_/n3 ) );
  XOR \ADD_/FAINST[54].FA_/U2  ( .A(b[54]), .B(\ADD_/c[54] ), .Z(
        \ADD_/FAINST[54].FA_/n2 ) );
  XOR \ADD_/FAINST[54].FA_/U1  ( .A(a[54]), .B(\ADD_/c[54] ), .Z(
        \ADD_/FAINST[54].FA_/n1 ) );
  XOR \ADD_/FAINST[53].FA_/U5  ( .A(\ADD_/FAINST[53].FA_/n3 ), .B(\ADD_/c[53] ), .Z(\ADD_/c[54] ) );
  XOR \ADD_/FAINST[53].FA_/U4  ( .A(\ADD_/FAINST[53].FA_/n1 ), .B(b[53]), .Z(
        c[53]) );
  AND \ADD_/FAINST[53].FA_/U3  ( .A(\ADD_/FAINST[53].FA_/n1 ), .B(
        \ADD_/FAINST[53].FA_/n2 ), .Z(\ADD_/FAINST[53].FA_/n3 ) );
  XOR \ADD_/FAINST[53].FA_/U2  ( .A(b[53]), .B(\ADD_/c[53] ), .Z(
        \ADD_/FAINST[53].FA_/n2 ) );
  XOR \ADD_/FAINST[53].FA_/U1  ( .A(a[53]), .B(\ADD_/c[53] ), .Z(
        \ADD_/FAINST[53].FA_/n1 ) );
  XOR \ADD_/FAINST[52].FA_/U5  ( .A(\ADD_/FAINST[52].FA_/n3 ), .B(\ADD_/c[52] ), .Z(\ADD_/c[53] ) );
  XOR \ADD_/FAINST[52].FA_/U4  ( .A(\ADD_/FAINST[52].FA_/n1 ), .B(b[52]), .Z(
        c[52]) );
  AND \ADD_/FAINST[52].FA_/U3  ( .A(\ADD_/FAINST[52].FA_/n1 ), .B(
        \ADD_/FAINST[52].FA_/n2 ), .Z(\ADD_/FAINST[52].FA_/n3 ) );
  XOR \ADD_/FAINST[52].FA_/U2  ( .A(b[52]), .B(\ADD_/c[52] ), .Z(
        \ADD_/FAINST[52].FA_/n2 ) );
  XOR \ADD_/FAINST[52].FA_/U1  ( .A(a[52]), .B(\ADD_/c[52] ), .Z(
        \ADD_/FAINST[52].FA_/n1 ) );
  XOR \ADD_/FAINST[51].FA_/U5  ( .A(\ADD_/FAINST[51].FA_/n3 ), .B(\ADD_/c[51] ), .Z(\ADD_/c[52] ) );
  XOR \ADD_/FAINST[51].FA_/U4  ( .A(\ADD_/FAINST[51].FA_/n1 ), .B(b[51]), .Z(
        c[51]) );
  AND \ADD_/FAINST[51].FA_/U3  ( .A(\ADD_/FAINST[51].FA_/n1 ), .B(
        \ADD_/FAINST[51].FA_/n2 ), .Z(\ADD_/FAINST[51].FA_/n3 ) );
  XOR \ADD_/FAINST[51].FA_/U2  ( .A(b[51]), .B(\ADD_/c[51] ), .Z(
        \ADD_/FAINST[51].FA_/n2 ) );
  XOR \ADD_/FAINST[51].FA_/U1  ( .A(a[51]), .B(\ADD_/c[51] ), .Z(
        \ADD_/FAINST[51].FA_/n1 ) );
  XOR \ADD_/FAINST[50].FA_/U5  ( .A(\ADD_/FAINST[50].FA_/n3 ), .B(\ADD_/c[50] ), .Z(\ADD_/c[51] ) );
  XOR \ADD_/FAINST[50].FA_/U4  ( .A(\ADD_/FAINST[50].FA_/n1 ), .B(b[50]), .Z(
        c[50]) );
  AND \ADD_/FAINST[50].FA_/U3  ( .A(\ADD_/FAINST[50].FA_/n1 ), .B(
        \ADD_/FAINST[50].FA_/n2 ), .Z(\ADD_/FAINST[50].FA_/n3 ) );
  XOR \ADD_/FAINST[50].FA_/U2  ( .A(b[50]), .B(\ADD_/c[50] ), .Z(
        \ADD_/FAINST[50].FA_/n2 ) );
  XOR \ADD_/FAINST[50].FA_/U1  ( .A(a[50]), .B(\ADD_/c[50] ), .Z(
        \ADD_/FAINST[50].FA_/n1 ) );
  XOR \ADD_/FAINST[49].FA_/U5  ( .A(\ADD_/FAINST[49].FA_/n3 ), .B(\ADD_/c[49] ), .Z(\ADD_/c[50] ) );
  XOR \ADD_/FAINST[49].FA_/U4  ( .A(\ADD_/FAINST[49].FA_/n1 ), .B(b[49]), .Z(
        c[49]) );
  AND \ADD_/FAINST[49].FA_/U3  ( .A(\ADD_/FAINST[49].FA_/n1 ), .B(
        \ADD_/FAINST[49].FA_/n2 ), .Z(\ADD_/FAINST[49].FA_/n3 ) );
  XOR \ADD_/FAINST[49].FA_/U2  ( .A(b[49]), .B(\ADD_/c[49] ), .Z(
        \ADD_/FAINST[49].FA_/n2 ) );
  XOR \ADD_/FAINST[49].FA_/U1  ( .A(a[49]), .B(\ADD_/c[49] ), .Z(
        \ADD_/FAINST[49].FA_/n1 ) );
  XOR \ADD_/FAINST[48].FA_/U5  ( .A(\ADD_/FAINST[48].FA_/n3 ), .B(\ADD_/c[48] ), .Z(\ADD_/c[49] ) );
  XOR \ADD_/FAINST[48].FA_/U4  ( .A(\ADD_/FAINST[48].FA_/n1 ), .B(b[48]), .Z(
        c[48]) );
  AND \ADD_/FAINST[48].FA_/U3  ( .A(\ADD_/FAINST[48].FA_/n1 ), .B(
        \ADD_/FAINST[48].FA_/n2 ), .Z(\ADD_/FAINST[48].FA_/n3 ) );
  XOR \ADD_/FAINST[48].FA_/U2  ( .A(b[48]), .B(\ADD_/c[48] ), .Z(
        \ADD_/FAINST[48].FA_/n2 ) );
  XOR \ADD_/FAINST[48].FA_/U1  ( .A(a[48]), .B(\ADD_/c[48] ), .Z(
        \ADD_/FAINST[48].FA_/n1 ) );
  XOR \ADD_/FAINST[47].FA_/U5  ( .A(\ADD_/FAINST[47].FA_/n3 ), .B(\ADD_/c[47] ), .Z(\ADD_/c[48] ) );
  XOR \ADD_/FAINST[47].FA_/U4  ( .A(\ADD_/FAINST[47].FA_/n1 ), .B(b[47]), .Z(
        c[47]) );
  AND \ADD_/FAINST[47].FA_/U3  ( .A(\ADD_/FAINST[47].FA_/n1 ), .B(
        \ADD_/FAINST[47].FA_/n2 ), .Z(\ADD_/FAINST[47].FA_/n3 ) );
  XOR \ADD_/FAINST[47].FA_/U2  ( .A(b[47]), .B(\ADD_/c[47] ), .Z(
        \ADD_/FAINST[47].FA_/n2 ) );
  XOR \ADD_/FAINST[47].FA_/U1  ( .A(a[47]), .B(\ADD_/c[47] ), .Z(
        \ADD_/FAINST[47].FA_/n1 ) );
  XOR \ADD_/FAINST[46].FA_/U5  ( .A(\ADD_/FAINST[46].FA_/n3 ), .B(\ADD_/c[46] ), .Z(\ADD_/c[47] ) );
  XOR \ADD_/FAINST[46].FA_/U4  ( .A(\ADD_/FAINST[46].FA_/n1 ), .B(b[46]), .Z(
        c[46]) );
  AND \ADD_/FAINST[46].FA_/U3  ( .A(\ADD_/FAINST[46].FA_/n1 ), .B(
        \ADD_/FAINST[46].FA_/n2 ), .Z(\ADD_/FAINST[46].FA_/n3 ) );
  XOR \ADD_/FAINST[46].FA_/U2  ( .A(b[46]), .B(\ADD_/c[46] ), .Z(
        \ADD_/FAINST[46].FA_/n2 ) );
  XOR \ADD_/FAINST[46].FA_/U1  ( .A(a[46]), .B(\ADD_/c[46] ), .Z(
        \ADD_/FAINST[46].FA_/n1 ) );
  XOR \ADD_/FAINST[45].FA_/U5  ( .A(\ADD_/FAINST[45].FA_/n3 ), .B(\ADD_/c[45] ), .Z(\ADD_/c[46] ) );
  XOR \ADD_/FAINST[45].FA_/U4  ( .A(\ADD_/FAINST[45].FA_/n1 ), .B(b[45]), .Z(
        c[45]) );
  AND \ADD_/FAINST[45].FA_/U3  ( .A(\ADD_/FAINST[45].FA_/n1 ), .B(
        \ADD_/FAINST[45].FA_/n2 ), .Z(\ADD_/FAINST[45].FA_/n3 ) );
  XOR \ADD_/FAINST[45].FA_/U2  ( .A(b[45]), .B(\ADD_/c[45] ), .Z(
        \ADD_/FAINST[45].FA_/n2 ) );
  XOR \ADD_/FAINST[45].FA_/U1  ( .A(a[45]), .B(\ADD_/c[45] ), .Z(
        \ADD_/FAINST[45].FA_/n1 ) );
  XOR \ADD_/FAINST[44].FA_/U5  ( .A(\ADD_/FAINST[44].FA_/n3 ), .B(\ADD_/c[44] ), .Z(\ADD_/c[45] ) );
  XOR \ADD_/FAINST[44].FA_/U4  ( .A(\ADD_/FAINST[44].FA_/n1 ), .B(b[44]), .Z(
        c[44]) );
  AND \ADD_/FAINST[44].FA_/U3  ( .A(\ADD_/FAINST[44].FA_/n1 ), .B(
        \ADD_/FAINST[44].FA_/n2 ), .Z(\ADD_/FAINST[44].FA_/n3 ) );
  XOR \ADD_/FAINST[44].FA_/U2  ( .A(b[44]), .B(\ADD_/c[44] ), .Z(
        \ADD_/FAINST[44].FA_/n2 ) );
  XOR \ADD_/FAINST[44].FA_/U1  ( .A(a[44]), .B(\ADD_/c[44] ), .Z(
        \ADD_/FAINST[44].FA_/n1 ) );
  XOR \ADD_/FAINST[43].FA_/U5  ( .A(\ADD_/FAINST[43].FA_/n3 ), .B(\ADD_/c[43] ), .Z(\ADD_/c[44] ) );
  XOR \ADD_/FAINST[43].FA_/U4  ( .A(\ADD_/FAINST[43].FA_/n1 ), .B(b[43]), .Z(
        c[43]) );
  AND \ADD_/FAINST[43].FA_/U3  ( .A(\ADD_/FAINST[43].FA_/n1 ), .B(
        \ADD_/FAINST[43].FA_/n2 ), .Z(\ADD_/FAINST[43].FA_/n3 ) );
  XOR \ADD_/FAINST[43].FA_/U2  ( .A(b[43]), .B(\ADD_/c[43] ), .Z(
        \ADD_/FAINST[43].FA_/n2 ) );
  XOR \ADD_/FAINST[43].FA_/U1  ( .A(a[43]), .B(\ADD_/c[43] ), .Z(
        \ADD_/FAINST[43].FA_/n1 ) );
  XOR \ADD_/FAINST[42].FA_/U5  ( .A(\ADD_/FAINST[42].FA_/n3 ), .B(\ADD_/c[42] ), .Z(\ADD_/c[43] ) );
  XOR \ADD_/FAINST[42].FA_/U4  ( .A(\ADD_/FAINST[42].FA_/n1 ), .B(b[42]), .Z(
        c[42]) );
  AND \ADD_/FAINST[42].FA_/U3  ( .A(\ADD_/FAINST[42].FA_/n1 ), .B(
        \ADD_/FAINST[42].FA_/n2 ), .Z(\ADD_/FAINST[42].FA_/n3 ) );
  XOR \ADD_/FAINST[42].FA_/U2  ( .A(b[42]), .B(\ADD_/c[42] ), .Z(
        \ADD_/FAINST[42].FA_/n2 ) );
  XOR \ADD_/FAINST[42].FA_/U1  ( .A(a[42]), .B(\ADD_/c[42] ), .Z(
        \ADD_/FAINST[42].FA_/n1 ) );
  XOR \ADD_/FAINST[41].FA_/U5  ( .A(\ADD_/FAINST[41].FA_/n3 ), .B(\ADD_/c[41] ), .Z(\ADD_/c[42] ) );
  XOR \ADD_/FAINST[41].FA_/U4  ( .A(\ADD_/FAINST[41].FA_/n1 ), .B(b[41]), .Z(
        c[41]) );
  AND \ADD_/FAINST[41].FA_/U3  ( .A(\ADD_/FAINST[41].FA_/n1 ), .B(
        \ADD_/FAINST[41].FA_/n2 ), .Z(\ADD_/FAINST[41].FA_/n3 ) );
  XOR \ADD_/FAINST[41].FA_/U2  ( .A(b[41]), .B(\ADD_/c[41] ), .Z(
        \ADD_/FAINST[41].FA_/n2 ) );
  XOR \ADD_/FAINST[41].FA_/U1  ( .A(a[41]), .B(\ADD_/c[41] ), .Z(
        \ADD_/FAINST[41].FA_/n1 ) );
  XOR \ADD_/FAINST[40].FA_/U5  ( .A(\ADD_/FAINST[40].FA_/n3 ), .B(\ADD_/c[40] ), .Z(\ADD_/c[41] ) );
  XOR \ADD_/FAINST[40].FA_/U4  ( .A(\ADD_/FAINST[40].FA_/n1 ), .B(b[40]), .Z(
        c[40]) );
  AND \ADD_/FAINST[40].FA_/U3  ( .A(\ADD_/FAINST[40].FA_/n1 ), .B(
        \ADD_/FAINST[40].FA_/n2 ), .Z(\ADD_/FAINST[40].FA_/n3 ) );
  XOR \ADD_/FAINST[40].FA_/U2  ( .A(b[40]), .B(\ADD_/c[40] ), .Z(
        \ADD_/FAINST[40].FA_/n2 ) );
  XOR \ADD_/FAINST[40].FA_/U1  ( .A(a[40]), .B(\ADD_/c[40] ), .Z(
        \ADD_/FAINST[40].FA_/n1 ) );
  XOR \ADD_/FAINST[39].FA_/U5  ( .A(\ADD_/FAINST[39].FA_/n3 ), .B(\ADD_/c[39] ), .Z(\ADD_/c[40] ) );
  XOR \ADD_/FAINST[39].FA_/U4  ( .A(\ADD_/FAINST[39].FA_/n1 ), .B(b[39]), .Z(
        c[39]) );
  AND \ADD_/FAINST[39].FA_/U3  ( .A(\ADD_/FAINST[39].FA_/n1 ), .B(
        \ADD_/FAINST[39].FA_/n2 ), .Z(\ADD_/FAINST[39].FA_/n3 ) );
  XOR \ADD_/FAINST[39].FA_/U2  ( .A(b[39]), .B(\ADD_/c[39] ), .Z(
        \ADD_/FAINST[39].FA_/n2 ) );
  XOR \ADD_/FAINST[39].FA_/U1  ( .A(a[39]), .B(\ADD_/c[39] ), .Z(
        \ADD_/FAINST[39].FA_/n1 ) );
  XOR \ADD_/FAINST[38].FA_/U5  ( .A(\ADD_/FAINST[38].FA_/n3 ), .B(\ADD_/c[38] ), .Z(\ADD_/c[39] ) );
  XOR \ADD_/FAINST[38].FA_/U4  ( .A(\ADD_/FAINST[38].FA_/n1 ), .B(b[38]), .Z(
        c[38]) );
  AND \ADD_/FAINST[38].FA_/U3  ( .A(\ADD_/FAINST[38].FA_/n1 ), .B(
        \ADD_/FAINST[38].FA_/n2 ), .Z(\ADD_/FAINST[38].FA_/n3 ) );
  XOR \ADD_/FAINST[38].FA_/U2  ( .A(b[38]), .B(\ADD_/c[38] ), .Z(
        \ADD_/FAINST[38].FA_/n2 ) );
  XOR \ADD_/FAINST[38].FA_/U1  ( .A(a[38]), .B(\ADD_/c[38] ), .Z(
        \ADD_/FAINST[38].FA_/n1 ) );
  XOR \ADD_/FAINST[37].FA_/U5  ( .A(\ADD_/FAINST[37].FA_/n3 ), .B(\ADD_/c[37] ), .Z(\ADD_/c[38] ) );
  XOR \ADD_/FAINST[37].FA_/U4  ( .A(\ADD_/FAINST[37].FA_/n1 ), .B(b[37]), .Z(
        c[37]) );
  AND \ADD_/FAINST[37].FA_/U3  ( .A(\ADD_/FAINST[37].FA_/n1 ), .B(
        \ADD_/FAINST[37].FA_/n2 ), .Z(\ADD_/FAINST[37].FA_/n3 ) );
  XOR \ADD_/FAINST[37].FA_/U2  ( .A(b[37]), .B(\ADD_/c[37] ), .Z(
        \ADD_/FAINST[37].FA_/n2 ) );
  XOR \ADD_/FAINST[37].FA_/U1  ( .A(a[37]), .B(\ADD_/c[37] ), .Z(
        \ADD_/FAINST[37].FA_/n1 ) );
  XOR \ADD_/FAINST[36].FA_/U5  ( .A(\ADD_/FAINST[36].FA_/n3 ), .B(\ADD_/c[36] ), .Z(\ADD_/c[37] ) );
  XOR \ADD_/FAINST[36].FA_/U4  ( .A(\ADD_/FAINST[36].FA_/n1 ), .B(b[36]), .Z(
        c[36]) );
  AND \ADD_/FAINST[36].FA_/U3  ( .A(\ADD_/FAINST[36].FA_/n1 ), .B(
        \ADD_/FAINST[36].FA_/n2 ), .Z(\ADD_/FAINST[36].FA_/n3 ) );
  XOR \ADD_/FAINST[36].FA_/U2  ( .A(b[36]), .B(\ADD_/c[36] ), .Z(
        \ADD_/FAINST[36].FA_/n2 ) );
  XOR \ADD_/FAINST[36].FA_/U1  ( .A(a[36]), .B(\ADD_/c[36] ), .Z(
        \ADD_/FAINST[36].FA_/n1 ) );
  XOR \ADD_/FAINST[35].FA_/U5  ( .A(\ADD_/FAINST[35].FA_/n3 ), .B(\ADD_/c[35] ), .Z(\ADD_/c[36] ) );
  XOR \ADD_/FAINST[35].FA_/U4  ( .A(\ADD_/FAINST[35].FA_/n1 ), .B(b[35]), .Z(
        c[35]) );
  AND \ADD_/FAINST[35].FA_/U3  ( .A(\ADD_/FAINST[35].FA_/n1 ), .B(
        \ADD_/FAINST[35].FA_/n2 ), .Z(\ADD_/FAINST[35].FA_/n3 ) );
  XOR \ADD_/FAINST[35].FA_/U2  ( .A(b[35]), .B(\ADD_/c[35] ), .Z(
        \ADD_/FAINST[35].FA_/n2 ) );
  XOR \ADD_/FAINST[35].FA_/U1  ( .A(a[35]), .B(\ADD_/c[35] ), .Z(
        \ADD_/FAINST[35].FA_/n1 ) );
  XOR \ADD_/FAINST[34].FA_/U5  ( .A(\ADD_/FAINST[34].FA_/n3 ), .B(\ADD_/c[34] ), .Z(\ADD_/c[35] ) );
  XOR \ADD_/FAINST[34].FA_/U4  ( .A(\ADD_/FAINST[34].FA_/n1 ), .B(b[34]), .Z(
        c[34]) );
  AND \ADD_/FAINST[34].FA_/U3  ( .A(\ADD_/FAINST[34].FA_/n1 ), .B(
        \ADD_/FAINST[34].FA_/n2 ), .Z(\ADD_/FAINST[34].FA_/n3 ) );
  XOR \ADD_/FAINST[34].FA_/U2  ( .A(b[34]), .B(\ADD_/c[34] ), .Z(
        \ADD_/FAINST[34].FA_/n2 ) );
  XOR \ADD_/FAINST[34].FA_/U1  ( .A(a[34]), .B(\ADD_/c[34] ), .Z(
        \ADD_/FAINST[34].FA_/n1 ) );
  XOR \ADD_/FAINST[33].FA_/U5  ( .A(\ADD_/FAINST[33].FA_/n3 ), .B(\ADD_/c[33] ), .Z(\ADD_/c[34] ) );
  XOR \ADD_/FAINST[33].FA_/U4  ( .A(\ADD_/FAINST[33].FA_/n1 ), .B(b[33]), .Z(
        c[33]) );
  AND \ADD_/FAINST[33].FA_/U3  ( .A(\ADD_/FAINST[33].FA_/n1 ), .B(
        \ADD_/FAINST[33].FA_/n2 ), .Z(\ADD_/FAINST[33].FA_/n3 ) );
  XOR \ADD_/FAINST[33].FA_/U2  ( .A(b[33]), .B(\ADD_/c[33] ), .Z(
        \ADD_/FAINST[33].FA_/n2 ) );
  XOR \ADD_/FAINST[33].FA_/U1  ( .A(a[33]), .B(\ADD_/c[33] ), .Z(
        \ADD_/FAINST[33].FA_/n1 ) );
  XOR \ADD_/FAINST[32].FA_/U5  ( .A(\ADD_/FAINST[32].FA_/n3 ), .B(\ADD_/c[32] ), .Z(\ADD_/c[33] ) );
  XOR \ADD_/FAINST[32].FA_/U4  ( .A(\ADD_/FAINST[32].FA_/n1 ), .B(b[32]), .Z(
        c[32]) );
  AND \ADD_/FAINST[32].FA_/U3  ( .A(\ADD_/FAINST[32].FA_/n1 ), .B(
        \ADD_/FAINST[32].FA_/n2 ), .Z(\ADD_/FAINST[32].FA_/n3 ) );
  XOR \ADD_/FAINST[32].FA_/U2  ( .A(b[32]), .B(\ADD_/c[32] ), .Z(
        \ADD_/FAINST[32].FA_/n2 ) );
  XOR \ADD_/FAINST[32].FA_/U1  ( .A(a[32]), .B(\ADD_/c[32] ), .Z(
        \ADD_/FAINST[32].FA_/n1 ) );
  XOR \ADD_/FAINST[31].FA_/U5  ( .A(\ADD_/FAINST[31].FA_/n3 ), .B(\ADD_/c[31] ), .Z(\ADD_/c[32] ) );
  XOR \ADD_/FAINST[31].FA_/U4  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(b[31]), .Z(
        c[31]) );
  AND \ADD_/FAINST[31].FA_/U3  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(
        \ADD_/FAINST[31].FA_/n2 ), .Z(\ADD_/FAINST[31].FA_/n3 ) );
  XOR \ADD_/FAINST[31].FA_/U2  ( .A(b[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n2 ) );
  XOR \ADD_/FAINST[31].FA_/U1  ( .A(a[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n1 ) );
  XOR \ADD_/FAINST[30].FA_/U5  ( .A(\ADD_/FAINST[30].FA_/n3 ), .B(\ADD_/c[30] ), .Z(\ADD_/c[31] ) );
  XOR \ADD_/FAINST[30].FA_/U4  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(b[30]), .Z(
        c[30]) );
  AND \ADD_/FAINST[30].FA_/U3  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(
        \ADD_/FAINST[30].FA_/n2 ), .Z(\ADD_/FAINST[30].FA_/n3 ) );
  XOR \ADD_/FAINST[30].FA_/U2  ( .A(b[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n2 ) );
  XOR \ADD_/FAINST[30].FA_/U1  ( .A(a[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n1 ) );
  XOR \ADD_/FAINST[29].FA_/U5  ( .A(\ADD_/FAINST[29].FA_/n3 ), .B(\ADD_/c[29] ), .Z(\ADD_/c[30] ) );
  XOR \ADD_/FAINST[29].FA_/U4  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(b[29]), .Z(
        c[29]) );
  AND \ADD_/FAINST[29].FA_/U3  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(
        \ADD_/FAINST[29].FA_/n2 ), .Z(\ADD_/FAINST[29].FA_/n3 ) );
  XOR \ADD_/FAINST[29].FA_/U2  ( .A(b[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n2 ) );
  XOR \ADD_/FAINST[29].FA_/U1  ( .A(a[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n1 ) );
  XOR \ADD_/FAINST[28].FA_/U5  ( .A(\ADD_/FAINST[28].FA_/n3 ), .B(\ADD_/c[28] ), .Z(\ADD_/c[29] ) );
  XOR \ADD_/FAINST[28].FA_/U4  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(b[28]), .Z(
        c[28]) );
  AND \ADD_/FAINST[28].FA_/U3  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(
        \ADD_/FAINST[28].FA_/n2 ), .Z(\ADD_/FAINST[28].FA_/n3 ) );
  XOR \ADD_/FAINST[28].FA_/U2  ( .A(b[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n2 ) );
  XOR \ADD_/FAINST[28].FA_/U1  ( .A(a[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n1 ) );
  XOR \ADD_/FAINST[27].FA_/U5  ( .A(\ADD_/FAINST[27].FA_/n3 ), .B(\ADD_/c[27] ), .Z(\ADD_/c[28] ) );
  XOR \ADD_/FAINST[27].FA_/U4  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(b[27]), .Z(
        c[27]) );
  AND \ADD_/FAINST[27].FA_/U3  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(
        \ADD_/FAINST[27].FA_/n2 ), .Z(\ADD_/FAINST[27].FA_/n3 ) );
  XOR \ADD_/FAINST[27].FA_/U2  ( .A(b[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n2 ) );
  XOR \ADD_/FAINST[27].FA_/U1  ( .A(a[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n1 ) );
  XOR \ADD_/FAINST[26].FA_/U5  ( .A(\ADD_/FAINST[26].FA_/n3 ), .B(\ADD_/c[26] ), .Z(\ADD_/c[27] ) );
  XOR \ADD_/FAINST[26].FA_/U4  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(b[26]), .Z(
        c[26]) );
  AND \ADD_/FAINST[26].FA_/U3  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(
        \ADD_/FAINST[26].FA_/n2 ), .Z(\ADD_/FAINST[26].FA_/n3 ) );
  XOR \ADD_/FAINST[26].FA_/U2  ( .A(b[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n2 ) );
  XOR \ADD_/FAINST[26].FA_/U1  ( .A(a[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n1 ) );
  XOR \ADD_/FAINST[25].FA_/U5  ( .A(\ADD_/FAINST[25].FA_/n3 ), .B(\ADD_/c[25] ), .Z(\ADD_/c[26] ) );
  XOR \ADD_/FAINST[25].FA_/U4  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(b[25]), .Z(
        c[25]) );
  AND \ADD_/FAINST[25].FA_/U3  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(
        \ADD_/FAINST[25].FA_/n2 ), .Z(\ADD_/FAINST[25].FA_/n3 ) );
  XOR \ADD_/FAINST[25].FA_/U2  ( .A(b[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n2 ) );
  XOR \ADD_/FAINST[25].FA_/U1  ( .A(a[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n1 ) );
  XOR \ADD_/FAINST[24].FA_/U5  ( .A(\ADD_/FAINST[24].FA_/n3 ), .B(\ADD_/c[24] ), .Z(\ADD_/c[25] ) );
  XOR \ADD_/FAINST[24].FA_/U4  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(b[24]), .Z(
        c[24]) );
  AND \ADD_/FAINST[24].FA_/U3  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(
        \ADD_/FAINST[24].FA_/n2 ), .Z(\ADD_/FAINST[24].FA_/n3 ) );
  XOR \ADD_/FAINST[24].FA_/U2  ( .A(b[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n2 ) );
  XOR \ADD_/FAINST[24].FA_/U1  ( .A(a[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n1 ) );
  XOR \ADD_/FAINST[23].FA_/U5  ( .A(\ADD_/FAINST[23].FA_/n3 ), .B(\ADD_/c[23] ), .Z(\ADD_/c[24] ) );
  XOR \ADD_/FAINST[23].FA_/U4  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(b[23]), .Z(
        c[23]) );
  AND \ADD_/FAINST[23].FA_/U3  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(
        \ADD_/FAINST[23].FA_/n2 ), .Z(\ADD_/FAINST[23].FA_/n3 ) );
  XOR \ADD_/FAINST[23].FA_/U2  ( .A(b[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n2 ) );
  XOR \ADD_/FAINST[23].FA_/U1  ( .A(a[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n1 ) );
  XOR \ADD_/FAINST[22].FA_/U5  ( .A(\ADD_/FAINST[22].FA_/n3 ), .B(\ADD_/c[22] ), .Z(\ADD_/c[23] ) );
  XOR \ADD_/FAINST[22].FA_/U4  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(b[22]), .Z(
        c[22]) );
  AND \ADD_/FAINST[22].FA_/U3  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(
        \ADD_/FAINST[22].FA_/n2 ), .Z(\ADD_/FAINST[22].FA_/n3 ) );
  XOR \ADD_/FAINST[22].FA_/U2  ( .A(b[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n2 ) );
  XOR \ADD_/FAINST[22].FA_/U1  ( .A(a[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n1 ) );
  XOR \ADD_/FAINST[21].FA_/U5  ( .A(\ADD_/FAINST[21].FA_/n3 ), .B(\ADD_/c[21] ), .Z(\ADD_/c[22] ) );
  XOR \ADD_/FAINST[21].FA_/U4  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(b[21]), .Z(
        c[21]) );
  AND \ADD_/FAINST[21].FA_/U3  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(
        \ADD_/FAINST[21].FA_/n2 ), .Z(\ADD_/FAINST[21].FA_/n3 ) );
  XOR \ADD_/FAINST[21].FA_/U2  ( .A(b[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n2 ) );
  XOR \ADD_/FAINST[21].FA_/U1  ( .A(a[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n1 ) );
  XOR \ADD_/FAINST[20].FA_/U5  ( .A(\ADD_/FAINST[20].FA_/n3 ), .B(\ADD_/c[20] ), .Z(\ADD_/c[21] ) );
  XOR \ADD_/FAINST[20].FA_/U4  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(b[20]), .Z(
        c[20]) );
  AND \ADD_/FAINST[20].FA_/U3  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(
        \ADD_/FAINST[20].FA_/n2 ), .Z(\ADD_/FAINST[20].FA_/n3 ) );
  XOR \ADD_/FAINST[20].FA_/U2  ( .A(b[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n2 ) );
  XOR \ADD_/FAINST[20].FA_/U1  ( .A(a[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n1 ) );
  XOR \ADD_/FAINST[19].FA_/U5  ( .A(\ADD_/FAINST[19].FA_/n3 ), .B(\ADD_/c[19] ), .Z(\ADD_/c[20] ) );
  XOR \ADD_/FAINST[19].FA_/U4  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(b[19]), .Z(
        c[19]) );
  AND \ADD_/FAINST[19].FA_/U3  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(
        \ADD_/FAINST[19].FA_/n2 ), .Z(\ADD_/FAINST[19].FA_/n3 ) );
  XOR \ADD_/FAINST[19].FA_/U2  ( .A(b[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n2 ) );
  XOR \ADD_/FAINST[19].FA_/U1  ( .A(a[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n1 ) );
  XOR \ADD_/FAINST[18].FA_/U5  ( .A(\ADD_/FAINST[18].FA_/n3 ), .B(\ADD_/c[18] ), .Z(\ADD_/c[19] ) );
  XOR \ADD_/FAINST[18].FA_/U4  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(b[18]), .Z(
        c[18]) );
  AND \ADD_/FAINST[18].FA_/U3  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(
        \ADD_/FAINST[18].FA_/n2 ), .Z(\ADD_/FAINST[18].FA_/n3 ) );
  XOR \ADD_/FAINST[18].FA_/U2  ( .A(b[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n2 ) );
  XOR \ADD_/FAINST[18].FA_/U1  ( .A(a[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n1 ) );
  XOR \ADD_/FAINST[17].FA_/U5  ( .A(\ADD_/FAINST[17].FA_/n3 ), .B(\ADD_/c[17] ), .Z(\ADD_/c[18] ) );
  XOR \ADD_/FAINST[17].FA_/U4  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(b[17]), .Z(
        c[17]) );
  AND \ADD_/FAINST[17].FA_/U3  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(
        \ADD_/FAINST[17].FA_/n2 ), .Z(\ADD_/FAINST[17].FA_/n3 ) );
  XOR \ADD_/FAINST[17].FA_/U2  ( .A(b[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n2 ) );
  XOR \ADD_/FAINST[17].FA_/U1  ( .A(a[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n1 ) );
  XOR \ADD_/FAINST[16].FA_/U5  ( .A(\ADD_/FAINST[16].FA_/n3 ), .B(\ADD_/c[16] ), .Z(\ADD_/c[17] ) );
  XOR \ADD_/FAINST[16].FA_/U4  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(b[16]), .Z(
        c[16]) );
  AND \ADD_/FAINST[16].FA_/U3  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(
        \ADD_/FAINST[16].FA_/n2 ), .Z(\ADD_/FAINST[16].FA_/n3 ) );
  XOR \ADD_/FAINST[16].FA_/U2  ( .A(b[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n2 ) );
  XOR \ADD_/FAINST[16].FA_/U1  ( .A(a[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n1 ) );
  XOR \ADD_/FAINST[15].FA_/U5  ( .A(\ADD_/FAINST[15].FA_/n3 ), .B(\ADD_/c[15] ), .Z(\ADD_/c[16] ) );
  XOR \ADD_/FAINST[15].FA_/U4  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(b[15]), .Z(
        c[15]) );
  AND \ADD_/FAINST[15].FA_/U3  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(
        \ADD_/FAINST[15].FA_/n2 ), .Z(\ADD_/FAINST[15].FA_/n3 ) );
  XOR \ADD_/FAINST[15].FA_/U2  ( .A(b[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n2 ) );
  XOR \ADD_/FAINST[15].FA_/U1  ( .A(a[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n1 ) );
  XOR \ADD_/FAINST[14].FA_/U5  ( .A(\ADD_/FAINST[14].FA_/n3 ), .B(\ADD_/c[14] ), .Z(\ADD_/c[15] ) );
  XOR \ADD_/FAINST[14].FA_/U4  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(b[14]), .Z(
        c[14]) );
  AND \ADD_/FAINST[14].FA_/U3  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(
        \ADD_/FAINST[14].FA_/n2 ), .Z(\ADD_/FAINST[14].FA_/n3 ) );
  XOR \ADD_/FAINST[14].FA_/U2  ( .A(b[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n2 ) );
  XOR \ADD_/FAINST[14].FA_/U1  ( .A(a[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n1 ) );
  XOR \ADD_/FAINST[13].FA_/U5  ( .A(\ADD_/FAINST[13].FA_/n3 ), .B(\ADD_/c[13] ), .Z(\ADD_/c[14] ) );
  XOR \ADD_/FAINST[13].FA_/U4  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(b[13]), .Z(
        c[13]) );
  AND \ADD_/FAINST[13].FA_/U3  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(
        \ADD_/FAINST[13].FA_/n2 ), .Z(\ADD_/FAINST[13].FA_/n3 ) );
  XOR \ADD_/FAINST[13].FA_/U2  ( .A(b[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n2 ) );
  XOR \ADD_/FAINST[13].FA_/U1  ( .A(a[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n1 ) );
  XOR \ADD_/FAINST[12].FA_/U5  ( .A(\ADD_/FAINST[12].FA_/n3 ), .B(\ADD_/c[12] ), .Z(\ADD_/c[13] ) );
  XOR \ADD_/FAINST[12].FA_/U4  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(b[12]), .Z(
        c[12]) );
  AND \ADD_/FAINST[12].FA_/U3  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(
        \ADD_/FAINST[12].FA_/n2 ), .Z(\ADD_/FAINST[12].FA_/n3 ) );
  XOR \ADD_/FAINST[12].FA_/U2  ( .A(b[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n2 ) );
  XOR \ADD_/FAINST[12].FA_/U1  ( .A(a[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n1 ) );
  XOR \ADD_/FAINST[11].FA_/U5  ( .A(\ADD_/FAINST[11].FA_/n3 ), .B(\ADD_/c[11] ), .Z(\ADD_/c[12] ) );
  XOR \ADD_/FAINST[11].FA_/U4  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(b[11]), .Z(
        c[11]) );
  AND \ADD_/FAINST[11].FA_/U3  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(
        \ADD_/FAINST[11].FA_/n2 ), .Z(\ADD_/FAINST[11].FA_/n3 ) );
  XOR \ADD_/FAINST[11].FA_/U2  ( .A(b[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n2 ) );
  XOR \ADD_/FAINST[11].FA_/U1  ( .A(a[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n1 ) );
  XOR \ADD_/FAINST[10].FA_/U5  ( .A(\ADD_/FAINST[10].FA_/n3 ), .B(\ADD_/c[10] ), .Z(\ADD_/c[11] ) );
  XOR \ADD_/FAINST[10].FA_/U4  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(b[10]), .Z(
        c[10]) );
  AND \ADD_/FAINST[10].FA_/U3  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(
        \ADD_/FAINST[10].FA_/n2 ), .Z(\ADD_/FAINST[10].FA_/n3 ) );
  XOR \ADD_/FAINST[10].FA_/U2  ( .A(b[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n2 ) );
  XOR \ADD_/FAINST[10].FA_/U1  ( .A(a[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n1 ) );
  XOR \ADD_/FAINST[9].FA_/U5  ( .A(\ADD_/FAINST[9].FA_/n3 ), .B(\ADD_/c[9] ), 
        .Z(\ADD_/c[10] ) );
  XOR \ADD_/FAINST[9].FA_/U4  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(b[9]), .Z(c[9]) );
  AND \ADD_/FAINST[9].FA_/U3  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(
        \ADD_/FAINST[9].FA_/n2 ), .Z(\ADD_/FAINST[9].FA_/n3 ) );
  XOR \ADD_/FAINST[9].FA_/U2  ( .A(b[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n2 ) );
  XOR \ADD_/FAINST[9].FA_/U1  ( .A(a[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n1 ) );
  XOR \ADD_/FAINST[8].FA_/U5  ( .A(\ADD_/FAINST[8].FA_/n3 ), .B(\ADD_/c[8] ), 
        .Z(\ADD_/c[9] ) );
  XOR \ADD_/FAINST[8].FA_/U4  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(b[8]), .Z(c[8]) );
  AND \ADD_/FAINST[8].FA_/U3  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(
        \ADD_/FAINST[8].FA_/n2 ), .Z(\ADD_/FAINST[8].FA_/n3 ) );
  XOR \ADD_/FAINST[8].FA_/U2  ( .A(b[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n2 ) );
  XOR \ADD_/FAINST[8].FA_/U1  ( .A(a[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n1 ) );
  XOR \ADD_/FAINST[7].FA_/U5  ( .A(\ADD_/FAINST[7].FA_/n3 ), .B(\ADD_/c[7] ), 
        .Z(\ADD_/c[8] ) );
  XOR \ADD_/FAINST[7].FA_/U4  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(b[7]), .Z(c[7]) );
  AND \ADD_/FAINST[7].FA_/U3  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(
        \ADD_/FAINST[7].FA_/n2 ), .Z(\ADD_/FAINST[7].FA_/n3 ) );
  XOR \ADD_/FAINST[7].FA_/U2  ( .A(b[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n2 ) );
  XOR \ADD_/FAINST[7].FA_/U1  ( .A(a[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n1 ) );
  XOR \ADD_/FAINST[6].FA_/U5  ( .A(\ADD_/FAINST[6].FA_/n3 ), .B(\ADD_/c[6] ), 
        .Z(\ADD_/c[7] ) );
  XOR \ADD_/FAINST[6].FA_/U4  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(b[6]), .Z(c[6]) );
  AND \ADD_/FAINST[6].FA_/U3  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(
        \ADD_/FAINST[6].FA_/n2 ), .Z(\ADD_/FAINST[6].FA_/n3 ) );
  XOR \ADD_/FAINST[6].FA_/U2  ( .A(b[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n2 ) );
  XOR \ADD_/FAINST[6].FA_/U1  ( .A(a[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n1 ) );
  XOR \ADD_/FAINST[5].FA_/U5  ( .A(\ADD_/FAINST[5].FA_/n3 ), .B(\ADD_/c[5] ), 
        .Z(\ADD_/c[6] ) );
  XOR \ADD_/FAINST[5].FA_/U4  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(b[5]), .Z(c[5]) );
  AND \ADD_/FAINST[5].FA_/U3  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(
        \ADD_/FAINST[5].FA_/n2 ), .Z(\ADD_/FAINST[5].FA_/n3 ) );
  XOR \ADD_/FAINST[5].FA_/U2  ( .A(b[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n2 ) );
  XOR \ADD_/FAINST[5].FA_/U1  ( .A(a[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n1 ) );
  XOR \ADD_/FAINST[4].FA_/U5  ( .A(\ADD_/FAINST[4].FA_/n3 ), .B(\ADD_/c[4] ), 
        .Z(\ADD_/c[5] ) );
  XOR \ADD_/FAINST[4].FA_/U4  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(b[4]), .Z(c[4]) );
  AND \ADD_/FAINST[4].FA_/U3  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(
        \ADD_/FAINST[4].FA_/n2 ), .Z(\ADD_/FAINST[4].FA_/n3 ) );
  XOR \ADD_/FAINST[4].FA_/U2  ( .A(b[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n2 ) );
  XOR \ADD_/FAINST[4].FA_/U1  ( .A(a[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n1 ) );
  XOR \ADD_/FAINST[3].FA_/U5  ( .A(\ADD_/FAINST[3].FA_/n3 ), .B(\ADD_/c[3] ), 
        .Z(\ADD_/c[4] ) );
  XOR \ADD_/FAINST[3].FA_/U4  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(b[3]), .Z(c[3]) );
  AND \ADD_/FAINST[3].FA_/U3  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(
        \ADD_/FAINST[3].FA_/n2 ), .Z(\ADD_/FAINST[3].FA_/n3 ) );
  XOR \ADD_/FAINST[3].FA_/U2  ( .A(b[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n2 ) );
  XOR \ADD_/FAINST[3].FA_/U1  ( .A(a[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n1 ) );
  XOR \ADD_/FAINST[2].FA_/U5  ( .A(\ADD_/FAINST[2].FA_/n3 ), .B(\ADD_/c[2] ), 
        .Z(\ADD_/c[3] ) );
  XOR \ADD_/FAINST[2].FA_/U4  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(b[2]), .Z(c[2]) );
  AND \ADD_/FAINST[2].FA_/U3  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(
        \ADD_/FAINST[2].FA_/n2 ), .Z(\ADD_/FAINST[2].FA_/n3 ) );
  XOR \ADD_/FAINST[2].FA_/U2  ( .A(b[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n2 ) );
  XOR \ADD_/FAINST[2].FA_/U1  ( .A(a[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n1 ) );
  XOR \ADD_/FAINST[1].FA_/U5  ( .A(\ADD_/FAINST[1].FA_/n3 ), .B(\ADD_/c[1] ), 
        .Z(\ADD_/c[2] ) );
  XOR \ADD_/FAINST[1].FA_/U4  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(b[1]), .Z(c[1]) );
  AND \ADD_/FAINST[1].FA_/U3  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(
        \ADD_/FAINST[1].FA_/n2 ), .Z(\ADD_/FAINST[1].FA_/n3 ) );
  XOR \ADD_/FAINST[1].FA_/U2  ( .A(b[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n2 ) );
  XOR \ADD_/FAINST[1].FA_/U1  ( .A(a[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n1 ) );
endmodule

