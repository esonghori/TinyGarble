
module first_nns_comb_W31_N128 ( q, DB, min_val_out );
  input [30:0] q;
  input [3967:0] DB;
  output [30:0] min_val_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950;

  XOR U3969 ( .A(DB[3946]), .B(n1), .Z(min_val_out[9]) );
  AND U3970 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3971 ( .A(n4), .B(n5), .Z(n3) );
  XOR U3972 ( .A(n6), .B(n7), .Z(n5) );
  IV U3973 ( .A(DB[3946]), .Z(n6) );
  AND U3974 ( .A(n8), .B(n9), .Z(n4) );
  XOR U3975 ( .A(n10), .B(n11), .Z(n9) );
  XOR U3976 ( .A(DB[3915]), .B(DB[3884]), .Z(n11) );
  AND U3977 ( .A(n12), .B(n13), .Z(n10) );
  XOR U3978 ( .A(n14), .B(n15), .Z(n13) );
  XOR U3979 ( .A(DB[3884]), .B(DB[3853]), .Z(n15) );
  AND U3980 ( .A(n16), .B(n17), .Z(n14) );
  XOR U3981 ( .A(n18), .B(n19), .Z(n17) );
  XOR U3982 ( .A(DB[3853]), .B(DB[3822]), .Z(n19) );
  AND U3983 ( .A(n20), .B(n21), .Z(n18) );
  XOR U3984 ( .A(n22), .B(n23), .Z(n21) );
  XOR U3985 ( .A(DB[3822]), .B(DB[3791]), .Z(n23) );
  AND U3986 ( .A(n24), .B(n25), .Z(n22) );
  XOR U3987 ( .A(n26), .B(n27), .Z(n25) );
  XOR U3988 ( .A(DB[3791]), .B(DB[3760]), .Z(n27) );
  AND U3989 ( .A(n28), .B(n29), .Z(n26) );
  XOR U3990 ( .A(n30), .B(n31), .Z(n29) );
  XOR U3991 ( .A(DB[3760]), .B(DB[3729]), .Z(n31) );
  AND U3992 ( .A(n32), .B(n33), .Z(n30) );
  XOR U3993 ( .A(n34), .B(n35), .Z(n33) );
  XOR U3994 ( .A(DB[3729]), .B(DB[3698]), .Z(n35) );
  AND U3995 ( .A(n36), .B(n37), .Z(n34) );
  XOR U3996 ( .A(n38), .B(n39), .Z(n37) );
  XOR U3997 ( .A(DB[3698]), .B(DB[3667]), .Z(n39) );
  AND U3998 ( .A(n40), .B(n41), .Z(n38) );
  XOR U3999 ( .A(n42), .B(n43), .Z(n41) );
  XOR U4000 ( .A(DB[3667]), .B(DB[3636]), .Z(n43) );
  AND U4001 ( .A(n44), .B(n45), .Z(n42) );
  XOR U4002 ( .A(n46), .B(n47), .Z(n45) );
  XOR U4003 ( .A(DB[3636]), .B(DB[3605]), .Z(n47) );
  AND U4004 ( .A(n48), .B(n49), .Z(n46) );
  XOR U4005 ( .A(n50), .B(n51), .Z(n49) );
  XOR U4006 ( .A(DB[3605]), .B(DB[3574]), .Z(n51) );
  AND U4007 ( .A(n52), .B(n53), .Z(n50) );
  XOR U4008 ( .A(n54), .B(n55), .Z(n53) );
  XOR U4009 ( .A(DB[3574]), .B(DB[3543]), .Z(n55) );
  AND U4010 ( .A(n56), .B(n57), .Z(n54) );
  XOR U4011 ( .A(n58), .B(n59), .Z(n57) );
  XOR U4012 ( .A(DB[3543]), .B(DB[3512]), .Z(n59) );
  AND U4013 ( .A(n60), .B(n61), .Z(n58) );
  XOR U4014 ( .A(n62), .B(n63), .Z(n61) );
  XOR U4015 ( .A(DB[3512]), .B(DB[3481]), .Z(n63) );
  AND U4016 ( .A(n64), .B(n65), .Z(n62) );
  XOR U4017 ( .A(n66), .B(n67), .Z(n65) );
  XOR U4018 ( .A(DB[3481]), .B(DB[3450]), .Z(n67) );
  AND U4019 ( .A(n68), .B(n69), .Z(n66) );
  XOR U4020 ( .A(n70), .B(n71), .Z(n69) );
  XOR U4021 ( .A(DB[3450]), .B(DB[3419]), .Z(n71) );
  AND U4022 ( .A(n72), .B(n73), .Z(n70) );
  XOR U4023 ( .A(n74), .B(n75), .Z(n73) );
  XOR U4024 ( .A(DB[3419]), .B(DB[3388]), .Z(n75) );
  AND U4025 ( .A(n76), .B(n77), .Z(n74) );
  XOR U4026 ( .A(n78), .B(n79), .Z(n77) );
  XOR U4027 ( .A(DB[3388]), .B(DB[3357]), .Z(n79) );
  AND U4028 ( .A(n80), .B(n81), .Z(n78) );
  XOR U4029 ( .A(n82), .B(n83), .Z(n81) );
  XOR U4030 ( .A(DB[3357]), .B(DB[3326]), .Z(n83) );
  AND U4031 ( .A(n84), .B(n85), .Z(n82) );
  XOR U4032 ( .A(n86), .B(n87), .Z(n85) );
  XOR U4033 ( .A(DB[3326]), .B(DB[3295]), .Z(n87) );
  AND U4034 ( .A(n88), .B(n89), .Z(n86) );
  XOR U4035 ( .A(n90), .B(n91), .Z(n89) );
  XOR U4036 ( .A(DB[3295]), .B(DB[3264]), .Z(n91) );
  AND U4037 ( .A(n92), .B(n93), .Z(n90) );
  XOR U4038 ( .A(n94), .B(n95), .Z(n93) );
  XOR U4039 ( .A(DB[3264]), .B(DB[3233]), .Z(n95) );
  AND U4040 ( .A(n96), .B(n97), .Z(n94) );
  XOR U4041 ( .A(n98), .B(n99), .Z(n97) );
  XOR U4042 ( .A(DB[3233]), .B(DB[3202]), .Z(n99) );
  AND U4043 ( .A(n100), .B(n101), .Z(n98) );
  XOR U4044 ( .A(n102), .B(n103), .Z(n101) );
  XOR U4045 ( .A(DB[3202]), .B(DB[3171]), .Z(n103) );
  AND U4046 ( .A(n104), .B(n105), .Z(n102) );
  XOR U4047 ( .A(n106), .B(n107), .Z(n105) );
  XOR U4048 ( .A(DB[3171]), .B(DB[3140]), .Z(n107) );
  AND U4049 ( .A(n108), .B(n109), .Z(n106) );
  XOR U4050 ( .A(n110), .B(n111), .Z(n109) );
  XOR U4051 ( .A(DB[3140]), .B(DB[3109]), .Z(n111) );
  AND U4052 ( .A(n112), .B(n113), .Z(n110) );
  XOR U4053 ( .A(n114), .B(n115), .Z(n113) );
  XOR U4054 ( .A(DB[3109]), .B(DB[3078]), .Z(n115) );
  AND U4055 ( .A(n116), .B(n117), .Z(n114) );
  XOR U4056 ( .A(n118), .B(n119), .Z(n117) );
  XOR U4057 ( .A(DB[3078]), .B(DB[3047]), .Z(n119) );
  AND U4058 ( .A(n120), .B(n121), .Z(n118) );
  XOR U4059 ( .A(n122), .B(n123), .Z(n121) );
  XOR U4060 ( .A(DB[3047]), .B(DB[3016]), .Z(n123) );
  AND U4061 ( .A(n124), .B(n125), .Z(n122) );
  XOR U4062 ( .A(n126), .B(n127), .Z(n125) );
  XOR U4063 ( .A(DB[3016]), .B(DB[2985]), .Z(n127) );
  AND U4064 ( .A(n128), .B(n129), .Z(n126) );
  XOR U4065 ( .A(n130), .B(n131), .Z(n129) );
  XOR U4066 ( .A(DB[2985]), .B(DB[2954]), .Z(n131) );
  AND U4067 ( .A(n132), .B(n133), .Z(n130) );
  XOR U4068 ( .A(n134), .B(n135), .Z(n133) );
  XOR U4069 ( .A(DB[2954]), .B(DB[2923]), .Z(n135) );
  AND U4070 ( .A(n136), .B(n137), .Z(n134) );
  XOR U4071 ( .A(n138), .B(n139), .Z(n137) );
  XOR U4072 ( .A(DB[2923]), .B(DB[2892]), .Z(n139) );
  AND U4073 ( .A(n140), .B(n141), .Z(n138) );
  XOR U4074 ( .A(n142), .B(n143), .Z(n141) );
  XOR U4075 ( .A(DB[2892]), .B(DB[2861]), .Z(n143) );
  AND U4076 ( .A(n144), .B(n145), .Z(n142) );
  XOR U4077 ( .A(n146), .B(n147), .Z(n145) );
  XOR U4078 ( .A(DB[2861]), .B(DB[2830]), .Z(n147) );
  AND U4079 ( .A(n148), .B(n149), .Z(n146) );
  XOR U4080 ( .A(n150), .B(n151), .Z(n149) );
  XOR U4081 ( .A(DB[2830]), .B(DB[2799]), .Z(n151) );
  AND U4082 ( .A(n152), .B(n153), .Z(n150) );
  XOR U4083 ( .A(n154), .B(n155), .Z(n153) );
  XOR U4084 ( .A(DB[2799]), .B(DB[2768]), .Z(n155) );
  AND U4085 ( .A(n156), .B(n157), .Z(n154) );
  XOR U4086 ( .A(n158), .B(n159), .Z(n157) );
  XOR U4087 ( .A(DB[2768]), .B(DB[2737]), .Z(n159) );
  AND U4088 ( .A(n160), .B(n161), .Z(n158) );
  XOR U4089 ( .A(n162), .B(n163), .Z(n161) );
  XOR U4090 ( .A(DB[2737]), .B(DB[2706]), .Z(n163) );
  AND U4091 ( .A(n164), .B(n165), .Z(n162) );
  XOR U4092 ( .A(n166), .B(n167), .Z(n165) );
  XOR U4093 ( .A(DB[2706]), .B(DB[2675]), .Z(n167) );
  AND U4094 ( .A(n168), .B(n169), .Z(n166) );
  XOR U4095 ( .A(n170), .B(n171), .Z(n169) );
  XOR U4096 ( .A(DB[2675]), .B(DB[2644]), .Z(n171) );
  AND U4097 ( .A(n172), .B(n173), .Z(n170) );
  XOR U4098 ( .A(n174), .B(n175), .Z(n173) );
  XOR U4099 ( .A(DB[2644]), .B(DB[2613]), .Z(n175) );
  AND U4100 ( .A(n176), .B(n177), .Z(n174) );
  XOR U4101 ( .A(n178), .B(n179), .Z(n177) );
  XOR U4102 ( .A(DB[2613]), .B(DB[2582]), .Z(n179) );
  AND U4103 ( .A(n180), .B(n181), .Z(n178) );
  XOR U4104 ( .A(n182), .B(n183), .Z(n181) );
  XOR U4105 ( .A(DB[2582]), .B(DB[2551]), .Z(n183) );
  AND U4106 ( .A(n184), .B(n185), .Z(n182) );
  XOR U4107 ( .A(n186), .B(n187), .Z(n185) );
  XOR U4108 ( .A(DB[2551]), .B(DB[2520]), .Z(n187) );
  AND U4109 ( .A(n188), .B(n189), .Z(n186) );
  XOR U4110 ( .A(n190), .B(n191), .Z(n189) );
  XOR U4111 ( .A(DB[2520]), .B(DB[2489]), .Z(n191) );
  AND U4112 ( .A(n192), .B(n193), .Z(n190) );
  XOR U4113 ( .A(n194), .B(n195), .Z(n193) );
  XOR U4114 ( .A(DB[2489]), .B(DB[2458]), .Z(n195) );
  AND U4115 ( .A(n196), .B(n197), .Z(n194) );
  XOR U4116 ( .A(n198), .B(n199), .Z(n197) );
  XOR U4117 ( .A(DB[2458]), .B(DB[2427]), .Z(n199) );
  AND U4118 ( .A(n200), .B(n201), .Z(n198) );
  XOR U4119 ( .A(n202), .B(n203), .Z(n201) );
  XOR U4120 ( .A(DB[2427]), .B(DB[2396]), .Z(n203) );
  AND U4121 ( .A(n204), .B(n205), .Z(n202) );
  XOR U4122 ( .A(n206), .B(n207), .Z(n205) );
  XOR U4123 ( .A(DB[2396]), .B(DB[2365]), .Z(n207) );
  AND U4124 ( .A(n208), .B(n209), .Z(n206) );
  XOR U4125 ( .A(n210), .B(n211), .Z(n209) );
  XOR U4126 ( .A(DB[2365]), .B(DB[2334]), .Z(n211) );
  AND U4127 ( .A(n212), .B(n213), .Z(n210) );
  XOR U4128 ( .A(n214), .B(n215), .Z(n213) );
  XOR U4129 ( .A(DB[2334]), .B(DB[2303]), .Z(n215) );
  AND U4130 ( .A(n216), .B(n217), .Z(n214) );
  XOR U4131 ( .A(n218), .B(n219), .Z(n217) );
  XOR U4132 ( .A(DB[2303]), .B(DB[2272]), .Z(n219) );
  AND U4133 ( .A(n220), .B(n221), .Z(n218) );
  XOR U4134 ( .A(n222), .B(n223), .Z(n221) );
  XOR U4135 ( .A(DB[2272]), .B(DB[2241]), .Z(n223) );
  AND U4136 ( .A(n224), .B(n225), .Z(n222) );
  XOR U4137 ( .A(n226), .B(n227), .Z(n225) );
  XOR U4138 ( .A(DB[2241]), .B(DB[2210]), .Z(n227) );
  AND U4139 ( .A(n228), .B(n229), .Z(n226) );
  XOR U4140 ( .A(n230), .B(n231), .Z(n229) );
  XOR U4141 ( .A(DB[2210]), .B(DB[2179]), .Z(n231) );
  AND U4142 ( .A(n232), .B(n233), .Z(n230) );
  XOR U4143 ( .A(n234), .B(n235), .Z(n233) );
  XOR U4144 ( .A(DB[2179]), .B(DB[2148]), .Z(n235) );
  AND U4145 ( .A(n236), .B(n237), .Z(n234) );
  XOR U4146 ( .A(n238), .B(n239), .Z(n237) );
  XOR U4147 ( .A(DB[2148]), .B(DB[2117]), .Z(n239) );
  AND U4148 ( .A(n240), .B(n241), .Z(n238) );
  XOR U4149 ( .A(n242), .B(n243), .Z(n241) );
  XOR U4150 ( .A(DB[2117]), .B(DB[2086]), .Z(n243) );
  AND U4151 ( .A(n244), .B(n245), .Z(n242) );
  XOR U4152 ( .A(n246), .B(n247), .Z(n245) );
  XOR U4153 ( .A(DB[2086]), .B(DB[2055]), .Z(n247) );
  AND U4154 ( .A(n248), .B(n249), .Z(n246) );
  XOR U4155 ( .A(n250), .B(n251), .Z(n249) );
  XOR U4156 ( .A(DB[2055]), .B(DB[2024]), .Z(n251) );
  AND U4157 ( .A(n252), .B(n253), .Z(n250) );
  XOR U4158 ( .A(n254), .B(n255), .Z(n253) );
  XOR U4159 ( .A(DB[2024]), .B(DB[1993]), .Z(n255) );
  AND U4160 ( .A(n256), .B(n257), .Z(n254) );
  XOR U4161 ( .A(n258), .B(n259), .Z(n257) );
  XOR U4162 ( .A(DB[1993]), .B(DB[1962]), .Z(n259) );
  AND U4163 ( .A(n260), .B(n261), .Z(n258) );
  XOR U4164 ( .A(n262), .B(n263), .Z(n261) );
  XOR U4165 ( .A(DB[1962]), .B(DB[1931]), .Z(n263) );
  AND U4166 ( .A(n264), .B(n265), .Z(n262) );
  XOR U4167 ( .A(n266), .B(n267), .Z(n265) );
  XOR U4168 ( .A(DB[1931]), .B(DB[1900]), .Z(n267) );
  AND U4169 ( .A(n268), .B(n269), .Z(n266) );
  XOR U4170 ( .A(n270), .B(n271), .Z(n269) );
  XOR U4171 ( .A(DB[1900]), .B(DB[1869]), .Z(n271) );
  AND U4172 ( .A(n272), .B(n273), .Z(n270) );
  XOR U4173 ( .A(n274), .B(n275), .Z(n273) );
  XOR U4174 ( .A(DB[1869]), .B(DB[1838]), .Z(n275) );
  AND U4175 ( .A(n276), .B(n277), .Z(n274) );
  XOR U4176 ( .A(n278), .B(n279), .Z(n277) );
  XOR U4177 ( .A(DB[1838]), .B(DB[1807]), .Z(n279) );
  AND U4178 ( .A(n280), .B(n281), .Z(n278) );
  XOR U4179 ( .A(n282), .B(n283), .Z(n281) );
  XOR U4180 ( .A(DB[1807]), .B(DB[1776]), .Z(n283) );
  AND U4181 ( .A(n284), .B(n285), .Z(n282) );
  XOR U4182 ( .A(n286), .B(n287), .Z(n285) );
  XOR U4183 ( .A(DB[1776]), .B(DB[1745]), .Z(n287) );
  AND U4184 ( .A(n288), .B(n289), .Z(n286) );
  XOR U4185 ( .A(n290), .B(n291), .Z(n289) );
  XOR U4186 ( .A(DB[1745]), .B(DB[1714]), .Z(n291) );
  AND U4187 ( .A(n292), .B(n293), .Z(n290) );
  XOR U4188 ( .A(n294), .B(n295), .Z(n293) );
  XOR U4189 ( .A(DB[1714]), .B(DB[1683]), .Z(n295) );
  AND U4190 ( .A(n296), .B(n297), .Z(n294) );
  XOR U4191 ( .A(n298), .B(n299), .Z(n297) );
  XOR U4192 ( .A(DB[1683]), .B(DB[1652]), .Z(n299) );
  AND U4193 ( .A(n300), .B(n301), .Z(n298) );
  XOR U4194 ( .A(n302), .B(n303), .Z(n301) );
  XOR U4195 ( .A(DB[1652]), .B(DB[1621]), .Z(n303) );
  AND U4196 ( .A(n304), .B(n305), .Z(n302) );
  XOR U4197 ( .A(n306), .B(n307), .Z(n305) );
  XOR U4198 ( .A(DB[1621]), .B(DB[1590]), .Z(n307) );
  AND U4199 ( .A(n308), .B(n309), .Z(n306) );
  XOR U4200 ( .A(n310), .B(n311), .Z(n309) );
  XOR U4201 ( .A(DB[1590]), .B(DB[1559]), .Z(n311) );
  AND U4202 ( .A(n312), .B(n313), .Z(n310) );
  XOR U4203 ( .A(n314), .B(n315), .Z(n313) );
  XOR U4204 ( .A(DB[1559]), .B(DB[1528]), .Z(n315) );
  AND U4205 ( .A(n316), .B(n317), .Z(n314) );
  XOR U4206 ( .A(n318), .B(n319), .Z(n317) );
  XOR U4207 ( .A(DB[1528]), .B(DB[1497]), .Z(n319) );
  AND U4208 ( .A(n320), .B(n321), .Z(n318) );
  XOR U4209 ( .A(n322), .B(n323), .Z(n321) );
  XOR U4210 ( .A(DB[1497]), .B(DB[1466]), .Z(n323) );
  AND U4211 ( .A(n324), .B(n325), .Z(n322) );
  XOR U4212 ( .A(n326), .B(n327), .Z(n325) );
  XOR U4213 ( .A(DB[1466]), .B(DB[1435]), .Z(n327) );
  AND U4214 ( .A(n328), .B(n329), .Z(n326) );
  XOR U4215 ( .A(n330), .B(n331), .Z(n329) );
  XOR U4216 ( .A(DB[1435]), .B(DB[1404]), .Z(n331) );
  AND U4217 ( .A(n332), .B(n333), .Z(n330) );
  XOR U4218 ( .A(n334), .B(n335), .Z(n333) );
  XOR U4219 ( .A(DB[1404]), .B(DB[1373]), .Z(n335) );
  AND U4220 ( .A(n336), .B(n337), .Z(n334) );
  XOR U4221 ( .A(n338), .B(n339), .Z(n337) );
  XOR U4222 ( .A(DB[1373]), .B(DB[1342]), .Z(n339) );
  AND U4223 ( .A(n340), .B(n341), .Z(n338) );
  XOR U4224 ( .A(n342), .B(n343), .Z(n341) );
  XOR U4225 ( .A(DB[1342]), .B(DB[1311]), .Z(n343) );
  AND U4226 ( .A(n344), .B(n345), .Z(n342) );
  XOR U4227 ( .A(n346), .B(n347), .Z(n345) );
  XOR U4228 ( .A(DB[1311]), .B(DB[1280]), .Z(n347) );
  AND U4229 ( .A(n348), .B(n349), .Z(n346) );
  XOR U4230 ( .A(n350), .B(n351), .Z(n349) );
  XOR U4231 ( .A(DB[1280]), .B(DB[1249]), .Z(n351) );
  AND U4232 ( .A(n352), .B(n353), .Z(n350) );
  XOR U4233 ( .A(n354), .B(n355), .Z(n353) );
  XOR U4234 ( .A(DB[1249]), .B(DB[1218]), .Z(n355) );
  AND U4235 ( .A(n356), .B(n357), .Z(n354) );
  XOR U4236 ( .A(n358), .B(n359), .Z(n357) );
  XOR U4237 ( .A(DB[1218]), .B(DB[1187]), .Z(n359) );
  AND U4238 ( .A(n360), .B(n361), .Z(n358) );
  XOR U4239 ( .A(n362), .B(n363), .Z(n361) );
  XOR U4240 ( .A(DB[1187]), .B(DB[1156]), .Z(n363) );
  AND U4241 ( .A(n364), .B(n365), .Z(n362) );
  XOR U4242 ( .A(n366), .B(n367), .Z(n365) );
  XOR U4243 ( .A(DB[1156]), .B(DB[1125]), .Z(n367) );
  AND U4244 ( .A(n368), .B(n369), .Z(n366) );
  XOR U4245 ( .A(n370), .B(n371), .Z(n369) );
  XOR U4246 ( .A(DB[1125]), .B(DB[1094]), .Z(n371) );
  AND U4247 ( .A(n372), .B(n373), .Z(n370) );
  XOR U4248 ( .A(n374), .B(n375), .Z(n373) );
  XOR U4249 ( .A(DB[1094]), .B(DB[1063]), .Z(n375) );
  AND U4250 ( .A(n376), .B(n377), .Z(n374) );
  XOR U4251 ( .A(n378), .B(n379), .Z(n377) );
  XOR U4252 ( .A(DB[1063]), .B(DB[1032]), .Z(n379) );
  AND U4253 ( .A(n380), .B(n381), .Z(n378) );
  XOR U4254 ( .A(n382), .B(n383), .Z(n381) );
  XOR U4255 ( .A(DB[1032]), .B(DB[1001]), .Z(n383) );
  AND U4256 ( .A(n384), .B(n385), .Z(n382) );
  XOR U4257 ( .A(n386), .B(n387), .Z(n385) );
  XOR U4258 ( .A(DB[970]), .B(DB[1001]), .Z(n387) );
  AND U4259 ( .A(n388), .B(n389), .Z(n386) );
  XOR U4260 ( .A(n390), .B(n391), .Z(n389) );
  XOR U4261 ( .A(DB[970]), .B(DB[939]), .Z(n391) );
  AND U4262 ( .A(n392), .B(n393), .Z(n390) );
  XOR U4263 ( .A(n394), .B(n395), .Z(n393) );
  XOR U4264 ( .A(DB[939]), .B(DB[908]), .Z(n395) );
  AND U4265 ( .A(n396), .B(n397), .Z(n394) );
  XOR U4266 ( .A(n398), .B(n399), .Z(n397) );
  XOR U4267 ( .A(DB[908]), .B(DB[877]), .Z(n399) );
  AND U4268 ( .A(n400), .B(n401), .Z(n398) );
  XOR U4269 ( .A(n402), .B(n403), .Z(n401) );
  XOR U4270 ( .A(DB[877]), .B(DB[846]), .Z(n403) );
  AND U4271 ( .A(n404), .B(n405), .Z(n402) );
  XOR U4272 ( .A(n406), .B(n407), .Z(n405) );
  XOR U4273 ( .A(DB[846]), .B(DB[815]), .Z(n407) );
  AND U4274 ( .A(n408), .B(n409), .Z(n406) );
  XOR U4275 ( .A(n410), .B(n411), .Z(n409) );
  XOR U4276 ( .A(DB[815]), .B(DB[784]), .Z(n411) );
  AND U4277 ( .A(n412), .B(n413), .Z(n410) );
  XOR U4278 ( .A(n414), .B(n415), .Z(n413) );
  XOR U4279 ( .A(DB[784]), .B(DB[753]), .Z(n415) );
  AND U4280 ( .A(n416), .B(n417), .Z(n414) );
  XOR U4281 ( .A(n418), .B(n419), .Z(n417) );
  XOR U4282 ( .A(DB[753]), .B(DB[722]), .Z(n419) );
  AND U4283 ( .A(n420), .B(n421), .Z(n418) );
  XOR U4284 ( .A(n422), .B(n423), .Z(n421) );
  XOR U4285 ( .A(DB[722]), .B(DB[691]), .Z(n423) );
  AND U4286 ( .A(n424), .B(n425), .Z(n422) );
  XOR U4287 ( .A(n426), .B(n427), .Z(n425) );
  XOR U4288 ( .A(DB[691]), .B(DB[660]), .Z(n427) );
  AND U4289 ( .A(n428), .B(n429), .Z(n426) );
  XOR U4290 ( .A(n430), .B(n431), .Z(n429) );
  XOR U4291 ( .A(DB[660]), .B(DB[629]), .Z(n431) );
  AND U4292 ( .A(n432), .B(n433), .Z(n430) );
  XOR U4293 ( .A(n434), .B(n435), .Z(n433) );
  XOR U4294 ( .A(DB[629]), .B(DB[598]), .Z(n435) );
  AND U4295 ( .A(n436), .B(n437), .Z(n434) );
  XOR U4296 ( .A(n438), .B(n439), .Z(n437) );
  XOR U4297 ( .A(DB[598]), .B(DB[567]), .Z(n439) );
  AND U4298 ( .A(n440), .B(n441), .Z(n438) );
  XOR U4299 ( .A(n442), .B(n443), .Z(n441) );
  XOR U4300 ( .A(DB[567]), .B(DB[536]), .Z(n443) );
  AND U4301 ( .A(n444), .B(n445), .Z(n442) );
  XOR U4302 ( .A(n446), .B(n447), .Z(n445) );
  XOR U4303 ( .A(DB[536]), .B(DB[505]), .Z(n447) );
  AND U4304 ( .A(n448), .B(n449), .Z(n446) );
  XOR U4305 ( .A(n450), .B(n451), .Z(n449) );
  XOR U4306 ( .A(DB[505]), .B(DB[474]), .Z(n451) );
  AND U4307 ( .A(n452), .B(n453), .Z(n450) );
  XOR U4308 ( .A(n454), .B(n455), .Z(n453) );
  XOR U4309 ( .A(DB[474]), .B(DB[443]), .Z(n455) );
  AND U4310 ( .A(n456), .B(n457), .Z(n454) );
  XOR U4311 ( .A(n458), .B(n459), .Z(n457) );
  XOR U4312 ( .A(DB[443]), .B(DB[412]), .Z(n459) );
  AND U4313 ( .A(n460), .B(n461), .Z(n458) );
  XOR U4314 ( .A(n462), .B(n463), .Z(n461) );
  XOR U4315 ( .A(DB[412]), .B(DB[381]), .Z(n463) );
  AND U4316 ( .A(n464), .B(n465), .Z(n462) );
  XOR U4317 ( .A(n466), .B(n467), .Z(n465) );
  XOR U4318 ( .A(DB[381]), .B(DB[350]), .Z(n467) );
  AND U4319 ( .A(n468), .B(n469), .Z(n466) );
  XOR U4320 ( .A(n470), .B(n471), .Z(n469) );
  XOR U4321 ( .A(DB[350]), .B(DB[319]), .Z(n471) );
  AND U4322 ( .A(n472), .B(n473), .Z(n470) );
  XOR U4323 ( .A(n474), .B(n475), .Z(n473) );
  XOR U4324 ( .A(DB[319]), .B(DB[288]), .Z(n475) );
  AND U4325 ( .A(n476), .B(n477), .Z(n474) );
  XOR U4326 ( .A(n478), .B(n479), .Z(n477) );
  XOR U4327 ( .A(DB[288]), .B(DB[257]), .Z(n479) );
  AND U4328 ( .A(n480), .B(n481), .Z(n478) );
  XOR U4329 ( .A(n482), .B(n483), .Z(n481) );
  XOR U4330 ( .A(DB[257]), .B(DB[226]), .Z(n483) );
  AND U4331 ( .A(n484), .B(n485), .Z(n482) );
  XOR U4332 ( .A(n486), .B(n487), .Z(n485) );
  XOR U4333 ( .A(DB[226]), .B(DB[195]), .Z(n487) );
  AND U4334 ( .A(n488), .B(n489), .Z(n486) );
  XOR U4335 ( .A(n490), .B(n491), .Z(n489) );
  XOR U4336 ( .A(DB[195]), .B(DB[164]), .Z(n491) );
  AND U4337 ( .A(n492), .B(n493), .Z(n490) );
  XOR U4338 ( .A(n494), .B(n495), .Z(n493) );
  XOR U4339 ( .A(DB[164]), .B(DB[133]), .Z(n495) );
  AND U4340 ( .A(n496), .B(n497), .Z(n494) );
  XOR U4341 ( .A(n498), .B(n499), .Z(n497) );
  XOR U4342 ( .A(DB[133]), .B(DB[102]), .Z(n499) );
  AND U4343 ( .A(n500), .B(n501), .Z(n498) );
  XOR U4344 ( .A(n502), .B(n503), .Z(n501) );
  XOR U4345 ( .A(DB[71]), .B(DB[102]), .Z(n503) );
  AND U4346 ( .A(n504), .B(n505), .Z(n502) );
  XOR U4347 ( .A(n506), .B(n507), .Z(n505) );
  XOR U4348 ( .A(DB[71]), .B(DB[40]), .Z(n507) );
  AND U4349 ( .A(n508), .B(n509), .Z(n506) );
  XOR U4350 ( .A(DB[9]), .B(DB[40]), .Z(n509) );
  XOR U4351 ( .A(DB[3945]), .B(n510), .Z(min_val_out[8]) );
  AND U4352 ( .A(n2), .B(n511), .Z(n510) );
  XOR U4353 ( .A(n512), .B(n513), .Z(n511) );
  XOR U4354 ( .A(DB[3945]), .B(DB[3914]), .Z(n513) );
  AND U4355 ( .A(n8), .B(n514), .Z(n512) );
  XOR U4356 ( .A(n515), .B(n516), .Z(n514) );
  XOR U4357 ( .A(DB[3914]), .B(DB[3883]), .Z(n516) );
  AND U4358 ( .A(n12), .B(n517), .Z(n515) );
  XOR U4359 ( .A(n518), .B(n519), .Z(n517) );
  XOR U4360 ( .A(DB[3883]), .B(DB[3852]), .Z(n519) );
  AND U4361 ( .A(n16), .B(n520), .Z(n518) );
  XOR U4362 ( .A(n521), .B(n522), .Z(n520) );
  XOR U4363 ( .A(DB[3852]), .B(DB[3821]), .Z(n522) );
  AND U4364 ( .A(n20), .B(n523), .Z(n521) );
  XOR U4365 ( .A(n524), .B(n525), .Z(n523) );
  XOR U4366 ( .A(DB[3821]), .B(DB[3790]), .Z(n525) );
  AND U4367 ( .A(n24), .B(n526), .Z(n524) );
  XOR U4368 ( .A(n527), .B(n528), .Z(n526) );
  XOR U4369 ( .A(DB[3790]), .B(DB[3759]), .Z(n528) );
  AND U4370 ( .A(n28), .B(n529), .Z(n527) );
  XOR U4371 ( .A(n530), .B(n531), .Z(n529) );
  XOR U4372 ( .A(DB[3759]), .B(DB[3728]), .Z(n531) );
  AND U4373 ( .A(n32), .B(n532), .Z(n530) );
  XOR U4374 ( .A(n533), .B(n534), .Z(n532) );
  XOR U4375 ( .A(DB[3728]), .B(DB[3697]), .Z(n534) );
  AND U4376 ( .A(n36), .B(n535), .Z(n533) );
  XOR U4377 ( .A(n536), .B(n537), .Z(n535) );
  XOR U4378 ( .A(DB[3697]), .B(DB[3666]), .Z(n537) );
  AND U4379 ( .A(n40), .B(n538), .Z(n536) );
  XOR U4380 ( .A(n539), .B(n540), .Z(n538) );
  XOR U4381 ( .A(DB[3666]), .B(DB[3635]), .Z(n540) );
  AND U4382 ( .A(n44), .B(n541), .Z(n539) );
  XOR U4383 ( .A(n542), .B(n543), .Z(n541) );
  XOR U4384 ( .A(DB[3635]), .B(DB[3604]), .Z(n543) );
  AND U4385 ( .A(n48), .B(n544), .Z(n542) );
  XOR U4386 ( .A(n545), .B(n546), .Z(n544) );
  XOR U4387 ( .A(DB[3604]), .B(DB[3573]), .Z(n546) );
  AND U4388 ( .A(n52), .B(n547), .Z(n545) );
  XOR U4389 ( .A(n548), .B(n549), .Z(n547) );
  XOR U4390 ( .A(DB[3573]), .B(DB[3542]), .Z(n549) );
  AND U4391 ( .A(n56), .B(n550), .Z(n548) );
  XOR U4392 ( .A(n551), .B(n552), .Z(n550) );
  XOR U4393 ( .A(DB[3542]), .B(DB[3511]), .Z(n552) );
  AND U4394 ( .A(n60), .B(n553), .Z(n551) );
  XOR U4395 ( .A(n554), .B(n555), .Z(n553) );
  XOR U4396 ( .A(DB[3511]), .B(DB[3480]), .Z(n555) );
  AND U4397 ( .A(n64), .B(n556), .Z(n554) );
  XOR U4398 ( .A(n557), .B(n558), .Z(n556) );
  XOR U4399 ( .A(DB[3480]), .B(DB[3449]), .Z(n558) );
  AND U4400 ( .A(n68), .B(n559), .Z(n557) );
  XOR U4401 ( .A(n560), .B(n561), .Z(n559) );
  XOR U4402 ( .A(DB[3449]), .B(DB[3418]), .Z(n561) );
  AND U4403 ( .A(n72), .B(n562), .Z(n560) );
  XOR U4404 ( .A(n563), .B(n564), .Z(n562) );
  XOR U4405 ( .A(DB[3418]), .B(DB[3387]), .Z(n564) );
  AND U4406 ( .A(n76), .B(n565), .Z(n563) );
  XOR U4407 ( .A(n566), .B(n567), .Z(n565) );
  XOR U4408 ( .A(DB[3387]), .B(DB[3356]), .Z(n567) );
  AND U4409 ( .A(n80), .B(n568), .Z(n566) );
  XOR U4410 ( .A(n569), .B(n570), .Z(n568) );
  XOR U4411 ( .A(DB[3356]), .B(DB[3325]), .Z(n570) );
  AND U4412 ( .A(n84), .B(n571), .Z(n569) );
  XOR U4413 ( .A(n572), .B(n573), .Z(n571) );
  XOR U4414 ( .A(DB[3325]), .B(DB[3294]), .Z(n573) );
  AND U4415 ( .A(n88), .B(n574), .Z(n572) );
  XOR U4416 ( .A(n575), .B(n576), .Z(n574) );
  XOR U4417 ( .A(DB[3294]), .B(DB[3263]), .Z(n576) );
  AND U4418 ( .A(n92), .B(n577), .Z(n575) );
  XOR U4419 ( .A(n578), .B(n579), .Z(n577) );
  XOR U4420 ( .A(DB[3263]), .B(DB[3232]), .Z(n579) );
  AND U4421 ( .A(n96), .B(n580), .Z(n578) );
  XOR U4422 ( .A(n581), .B(n582), .Z(n580) );
  XOR U4423 ( .A(DB[3232]), .B(DB[3201]), .Z(n582) );
  AND U4424 ( .A(n100), .B(n583), .Z(n581) );
  XOR U4425 ( .A(n584), .B(n585), .Z(n583) );
  XOR U4426 ( .A(DB[3201]), .B(DB[3170]), .Z(n585) );
  AND U4427 ( .A(n104), .B(n586), .Z(n584) );
  XOR U4428 ( .A(n587), .B(n588), .Z(n586) );
  XOR U4429 ( .A(DB[3170]), .B(DB[3139]), .Z(n588) );
  AND U4430 ( .A(n108), .B(n589), .Z(n587) );
  XOR U4431 ( .A(n590), .B(n591), .Z(n589) );
  XOR U4432 ( .A(DB[3139]), .B(DB[3108]), .Z(n591) );
  AND U4433 ( .A(n112), .B(n592), .Z(n590) );
  XOR U4434 ( .A(n593), .B(n594), .Z(n592) );
  XOR U4435 ( .A(DB[3108]), .B(DB[3077]), .Z(n594) );
  AND U4436 ( .A(n116), .B(n595), .Z(n593) );
  XOR U4437 ( .A(n596), .B(n597), .Z(n595) );
  XOR U4438 ( .A(DB[3077]), .B(DB[3046]), .Z(n597) );
  AND U4439 ( .A(n120), .B(n598), .Z(n596) );
  XOR U4440 ( .A(n599), .B(n600), .Z(n598) );
  XOR U4441 ( .A(DB[3046]), .B(DB[3015]), .Z(n600) );
  AND U4442 ( .A(n124), .B(n601), .Z(n599) );
  XOR U4443 ( .A(n602), .B(n603), .Z(n601) );
  XOR U4444 ( .A(DB[3015]), .B(DB[2984]), .Z(n603) );
  AND U4445 ( .A(n128), .B(n604), .Z(n602) );
  XOR U4446 ( .A(n605), .B(n606), .Z(n604) );
  XOR U4447 ( .A(DB[2984]), .B(DB[2953]), .Z(n606) );
  AND U4448 ( .A(n132), .B(n607), .Z(n605) );
  XOR U4449 ( .A(n608), .B(n609), .Z(n607) );
  XOR U4450 ( .A(DB[2953]), .B(DB[2922]), .Z(n609) );
  AND U4451 ( .A(n136), .B(n610), .Z(n608) );
  XOR U4452 ( .A(n611), .B(n612), .Z(n610) );
  XOR U4453 ( .A(DB[2922]), .B(DB[2891]), .Z(n612) );
  AND U4454 ( .A(n140), .B(n613), .Z(n611) );
  XOR U4455 ( .A(n614), .B(n615), .Z(n613) );
  XOR U4456 ( .A(DB[2891]), .B(DB[2860]), .Z(n615) );
  AND U4457 ( .A(n144), .B(n616), .Z(n614) );
  XOR U4458 ( .A(n617), .B(n618), .Z(n616) );
  XOR U4459 ( .A(DB[2860]), .B(DB[2829]), .Z(n618) );
  AND U4460 ( .A(n148), .B(n619), .Z(n617) );
  XOR U4461 ( .A(n620), .B(n621), .Z(n619) );
  XOR U4462 ( .A(DB[2829]), .B(DB[2798]), .Z(n621) );
  AND U4463 ( .A(n152), .B(n622), .Z(n620) );
  XOR U4464 ( .A(n623), .B(n624), .Z(n622) );
  XOR U4465 ( .A(DB[2798]), .B(DB[2767]), .Z(n624) );
  AND U4466 ( .A(n156), .B(n625), .Z(n623) );
  XOR U4467 ( .A(n626), .B(n627), .Z(n625) );
  XOR U4468 ( .A(DB[2767]), .B(DB[2736]), .Z(n627) );
  AND U4469 ( .A(n160), .B(n628), .Z(n626) );
  XOR U4470 ( .A(n629), .B(n630), .Z(n628) );
  XOR U4471 ( .A(DB[2736]), .B(DB[2705]), .Z(n630) );
  AND U4472 ( .A(n164), .B(n631), .Z(n629) );
  XOR U4473 ( .A(n632), .B(n633), .Z(n631) );
  XOR U4474 ( .A(DB[2705]), .B(DB[2674]), .Z(n633) );
  AND U4475 ( .A(n168), .B(n634), .Z(n632) );
  XOR U4476 ( .A(n635), .B(n636), .Z(n634) );
  XOR U4477 ( .A(DB[2674]), .B(DB[2643]), .Z(n636) );
  AND U4478 ( .A(n172), .B(n637), .Z(n635) );
  XOR U4479 ( .A(n638), .B(n639), .Z(n637) );
  XOR U4480 ( .A(DB[2643]), .B(DB[2612]), .Z(n639) );
  AND U4481 ( .A(n176), .B(n640), .Z(n638) );
  XOR U4482 ( .A(n641), .B(n642), .Z(n640) );
  XOR U4483 ( .A(DB[2612]), .B(DB[2581]), .Z(n642) );
  AND U4484 ( .A(n180), .B(n643), .Z(n641) );
  XOR U4485 ( .A(n644), .B(n645), .Z(n643) );
  XOR U4486 ( .A(DB[2581]), .B(DB[2550]), .Z(n645) );
  AND U4487 ( .A(n184), .B(n646), .Z(n644) );
  XOR U4488 ( .A(n647), .B(n648), .Z(n646) );
  XOR U4489 ( .A(DB[2550]), .B(DB[2519]), .Z(n648) );
  AND U4490 ( .A(n188), .B(n649), .Z(n647) );
  XOR U4491 ( .A(n650), .B(n651), .Z(n649) );
  XOR U4492 ( .A(DB[2519]), .B(DB[2488]), .Z(n651) );
  AND U4493 ( .A(n192), .B(n652), .Z(n650) );
  XOR U4494 ( .A(n653), .B(n654), .Z(n652) );
  XOR U4495 ( .A(DB[2488]), .B(DB[2457]), .Z(n654) );
  AND U4496 ( .A(n196), .B(n655), .Z(n653) );
  XOR U4497 ( .A(n656), .B(n657), .Z(n655) );
  XOR U4498 ( .A(DB[2457]), .B(DB[2426]), .Z(n657) );
  AND U4499 ( .A(n200), .B(n658), .Z(n656) );
  XOR U4500 ( .A(n659), .B(n660), .Z(n658) );
  XOR U4501 ( .A(DB[2426]), .B(DB[2395]), .Z(n660) );
  AND U4502 ( .A(n204), .B(n661), .Z(n659) );
  XOR U4503 ( .A(n662), .B(n663), .Z(n661) );
  XOR U4504 ( .A(DB[2395]), .B(DB[2364]), .Z(n663) );
  AND U4505 ( .A(n208), .B(n664), .Z(n662) );
  XOR U4506 ( .A(n665), .B(n666), .Z(n664) );
  XOR U4507 ( .A(DB[2364]), .B(DB[2333]), .Z(n666) );
  AND U4508 ( .A(n212), .B(n667), .Z(n665) );
  XOR U4509 ( .A(n668), .B(n669), .Z(n667) );
  XOR U4510 ( .A(DB[2333]), .B(DB[2302]), .Z(n669) );
  AND U4511 ( .A(n216), .B(n670), .Z(n668) );
  XOR U4512 ( .A(n671), .B(n672), .Z(n670) );
  XOR U4513 ( .A(DB[2302]), .B(DB[2271]), .Z(n672) );
  AND U4514 ( .A(n220), .B(n673), .Z(n671) );
  XOR U4515 ( .A(n674), .B(n675), .Z(n673) );
  XOR U4516 ( .A(DB[2271]), .B(DB[2240]), .Z(n675) );
  AND U4517 ( .A(n224), .B(n676), .Z(n674) );
  XOR U4518 ( .A(n677), .B(n678), .Z(n676) );
  XOR U4519 ( .A(DB[2240]), .B(DB[2209]), .Z(n678) );
  AND U4520 ( .A(n228), .B(n679), .Z(n677) );
  XOR U4521 ( .A(n680), .B(n681), .Z(n679) );
  XOR U4522 ( .A(DB[2209]), .B(DB[2178]), .Z(n681) );
  AND U4523 ( .A(n232), .B(n682), .Z(n680) );
  XOR U4524 ( .A(n683), .B(n684), .Z(n682) );
  XOR U4525 ( .A(DB[2178]), .B(DB[2147]), .Z(n684) );
  AND U4526 ( .A(n236), .B(n685), .Z(n683) );
  XOR U4527 ( .A(n686), .B(n687), .Z(n685) );
  XOR U4528 ( .A(DB[2147]), .B(DB[2116]), .Z(n687) );
  AND U4529 ( .A(n240), .B(n688), .Z(n686) );
  XOR U4530 ( .A(n689), .B(n690), .Z(n688) );
  XOR U4531 ( .A(DB[2116]), .B(DB[2085]), .Z(n690) );
  AND U4532 ( .A(n244), .B(n691), .Z(n689) );
  XOR U4533 ( .A(n692), .B(n693), .Z(n691) );
  XOR U4534 ( .A(DB[2085]), .B(DB[2054]), .Z(n693) );
  AND U4535 ( .A(n248), .B(n694), .Z(n692) );
  XOR U4536 ( .A(n695), .B(n696), .Z(n694) );
  XOR U4537 ( .A(DB[2054]), .B(DB[2023]), .Z(n696) );
  AND U4538 ( .A(n252), .B(n697), .Z(n695) );
  XOR U4539 ( .A(n698), .B(n699), .Z(n697) );
  XOR U4540 ( .A(DB[2023]), .B(DB[1992]), .Z(n699) );
  AND U4541 ( .A(n256), .B(n700), .Z(n698) );
  XOR U4542 ( .A(n701), .B(n702), .Z(n700) );
  XOR U4543 ( .A(DB[1992]), .B(DB[1961]), .Z(n702) );
  AND U4544 ( .A(n260), .B(n703), .Z(n701) );
  XOR U4545 ( .A(n704), .B(n705), .Z(n703) );
  XOR U4546 ( .A(DB[1961]), .B(DB[1930]), .Z(n705) );
  AND U4547 ( .A(n264), .B(n706), .Z(n704) );
  XOR U4548 ( .A(n707), .B(n708), .Z(n706) );
  XOR U4549 ( .A(DB[1930]), .B(DB[1899]), .Z(n708) );
  AND U4550 ( .A(n268), .B(n709), .Z(n707) );
  XOR U4551 ( .A(n710), .B(n711), .Z(n709) );
  XOR U4552 ( .A(DB[1899]), .B(DB[1868]), .Z(n711) );
  AND U4553 ( .A(n272), .B(n712), .Z(n710) );
  XOR U4554 ( .A(n713), .B(n714), .Z(n712) );
  XOR U4555 ( .A(DB[1868]), .B(DB[1837]), .Z(n714) );
  AND U4556 ( .A(n276), .B(n715), .Z(n713) );
  XOR U4557 ( .A(n716), .B(n717), .Z(n715) );
  XOR U4558 ( .A(DB[1837]), .B(DB[1806]), .Z(n717) );
  AND U4559 ( .A(n280), .B(n718), .Z(n716) );
  XOR U4560 ( .A(n719), .B(n720), .Z(n718) );
  XOR U4561 ( .A(DB[1806]), .B(DB[1775]), .Z(n720) );
  AND U4562 ( .A(n284), .B(n721), .Z(n719) );
  XOR U4563 ( .A(n722), .B(n723), .Z(n721) );
  XOR U4564 ( .A(DB[1775]), .B(DB[1744]), .Z(n723) );
  AND U4565 ( .A(n288), .B(n724), .Z(n722) );
  XOR U4566 ( .A(n725), .B(n726), .Z(n724) );
  XOR U4567 ( .A(DB[1744]), .B(DB[1713]), .Z(n726) );
  AND U4568 ( .A(n292), .B(n727), .Z(n725) );
  XOR U4569 ( .A(n728), .B(n729), .Z(n727) );
  XOR U4570 ( .A(DB[1713]), .B(DB[1682]), .Z(n729) );
  AND U4571 ( .A(n296), .B(n730), .Z(n728) );
  XOR U4572 ( .A(n731), .B(n732), .Z(n730) );
  XOR U4573 ( .A(DB[1682]), .B(DB[1651]), .Z(n732) );
  AND U4574 ( .A(n300), .B(n733), .Z(n731) );
  XOR U4575 ( .A(n734), .B(n735), .Z(n733) );
  XOR U4576 ( .A(DB[1651]), .B(DB[1620]), .Z(n735) );
  AND U4577 ( .A(n304), .B(n736), .Z(n734) );
  XOR U4578 ( .A(n737), .B(n738), .Z(n736) );
  XOR U4579 ( .A(DB[1620]), .B(DB[1589]), .Z(n738) );
  AND U4580 ( .A(n308), .B(n739), .Z(n737) );
  XOR U4581 ( .A(n740), .B(n741), .Z(n739) );
  XOR U4582 ( .A(DB[1589]), .B(DB[1558]), .Z(n741) );
  AND U4583 ( .A(n312), .B(n742), .Z(n740) );
  XOR U4584 ( .A(n743), .B(n744), .Z(n742) );
  XOR U4585 ( .A(DB[1558]), .B(DB[1527]), .Z(n744) );
  AND U4586 ( .A(n316), .B(n745), .Z(n743) );
  XOR U4587 ( .A(n746), .B(n747), .Z(n745) );
  XOR U4588 ( .A(DB[1527]), .B(DB[1496]), .Z(n747) );
  AND U4589 ( .A(n320), .B(n748), .Z(n746) );
  XOR U4590 ( .A(n749), .B(n750), .Z(n748) );
  XOR U4591 ( .A(DB[1496]), .B(DB[1465]), .Z(n750) );
  AND U4592 ( .A(n324), .B(n751), .Z(n749) );
  XOR U4593 ( .A(n752), .B(n753), .Z(n751) );
  XOR U4594 ( .A(DB[1465]), .B(DB[1434]), .Z(n753) );
  AND U4595 ( .A(n328), .B(n754), .Z(n752) );
  XOR U4596 ( .A(n755), .B(n756), .Z(n754) );
  XOR U4597 ( .A(DB[1434]), .B(DB[1403]), .Z(n756) );
  AND U4598 ( .A(n332), .B(n757), .Z(n755) );
  XOR U4599 ( .A(n758), .B(n759), .Z(n757) );
  XOR U4600 ( .A(DB[1403]), .B(DB[1372]), .Z(n759) );
  AND U4601 ( .A(n336), .B(n760), .Z(n758) );
  XOR U4602 ( .A(n761), .B(n762), .Z(n760) );
  XOR U4603 ( .A(DB[1372]), .B(DB[1341]), .Z(n762) );
  AND U4604 ( .A(n340), .B(n763), .Z(n761) );
  XOR U4605 ( .A(n764), .B(n765), .Z(n763) );
  XOR U4606 ( .A(DB[1341]), .B(DB[1310]), .Z(n765) );
  AND U4607 ( .A(n344), .B(n766), .Z(n764) );
  XOR U4608 ( .A(n767), .B(n768), .Z(n766) );
  XOR U4609 ( .A(DB[1310]), .B(DB[1279]), .Z(n768) );
  AND U4610 ( .A(n348), .B(n769), .Z(n767) );
  XOR U4611 ( .A(n770), .B(n771), .Z(n769) );
  XOR U4612 ( .A(DB[1279]), .B(DB[1248]), .Z(n771) );
  AND U4613 ( .A(n352), .B(n772), .Z(n770) );
  XOR U4614 ( .A(n773), .B(n774), .Z(n772) );
  XOR U4615 ( .A(DB[1248]), .B(DB[1217]), .Z(n774) );
  AND U4616 ( .A(n356), .B(n775), .Z(n773) );
  XOR U4617 ( .A(n776), .B(n777), .Z(n775) );
  XOR U4618 ( .A(DB[1217]), .B(DB[1186]), .Z(n777) );
  AND U4619 ( .A(n360), .B(n778), .Z(n776) );
  XOR U4620 ( .A(n779), .B(n780), .Z(n778) );
  XOR U4621 ( .A(DB[1186]), .B(DB[1155]), .Z(n780) );
  AND U4622 ( .A(n364), .B(n781), .Z(n779) );
  XOR U4623 ( .A(n782), .B(n783), .Z(n781) );
  XOR U4624 ( .A(DB[1155]), .B(DB[1124]), .Z(n783) );
  AND U4625 ( .A(n368), .B(n784), .Z(n782) );
  XOR U4626 ( .A(n785), .B(n786), .Z(n784) );
  XOR U4627 ( .A(DB[1124]), .B(DB[1093]), .Z(n786) );
  AND U4628 ( .A(n372), .B(n787), .Z(n785) );
  XOR U4629 ( .A(n788), .B(n789), .Z(n787) );
  XOR U4630 ( .A(DB[1093]), .B(DB[1062]), .Z(n789) );
  AND U4631 ( .A(n376), .B(n790), .Z(n788) );
  XOR U4632 ( .A(n791), .B(n792), .Z(n790) );
  XOR U4633 ( .A(DB[1062]), .B(DB[1031]), .Z(n792) );
  AND U4634 ( .A(n380), .B(n793), .Z(n791) );
  XOR U4635 ( .A(n794), .B(n795), .Z(n793) );
  XOR U4636 ( .A(DB[1031]), .B(DB[1000]), .Z(n795) );
  AND U4637 ( .A(n384), .B(n796), .Z(n794) );
  XOR U4638 ( .A(n797), .B(n798), .Z(n796) );
  XOR U4639 ( .A(DB[969]), .B(DB[1000]), .Z(n798) );
  AND U4640 ( .A(n388), .B(n799), .Z(n797) );
  XOR U4641 ( .A(n800), .B(n801), .Z(n799) );
  XOR U4642 ( .A(DB[969]), .B(DB[938]), .Z(n801) );
  AND U4643 ( .A(n392), .B(n802), .Z(n800) );
  XOR U4644 ( .A(n803), .B(n804), .Z(n802) );
  XOR U4645 ( .A(DB[938]), .B(DB[907]), .Z(n804) );
  AND U4646 ( .A(n396), .B(n805), .Z(n803) );
  XOR U4647 ( .A(n806), .B(n807), .Z(n805) );
  XOR U4648 ( .A(DB[907]), .B(DB[876]), .Z(n807) );
  AND U4649 ( .A(n400), .B(n808), .Z(n806) );
  XOR U4650 ( .A(n809), .B(n810), .Z(n808) );
  XOR U4651 ( .A(DB[876]), .B(DB[845]), .Z(n810) );
  AND U4652 ( .A(n404), .B(n811), .Z(n809) );
  XOR U4653 ( .A(n812), .B(n813), .Z(n811) );
  XOR U4654 ( .A(DB[845]), .B(DB[814]), .Z(n813) );
  AND U4655 ( .A(n408), .B(n814), .Z(n812) );
  XOR U4656 ( .A(n815), .B(n816), .Z(n814) );
  XOR U4657 ( .A(DB[814]), .B(DB[783]), .Z(n816) );
  AND U4658 ( .A(n412), .B(n817), .Z(n815) );
  XOR U4659 ( .A(n818), .B(n819), .Z(n817) );
  XOR U4660 ( .A(DB[783]), .B(DB[752]), .Z(n819) );
  AND U4661 ( .A(n416), .B(n820), .Z(n818) );
  XOR U4662 ( .A(n821), .B(n822), .Z(n820) );
  XOR U4663 ( .A(DB[752]), .B(DB[721]), .Z(n822) );
  AND U4664 ( .A(n420), .B(n823), .Z(n821) );
  XOR U4665 ( .A(n824), .B(n825), .Z(n823) );
  XOR U4666 ( .A(DB[721]), .B(DB[690]), .Z(n825) );
  AND U4667 ( .A(n424), .B(n826), .Z(n824) );
  XOR U4668 ( .A(n827), .B(n828), .Z(n826) );
  XOR U4669 ( .A(DB[690]), .B(DB[659]), .Z(n828) );
  AND U4670 ( .A(n428), .B(n829), .Z(n827) );
  XOR U4671 ( .A(n830), .B(n831), .Z(n829) );
  XOR U4672 ( .A(DB[659]), .B(DB[628]), .Z(n831) );
  AND U4673 ( .A(n432), .B(n832), .Z(n830) );
  XOR U4674 ( .A(n833), .B(n834), .Z(n832) );
  XOR U4675 ( .A(DB[628]), .B(DB[597]), .Z(n834) );
  AND U4676 ( .A(n436), .B(n835), .Z(n833) );
  XOR U4677 ( .A(n836), .B(n837), .Z(n835) );
  XOR U4678 ( .A(DB[597]), .B(DB[566]), .Z(n837) );
  AND U4679 ( .A(n440), .B(n838), .Z(n836) );
  XOR U4680 ( .A(n839), .B(n840), .Z(n838) );
  XOR U4681 ( .A(DB[566]), .B(DB[535]), .Z(n840) );
  AND U4682 ( .A(n444), .B(n841), .Z(n839) );
  XOR U4683 ( .A(n842), .B(n843), .Z(n841) );
  XOR U4684 ( .A(DB[535]), .B(DB[504]), .Z(n843) );
  AND U4685 ( .A(n448), .B(n844), .Z(n842) );
  XOR U4686 ( .A(n845), .B(n846), .Z(n844) );
  XOR U4687 ( .A(DB[504]), .B(DB[473]), .Z(n846) );
  AND U4688 ( .A(n452), .B(n847), .Z(n845) );
  XOR U4689 ( .A(n848), .B(n849), .Z(n847) );
  XOR U4690 ( .A(DB[473]), .B(DB[442]), .Z(n849) );
  AND U4691 ( .A(n456), .B(n850), .Z(n848) );
  XOR U4692 ( .A(n851), .B(n852), .Z(n850) );
  XOR U4693 ( .A(DB[442]), .B(DB[411]), .Z(n852) );
  AND U4694 ( .A(n460), .B(n853), .Z(n851) );
  XOR U4695 ( .A(n854), .B(n855), .Z(n853) );
  XOR U4696 ( .A(DB[411]), .B(DB[380]), .Z(n855) );
  AND U4697 ( .A(n464), .B(n856), .Z(n854) );
  XOR U4698 ( .A(n857), .B(n858), .Z(n856) );
  XOR U4699 ( .A(DB[380]), .B(DB[349]), .Z(n858) );
  AND U4700 ( .A(n468), .B(n859), .Z(n857) );
  XOR U4701 ( .A(n860), .B(n861), .Z(n859) );
  XOR U4702 ( .A(DB[349]), .B(DB[318]), .Z(n861) );
  AND U4703 ( .A(n472), .B(n862), .Z(n860) );
  XOR U4704 ( .A(n863), .B(n864), .Z(n862) );
  XOR U4705 ( .A(DB[318]), .B(DB[287]), .Z(n864) );
  AND U4706 ( .A(n476), .B(n865), .Z(n863) );
  XOR U4707 ( .A(n866), .B(n867), .Z(n865) );
  XOR U4708 ( .A(DB[287]), .B(DB[256]), .Z(n867) );
  AND U4709 ( .A(n480), .B(n868), .Z(n866) );
  XOR U4710 ( .A(n869), .B(n870), .Z(n868) );
  XOR U4711 ( .A(DB[256]), .B(DB[225]), .Z(n870) );
  AND U4712 ( .A(n484), .B(n871), .Z(n869) );
  XOR U4713 ( .A(n872), .B(n873), .Z(n871) );
  XOR U4714 ( .A(DB[225]), .B(DB[194]), .Z(n873) );
  AND U4715 ( .A(n488), .B(n874), .Z(n872) );
  XOR U4716 ( .A(n875), .B(n876), .Z(n874) );
  XOR U4717 ( .A(DB[194]), .B(DB[163]), .Z(n876) );
  AND U4718 ( .A(n492), .B(n877), .Z(n875) );
  XOR U4719 ( .A(n878), .B(n879), .Z(n877) );
  XOR U4720 ( .A(DB[163]), .B(DB[132]), .Z(n879) );
  AND U4721 ( .A(n496), .B(n880), .Z(n878) );
  XOR U4722 ( .A(n881), .B(n882), .Z(n880) );
  XOR U4723 ( .A(DB[132]), .B(DB[101]), .Z(n882) );
  AND U4724 ( .A(n500), .B(n883), .Z(n881) );
  XOR U4725 ( .A(n884), .B(n885), .Z(n883) );
  XOR U4726 ( .A(DB[70]), .B(DB[101]), .Z(n885) );
  AND U4727 ( .A(n504), .B(n886), .Z(n884) );
  XOR U4728 ( .A(n887), .B(n888), .Z(n886) );
  XOR U4729 ( .A(DB[70]), .B(DB[39]), .Z(n888) );
  AND U4730 ( .A(n508), .B(n889), .Z(n887) );
  XOR U4731 ( .A(DB[8]), .B(DB[39]), .Z(n889) );
  XOR U4732 ( .A(DB[3944]), .B(n890), .Z(min_val_out[7]) );
  AND U4733 ( .A(n2), .B(n891), .Z(n890) );
  XOR U4734 ( .A(n892), .B(n893), .Z(n891) );
  XOR U4735 ( .A(DB[3944]), .B(DB[3913]), .Z(n893) );
  AND U4736 ( .A(n8), .B(n894), .Z(n892) );
  XOR U4737 ( .A(n895), .B(n896), .Z(n894) );
  XOR U4738 ( .A(DB[3913]), .B(DB[3882]), .Z(n896) );
  AND U4739 ( .A(n12), .B(n897), .Z(n895) );
  XOR U4740 ( .A(n898), .B(n899), .Z(n897) );
  XOR U4741 ( .A(DB[3882]), .B(DB[3851]), .Z(n899) );
  AND U4742 ( .A(n16), .B(n900), .Z(n898) );
  XOR U4743 ( .A(n901), .B(n902), .Z(n900) );
  XOR U4744 ( .A(DB[3851]), .B(DB[3820]), .Z(n902) );
  AND U4745 ( .A(n20), .B(n903), .Z(n901) );
  XOR U4746 ( .A(n904), .B(n905), .Z(n903) );
  XOR U4747 ( .A(DB[3820]), .B(DB[3789]), .Z(n905) );
  AND U4748 ( .A(n24), .B(n906), .Z(n904) );
  XOR U4749 ( .A(n907), .B(n908), .Z(n906) );
  XOR U4750 ( .A(DB[3789]), .B(DB[3758]), .Z(n908) );
  AND U4751 ( .A(n28), .B(n909), .Z(n907) );
  XOR U4752 ( .A(n910), .B(n911), .Z(n909) );
  XOR U4753 ( .A(DB[3758]), .B(DB[3727]), .Z(n911) );
  AND U4754 ( .A(n32), .B(n912), .Z(n910) );
  XOR U4755 ( .A(n913), .B(n914), .Z(n912) );
  XOR U4756 ( .A(DB[3727]), .B(DB[3696]), .Z(n914) );
  AND U4757 ( .A(n36), .B(n915), .Z(n913) );
  XOR U4758 ( .A(n916), .B(n917), .Z(n915) );
  XOR U4759 ( .A(DB[3696]), .B(DB[3665]), .Z(n917) );
  AND U4760 ( .A(n40), .B(n918), .Z(n916) );
  XOR U4761 ( .A(n919), .B(n920), .Z(n918) );
  XOR U4762 ( .A(DB[3665]), .B(DB[3634]), .Z(n920) );
  AND U4763 ( .A(n44), .B(n921), .Z(n919) );
  XOR U4764 ( .A(n922), .B(n923), .Z(n921) );
  XOR U4765 ( .A(DB[3634]), .B(DB[3603]), .Z(n923) );
  AND U4766 ( .A(n48), .B(n924), .Z(n922) );
  XOR U4767 ( .A(n925), .B(n926), .Z(n924) );
  XOR U4768 ( .A(DB[3603]), .B(DB[3572]), .Z(n926) );
  AND U4769 ( .A(n52), .B(n927), .Z(n925) );
  XOR U4770 ( .A(n928), .B(n929), .Z(n927) );
  XOR U4771 ( .A(DB[3572]), .B(DB[3541]), .Z(n929) );
  AND U4772 ( .A(n56), .B(n930), .Z(n928) );
  XOR U4773 ( .A(n931), .B(n932), .Z(n930) );
  XOR U4774 ( .A(DB[3541]), .B(DB[3510]), .Z(n932) );
  AND U4775 ( .A(n60), .B(n933), .Z(n931) );
  XOR U4776 ( .A(n934), .B(n935), .Z(n933) );
  XOR U4777 ( .A(DB[3510]), .B(DB[3479]), .Z(n935) );
  AND U4778 ( .A(n64), .B(n936), .Z(n934) );
  XOR U4779 ( .A(n937), .B(n938), .Z(n936) );
  XOR U4780 ( .A(DB[3479]), .B(DB[3448]), .Z(n938) );
  AND U4781 ( .A(n68), .B(n939), .Z(n937) );
  XOR U4782 ( .A(n940), .B(n941), .Z(n939) );
  XOR U4783 ( .A(DB[3448]), .B(DB[3417]), .Z(n941) );
  AND U4784 ( .A(n72), .B(n942), .Z(n940) );
  XOR U4785 ( .A(n943), .B(n944), .Z(n942) );
  XOR U4786 ( .A(DB[3417]), .B(DB[3386]), .Z(n944) );
  AND U4787 ( .A(n76), .B(n945), .Z(n943) );
  XOR U4788 ( .A(n946), .B(n947), .Z(n945) );
  XOR U4789 ( .A(DB[3386]), .B(DB[3355]), .Z(n947) );
  AND U4790 ( .A(n80), .B(n948), .Z(n946) );
  XOR U4791 ( .A(n949), .B(n950), .Z(n948) );
  XOR U4792 ( .A(DB[3355]), .B(DB[3324]), .Z(n950) );
  AND U4793 ( .A(n84), .B(n951), .Z(n949) );
  XOR U4794 ( .A(n952), .B(n953), .Z(n951) );
  XOR U4795 ( .A(DB[3324]), .B(DB[3293]), .Z(n953) );
  AND U4796 ( .A(n88), .B(n954), .Z(n952) );
  XOR U4797 ( .A(n955), .B(n956), .Z(n954) );
  XOR U4798 ( .A(DB[3293]), .B(DB[3262]), .Z(n956) );
  AND U4799 ( .A(n92), .B(n957), .Z(n955) );
  XOR U4800 ( .A(n958), .B(n959), .Z(n957) );
  XOR U4801 ( .A(DB[3262]), .B(DB[3231]), .Z(n959) );
  AND U4802 ( .A(n96), .B(n960), .Z(n958) );
  XOR U4803 ( .A(n961), .B(n962), .Z(n960) );
  XOR U4804 ( .A(DB[3231]), .B(DB[3200]), .Z(n962) );
  AND U4805 ( .A(n100), .B(n963), .Z(n961) );
  XOR U4806 ( .A(n964), .B(n965), .Z(n963) );
  XOR U4807 ( .A(DB[3200]), .B(DB[3169]), .Z(n965) );
  AND U4808 ( .A(n104), .B(n966), .Z(n964) );
  XOR U4809 ( .A(n967), .B(n968), .Z(n966) );
  XOR U4810 ( .A(DB[3169]), .B(DB[3138]), .Z(n968) );
  AND U4811 ( .A(n108), .B(n969), .Z(n967) );
  XOR U4812 ( .A(n970), .B(n971), .Z(n969) );
  XOR U4813 ( .A(DB[3138]), .B(DB[3107]), .Z(n971) );
  AND U4814 ( .A(n112), .B(n972), .Z(n970) );
  XOR U4815 ( .A(n973), .B(n974), .Z(n972) );
  XOR U4816 ( .A(DB[3107]), .B(DB[3076]), .Z(n974) );
  AND U4817 ( .A(n116), .B(n975), .Z(n973) );
  XOR U4818 ( .A(n976), .B(n977), .Z(n975) );
  XOR U4819 ( .A(DB[3076]), .B(DB[3045]), .Z(n977) );
  AND U4820 ( .A(n120), .B(n978), .Z(n976) );
  XOR U4821 ( .A(n979), .B(n980), .Z(n978) );
  XOR U4822 ( .A(DB[3045]), .B(DB[3014]), .Z(n980) );
  AND U4823 ( .A(n124), .B(n981), .Z(n979) );
  XOR U4824 ( .A(n982), .B(n983), .Z(n981) );
  XOR U4825 ( .A(DB[3014]), .B(DB[2983]), .Z(n983) );
  AND U4826 ( .A(n128), .B(n984), .Z(n982) );
  XOR U4827 ( .A(n985), .B(n986), .Z(n984) );
  XOR U4828 ( .A(DB[2983]), .B(DB[2952]), .Z(n986) );
  AND U4829 ( .A(n132), .B(n987), .Z(n985) );
  XOR U4830 ( .A(n988), .B(n989), .Z(n987) );
  XOR U4831 ( .A(DB[2952]), .B(DB[2921]), .Z(n989) );
  AND U4832 ( .A(n136), .B(n990), .Z(n988) );
  XOR U4833 ( .A(n991), .B(n992), .Z(n990) );
  XOR U4834 ( .A(DB[2921]), .B(DB[2890]), .Z(n992) );
  AND U4835 ( .A(n140), .B(n993), .Z(n991) );
  XOR U4836 ( .A(n994), .B(n995), .Z(n993) );
  XOR U4837 ( .A(DB[2890]), .B(DB[2859]), .Z(n995) );
  AND U4838 ( .A(n144), .B(n996), .Z(n994) );
  XOR U4839 ( .A(n997), .B(n998), .Z(n996) );
  XOR U4840 ( .A(DB[2859]), .B(DB[2828]), .Z(n998) );
  AND U4841 ( .A(n148), .B(n999), .Z(n997) );
  XOR U4842 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U4843 ( .A(DB[2828]), .B(DB[2797]), .Z(n1001) );
  AND U4844 ( .A(n152), .B(n1002), .Z(n1000) );
  XOR U4845 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR U4846 ( .A(DB[2797]), .B(DB[2766]), .Z(n1004) );
  AND U4847 ( .A(n156), .B(n1005), .Z(n1003) );
  XOR U4848 ( .A(n1006), .B(n1007), .Z(n1005) );
  XOR U4849 ( .A(DB[2766]), .B(DB[2735]), .Z(n1007) );
  AND U4850 ( .A(n160), .B(n1008), .Z(n1006) );
  XOR U4851 ( .A(n1009), .B(n1010), .Z(n1008) );
  XOR U4852 ( .A(DB[2735]), .B(DB[2704]), .Z(n1010) );
  AND U4853 ( .A(n164), .B(n1011), .Z(n1009) );
  XOR U4854 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR U4855 ( .A(DB[2704]), .B(DB[2673]), .Z(n1013) );
  AND U4856 ( .A(n168), .B(n1014), .Z(n1012) );
  XOR U4857 ( .A(n1015), .B(n1016), .Z(n1014) );
  XOR U4858 ( .A(DB[2673]), .B(DB[2642]), .Z(n1016) );
  AND U4859 ( .A(n172), .B(n1017), .Z(n1015) );
  XOR U4860 ( .A(n1018), .B(n1019), .Z(n1017) );
  XOR U4861 ( .A(DB[2642]), .B(DB[2611]), .Z(n1019) );
  AND U4862 ( .A(n176), .B(n1020), .Z(n1018) );
  XOR U4863 ( .A(n1021), .B(n1022), .Z(n1020) );
  XOR U4864 ( .A(DB[2611]), .B(DB[2580]), .Z(n1022) );
  AND U4865 ( .A(n180), .B(n1023), .Z(n1021) );
  XOR U4866 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U4867 ( .A(DB[2580]), .B(DB[2549]), .Z(n1025) );
  AND U4868 ( .A(n184), .B(n1026), .Z(n1024) );
  XOR U4869 ( .A(n1027), .B(n1028), .Z(n1026) );
  XOR U4870 ( .A(DB[2549]), .B(DB[2518]), .Z(n1028) );
  AND U4871 ( .A(n188), .B(n1029), .Z(n1027) );
  XOR U4872 ( .A(n1030), .B(n1031), .Z(n1029) );
  XOR U4873 ( .A(DB[2518]), .B(DB[2487]), .Z(n1031) );
  AND U4874 ( .A(n192), .B(n1032), .Z(n1030) );
  XOR U4875 ( .A(n1033), .B(n1034), .Z(n1032) );
  XOR U4876 ( .A(DB[2487]), .B(DB[2456]), .Z(n1034) );
  AND U4877 ( .A(n196), .B(n1035), .Z(n1033) );
  XOR U4878 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR U4879 ( .A(DB[2456]), .B(DB[2425]), .Z(n1037) );
  AND U4880 ( .A(n200), .B(n1038), .Z(n1036) );
  XOR U4881 ( .A(n1039), .B(n1040), .Z(n1038) );
  XOR U4882 ( .A(DB[2425]), .B(DB[2394]), .Z(n1040) );
  AND U4883 ( .A(n204), .B(n1041), .Z(n1039) );
  XOR U4884 ( .A(n1042), .B(n1043), .Z(n1041) );
  XOR U4885 ( .A(DB[2394]), .B(DB[2363]), .Z(n1043) );
  AND U4886 ( .A(n208), .B(n1044), .Z(n1042) );
  XOR U4887 ( .A(n1045), .B(n1046), .Z(n1044) );
  XOR U4888 ( .A(DB[2363]), .B(DB[2332]), .Z(n1046) );
  AND U4889 ( .A(n212), .B(n1047), .Z(n1045) );
  XOR U4890 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U4891 ( .A(DB[2332]), .B(DB[2301]), .Z(n1049) );
  AND U4892 ( .A(n216), .B(n1050), .Z(n1048) );
  XOR U4893 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U4894 ( .A(DB[2301]), .B(DB[2270]), .Z(n1052) );
  AND U4895 ( .A(n220), .B(n1053), .Z(n1051) );
  XOR U4896 ( .A(n1054), .B(n1055), .Z(n1053) );
  XOR U4897 ( .A(DB[2270]), .B(DB[2239]), .Z(n1055) );
  AND U4898 ( .A(n224), .B(n1056), .Z(n1054) );
  XOR U4899 ( .A(n1057), .B(n1058), .Z(n1056) );
  XOR U4900 ( .A(DB[2239]), .B(DB[2208]), .Z(n1058) );
  AND U4901 ( .A(n228), .B(n1059), .Z(n1057) );
  XOR U4902 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR U4903 ( .A(DB[2208]), .B(DB[2177]), .Z(n1061) );
  AND U4904 ( .A(n232), .B(n1062), .Z(n1060) );
  XOR U4905 ( .A(n1063), .B(n1064), .Z(n1062) );
  XOR U4906 ( .A(DB[2177]), .B(DB[2146]), .Z(n1064) );
  AND U4907 ( .A(n236), .B(n1065), .Z(n1063) );
  XOR U4908 ( .A(n1066), .B(n1067), .Z(n1065) );
  XOR U4909 ( .A(DB[2146]), .B(DB[2115]), .Z(n1067) );
  AND U4910 ( .A(n240), .B(n1068), .Z(n1066) );
  XOR U4911 ( .A(n1069), .B(n1070), .Z(n1068) );
  XOR U4912 ( .A(DB[2115]), .B(DB[2084]), .Z(n1070) );
  AND U4913 ( .A(n244), .B(n1071), .Z(n1069) );
  XOR U4914 ( .A(n1072), .B(n1073), .Z(n1071) );
  XOR U4915 ( .A(DB[2084]), .B(DB[2053]), .Z(n1073) );
  AND U4916 ( .A(n248), .B(n1074), .Z(n1072) );
  XOR U4917 ( .A(n1075), .B(n1076), .Z(n1074) );
  XOR U4918 ( .A(DB[2053]), .B(DB[2022]), .Z(n1076) );
  AND U4919 ( .A(n252), .B(n1077), .Z(n1075) );
  XOR U4920 ( .A(n1078), .B(n1079), .Z(n1077) );
  XOR U4921 ( .A(DB[2022]), .B(DB[1991]), .Z(n1079) );
  AND U4922 ( .A(n256), .B(n1080), .Z(n1078) );
  XOR U4923 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR U4924 ( .A(DB[1991]), .B(DB[1960]), .Z(n1082) );
  AND U4925 ( .A(n260), .B(n1083), .Z(n1081) );
  XOR U4926 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U4927 ( .A(DB[1960]), .B(DB[1929]), .Z(n1085) );
  AND U4928 ( .A(n264), .B(n1086), .Z(n1084) );
  XOR U4929 ( .A(n1087), .B(n1088), .Z(n1086) );
  XOR U4930 ( .A(DB[1929]), .B(DB[1898]), .Z(n1088) );
  AND U4931 ( .A(n268), .B(n1089), .Z(n1087) );
  XOR U4932 ( .A(n1090), .B(n1091), .Z(n1089) );
  XOR U4933 ( .A(DB[1898]), .B(DB[1867]), .Z(n1091) );
  AND U4934 ( .A(n272), .B(n1092), .Z(n1090) );
  XOR U4935 ( .A(n1093), .B(n1094), .Z(n1092) );
  XOR U4936 ( .A(DB[1867]), .B(DB[1836]), .Z(n1094) );
  AND U4937 ( .A(n276), .B(n1095), .Z(n1093) );
  XOR U4938 ( .A(n1096), .B(n1097), .Z(n1095) );
  XOR U4939 ( .A(DB[1836]), .B(DB[1805]), .Z(n1097) );
  AND U4940 ( .A(n280), .B(n1098), .Z(n1096) );
  XOR U4941 ( .A(n1099), .B(n1100), .Z(n1098) );
  XOR U4942 ( .A(DB[1805]), .B(DB[1774]), .Z(n1100) );
  AND U4943 ( .A(n284), .B(n1101), .Z(n1099) );
  XOR U4944 ( .A(n1102), .B(n1103), .Z(n1101) );
  XOR U4945 ( .A(DB[1774]), .B(DB[1743]), .Z(n1103) );
  AND U4946 ( .A(n288), .B(n1104), .Z(n1102) );
  XOR U4947 ( .A(n1105), .B(n1106), .Z(n1104) );
  XOR U4948 ( .A(DB[1743]), .B(DB[1712]), .Z(n1106) );
  AND U4949 ( .A(n292), .B(n1107), .Z(n1105) );
  XOR U4950 ( .A(n1108), .B(n1109), .Z(n1107) );
  XOR U4951 ( .A(DB[1712]), .B(DB[1681]), .Z(n1109) );
  AND U4952 ( .A(n296), .B(n1110), .Z(n1108) );
  XOR U4953 ( .A(n1111), .B(n1112), .Z(n1110) );
  XOR U4954 ( .A(DB[1681]), .B(DB[1650]), .Z(n1112) );
  AND U4955 ( .A(n300), .B(n1113), .Z(n1111) );
  XOR U4956 ( .A(n1114), .B(n1115), .Z(n1113) );
  XOR U4957 ( .A(DB[1650]), .B(DB[1619]), .Z(n1115) );
  AND U4958 ( .A(n304), .B(n1116), .Z(n1114) );
  XOR U4959 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U4960 ( .A(DB[1619]), .B(DB[1588]), .Z(n1118) );
  AND U4961 ( .A(n308), .B(n1119), .Z(n1117) );
  XOR U4962 ( .A(n1120), .B(n1121), .Z(n1119) );
  XOR U4963 ( .A(DB[1588]), .B(DB[1557]), .Z(n1121) );
  AND U4964 ( .A(n312), .B(n1122), .Z(n1120) );
  XOR U4965 ( .A(n1123), .B(n1124), .Z(n1122) );
  XOR U4966 ( .A(DB[1557]), .B(DB[1526]), .Z(n1124) );
  AND U4967 ( .A(n316), .B(n1125), .Z(n1123) );
  XOR U4968 ( .A(n1126), .B(n1127), .Z(n1125) );
  XOR U4969 ( .A(DB[1526]), .B(DB[1495]), .Z(n1127) );
  AND U4970 ( .A(n320), .B(n1128), .Z(n1126) );
  XOR U4971 ( .A(n1129), .B(n1130), .Z(n1128) );
  XOR U4972 ( .A(DB[1495]), .B(DB[1464]), .Z(n1130) );
  AND U4973 ( .A(n324), .B(n1131), .Z(n1129) );
  XOR U4974 ( .A(n1132), .B(n1133), .Z(n1131) );
  XOR U4975 ( .A(DB[1464]), .B(DB[1433]), .Z(n1133) );
  AND U4976 ( .A(n328), .B(n1134), .Z(n1132) );
  XOR U4977 ( .A(n1135), .B(n1136), .Z(n1134) );
  XOR U4978 ( .A(DB[1433]), .B(DB[1402]), .Z(n1136) );
  AND U4979 ( .A(n332), .B(n1137), .Z(n1135) );
  XOR U4980 ( .A(n1138), .B(n1139), .Z(n1137) );
  XOR U4981 ( .A(DB[1402]), .B(DB[1371]), .Z(n1139) );
  AND U4982 ( .A(n336), .B(n1140), .Z(n1138) );
  XOR U4983 ( .A(n1141), .B(n1142), .Z(n1140) );
  XOR U4984 ( .A(DB[1371]), .B(DB[1340]), .Z(n1142) );
  AND U4985 ( .A(n340), .B(n1143), .Z(n1141) );
  XOR U4986 ( .A(n1144), .B(n1145), .Z(n1143) );
  XOR U4987 ( .A(DB[1340]), .B(DB[1309]), .Z(n1145) );
  AND U4988 ( .A(n344), .B(n1146), .Z(n1144) );
  XOR U4989 ( .A(n1147), .B(n1148), .Z(n1146) );
  XOR U4990 ( .A(DB[1309]), .B(DB[1278]), .Z(n1148) );
  AND U4991 ( .A(n348), .B(n1149), .Z(n1147) );
  XOR U4992 ( .A(n1150), .B(n1151), .Z(n1149) );
  XOR U4993 ( .A(DB[1278]), .B(DB[1247]), .Z(n1151) );
  AND U4994 ( .A(n352), .B(n1152), .Z(n1150) );
  XOR U4995 ( .A(n1153), .B(n1154), .Z(n1152) );
  XOR U4996 ( .A(DB[1247]), .B(DB[1216]), .Z(n1154) );
  AND U4997 ( .A(n356), .B(n1155), .Z(n1153) );
  XOR U4998 ( .A(n1156), .B(n1157), .Z(n1155) );
  XOR U4999 ( .A(DB[1216]), .B(DB[1185]), .Z(n1157) );
  AND U5000 ( .A(n360), .B(n1158), .Z(n1156) );
  XOR U5001 ( .A(n1159), .B(n1160), .Z(n1158) );
  XOR U5002 ( .A(DB[1185]), .B(DB[1154]), .Z(n1160) );
  AND U5003 ( .A(n364), .B(n1161), .Z(n1159) );
  XOR U5004 ( .A(n1162), .B(n1163), .Z(n1161) );
  XOR U5005 ( .A(DB[1154]), .B(DB[1123]), .Z(n1163) );
  AND U5006 ( .A(n368), .B(n1164), .Z(n1162) );
  XOR U5007 ( .A(n1165), .B(n1166), .Z(n1164) );
  XOR U5008 ( .A(DB[1123]), .B(DB[1092]), .Z(n1166) );
  AND U5009 ( .A(n372), .B(n1167), .Z(n1165) );
  XOR U5010 ( .A(n1168), .B(n1169), .Z(n1167) );
  XOR U5011 ( .A(DB[1092]), .B(DB[1061]), .Z(n1169) );
  AND U5012 ( .A(n376), .B(n1170), .Z(n1168) );
  XOR U5013 ( .A(n1171), .B(n1172), .Z(n1170) );
  XOR U5014 ( .A(DB[1061]), .B(DB[1030]), .Z(n1172) );
  AND U5015 ( .A(n380), .B(n1173), .Z(n1171) );
  XOR U5016 ( .A(n1174), .B(n1175), .Z(n1173) );
  XOR U5017 ( .A(DB[999]), .B(DB[1030]), .Z(n1175) );
  AND U5018 ( .A(n384), .B(n1176), .Z(n1174) );
  XOR U5019 ( .A(n1177), .B(n1178), .Z(n1176) );
  XOR U5020 ( .A(DB[999]), .B(DB[968]), .Z(n1178) );
  AND U5021 ( .A(n388), .B(n1179), .Z(n1177) );
  XOR U5022 ( .A(n1180), .B(n1181), .Z(n1179) );
  XOR U5023 ( .A(DB[968]), .B(DB[937]), .Z(n1181) );
  AND U5024 ( .A(n392), .B(n1182), .Z(n1180) );
  XOR U5025 ( .A(n1183), .B(n1184), .Z(n1182) );
  XOR U5026 ( .A(DB[937]), .B(DB[906]), .Z(n1184) );
  AND U5027 ( .A(n396), .B(n1185), .Z(n1183) );
  XOR U5028 ( .A(n1186), .B(n1187), .Z(n1185) );
  XOR U5029 ( .A(DB[906]), .B(DB[875]), .Z(n1187) );
  AND U5030 ( .A(n400), .B(n1188), .Z(n1186) );
  XOR U5031 ( .A(n1189), .B(n1190), .Z(n1188) );
  XOR U5032 ( .A(DB[875]), .B(DB[844]), .Z(n1190) );
  AND U5033 ( .A(n404), .B(n1191), .Z(n1189) );
  XOR U5034 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U5035 ( .A(DB[844]), .B(DB[813]), .Z(n1193) );
  AND U5036 ( .A(n408), .B(n1194), .Z(n1192) );
  XOR U5037 ( .A(n1195), .B(n1196), .Z(n1194) );
  XOR U5038 ( .A(DB[813]), .B(DB[782]), .Z(n1196) );
  AND U5039 ( .A(n412), .B(n1197), .Z(n1195) );
  XOR U5040 ( .A(n1198), .B(n1199), .Z(n1197) );
  XOR U5041 ( .A(DB[782]), .B(DB[751]), .Z(n1199) );
  AND U5042 ( .A(n416), .B(n1200), .Z(n1198) );
  XOR U5043 ( .A(n1201), .B(n1202), .Z(n1200) );
  XOR U5044 ( .A(DB[751]), .B(DB[720]), .Z(n1202) );
  AND U5045 ( .A(n420), .B(n1203), .Z(n1201) );
  XOR U5046 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U5047 ( .A(DB[720]), .B(DB[689]), .Z(n1205) );
  AND U5048 ( .A(n424), .B(n1206), .Z(n1204) );
  XOR U5049 ( .A(n1207), .B(n1208), .Z(n1206) );
  XOR U5050 ( .A(DB[689]), .B(DB[658]), .Z(n1208) );
  AND U5051 ( .A(n428), .B(n1209), .Z(n1207) );
  XOR U5052 ( .A(n1210), .B(n1211), .Z(n1209) );
  XOR U5053 ( .A(DB[658]), .B(DB[627]), .Z(n1211) );
  AND U5054 ( .A(n432), .B(n1212), .Z(n1210) );
  XOR U5055 ( .A(n1213), .B(n1214), .Z(n1212) );
  XOR U5056 ( .A(DB[627]), .B(DB[596]), .Z(n1214) );
  AND U5057 ( .A(n436), .B(n1215), .Z(n1213) );
  XOR U5058 ( .A(n1216), .B(n1217), .Z(n1215) );
  XOR U5059 ( .A(DB[596]), .B(DB[565]), .Z(n1217) );
  AND U5060 ( .A(n440), .B(n1218), .Z(n1216) );
  XOR U5061 ( .A(n1219), .B(n1220), .Z(n1218) );
  XOR U5062 ( .A(DB[565]), .B(DB[534]), .Z(n1220) );
  AND U5063 ( .A(n444), .B(n1221), .Z(n1219) );
  XOR U5064 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U5065 ( .A(DB[534]), .B(DB[503]), .Z(n1223) );
  AND U5066 ( .A(n448), .B(n1224), .Z(n1222) );
  XOR U5067 ( .A(n1225), .B(n1226), .Z(n1224) );
  XOR U5068 ( .A(DB[503]), .B(DB[472]), .Z(n1226) );
  AND U5069 ( .A(n452), .B(n1227), .Z(n1225) );
  XOR U5070 ( .A(n1228), .B(n1229), .Z(n1227) );
  XOR U5071 ( .A(DB[472]), .B(DB[441]), .Z(n1229) );
  AND U5072 ( .A(n456), .B(n1230), .Z(n1228) );
  XOR U5073 ( .A(n1231), .B(n1232), .Z(n1230) );
  XOR U5074 ( .A(DB[441]), .B(DB[410]), .Z(n1232) );
  AND U5075 ( .A(n460), .B(n1233), .Z(n1231) );
  XOR U5076 ( .A(n1234), .B(n1235), .Z(n1233) );
  XOR U5077 ( .A(DB[410]), .B(DB[379]), .Z(n1235) );
  AND U5078 ( .A(n464), .B(n1236), .Z(n1234) );
  XOR U5079 ( .A(n1237), .B(n1238), .Z(n1236) );
  XOR U5080 ( .A(DB[379]), .B(DB[348]), .Z(n1238) );
  AND U5081 ( .A(n468), .B(n1239), .Z(n1237) );
  XOR U5082 ( .A(n1240), .B(n1241), .Z(n1239) );
  XOR U5083 ( .A(DB[348]), .B(DB[317]), .Z(n1241) );
  AND U5084 ( .A(n472), .B(n1242), .Z(n1240) );
  XOR U5085 ( .A(n1243), .B(n1244), .Z(n1242) );
  XOR U5086 ( .A(DB[317]), .B(DB[286]), .Z(n1244) );
  AND U5087 ( .A(n476), .B(n1245), .Z(n1243) );
  XOR U5088 ( .A(n1246), .B(n1247), .Z(n1245) );
  XOR U5089 ( .A(DB[286]), .B(DB[255]), .Z(n1247) );
  AND U5090 ( .A(n480), .B(n1248), .Z(n1246) );
  XOR U5091 ( .A(n1249), .B(n1250), .Z(n1248) );
  XOR U5092 ( .A(DB[255]), .B(DB[224]), .Z(n1250) );
  AND U5093 ( .A(n484), .B(n1251), .Z(n1249) );
  XOR U5094 ( .A(n1252), .B(n1253), .Z(n1251) );
  XOR U5095 ( .A(DB[224]), .B(DB[193]), .Z(n1253) );
  AND U5096 ( .A(n488), .B(n1254), .Z(n1252) );
  XOR U5097 ( .A(n1255), .B(n1256), .Z(n1254) );
  XOR U5098 ( .A(DB[193]), .B(DB[162]), .Z(n1256) );
  AND U5099 ( .A(n492), .B(n1257), .Z(n1255) );
  XOR U5100 ( .A(n1258), .B(n1259), .Z(n1257) );
  XOR U5101 ( .A(DB[162]), .B(DB[131]), .Z(n1259) );
  AND U5102 ( .A(n496), .B(n1260), .Z(n1258) );
  XOR U5103 ( .A(n1261), .B(n1262), .Z(n1260) );
  XOR U5104 ( .A(DB[131]), .B(DB[100]), .Z(n1262) );
  AND U5105 ( .A(n500), .B(n1263), .Z(n1261) );
  XOR U5106 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U5107 ( .A(DB[69]), .B(DB[100]), .Z(n1265) );
  AND U5108 ( .A(n504), .B(n1266), .Z(n1264) );
  XOR U5109 ( .A(n1267), .B(n1268), .Z(n1266) );
  XOR U5110 ( .A(DB[69]), .B(DB[38]), .Z(n1268) );
  AND U5111 ( .A(n508), .B(n1269), .Z(n1267) );
  XOR U5112 ( .A(DB[7]), .B(DB[38]), .Z(n1269) );
  XOR U5113 ( .A(DB[3943]), .B(n1270), .Z(min_val_out[6]) );
  AND U5114 ( .A(n2), .B(n1271), .Z(n1270) );
  XOR U5115 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U5116 ( .A(DB[3943]), .B(DB[3912]), .Z(n1273) );
  AND U5117 ( .A(n8), .B(n1274), .Z(n1272) );
  XOR U5118 ( .A(n1275), .B(n1276), .Z(n1274) );
  XOR U5119 ( .A(DB[3912]), .B(DB[3881]), .Z(n1276) );
  AND U5120 ( .A(n12), .B(n1277), .Z(n1275) );
  XOR U5121 ( .A(n1278), .B(n1279), .Z(n1277) );
  XOR U5122 ( .A(DB[3881]), .B(DB[3850]), .Z(n1279) );
  AND U5123 ( .A(n16), .B(n1280), .Z(n1278) );
  XOR U5124 ( .A(n1281), .B(n1282), .Z(n1280) );
  XOR U5125 ( .A(DB[3850]), .B(DB[3819]), .Z(n1282) );
  AND U5126 ( .A(n20), .B(n1283), .Z(n1281) );
  XOR U5127 ( .A(n1284), .B(n1285), .Z(n1283) );
  XOR U5128 ( .A(DB[3819]), .B(DB[3788]), .Z(n1285) );
  AND U5129 ( .A(n24), .B(n1286), .Z(n1284) );
  XOR U5130 ( .A(n1287), .B(n1288), .Z(n1286) );
  XOR U5131 ( .A(DB[3788]), .B(DB[3757]), .Z(n1288) );
  AND U5132 ( .A(n28), .B(n1289), .Z(n1287) );
  XOR U5133 ( .A(n1290), .B(n1291), .Z(n1289) );
  XOR U5134 ( .A(DB[3757]), .B(DB[3726]), .Z(n1291) );
  AND U5135 ( .A(n32), .B(n1292), .Z(n1290) );
  XOR U5136 ( .A(n1293), .B(n1294), .Z(n1292) );
  XOR U5137 ( .A(DB[3726]), .B(DB[3695]), .Z(n1294) );
  AND U5138 ( .A(n36), .B(n1295), .Z(n1293) );
  XOR U5139 ( .A(n1296), .B(n1297), .Z(n1295) );
  XOR U5140 ( .A(DB[3695]), .B(DB[3664]), .Z(n1297) );
  AND U5141 ( .A(n40), .B(n1298), .Z(n1296) );
  XOR U5142 ( .A(n1299), .B(n1300), .Z(n1298) );
  XOR U5143 ( .A(DB[3664]), .B(DB[3633]), .Z(n1300) );
  AND U5144 ( .A(n44), .B(n1301), .Z(n1299) );
  XOR U5145 ( .A(n1302), .B(n1303), .Z(n1301) );
  XOR U5146 ( .A(DB[3633]), .B(DB[3602]), .Z(n1303) );
  AND U5147 ( .A(n48), .B(n1304), .Z(n1302) );
  XOR U5148 ( .A(n1305), .B(n1306), .Z(n1304) );
  XOR U5149 ( .A(DB[3602]), .B(DB[3571]), .Z(n1306) );
  AND U5150 ( .A(n52), .B(n1307), .Z(n1305) );
  XOR U5151 ( .A(n1308), .B(n1309), .Z(n1307) );
  XOR U5152 ( .A(DB[3571]), .B(DB[3540]), .Z(n1309) );
  AND U5153 ( .A(n56), .B(n1310), .Z(n1308) );
  XOR U5154 ( .A(n1311), .B(n1312), .Z(n1310) );
  XOR U5155 ( .A(DB[3540]), .B(DB[3509]), .Z(n1312) );
  AND U5156 ( .A(n60), .B(n1313), .Z(n1311) );
  XOR U5157 ( .A(n1314), .B(n1315), .Z(n1313) );
  XOR U5158 ( .A(DB[3509]), .B(DB[3478]), .Z(n1315) );
  AND U5159 ( .A(n64), .B(n1316), .Z(n1314) );
  XOR U5160 ( .A(n1317), .B(n1318), .Z(n1316) );
  XOR U5161 ( .A(DB[3478]), .B(DB[3447]), .Z(n1318) );
  AND U5162 ( .A(n68), .B(n1319), .Z(n1317) );
  XOR U5163 ( .A(n1320), .B(n1321), .Z(n1319) );
  XOR U5164 ( .A(DB[3447]), .B(DB[3416]), .Z(n1321) );
  AND U5165 ( .A(n72), .B(n1322), .Z(n1320) );
  XOR U5166 ( .A(n1323), .B(n1324), .Z(n1322) );
  XOR U5167 ( .A(DB[3416]), .B(DB[3385]), .Z(n1324) );
  AND U5168 ( .A(n76), .B(n1325), .Z(n1323) );
  XOR U5169 ( .A(n1326), .B(n1327), .Z(n1325) );
  XOR U5170 ( .A(DB[3385]), .B(DB[3354]), .Z(n1327) );
  AND U5171 ( .A(n80), .B(n1328), .Z(n1326) );
  XOR U5172 ( .A(n1329), .B(n1330), .Z(n1328) );
  XOR U5173 ( .A(DB[3354]), .B(DB[3323]), .Z(n1330) );
  AND U5174 ( .A(n84), .B(n1331), .Z(n1329) );
  XOR U5175 ( .A(n1332), .B(n1333), .Z(n1331) );
  XOR U5176 ( .A(DB[3323]), .B(DB[3292]), .Z(n1333) );
  AND U5177 ( .A(n88), .B(n1334), .Z(n1332) );
  XOR U5178 ( .A(n1335), .B(n1336), .Z(n1334) );
  XOR U5179 ( .A(DB[3292]), .B(DB[3261]), .Z(n1336) );
  AND U5180 ( .A(n92), .B(n1337), .Z(n1335) );
  XOR U5181 ( .A(n1338), .B(n1339), .Z(n1337) );
  XOR U5182 ( .A(DB[3261]), .B(DB[3230]), .Z(n1339) );
  AND U5183 ( .A(n96), .B(n1340), .Z(n1338) );
  XOR U5184 ( .A(n1341), .B(n1342), .Z(n1340) );
  XOR U5185 ( .A(DB[3230]), .B(DB[3199]), .Z(n1342) );
  AND U5186 ( .A(n100), .B(n1343), .Z(n1341) );
  XOR U5187 ( .A(n1344), .B(n1345), .Z(n1343) );
  XOR U5188 ( .A(DB[3199]), .B(DB[3168]), .Z(n1345) );
  AND U5189 ( .A(n104), .B(n1346), .Z(n1344) );
  XOR U5190 ( .A(n1347), .B(n1348), .Z(n1346) );
  XOR U5191 ( .A(DB[3168]), .B(DB[3137]), .Z(n1348) );
  AND U5192 ( .A(n108), .B(n1349), .Z(n1347) );
  XOR U5193 ( .A(n1350), .B(n1351), .Z(n1349) );
  XOR U5194 ( .A(DB[3137]), .B(DB[3106]), .Z(n1351) );
  AND U5195 ( .A(n112), .B(n1352), .Z(n1350) );
  XOR U5196 ( .A(n1353), .B(n1354), .Z(n1352) );
  XOR U5197 ( .A(DB[3106]), .B(DB[3075]), .Z(n1354) );
  AND U5198 ( .A(n116), .B(n1355), .Z(n1353) );
  XOR U5199 ( .A(n1356), .B(n1357), .Z(n1355) );
  XOR U5200 ( .A(DB[3075]), .B(DB[3044]), .Z(n1357) );
  AND U5201 ( .A(n120), .B(n1358), .Z(n1356) );
  XOR U5202 ( .A(n1359), .B(n1360), .Z(n1358) );
  XOR U5203 ( .A(DB[3044]), .B(DB[3013]), .Z(n1360) );
  AND U5204 ( .A(n124), .B(n1361), .Z(n1359) );
  XOR U5205 ( .A(n1362), .B(n1363), .Z(n1361) );
  XOR U5206 ( .A(DB[3013]), .B(DB[2982]), .Z(n1363) );
  AND U5207 ( .A(n128), .B(n1364), .Z(n1362) );
  XOR U5208 ( .A(n1365), .B(n1366), .Z(n1364) );
  XOR U5209 ( .A(DB[2982]), .B(DB[2951]), .Z(n1366) );
  AND U5210 ( .A(n132), .B(n1367), .Z(n1365) );
  XOR U5211 ( .A(n1368), .B(n1369), .Z(n1367) );
  XOR U5212 ( .A(DB[2951]), .B(DB[2920]), .Z(n1369) );
  AND U5213 ( .A(n136), .B(n1370), .Z(n1368) );
  XOR U5214 ( .A(n1371), .B(n1372), .Z(n1370) );
  XOR U5215 ( .A(DB[2920]), .B(DB[2889]), .Z(n1372) );
  AND U5216 ( .A(n140), .B(n1373), .Z(n1371) );
  XOR U5217 ( .A(n1374), .B(n1375), .Z(n1373) );
  XOR U5218 ( .A(DB[2889]), .B(DB[2858]), .Z(n1375) );
  AND U5219 ( .A(n144), .B(n1376), .Z(n1374) );
  XOR U5220 ( .A(n1377), .B(n1378), .Z(n1376) );
  XOR U5221 ( .A(DB[2858]), .B(DB[2827]), .Z(n1378) );
  AND U5222 ( .A(n148), .B(n1379), .Z(n1377) );
  XOR U5223 ( .A(n1380), .B(n1381), .Z(n1379) );
  XOR U5224 ( .A(DB[2827]), .B(DB[2796]), .Z(n1381) );
  AND U5225 ( .A(n152), .B(n1382), .Z(n1380) );
  XOR U5226 ( .A(n1383), .B(n1384), .Z(n1382) );
  XOR U5227 ( .A(DB[2796]), .B(DB[2765]), .Z(n1384) );
  AND U5228 ( .A(n156), .B(n1385), .Z(n1383) );
  XOR U5229 ( .A(n1386), .B(n1387), .Z(n1385) );
  XOR U5230 ( .A(DB[2765]), .B(DB[2734]), .Z(n1387) );
  AND U5231 ( .A(n160), .B(n1388), .Z(n1386) );
  XOR U5232 ( .A(n1389), .B(n1390), .Z(n1388) );
  XOR U5233 ( .A(DB[2734]), .B(DB[2703]), .Z(n1390) );
  AND U5234 ( .A(n164), .B(n1391), .Z(n1389) );
  XOR U5235 ( .A(n1392), .B(n1393), .Z(n1391) );
  XOR U5236 ( .A(DB[2703]), .B(DB[2672]), .Z(n1393) );
  AND U5237 ( .A(n168), .B(n1394), .Z(n1392) );
  XOR U5238 ( .A(n1395), .B(n1396), .Z(n1394) );
  XOR U5239 ( .A(DB[2672]), .B(DB[2641]), .Z(n1396) );
  AND U5240 ( .A(n172), .B(n1397), .Z(n1395) );
  XOR U5241 ( .A(n1398), .B(n1399), .Z(n1397) );
  XOR U5242 ( .A(DB[2641]), .B(DB[2610]), .Z(n1399) );
  AND U5243 ( .A(n176), .B(n1400), .Z(n1398) );
  XOR U5244 ( .A(n1401), .B(n1402), .Z(n1400) );
  XOR U5245 ( .A(DB[2610]), .B(DB[2579]), .Z(n1402) );
  AND U5246 ( .A(n180), .B(n1403), .Z(n1401) );
  XOR U5247 ( .A(n1404), .B(n1405), .Z(n1403) );
  XOR U5248 ( .A(DB[2579]), .B(DB[2548]), .Z(n1405) );
  AND U5249 ( .A(n184), .B(n1406), .Z(n1404) );
  XOR U5250 ( .A(n1407), .B(n1408), .Z(n1406) );
  XOR U5251 ( .A(DB[2548]), .B(DB[2517]), .Z(n1408) );
  AND U5252 ( .A(n188), .B(n1409), .Z(n1407) );
  XOR U5253 ( .A(n1410), .B(n1411), .Z(n1409) );
  XOR U5254 ( .A(DB[2517]), .B(DB[2486]), .Z(n1411) );
  AND U5255 ( .A(n192), .B(n1412), .Z(n1410) );
  XOR U5256 ( .A(n1413), .B(n1414), .Z(n1412) );
  XOR U5257 ( .A(DB[2486]), .B(DB[2455]), .Z(n1414) );
  AND U5258 ( .A(n196), .B(n1415), .Z(n1413) );
  XOR U5259 ( .A(n1416), .B(n1417), .Z(n1415) );
  XOR U5260 ( .A(DB[2455]), .B(DB[2424]), .Z(n1417) );
  AND U5261 ( .A(n200), .B(n1418), .Z(n1416) );
  XOR U5262 ( .A(n1419), .B(n1420), .Z(n1418) );
  XOR U5263 ( .A(DB[2424]), .B(DB[2393]), .Z(n1420) );
  AND U5264 ( .A(n204), .B(n1421), .Z(n1419) );
  XOR U5265 ( .A(n1422), .B(n1423), .Z(n1421) );
  XOR U5266 ( .A(DB[2393]), .B(DB[2362]), .Z(n1423) );
  AND U5267 ( .A(n208), .B(n1424), .Z(n1422) );
  XOR U5268 ( .A(n1425), .B(n1426), .Z(n1424) );
  XOR U5269 ( .A(DB[2362]), .B(DB[2331]), .Z(n1426) );
  AND U5270 ( .A(n212), .B(n1427), .Z(n1425) );
  XOR U5271 ( .A(n1428), .B(n1429), .Z(n1427) );
  XOR U5272 ( .A(DB[2331]), .B(DB[2300]), .Z(n1429) );
  AND U5273 ( .A(n216), .B(n1430), .Z(n1428) );
  XOR U5274 ( .A(n1431), .B(n1432), .Z(n1430) );
  XOR U5275 ( .A(DB[2300]), .B(DB[2269]), .Z(n1432) );
  AND U5276 ( .A(n220), .B(n1433), .Z(n1431) );
  XOR U5277 ( .A(n1434), .B(n1435), .Z(n1433) );
  XOR U5278 ( .A(DB[2269]), .B(DB[2238]), .Z(n1435) );
  AND U5279 ( .A(n224), .B(n1436), .Z(n1434) );
  XOR U5280 ( .A(n1437), .B(n1438), .Z(n1436) );
  XOR U5281 ( .A(DB[2238]), .B(DB[2207]), .Z(n1438) );
  AND U5282 ( .A(n228), .B(n1439), .Z(n1437) );
  XOR U5283 ( .A(n1440), .B(n1441), .Z(n1439) );
  XOR U5284 ( .A(DB[2207]), .B(DB[2176]), .Z(n1441) );
  AND U5285 ( .A(n232), .B(n1442), .Z(n1440) );
  XOR U5286 ( .A(n1443), .B(n1444), .Z(n1442) );
  XOR U5287 ( .A(DB[2176]), .B(DB[2145]), .Z(n1444) );
  AND U5288 ( .A(n236), .B(n1445), .Z(n1443) );
  XOR U5289 ( .A(n1446), .B(n1447), .Z(n1445) );
  XOR U5290 ( .A(DB[2145]), .B(DB[2114]), .Z(n1447) );
  AND U5291 ( .A(n240), .B(n1448), .Z(n1446) );
  XOR U5292 ( .A(n1449), .B(n1450), .Z(n1448) );
  XOR U5293 ( .A(DB[2114]), .B(DB[2083]), .Z(n1450) );
  AND U5294 ( .A(n244), .B(n1451), .Z(n1449) );
  XOR U5295 ( .A(n1452), .B(n1453), .Z(n1451) );
  XOR U5296 ( .A(DB[2083]), .B(DB[2052]), .Z(n1453) );
  AND U5297 ( .A(n248), .B(n1454), .Z(n1452) );
  XOR U5298 ( .A(n1455), .B(n1456), .Z(n1454) );
  XOR U5299 ( .A(DB[2052]), .B(DB[2021]), .Z(n1456) );
  AND U5300 ( .A(n252), .B(n1457), .Z(n1455) );
  XOR U5301 ( .A(n1458), .B(n1459), .Z(n1457) );
  XOR U5302 ( .A(DB[2021]), .B(DB[1990]), .Z(n1459) );
  AND U5303 ( .A(n256), .B(n1460), .Z(n1458) );
  XOR U5304 ( .A(n1461), .B(n1462), .Z(n1460) );
  XOR U5305 ( .A(DB[1990]), .B(DB[1959]), .Z(n1462) );
  AND U5306 ( .A(n260), .B(n1463), .Z(n1461) );
  XOR U5307 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U5308 ( .A(DB[1959]), .B(DB[1928]), .Z(n1465) );
  AND U5309 ( .A(n264), .B(n1466), .Z(n1464) );
  XOR U5310 ( .A(n1467), .B(n1468), .Z(n1466) );
  XOR U5311 ( .A(DB[1928]), .B(DB[1897]), .Z(n1468) );
  AND U5312 ( .A(n268), .B(n1469), .Z(n1467) );
  XOR U5313 ( .A(n1470), .B(n1471), .Z(n1469) );
  XOR U5314 ( .A(DB[1897]), .B(DB[1866]), .Z(n1471) );
  AND U5315 ( .A(n272), .B(n1472), .Z(n1470) );
  XOR U5316 ( .A(n1473), .B(n1474), .Z(n1472) );
  XOR U5317 ( .A(DB[1866]), .B(DB[1835]), .Z(n1474) );
  AND U5318 ( .A(n276), .B(n1475), .Z(n1473) );
  XOR U5319 ( .A(n1476), .B(n1477), .Z(n1475) );
  XOR U5320 ( .A(DB[1835]), .B(DB[1804]), .Z(n1477) );
  AND U5321 ( .A(n280), .B(n1478), .Z(n1476) );
  XOR U5322 ( .A(n1479), .B(n1480), .Z(n1478) );
  XOR U5323 ( .A(DB[1804]), .B(DB[1773]), .Z(n1480) );
  AND U5324 ( .A(n284), .B(n1481), .Z(n1479) );
  XOR U5325 ( .A(n1482), .B(n1483), .Z(n1481) );
  XOR U5326 ( .A(DB[1773]), .B(DB[1742]), .Z(n1483) );
  AND U5327 ( .A(n288), .B(n1484), .Z(n1482) );
  XOR U5328 ( .A(n1485), .B(n1486), .Z(n1484) );
  XOR U5329 ( .A(DB[1742]), .B(DB[1711]), .Z(n1486) );
  AND U5330 ( .A(n292), .B(n1487), .Z(n1485) );
  XOR U5331 ( .A(n1488), .B(n1489), .Z(n1487) );
  XOR U5332 ( .A(DB[1711]), .B(DB[1680]), .Z(n1489) );
  AND U5333 ( .A(n296), .B(n1490), .Z(n1488) );
  XOR U5334 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U5335 ( .A(DB[1680]), .B(DB[1649]), .Z(n1492) );
  AND U5336 ( .A(n300), .B(n1493), .Z(n1491) );
  XOR U5337 ( .A(n1494), .B(n1495), .Z(n1493) );
  XOR U5338 ( .A(DB[1649]), .B(DB[1618]), .Z(n1495) );
  AND U5339 ( .A(n304), .B(n1496), .Z(n1494) );
  XOR U5340 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR U5341 ( .A(DB[1618]), .B(DB[1587]), .Z(n1498) );
  AND U5342 ( .A(n308), .B(n1499), .Z(n1497) );
  XOR U5343 ( .A(n1500), .B(n1501), .Z(n1499) );
  XOR U5344 ( .A(DB[1587]), .B(DB[1556]), .Z(n1501) );
  AND U5345 ( .A(n312), .B(n1502), .Z(n1500) );
  XOR U5346 ( .A(n1503), .B(n1504), .Z(n1502) );
  XOR U5347 ( .A(DB[1556]), .B(DB[1525]), .Z(n1504) );
  AND U5348 ( .A(n316), .B(n1505), .Z(n1503) );
  XOR U5349 ( .A(n1506), .B(n1507), .Z(n1505) );
  XOR U5350 ( .A(DB[1525]), .B(DB[1494]), .Z(n1507) );
  AND U5351 ( .A(n320), .B(n1508), .Z(n1506) );
  XOR U5352 ( .A(n1509), .B(n1510), .Z(n1508) );
  XOR U5353 ( .A(DB[1494]), .B(DB[1463]), .Z(n1510) );
  AND U5354 ( .A(n324), .B(n1511), .Z(n1509) );
  XOR U5355 ( .A(n1512), .B(n1513), .Z(n1511) );
  XOR U5356 ( .A(DB[1463]), .B(DB[1432]), .Z(n1513) );
  AND U5357 ( .A(n328), .B(n1514), .Z(n1512) );
  XOR U5358 ( .A(n1515), .B(n1516), .Z(n1514) );
  XOR U5359 ( .A(DB[1432]), .B(DB[1401]), .Z(n1516) );
  AND U5360 ( .A(n332), .B(n1517), .Z(n1515) );
  XOR U5361 ( .A(n1518), .B(n1519), .Z(n1517) );
  XOR U5362 ( .A(DB[1401]), .B(DB[1370]), .Z(n1519) );
  AND U5363 ( .A(n336), .B(n1520), .Z(n1518) );
  XOR U5364 ( .A(n1521), .B(n1522), .Z(n1520) );
  XOR U5365 ( .A(DB[1370]), .B(DB[1339]), .Z(n1522) );
  AND U5366 ( .A(n340), .B(n1523), .Z(n1521) );
  XOR U5367 ( .A(n1524), .B(n1525), .Z(n1523) );
  XOR U5368 ( .A(DB[1339]), .B(DB[1308]), .Z(n1525) );
  AND U5369 ( .A(n344), .B(n1526), .Z(n1524) );
  XOR U5370 ( .A(n1527), .B(n1528), .Z(n1526) );
  XOR U5371 ( .A(DB[1308]), .B(DB[1277]), .Z(n1528) );
  AND U5372 ( .A(n348), .B(n1529), .Z(n1527) );
  XOR U5373 ( .A(n1530), .B(n1531), .Z(n1529) );
  XOR U5374 ( .A(DB[1277]), .B(DB[1246]), .Z(n1531) );
  AND U5375 ( .A(n352), .B(n1532), .Z(n1530) );
  XOR U5376 ( .A(n1533), .B(n1534), .Z(n1532) );
  XOR U5377 ( .A(DB[1246]), .B(DB[1215]), .Z(n1534) );
  AND U5378 ( .A(n356), .B(n1535), .Z(n1533) );
  XOR U5379 ( .A(n1536), .B(n1537), .Z(n1535) );
  XOR U5380 ( .A(DB[1215]), .B(DB[1184]), .Z(n1537) );
  AND U5381 ( .A(n360), .B(n1538), .Z(n1536) );
  XOR U5382 ( .A(n1539), .B(n1540), .Z(n1538) );
  XOR U5383 ( .A(DB[1184]), .B(DB[1153]), .Z(n1540) );
  AND U5384 ( .A(n364), .B(n1541), .Z(n1539) );
  XOR U5385 ( .A(n1542), .B(n1543), .Z(n1541) );
  XOR U5386 ( .A(DB[1153]), .B(DB[1122]), .Z(n1543) );
  AND U5387 ( .A(n368), .B(n1544), .Z(n1542) );
  XOR U5388 ( .A(n1545), .B(n1546), .Z(n1544) );
  XOR U5389 ( .A(DB[1122]), .B(DB[1091]), .Z(n1546) );
  AND U5390 ( .A(n372), .B(n1547), .Z(n1545) );
  XOR U5391 ( .A(n1548), .B(n1549), .Z(n1547) );
  XOR U5392 ( .A(DB[1091]), .B(DB[1060]), .Z(n1549) );
  AND U5393 ( .A(n376), .B(n1550), .Z(n1548) );
  XOR U5394 ( .A(n1551), .B(n1552), .Z(n1550) );
  XOR U5395 ( .A(DB[1060]), .B(DB[1029]), .Z(n1552) );
  AND U5396 ( .A(n380), .B(n1553), .Z(n1551) );
  XOR U5397 ( .A(n1554), .B(n1555), .Z(n1553) );
  XOR U5398 ( .A(DB[998]), .B(DB[1029]), .Z(n1555) );
  AND U5399 ( .A(n384), .B(n1556), .Z(n1554) );
  XOR U5400 ( .A(n1557), .B(n1558), .Z(n1556) );
  XOR U5401 ( .A(DB[998]), .B(DB[967]), .Z(n1558) );
  AND U5402 ( .A(n388), .B(n1559), .Z(n1557) );
  XOR U5403 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U5404 ( .A(DB[967]), .B(DB[936]), .Z(n1561) );
  AND U5405 ( .A(n392), .B(n1562), .Z(n1560) );
  XOR U5406 ( .A(n1563), .B(n1564), .Z(n1562) );
  XOR U5407 ( .A(DB[936]), .B(DB[905]), .Z(n1564) );
  AND U5408 ( .A(n396), .B(n1565), .Z(n1563) );
  XOR U5409 ( .A(n1566), .B(n1567), .Z(n1565) );
  XOR U5410 ( .A(DB[905]), .B(DB[874]), .Z(n1567) );
  AND U5411 ( .A(n400), .B(n1568), .Z(n1566) );
  XOR U5412 ( .A(n1569), .B(n1570), .Z(n1568) );
  XOR U5413 ( .A(DB[874]), .B(DB[843]), .Z(n1570) );
  AND U5414 ( .A(n404), .B(n1571), .Z(n1569) );
  XOR U5415 ( .A(n1572), .B(n1573), .Z(n1571) );
  XOR U5416 ( .A(DB[843]), .B(DB[812]), .Z(n1573) );
  AND U5417 ( .A(n408), .B(n1574), .Z(n1572) );
  XOR U5418 ( .A(n1575), .B(n1576), .Z(n1574) );
  XOR U5419 ( .A(DB[812]), .B(DB[781]), .Z(n1576) );
  AND U5420 ( .A(n412), .B(n1577), .Z(n1575) );
  XOR U5421 ( .A(n1578), .B(n1579), .Z(n1577) );
  XOR U5422 ( .A(DB[781]), .B(DB[750]), .Z(n1579) );
  AND U5423 ( .A(n416), .B(n1580), .Z(n1578) );
  XOR U5424 ( .A(n1581), .B(n1582), .Z(n1580) );
  XOR U5425 ( .A(DB[750]), .B(DB[719]), .Z(n1582) );
  AND U5426 ( .A(n420), .B(n1583), .Z(n1581) );
  XOR U5427 ( .A(n1584), .B(n1585), .Z(n1583) );
  XOR U5428 ( .A(DB[719]), .B(DB[688]), .Z(n1585) );
  AND U5429 ( .A(n424), .B(n1586), .Z(n1584) );
  XOR U5430 ( .A(n1587), .B(n1588), .Z(n1586) );
  XOR U5431 ( .A(DB[688]), .B(DB[657]), .Z(n1588) );
  AND U5432 ( .A(n428), .B(n1589), .Z(n1587) );
  XOR U5433 ( .A(n1590), .B(n1591), .Z(n1589) );
  XOR U5434 ( .A(DB[657]), .B(DB[626]), .Z(n1591) );
  AND U5435 ( .A(n432), .B(n1592), .Z(n1590) );
  XOR U5436 ( .A(n1593), .B(n1594), .Z(n1592) );
  XOR U5437 ( .A(DB[626]), .B(DB[595]), .Z(n1594) );
  AND U5438 ( .A(n436), .B(n1595), .Z(n1593) );
  XOR U5439 ( .A(n1596), .B(n1597), .Z(n1595) );
  XOR U5440 ( .A(DB[595]), .B(DB[564]), .Z(n1597) );
  AND U5441 ( .A(n440), .B(n1598), .Z(n1596) );
  XOR U5442 ( .A(n1599), .B(n1600), .Z(n1598) );
  XOR U5443 ( .A(DB[564]), .B(DB[533]), .Z(n1600) );
  AND U5444 ( .A(n444), .B(n1601), .Z(n1599) );
  XOR U5445 ( .A(n1602), .B(n1603), .Z(n1601) );
  XOR U5446 ( .A(DB[533]), .B(DB[502]), .Z(n1603) );
  AND U5447 ( .A(n448), .B(n1604), .Z(n1602) );
  XOR U5448 ( .A(n1605), .B(n1606), .Z(n1604) );
  XOR U5449 ( .A(DB[502]), .B(DB[471]), .Z(n1606) );
  AND U5450 ( .A(n452), .B(n1607), .Z(n1605) );
  XOR U5451 ( .A(n1608), .B(n1609), .Z(n1607) );
  XOR U5452 ( .A(DB[471]), .B(DB[440]), .Z(n1609) );
  AND U5453 ( .A(n456), .B(n1610), .Z(n1608) );
  XOR U5454 ( .A(n1611), .B(n1612), .Z(n1610) );
  XOR U5455 ( .A(DB[440]), .B(DB[409]), .Z(n1612) );
  AND U5456 ( .A(n460), .B(n1613), .Z(n1611) );
  XOR U5457 ( .A(n1614), .B(n1615), .Z(n1613) );
  XOR U5458 ( .A(DB[409]), .B(DB[378]), .Z(n1615) );
  AND U5459 ( .A(n464), .B(n1616), .Z(n1614) );
  XOR U5460 ( .A(n1617), .B(n1618), .Z(n1616) );
  XOR U5461 ( .A(DB[378]), .B(DB[347]), .Z(n1618) );
  AND U5462 ( .A(n468), .B(n1619), .Z(n1617) );
  XOR U5463 ( .A(n1620), .B(n1621), .Z(n1619) );
  XOR U5464 ( .A(DB[347]), .B(DB[316]), .Z(n1621) );
  AND U5465 ( .A(n472), .B(n1622), .Z(n1620) );
  XOR U5466 ( .A(n1623), .B(n1624), .Z(n1622) );
  XOR U5467 ( .A(DB[316]), .B(DB[285]), .Z(n1624) );
  AND U5468 ( .A(n476), .B(n1625), .Z(n1623) );
  XOR U5469 ( .A(n1626), .B(n1627), .Z(n1625) );
  XOR U5470 ( .A(DB[285]), .B(DB[254]), .Z(n1627) );
  AND U5471 ( .A(n480), .B(n1628), .Z(n1626) );
  XOR U5472 ( .A(n1629), .B(n1630), .Z(n1628) );
  XOR U5473 ( .A(DB[254]), .B(DB[223]), .Z(n1630) );
  AND U5474 ( .A(n484), .B(n1631), .Z(n1629) );
  XOR U5475 ( .A(n1632), .B(n1633), .Z(n1631) );
  XOR U5476 ( .A(DB[223]), .B(DB[192]), .Z(n1633) );
  AND U5477 ( .A(n488), .B(n1634), .Z(n1632) );
  XOR U5478 ( .A(n1635), .B(n1636), .Z(n1634) );
  XOR U5479 ( .A(DB[192]), .B(DB[161]), .Z(n1636) );
  AND U5480 ( .A(n492), .B(n1637), .Z(n1635) );
  XOR U5481 ( .A(n1638), .B(n1639), .Z(n1637) );
  XOR U5482 ( .A(DB[161]), .B(DB[130]), .Z(n1639) );
  AND U5483 ( .A(n496), .B(n1640), .Z(n1638) );
  XOR U5484 ( .A(n1641), .B(n1642), .Z(n1640) );
  XOR U5485 ( .A(DB[99]), .B(DB[130]), .Z(n1642) );
  AND U5486 ( .A(n500), .B(n1643), .Z(n1641) );
  XOR U5487 ( .A(n1644), .B(n1645), .Z(n1643) );
  XOR U5488 ( .A(DB[99]), .B(DB[68]), .Z(n1645) );
  AND U5489 ( .A(n504), .B(n1646), .Z(n1644) );
  XOR U5490 ( .A(n1647), .B(n1648), .Z(n1646) );
  XOR U5491 ( .A(DB[68]), .B(DB[37]), .Z(n1648) );
  AND U5492 ( .A(n508), .B(n1649), .Z(n1647) );
  XOR U5493 ( .A(DB[6]), .B(DB[37]), .Z(n1649) );
  XOR U5494 ( .A(DB[3942]), .B(n1650), .Z(min_val_out[5]) );
  AND U5495 ( .A(n2), .B(n1651), .Z(n1650) );
  XOR U5496 ( .A(n1652), .B(n1653), .Z(n1651) );
  XOR U5497 ( .A(DB[3942]), .B(DB[3911]), .Z(n1653) );
  AND U5498 ( .A(n8), .B(n1654), .Z(n1652) );
  XOR U5499 ( .A(n1655), .B(n1656), .Z(n1654) );
  XOR U5500 ( .A(DB[3911]), .B(DB[3880]), .Z(n1656) );
  AND U5501 ( .A(n12), .B(n1657), .Z(n1655) );
  XOR U5502 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U5503 ( .A(DB[3880]), .B(DB[3849]), .Z(n1659) );
  AND U5504 ( .A(n16), .B(n1660), .Z(n1658) );
  XOR U5505 ( .A(n1661), .B(n1662), .Z(n1660) );
  XOR U5506 ( .A(DB[3849]), .B(DB[3818]), .Z(n1662) );
  AND U5507 ( .A(n20), .B(n1663), .Z(n1661) );
  XOR U5508 ( .A(n1664), .B(n1665), .Z(n1663) );
  XOR U5509 ( .A(DB[3818]), .B(DB[3787]), .Z(n1665) );
  AND U5510 ( .A(n24), .B(n1666), .Z(n1664) );
  XOR U5511 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U5512 ( .A(DB[3787]), .B(DB[3756]), .Z(n1668) );
  AND U5513 ( .A(n28), .B(n1669), .Z(n1667) );
  XOR U5514 ( .A(n1670), .B(n1671), .Z(n1669) );
  XOR U5515 ( .A(DB[3756]), .B(DB[3725]), .Z(n1671) );
  AND U5516 ( .A(n32), .B(n1672), .Z(n1670) );
  XOR U5517 ( .A(n1673), .B(n1674), .Z(n1672) );
  XOR U5518 ( .A(DB[3725]), .B(DB[3694]), .Z(n1674) );
  AND U5519 ( .A(n36), .B(n1675), .Z(n1673) );
  XOR U5520 ( .A(n1676), .B(n1677), .Z(n1675) );
  XOR U5521 ( .A(DB[3694]), .B(DB[3663]), .Z(n1677) );
  AND U5522 ( .A(n40), .B(n1678), .Z(n1676) );
  XOR U5523 ( .A(n1679), .B(n1680), .Z(n1678) );
  XOR U5524 ( .A(DB[3663]), .B(DB[3632]), .Z(n1680) );
  AND U5525 ( .A(n44), .B(n1681), .Z(n1679) );
  XOR U5526 ( .A(n1682), .B(n1683), .Z(n1681) );
  XOR U5527 ( .A(DB[3632]), .B(DB[3601]), .Z(n1683) );
  AND U5528 ( .A(n48), .B(n1684), .Z(n1682) );
  XOR U5529 ( .A(n1685), .B(n1686), .Z(n1684) );
  XOR U5530 ( .A(DB[3601]), .B(DB[3570]), .Z(n1686) );
  AND U5531 ( .A(n52), .B(n1687), .Z(n1685) );
  XOR U5532 ( .A(n1688), .B(n1689), .Z(n1687) );
  XOR U5533 ( .A(DB[3570]), .B(DB[3539]), .Z(n1689) );
  AND U5534 ( .A(n56), .B(n1690), .Z(n1688) );
  XOR U5535 ( .A(n1691), .B(n1692), .Z(n1690) );
  XOR U5536 ( .A(DB[3539]), .B(DB[3508]), .Z(n1692) );
  AND U5537 ( .A(n60), .B(n1693), .Z(n1691) );
  XOR U5538 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U5539 ( .A(DB[3508]), .B(DB[3477]), .Z(n1695) );
  AND U5540 ( .A(n64), .B(n1696), .Z(n1694) );
  XOR U5541 ( .A(n1697), .B(n1698), .Z(n1696) );
  XOR U5542 ( .A(DB[3477]), .B(DB[3446]), .Z(n1698) );
  AND U5543 ( .A(n68), .B(n1699), .Z(n1697) );
  XOR U5544 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U5545 ( .A(DB[3446]), .B(DB[3415]), .Z(n1701) );
  AND U5546 ( .A(n72), .B(n1702), .Z(n1700) );
  XOR U5547 ( .A(n1703), .B(n1704), .Z(n1702) );
  XOR U5548 ( .A(DB[3415]), .B(DB[3384]), .Z(n1704) );
  AND U5549 ( .A(n76), .B(n1705), .Z(n1703) );
  XOR U5550 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U5551 ( .A(DB[3384]), .B(DB[3353]), .Z(n1707) );
  AND U5552 ( .A(n80), .B(n1708), .Z(n1706) );
  XOR U5553 ( .A(n1709), .B(n1710), .Z(n1708) );
  XOR U5554 ( .A(DB[3353]), .B(DB[3322]), .Z(n1710) );
  AND U5555 ( .A(n84), .B(n1711), .Z(n1709) );
  XOR U5556 ( .A(n1712), .B(n1713), .Z(n1711) );
  XOR U5557 ( .A(DB[3322]), .B(DB[3291]), .Z(n1713) );
  AND U5558 ( .A(n88), .B(n1714), .Z(n1712) );
  XOR U5559 ( .A(n1715), .B(n1716), .Z(n1714) );
  XOR U5560 ( .A(DB[3291]), .B(DB[3260]), .Z(n1716) );
  AND U5561 ( .A(n92), .B(n1717), .Z(n1715) );
  XOR U5562 ( .A(n1718), .B(n1719), .Z(n1717) );
  XOR U5563 ( .A(DB[3260]), .B(DB[3229]), .Z(n1719) );
  AND U5564 ( .A(n96), .B(n1720), .Z(n1718) );
  XOR U5565 ( .A(n1721), .B(n1722), .Z(n1720) );
  XOR U5566 ( .A(DB[3229]), .B(DB[3198]), .Z(n1722) );
  AND U5567 ( .A(n100), .B(n1723), .Z(n1721) );
  XOR U5568 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U5569 ( .A(DB[3198]), .B(DB[3167]), .Z(n1725) );
  AND U5570 ( .A(n104), .B(n1726), .Z(n1724) );
  XOR U5571 ( .A(n1727), .B(n1728), .Z(n1726) );
  XOR U5572 ( .A(DB[3167]), .B(DB[3136]), .Z(n1728) );
  AND U5573 ( .A(n108), .B(n1729), .Z(n1727) );
  XOR U5574 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U5575 ( .A(DB[3136]), .B(DB[3105]), .Z(n1731) );
  AND U5576 ( .A(n112), .B(n1732), .Z(n1730) );
  XOR U5577 ( .A(n1733), .B(n1734), .Z(n1732) );
  XOR U5578 ( .A(DB[3105]), .B(DB[3074]), .Z(n1734) );
  AND U5579 ( .A(n116), .B(n1735), .Z(n1733) );
  XOR U5580 ( .A(n1736), .B(n1737), .Z(n1735) );
  XOR U5581 ( .A(DB[3074]), .B(DB[3043]), .Z(n1737) );
  AND U5582 ( .A(n120), .B(n1738), .Z(n1736) );
  XOR U5583 ( .A(n1739), .B(n1740), .Z(n1738) );
  XOR U5584 ( .A(DB[3043]), .B(DB[3012]), .Z(n1740) );
  AND U5585 ( .A(n124), .B(n1741), .Z(n1739) );
  XOR U5586 ( .A(n1742), .B(n1743), .Z(n1741) );
  XOR U5587 ( .A(DB[3012]), .B(DB[2981]), .Z(n1743) );
  AND U5588 ( .A(n128), .B(n1744), .Z(n1742) );
  XOR U5589 ( .A(n1745), .B(n1746), .Z(n1744) );
  XOR U5590 ( .A(DB[2981]), .B(DB[2950]), .Z(n1746) );
  AND U5591 ( .A(n132), .B(n1747), .Z(n1745) );
  XOR U5592 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U5593 ( .A(DB[2950]), .B(DB[2919]), .Z(n1749) );
  AND U5594 ( .A(n136), .B(n1750), .Z(n1748) );
  XOR U5595 ( .A(n1751), .B(n1752), .Z(n1750) );
  XOR U5596 ( .A(DB[2919]), .B(DB[2888]), .Z(n1752) );
  AND U5597 ( .A(n140), .B(n1753), .Z(n1751) );
  XOR U5598 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U5599 ( .A(DB[2888]), .B(DB[2857]), .Z(n1755) );
  AND U5600 ( .A(n144), .B(n1756), .Z(n1754) );
  XOR U5601 ( .A(n1757), .B(n1758), .Z(n1756) );
  XOR U5602 ( .A(DB[2857]), .B(DB[2826]), .Z(n1758) );
  AND U5603 ( .A(n148), .B(n1759), .Z(n1757) );
  XOR U5604 ( .A(n1760), .B(n1761), .Z(n1759) );
  XOR U5605 ( .A(DB[2826]), .B(DB[2795]), .Z(n1761) );
  AND U5606 ( .A(n152), .B(n1762), .Z(n1760) );
  XOR U5607 ( .A(n1763), .B(n1764), .Z(n1762) );
  XOR U5608 ( .A(DB[2795]), .B(DB[2764]), .Z(n1764) );
  AND U5609 ( .A(n156), .B(n1765), .Z(n1763) );
  XOR U5610 ( .A(n1766), .B(n1767), .Z(n1765) );
  XOR U5611 ( .A(DB[2764]), .B(DB[2733]), .Z(n1767) );
  AND U5612 ( .A(n160), .B(n1768), .Z(n1766) );
  XOR U5613 ( .A(n1769), .B(n1770), .Z(n1768) );
  XOR U5614 ( .A(DB[2733]), .B(DB[2702]), .Z(n1770) );
  AND U5615 ( .A(n164), .B(n1771), .Z(n1769) );
  XOR U5616 ( .A(n1772), .B(n1773), .Z(n1771) );
  XOR U5617 ( .A(DB[2702]), .B(DB[2671]), .Z(n1773) );
  AND U5618 ( .A(n168), .B(n1774), .Z(n1772) );
  XOR U5619 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U5620 ( .A(DB[2671]), .B(DB[2640]), .Z(n1776) );
  AND U5621 ( .A(n172), .B(n1777), .Z(n1775) );
  XOR U5622 ( .A(n1778), .B(n1779), .Z(n1777) );
  XOR U5623 ( .A(DB[2640]), .B(DB[2609]), .Z(n1779) );
  AND U5624 ( .A(n176), .B(n1780), .Z(n1778) );
  XOR U5625 ( .A(n1781), .B(n1782), .Z(n1780) );
  XOR U5626 ( .A(DB[2609]), .B(DB[2578]), .Z(n1782) );
  AND U5627 ( .A(n180), .B(n1783), .Z(n1781) );
  XOR U5628 ( .A(n1784), .B(n1785), .Z(n1783) );
  XOR U5629 ( .A(DB[2578]), .B(DB[2547]), .Z(n1785) );
  AND U5630 ( .A(n184), .B(n1786), .Z(n1784) );
  XOR U5631 ( .A(n1787), .B(n1788), .Z(n1786) );
  XOR U5632 ( .A(DB[2547]), .B(DB[2516]), .Z(n1788) );
  AND U5633 ( .A(n188), .B(n1789), .Z(n1787) );
  XOR U5634 ( .A(n1790), .B(n1791), .Z(n1789) );
  XOR U5635 ( .A(DB[2516]), .B(DB[2485]), .Z(n1791) );
  AND U5636 ( .A(n192), .B(n1792), .Z(n1790) );
  XOR U5637 ( .A(n1793), .B(n1794), .Z(n1792) );
  XOR U5638 ( .A(DB[2485]), .B(DB[2454]), .Z(n1794) );
  AND U5639 ( .A(n196), .B(n1795), .Z(n1793) );
  XOR U5640 ( .A(n1796), .B(n1797), .Z(n1795) );
  XOR U5641 ( .A(DB[2454]), .B(DB[2423]), .Z(n1797) );
  AND U5642 ( .A(n200), .B(n1798), .Z(n1796) );
  XOR U5643 ( .A(n1799), .B(n1800), .Z(n1798) );
  XOR U5644 ( .A(DB[2423]), .B(DB[2392]), .Z(n1800) );
  AND U5645 ( .A(n204), .B(n1801), .Z(n1799) );
  XOR U5646 ( .A(n1802), .B(n1803), .Z(n1801) );
  XOR U5647 ( .A(DB[2392]), .B(DB[2361]), .Z(n1803) );
  AND U5648 ( .A(n208), .B(n1804), .Z(n1802) );
  XOR U5649 ( .A(n1805), .B(n1806), .Z(n1804) );
  XOR U5650 ( .A(DB[2361]), .B(DB[2330]), .Z(n1806) );
  AND U5651 ( .A(n212), .B(n1807), .Z(n1805) );
  XOR U5652 ( .A(n1808), .B(n1809), .Z(n1807) );
  XOR U5653 ( .A(DB[2330]), .B(DB[2299]), .Z(n1809) );
  AND U5654 ( .A(n216), .B(n1810), .Z(n1808) );
  XOR U5655 ( .A(n1811), .B(n1812), .Z(n1810) );
  XOR U5656 ( .A(DB[2299]), .B(DB[2268]), .Z(n1812) );
  AND U5657 ( .A(n220), .B(n1813), .Z(n1811) );
  XOR U5658 ( .A(n1814), .B(n1815), .Z(n1813) );
  XOR U5659 ( .A(DB[2268]), .B(DB[2237]), .Z(n1815) );
  AND U5660 ( .A(n224), .B(n1816), .Z(n1814) );
  XOR U5661 ( .A(n1817), .B(n1818), .Z(n1816) );
  XOR U5662 ( .A(DB[2237]), .B(DB[2206]), .Z(n1818) );
  AND U5663 ( .A(n228), .B(n1819), .Z(n1817) );
  XOR U5664 ( .A(n1820), .B(n1821), .Z(n1819) );
  XOR U5665 ( .A(DB[2206]), .B(DB[2175]), .Z(n1821) );
  AND U5666 ( .A(n232), .B(n1822), .Z(n1820) );
  XOR U5667 ( .A(n1823), .B(n1824), .Z(n1822) );
  XOR U5668 ( .A(DB[2175]), .B(DB[2144]), .Z(n1824) );
  AND U5669 ( .A(n236), .B(n1825), .Z(n1823) );
  XOR U5670 ( .A(n1826), .B(n1827), .Z(n1825) );
  XOR U5671 ( .A(DB[2144]), .B(DB[2113]), .Z(n1827) );
  AND U5672 ( .A(n240), .B(n1828), .Z(n1826) );
  XOR U5673 ( .A(n1829), .B(n1830), .Z(n1828) );
  XOR U5674 ( .A(DB[2113]), .B(DB[2082]), .Z(n1830) );
  AND U5675 ( .A(n244), .B(n1831), .Z(n1829) );
  XOR U5676 ( .A(n1832), .B(n1833), .Z(n1831) );
  XOR U5677 ( .A(DB[2082]), .B(DB[2051]), .Z(n1833) );
  AND U5678 ( .A(n248), .B(n1834), .Z(n1832) );
  XOR U5679 ( .A(n1835), .B(n1836), .Z(n1834) );
  XOR U5680 ( .A(DB[2051]), .B(DB[2020]), .Z(n1836) );
  AND U5681 ( .A(n252), .B(n1837), .Z(n1835) );
  XOR U5682 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U5683 ( .A(DB[2020]), .B(DB[1989]), .Z(n1839) );
  AND U5684 ( .A(n256), .B(n1840), .Z(n1838) );
  XOR U5685 ( .A(n1841), .B(n1842), .Z(n1840) );
  XOR U5686 ( .A(DB[1989]), .B(DB[1958]), .Z(n1842) );
  AND U5687 ( .A(n260), .B(n1843), .Z(n1841) );
  XOR U5688 ( .A(n1844), .B(n1845), .Z(n1843) );
  XOR U5689 ( .A(DB[1958]), .B(DB[1927]), .Z(n1845) );
  AND U5690 ( .A(n264), .B(n1846), .Z(n1844) );
  XOR U5691 ( .A(n1847), .B(n1848), .Z(n1846) );
  XOR U5692 ( .A(DB[1927]), .B(DB[1896]), .Z(n1848) );
  AND U5693 ( .A(n268), .B(n1849), .Z(n1847) );
  XOR U5694 ( .A(n1850), .B(n1851), .Z(n1849) );
  XOR U5695 ( .A(DB[1896]), .B(DB[1865]), .Z(n1851) );
  AND U5696 ( .A(n272), .B(n1852), .Z(n1850) );
  XOR U5697 ( .A(n1853), .B(n1854), .Z(n1852) );
  XOR U5698 ( .A(DB[1865]), .B(DB[1834]), .Z(n1854) );
  AND U5699 ( .A(n276), .B(n1855), .Z(n1853) );
  XOR U5700 ( .A(n1856), .B(n1857), .Z(n1855) );
  XOR U5701 ( .A(DB[1834]), .B(DB[1803]), .Z(n1857) );
  AND U5702 ( .A(n280), .B(n1858), .Z(n1856) );
  XOR U5703 ( .A(n1859), .B(n1860), .Z(n1858) );
  XOR U5704 ( .A(DB[1803]), .B(DB[1772]), .Z(n1860) );
  AND U5705 ( .A(n284), .B(n1861), .Z(n1859) );
  XOR U5706 ( .A(n1862), .B(n1863), .Z(n1861) );
  XOR U5707 ( .A(DB[1772]), .B(DB[1741]), .Z(n1863) );
  AND U5708 ( .A(n288), .B(n1864), .Z(n1862) );
  XOR U5709 ( .A(n1865), .B(n1866), .Z(n1864) );
  XOR U5710 ( .A(DB[1741]), .B(DB[1710]), .Z(n1866) );
  AND U5711 ( .A(n292), .B(n1867), .Z(n1865) );
  XOR U5712 ( .A(n1868), .B(n1869), .Z(n1867) );
  XOR U5713 ( .A(DB[1710]), .B(DB[1679]), .Z(n1869) );
  AND U5714 ( .A(n296), .B(n1870), .Z(n1868) );
  XOR U5715 ( .A(n1871), .B(n1872), .Z(n1870) );
  XOR U5716 ( .A(DB[1679]), .B(DB[1648]), .Z(n1872) );
  AND U5717 ( .A(n300), .B(n1873), .Z(n1871) );
  XOR U5718 ( .A(n1874), .B(n1875), .Z(n1873) );
  XOR U5719 ( .A(DB[1648]), .B(DB[1617]), .Z(n1875) );
  AND U5720 ( .A(n304), .B(n1876), .Z(n1874) );
  XOR U5721 ( .A(n1877), .B(n1878), .Z(n1876) );
  XOR U5722 ( .A(DB[1617]), .B(DB[1586]), .Z(n1878) );
  AND U5723 ( .A(n308), .B(n1879), .Z(n1877) );
  XOR U5724 ( .A(n1880), .B(n1881), .Z(n1879) );
  XOR U5725 ( .A(DB[1586]), .B(DB[1555]), .Z(n1881) );
  AND U5726 ( .A(n312), .B(n1882), .Z(n1880) );
  XOR U5727 ( .A(n1883), .B(n1884), .Z(n1882) );
  XOR U5728 ( .A(DB[1555]), .B(DB[1524]), .Z(n1884) );
  AND U5729 ( .A(n316), .B(n1885), .Z(n1883) );
  XOR U5730 ( .A(n1886), .B(n1887), .Z(n1885) );
  XOR U5731 ( .A(DB[1524]), .B(DB[1493]), .Z(n1887) );
  AND U5732 ( .A(n320), .B(n1888), .Z(n1886) );
  XOR U5733 ( .A(n1889), .B(n1890), .Z(n1888) );
  XOR U5734 ( .A(DB[1493]), .B(DB[1462]), .Z(n1890) );
  AND U5735 ( .A(n324), .B(n1891), .Z(n1889) );
  XOR U5736 ( .A(n1892), .B(n1893), .Z(n1891) );
  XOR U5737 ( .A(DB[1462]), .B(DB[1431]), .Z(n1893) );
  AND U5738 ( .A(n328), .B(n1894), .Z(n1892) );
  XOR U5739 ( .A(n1895), .B(n1896), .Z(n1894) );
  XOR U5740 ( .A(DB[1431]), .B(DB[1400]), .Z(n1896) );
  AND U5741 ( .A(n332), .B(n1897), .Z(n1895) );
  XOR U5742 ( .A(n1898), .B(n1899), .Z(n1897) );
  XOR U5743 ( .A(DB[1400]), .B(DB[1369]), .Z(n1899) );
  AND U5744 ( .A(n336), .B(n1900), .Z(n1898) );
  XOR U5745 ( .A(n1901), .B(n1902), .Z(n1900) );
  XOR U5746 ( .A(DB[1369]), .B(DB[1338]), .Z(n1902) );
  AND U5747 ( .A(n340), .B(n1903), .Z(n1901) );
  XOR U5748 ( .A(n1904), .B(n1905), .Z(n1903) );
  XOR U5749 ( .A(DB[1338]), .B(DB[1307]), .Z(n1905) );
  AND U5750 ( .A(n344), .B(n1906), .Z(n1904) );
  XOR U5751 ( .A(n1907), .B(n1908), .Z(n1906) );
  XOR U5752 ( .A(DB[1307]), .B(DB[1276]), .Z(n1908) );
  AND U5753 ( .A(n348), .B(n1909), .Z(n1907) );
  XOR U5754 ( .A(n1910), .B(n1911), .Z(n1909) );
  XOR U5755 ( .A(DB[1276]), .B(DB[1245]), .Z(n1911) );
  AND U5756 ( .A(n352), .B(n1912), .Z(n1910) );
  XOR U5757 ( .A(n1913), .B(n1914), .Z(n1912) );
  XOR U5758 ( .A(DB[1245]), .B(DB[1214]), .Z(n1914) );
  AND U5759 ( .A(n356), .B(n1915), .Z(n1913) );
  XOR U5760 ( .A(n1916), .B(n1917), .Z(n1915) );
  XOR U5761 ( .A(DB[1214]), .B(DB[1183]), .Z(n1917) );
  AND U5762 ( .A(n360), .B(n1918), .Z(n1916) );
  XOR U5763 ( .A(n1919), .B(n1920), .Z(n1918) );
  XOR U5764 ( .A(DB[1183]), .B(DB[1152]), .Z(n1920) );
  AND U5765 ( .A(n364), .B(n1921), .Z(n1919) );
  XOR U5766 ( .A(n1922), .B(n1923), .Z(n1921) );
  XOR U5767 ( .A(DB[1152]), .B(DB[1121]), .Z(n1923) );
  AND U5768 ( .A(n368), .B(n1924), .Z(n1922) );
  XOR U5769 ( .A(n1925), .B(n1926), .Z(n1924) );
  XOR U5770 ( .A(DB[1121]), .B(DB[1090]), .Z(n1926) );
  AND U5771 ( .A(n372), .B(n1927), .Z(n1925) );
  XOR U5772 ( .A(n1928), .B(n1929), .Z(n1927) );
  XOR U5773 ( .A(DB[1090]), .B(DB[1059]), .Z(n1929) );
  AND U5774 ( .A(n376), .B(n1930), .Z(n1928) );
  XOR U5775 ( .A(n1931), .B(n1932), .Z(n1930) );
  XOR U5776 ( .A(DB[1059]), .B(DB[1028]), .Z(n1932) );
  AND U5777 ( .A(n380), .B(n1933), .Z(n1931) );
  XOR U5778 ( .A(n1934), .B(n1935), .Z(n1933) );
  XOR U5779 ( .A(DB[997]), .B(DB[1028]), .Z(n1935) );
  AND U5780 ( .A(n384), .B(n1936), .Z(n1934) );
  XOR U5781 ( .A(n1937), .B(n1938), .Z(n1936) );
  XOR U5782 ( .A(DB[997]), .B(DB[966]), .Z(n1938) );
  AND U5783 ( .A(n388), .B(n1939), .Z(n1937) );
  XOR U5784 ( .A(n1940), .B(n1941), .Z(n1939) );
  XOR U5785 ( .A(DB[966]), .B(DB[935]), .Z(n1941) );
  AND U5786 ( .A(n392), .B(n1942), .Z(n1940) );
  XOR U5787 ( .A(n1943), .B(n1944), .Z(n1942) );
  XOR U5788 ( .A(DB[935]), .B(DB[904]), .Z(n1944) );
  AND U5789 ( .A(n396), .B(n1945), .Z(n1943) );
  XOR U5790 ( .A(n1946), .B(n1947), .Z(n1945) );
  XOR U5791 ( .A(DB[904]), .B(DB[873]), .Z(n1947) );
  AND U5792 ( .A(n400), .B(n1948), .Z(n1946) );
  XOR U5793 ( .A(n1949), .B(n1950), .Z(n1948) );
  XOR U5794 ( .A(DB[873]), .B(DB[842]), .Z(n1950) );
  AND U5795 ( .A(n404), .B(n1951), .Z(n1949) );
  XOR U5796 ( .A(n1952), .B(n1953), .Z(n1951) );
  XOR U5797 ( .A(DB[842]), .B(DB[811]), .Z(n1953) );
  AND U5798 ( .A(n408), .B(n1954), .Z(n1952) );
  XOR U5799 ( .A(n1955), .B(n1956), .Z(n1954) );
  XOR U5800 ( .A(DB[811]), .B(DB[780]), .Z(n1956) );
  AND U5801 ( .A(n412), .B(n1957), .Z(n1955) );
  XOR U5802 ( .A(n1958), .B(n1959), .Z(n1957) );
  XOR U5803 ( .A(DB[780]), .B(DB[749]), .Z(n1959) );
  AND U5804 ( .A(n416), .B(n1960), .Z(n1958) );
  XOR U5805 ( .A(n1961), .B(n1962), .Z(n1960) );
  XOR U5806 ( .A(DB[749]), .B(DB[718]), .Z(n1962) );
  AND U5807 ( .A(n420), .B(n1963), .Z(n1961) );
  XOR U5808 ( .A(n1964), .B(n1965), .Z(n1963) );
  XOR U5809 ( .A(DB[718]), .B(DB[687]), .Z(n1965) );
  AND U5810 ( .A(n424), .B(n1966), .Z(n1964) );
  XOR U5811 ( .A(n1967), .B(n1968), .Z(n1966) );
  XOR U5812 ( .A(DB[687]), .B(DB[656]), .Z(n1968) );
  AND U5813 ( .A(n428), .B(n1969), .Z(n1967) );
  XOR U5814 ( .A(n1970), .B(n1971), .Z(n1969) );
  XOR U5815 ( .A(DB[656]), .B(DB[625]), .Z(n1971) );
  AND U5816 ( .A(n432), .B(n1972), .Z(n1970) );
  XOR U5817 ( .A(n1973), .B(n1974), .Z(n1972) );
  XOR U5818 ( .A(DB[625]), .B(DB[594]), .Z(n1974) );
  AND U5819 ( .A(n436), .B(n1975), .Z(n1973) );
  XOR U5820 ( .A(n1976), .B(n1977), .Z(n1975) );
  XOR U5821 ( .A(DB[594]), .B(DB[563]), .Z(n1977) );
  AND U5822 ( .A(n440), .B(n1978), .Z(n1976) );
  XOR U5823 ( .A(n1979), .B(n1980), .Z(n1978) );
  XOR U5824 ( .A(DB[563]), .B(DB[532]), .Z(n1980) );
  AND U5825 ( .A(n444), .B(n1981), .Z(n1979) );
  XOR U5826 ( .A(n1982), .B(n1983), .Z(n1981) );
  XOR U5827 ( .A(DB[532]), .B(DB[501]), .Z(n1983) );
  AND U5828 ( .A(n448), .B(n1984), .Z(n1982) );
  XOR U5829 ( .A(n1985), .B(n1986), .Z(n1984) );
  XOR U5830 ( .A(DB[501]), .B(DB[470]), .Z(n1986) );
  AND U5831 ( .A(n452), .B(n1987), .Z(n1985) );
  XOR U5832 ( .A(n1988), .B(n1989), .Z(n1987) );
  XOR U5833 ( .A(DB[470]), .B(DB[439]), .Z(n1989) );
  AND U5834 ( .A(n456), .B(n1990), .Z(n1988) );
  XOR U5835 ( .A(n1991), .B(n1992), .Z(n1990) );
  XOR U5836 ( .A(DB[439]), .B(DB[408]), .Z(n1992) );
  AND U5837 ( .A(n460), .B(n1993), .Z(n1991) );
  XOR U5838 ( .A(n1994), .B(n1995), .Z(n1993) );
  XOR U5839 ( .A(DB[408]), .B(DB[377]), .Z(n1995) );
  AND U5840 ( .A(n464), .B(n1996), .Z(n1994) );
  XOR U5841 ( .A(n1997), .B(n1998), .Z(n1996) );
  XOR U5842 ( .A(DB[377]), .B(DB[346]), .Z(n1998) );
  AND U5843 ( .A(n468), .B(n1999), .Z(n1997) );
  XOR U5844 ( .A(n2000), .B(n2001), .Z(n1999) );
  XOR U5845 ( .A(DB[346]), .B(DB[315]), .Z(n2001) );
  AND U5846 ( .A(n472), .B(n2002), .Z(n2000) );
  XOR U5847 ( .A(n2003), .B(n2004), .Z(n2002) );
  XOR U5848 ( .A(DB[315]), .B(DB[284]), .Z(n2004) );
  AND U5849 ( .A(n476), .B(n2005), .Z(n2003) );
  XOR U5850 ( .A(n2006), .B(n2007), .Z(n2005) );
  XOR U5851 ( .A(DB[284]), .B(DB[253]), .Z(n2007) );
  AND U5852 ( .A(n480), .B(n2008), .Z(n2006) );
  XOR U5853 ( .A(n2009), .B(n2010), .Z(n2008) );
  XOR U5854 ( .A(DB[253]), .B(DB[222]), .Z(n2010) );
  AND U5855 ( .A(n484), .B(n2011), .Z(n2009) );
  XOR U5856 ( .A(n2012), .B(n2013), .Z(n2011) );
  XOR U5857 ( .A(DB[222]), .B(DB[191]), .Z(n2013) );
  AND U5858 ( .A(n488), .B(n2014), .Z(n2012) );
  XOR U5859 ( .A(n2015), .B(n2016), .Z(n2014) );
  XOR U5860 ( .A(DB[191]), .B(DB[160]), .Z(n2016) );
  AND U5861 ( .A(n492), .B(n2017), .Z(n2015) );
  XOR U5862 ( .A(n2018), .B(n2019), .Z(n2017) );
  XOR U5863 ( .A(DB[160]), .B(DB[129]), .Z(n2019) );
  AND U5864 ( .A(n496), .B(n2020), .Z(n2018) );
  XOR U5865 ( .A(n2021), .B(n2022), .Z(n2020) );
  XOR U5866 ( .A(DB[98]), .B(DB[129]), .Z(n2022) );
  AND U5867 ( .A(n500), .B(n2023), .Z(n2021) );
  XOR U5868 ( .A(n2024), .B(n2025), .Z(n2023) );
  XOR U5869 ( .A(DB[98]), .B(DB[67]), .Z(n2025) );
  AND U5870 ( .A(n504), .B(n2026), .Z(n2024) );
  XOR U5871 ( .A(n2027), .B(n2028), .Z(n2026) );
  XOR U5872 ( .A(DB[67]), .B(DB[36]), .Z(n2028) );
  AND U5873 ( .A(n508), .B(n2029), .Z(n2027) );
  XOR U5874 ( .A(DB[5]), .B(DB[36]), .Z(n2029) );
  XOR U5875 ( .A(DB[3941]), .B(n2030), .Z(min_val_out[4]) );
  AND U5876 ( .A(n2), .B(n2031), .Z(n2030) );
  XOR U5877 ( .A(n2032), .B(n2033), .Z(n2031) );
  XOR U5878 ( .A(DB[3941]), .B(DB[3910]), .Z(n2033) );
  AND U5879 ( .A(n8), .B(n2034), .Z(n2032) );
  XOR U5880 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U5881 ( .A(DB[3910]), .B(DB[3879]), .Z(n2036) );
  AND U5882 ( .A(n12), .B(n2037), .Z(n2035) );
  XOR U5883 ( .A(n2038), .B(n2039), .Z(n2037) );
  XOR U5884 ( .A(DB[3879]), .B(DB[3848]), .Z(n2039) );
  AND U5885 ( .A(n16), .B(n2040), .Z(n2038) );
  XOR U5886 ( .A(n2041), .B(n2042), .Z(n2040) );
  XOR U5887 ( .A(DB[3848]), .B(DB[3817]), .Z(n2042) );
  AND U5888 ( .A(n20), .B(n2043), .Z(n2041) );
  XOR U5889 ( .A(n2044), .B(n2045), .Z(n2043) );
  XOR U5890 ( .A(DB[3817]), .B(DB[3786]), .Z(n2045) );
  AND U5891 ( .A(n24), .B(n2046), .Z(n2044) );
  XOR U5892 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U5893 ( .A(DB[3786]), .B(DB[3755]), .Z(n2048) );
  AND U5894 ( .A(n28), .B(n2049), .Z(n2047) );
  XOR U5895 ( .A(n2050), .B(n2051), .Z(n2049) );
  XOR U5896 ( .A(DB[3755]), .B(DB[3724]), .Z(n2051) );
  AND U5897 ( .A(n32), .B(n2052), .Z(n2050) );
  XOR U5898 ( .A(n2053), .B(n2054), .Z(n2052) );
  XOR U5899 ( .A(DB[3724]), .B(DB[3693]), .Z(n2054) );
  AND U5900 ( .A(n36), .B(n2055), .Z(n2053) );
  XOR U5901 ( .A(n2056), .B(n2057), .Z(n2055) );
  XOR U5902 ( .A(DB[3693]), .B(DB[3662]), .Z(n2057) );
  AND U5903 ( .A(n40), .B(n2058), .Z(n2056) );
  XOR U5904 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U5905 ( .A(DB[3662]), .B(DB[3631]), .Z(n2060) );
  AND U5906 ( .A(n44), .B(n2061), .Z(n2059) );
  XOR U5907 ( .A(n2062), .B(n2063), .Z(n2061) );
  XOR U5908 ( .A(DB[3631]), .B(DB[3600]), .Z(n2063) );
  AND U5909 ( .A(n48), .B(n2064), .Z(n2062) );
  XOR U5910 ( .A(n2065), .B(n2066), .Z(n2064) );
  XOR U5911 ( .A(DB[3600]), .B(DB[3569]), .Z(n2066) );
  AND U5912 ( .A(n52), .B(n2067), .Z(n2065) );
  XOR U5913 ( .A(n2068), .B(n2069), .Z(n2067) );
  XOR U5914 ( .A(DB[3569]), .B(DB[3538]), .Z(n2069) );
  AND U5915 ( .A(n56), .B(n2070), .Z(n2068) );
  XOR U5916 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U5917 ( .A(DB[3538]), .B(DB[3507]), .Z(n2072) );
  AND U5918 ( .A(n60), .B(n2073), .Z(n2071) );
  XOR U5919 ( .A(n2074), .B(n2075), .Z(n2073) );
  XOR U5920 ( .A(DB[3507]), .B(DB[3476]), .Z(n2075) );
  AND U5921 ( .A(n64), .B(n2076), .Z(n2074) );
  XOR U5922 ( .A(n2077), .B(n2078), .Z(n2076) );
  XOR U5923 ( .A(DB[3476]), .B(DB[3445]), .Z(n2078) );
  AND U5924 ( .A(n68), .B(n2079), .Z(n2077) );
  XOR U5925 ( .A(n2080), .B(n2081), .Z(n2079) );
  XOR U5926 ( .A(DB[3445]), .B(DB[3414]), .Z(n2081) );
  AND U5927 ( .A(n72), .B(n2082), .Z(n2080) );
  XOR U5928 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U5929 ( .A(DB[3414]), .B(DB[3383]), .Z(n2084) );
  AND U5930 ( .A(n76), .B(n2085), .Z(n2083) );
  XOR U5931 ( .A(n2086), .B(n2087), .Z(n2085) );
  XOR U5932 ( .A(DB[3383]), .B(DB[3352]), .Z(n2087) );
  AND U5933 ( .A(n80), .B(n2088), .Z(n2086) );
  XOR U5934 ( .A(n2089), .B(n2090), .Z(n2088) );
  XOR U5935 ( .A(DB[3352]), .B(DB[3321]), .Z(n2090) );
  AND U5936 ( .A(n84), .B(n2091), .Z(n2089) );
  XOR U5937 ( .A(n2092), .B(n2093), .Z(n2091) );
  XOR U5938 ( .A(DB[3321]), .B(DB[3290]), .Z(n2093) );
  AND U5939 ( .A(n88), .B(n2094), .Z(n2092) );
  XOR U5940 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U5941 ( .A(DB[3290]), .B(DB[3259]), .Z(n2096) );
  AND U5942 ( .A(n92), .B(n2097), .Z(n2095) );
  XOR U5943 ( .A(n2098), .B(n2099), .Z(n2097) );
  XOR U5944 ( .A(DB[3259]), .B(DB[3228]), .Z(n2099) );
  AND U5945 ( .A(n96), .B(n2100), .Z(n2098) );
  XOR U5946 ( .A(n2101), .B(n2102), .Z(n2100) );
  XOR U5947 ( .A(DB[3228]), .B(DB[3197]), .Z(n2102) );
  AND U5948 ( .A(n100), .B(n2103), .Z(n2101) );
  XOR U5949 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR U5950 ( .A(DB[3197]), .B(DB[3166]), .Z(n2105) );
  AND U5951 ( .A(n104), .B(n2106), .Z(n2104) );
  XOR U5952 ( .A(n2107), .B(n2108), .Z(n2106) );
  XOR U5953 ( .A(DB[3166]), .B(DB[3135]), .Z(n2108) );
  AND U5954 ( .A(n108), .B(n2109), .Z(n2107) );
  XOR U5955 ( .A(n2110), .B(n2111), .Z(n2109) );
  XOR U5956 ( .A(DB[3135]), .B(DB[3104]), .Z(n2111) );
  AND U5957 ( .A(n112), .B(n2112), .Z(n2110) );
  XOR U5958 ( .A(n2113), .B(n2114), .Z(n2112) );
  XOR U5959 ( .A(DB[3104]), .B(DB[3073]), .Z(n2114) );
  AND U5960 ( .A(n116), .B(n2115), .Z(n2113) );
  XOR U5961 ( .A(n2116), .B(n2117), .Z(n2115) );
  XOR U5962 ( .A(DB[3073]), .B(DB[3042]), .Z(n2117) );
  AND U5963 ( .A(n120), .B(n2118), .Z(n2116) );
  XOR U5964 ( .A(n2119), .B(n2120), .Z(n2118) );
  XOR U5965 ( .A(DB[3042]), .B(DB[3011]), .Z(n2120) );
  AND U5966 ( .A(n124), .B(n2121), .Z(n2119) );
  XOR U5967 ( .A(n2122), .B(n2123), .Z(n2121) );
  XOR U5968 ( .A(DB[3011]), .B(DB[2980]), .Z(n2123) );
  AND U5969 ( .A(n128), .B(n2124), .Z(n2122) );
  XOR U5970 ( .A(n2125), .B(n2126), .Z(n2124) );
  XOR U5971 ( .A(DB[2980]), .B(DB[2949]), .Z(n2126) );
  AND U5972 ( .A(n132), .B(n2127), .Z(n2125) );
  XOR U5973 ( .A(n2128), .B(n2129), .Z(n2127) );
  XOR U5974 ( .A(DB[2949]), .B(DB[2918]), .Z(n2129) );
  AND U5975 ( .A(n136), .B(n2130), .Z(n2128) );
  XOR U5976 ( .A(n2131), .B(n2132), .Z(n2130) );
  XOR U5977 ( .A(DB[2918]), .B(DB[2887]), .Z(n2132) );
  AND U5978 ( .A(n140), .B(n2133), .Z(n2131) );
  XOR U5979 ( .A(n2134), .B(n2135), .Z(n2133) );
  XOR U5980 ( .A(DB[2887]), .B(DB[2856]), .Z(n2135) );
  AND U5981 ( .A(n144), .B(n2136), .Z(n2134) );
  XOR U5982 ( .A(n2137), .B(n2138), .Z(n2136) );
  XOR U5983 ( .A(DB[2856]), .B(DB[2825]), .Z(n2138) );
  AND U5984 ( .A(n148), .B(n2139), .Z(n2137) );
  XOR U5985 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U5986 ( .A(DB[2825]), .B(DB[2794]), .Z(n2141) );
  AND U5987 ( .A(n152), .B(n2142), .Z(n2140) );
  XOR U5988 ( .A(n2143), .B(n2144), .Z(n2142) );
  XOR U5989 ( .A(DB[2794]), .B(DB[2763]), .Z(n2144) );
  AND U5990 ( .A(n156), .B(n2145), .Z(n2143) );
  XOR U5991 ( .A(n2146), .B(n2147), .Z(n2145) );
  XOR U5992 ( .A(DB[2763]), .B(DB[2732]), .Z(n2147) );
  AND U5993 ( .A(n160), .B(n2148), .Z(n2146) );
  XOR U5994 ( .A(n2149), .B(n2150), .Z(n2148) );
  XOR U5995 ( .A(DB[2732]), .B(DB[2701]), .Z(n2150) );
  AND U5996 ( .A(n164), .B(n2151), .Z(n2149) );
  XOR U5997 ( .A(n2152), .B(n2153), .Z(n2151) );
  XOR U5998 ( .A(DB[2701]), .B(DB[2670]), .Z(n2153) );
  AND U5999 ( .A(n168), .B(n2154), .Z(n2152) );
  XOR U6000 ( .A(n2155), .B(n2156), .Z(n2154) );
  XOR U6001 ( .A(DB[2670]), .B(DB[2639]), .Z(n2156) );
  AND U6002 ( .A(n172), .B(n2157), .Z(n2155) );
  XOR U6003 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U6004 ( .A(DB[2639]), .B(DB[2608]), .Z(n2159) );
  AND U6005 ( .A(n176), .B(n2160), .Z(n2158) );
  XOR U6006 ( .A(n2161), .B(n2162), .Z(n2160) );
  XOR U6007 ( .A(DB[2608]), .B(DB[2577]), .Z(n2162) );
  AND U6008 ( .A(n180), .B(n2163), .Z(n2161) );
  XOR U6009 ( .A(n2164), .B(n2165), .Z(n2163) );
  XOR U6010 ( .A(DB[2577]), .B(DB[2546]), .Z(n2165) );
  AND U6011 ( .A(n184), .B(n2166), .Z(n2164) );
  XOR U6012 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U6013 ( .A(DB[2546]), .B(DB[2515]), .Z(n2168) );
  AND U6014 ( .A(n188), .B(n2169), .Z(n2167) );
  XOR U6015 ( .A(n2170), .B(n2171), .Z(n2169) );
  XOR U6016 ( .A(DB[2515]), .B(DB[2484]), .Z(n2171) );
  AND U6017 ( .A(n192), .B(n2172), .Z(n2170) );
  XOR U6018 ( .A(n2173), .B(n2174), .Z(n2172) );
  XOR U6019 ( .A(DB[2484]), .B(DB[2453]), .Z(n2174) );
  AND U6020 ( .A(n196), .B(n2175), .Z(n2173) );
  XOR U6021 ( .A(n2176), .B(n2177), .Z(n2175) );
  XOR U6022 ( .A(DB[2453]), .B(DB[2422]), .Z(n2177) );
  AND U6023 ( .A(n200), .B(n2178), .Z(n2176) );
  XOR U6024 ( .A(n2179), .B(n2180), .Z(n2178) );
  XOR U6025 ( .A(DB[2422]), .B(DB[2391]), .Z(n2180) );
  AND U6026 ( .A(n204), .B(n2181), .Z(n2179) );
  XOR U6027 ( .A(n2182), .B(n2183), .Z(n2181) );
  XOR U6028 ( .A(DB[2391]), .B(DB[2360]), .Z(n2183) );
  AND U6029 ( .A(n208), .B(n2184), .Z(n2182) );
  XOR U6030 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U6031 ( .A(DB[2360]), .B(DB[2329]), .Z(n2186) );
  AND U6032 ( .A(n212), .B(n2187), .Z(n2185) );
  XOR U6033 ( .A(n2188), .B(n2189), .Z(n2187) );
  XOR U6034 ( .A(DB[2329]), .B(DB[2298]), .Z(n2189) );
  AND U6035 ( .A(n216), .B(n2190), .Z(n2188) );
  XOR U6036 ( .A(n2191), .B(n2192), .Z(n2190) );
  XOR U6037 ( .A(DB[2298]), .B(DB[2267]), .Z(n2192) );
  AND U6038 ( .A(n220), .B(n2193), .Z(n2191) );
  XOR U6039 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U6040 ( .A(DB[2267]), .B(DB[2236]), .Z(n2195) );
  AND U6041 ( .A(n224), .B(n2196), .Z(n2194) );
  XOR U6042 ( .A(n2197), .B(n2198), .Z(n2196) );
  XOR U6043 ( .A(DB[2236]), .B(DB[2205]), .Z(n2198) );
  AND U6044 ( .A(n228), .B(n2199), .Z(n2197) );
  XOR U6045 ( .A(n2200), .B(n2201), .Z(n2199) );
  XOR U6046 ( .A(DB[2205]), .B(DB[2174]), .Z(n2201) );
  AND U6047 ( .A(n232), .B(n2202), .Z(n2200) );
  XOR U6048 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR U6049 ( .A(DB[2174]), .B(DB[2143]), .Z(n2204) );
  AND U6050 ( .A(n236), .B(n2205), .Z(n2203) );
  XOR U6051 ( .A(n2206), .B(n2207), .Z(n2205) );
  XOR U6052 ( .A(DB[2143]), .B(DB[2112]), .Z(n2207) );
  AND U6053 ( .A(n240), .B(n2208), .Z(n2206) );
  XOR U6054 ( .A(n2209), .B(n2210), .Z(n2208) );
  XOR U6055 ( .A(DB[2112]), .B(DB[2081]), .Z(n2210) );
  AND U6056 ( .A(n244), .B(n2211), .Z(n2209) );
  XOR U6057 ( .A(n2212), .B(n2213), .Z(n2211) );
  XOR U6058 ( .A(DB[2081]), .B(DB[2050]), .Z(n2213) );
  AND U6059 ( .A(n248), .B(n2214), .Z(n2212) );
  XOR U6060 ( .A(n2215), .B(n2216), .Z(n2214) );
  XOR U6061 ( .A(DB[2050]), .B(DB[2019]), .Z(n2216) );
  AND U6062 ( .A(n252), .B(n2217), .Z(n2215) );
  XOR U6063 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U6064 ( .A(DB[2019]), .B(DB[1988]), .Z(n2219) );
  AND U6065 ( .A(n256), .B(n2220), .Z(n2218) );
  XOR U6066 ( .A(n2221), .B(n2222), .Z(n2220) );
  XOR U6067 ( .A(DB[1988]), .B(DB[1957]), .Z(n2222) );
  AND U6068 ( .A(n260), .B(n2223), .Z(n2221) );
  XOR U6069 ( .A(n2224), .B(n2225), .Z(n2223) );
  XOR U6070 ( .A(DB[1957]), .B(DB[1926]), .Z(n2225) );
  AND U6071 ( .A(n264), .B(n2226), .Z(n2224) );
  XOR U6072 ( .A(n2227), .B(n2228), .Z(n2226) );
  XOR U6073 ( .A(DB[1926]), .B(DB[1895]), .Z(n2228) );
  AND U6074 ( .A(n268), .B(n2229), .Z(n2227) );
  XOR U6075 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U6076 ( .A(DB[1895]), .B(DB[1864]), .Z(n2231) );
  AND U6077 ( .A(n272), .B(n2232), .Z(n2230) );
  XOR U6078 ( .A(n2233), .B(n2234), .Z(n2232) );
  XOR U6079 ( .A(DB[1864]), .B(DB[1833]), .Z(n2234) );
  AND U6080 ( .A(n276), .B(n2235), .Z(n2233) );
  XOR U6081 ( .A(n2236), .B(n2237), .Z(n2235) );
  XOR U6082 ( .A(DB[1833]), .B(DB[1802]), .Z(n2237) );
  AND U6083 ( .A(n280), .B(n2238), .Z(n2236) );
  XOR U6084 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U6085 ( .A(DB[1802]), .B(DB[1771]), .Z(n2240) );
  AND U6086 ( .A(n284), .B(n2241), .Z(n2239) );
  XOR U6087 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U6088 ( .A(DB[1771]), .B(DB[1740]), .Z(n2243) );
  AND U6089 ( .A(n288), .B(n2244), .Z(n2242) );
  XOR U6090 ( .A(n2245), .B(n2246), .Z(n2244) );
  XOR U6091 ( .A(DB[1740]), .B(DB[1709]), .Z(n2246) );
  AND U6092 ( .A(n292), .B(n2247), .Z(n2245) );
  XOR U6093 ( .A(n2248), .B(n2249), .Z(n2247) );
  XOR U6094 ( .A(DB[1709]), .B(DB[1678]), .Z(n2249) );
  AND U6095 ( .A(n296), .B(n2250), .Z(n2248) );
  XOR U6096 ( .A(n2251), .B(n2252), .Z(n2250) );
  XOR U6097 ( .A(DB[1678]), .B(DB[1647]), .Z(n2252) );
  AND U6098 ( .A(n300), .B(n2253), .Z(n2251) );
  XOR U6099 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR U6100 ( .A(DB[1647]), .B(DB[1616]), .Z(n2255) );
  AND U6101 ( .A(n304), .B(n2256), .Z(n2254) );
  XOR U6102 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U6103 ( .A(DB[1616]), .B(DB[1585]), .Z(n2258) );
  AND U6104 ( .A(n308), .B(n2259), .Z(n2257) );
  XOR U6105 ( .A(n2260), .B(n2261), .Z(n2259) );
  XOR U6106 ( .A(DB[1585]), .B(DB[1554]), .Z(n2261) );
  AND U6107 ( .A(n312), .B(n2262), .Z(n2260) );
  XOR U6108 ( .A(n2263), .B(n2264), .Z(n2262) );
  XOR U6109 ( .A(DB[1554]), .B(DB[1523]), .Z(n2264) );
  AND U6110 ( .A(n316), .B(n2265), .Z(n2263) );
  XOR U6111 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U6112 ( .A(DB[1523]), .B(DB[1492]), .Z(n2267) );
  AND U6113 ( .A(n320), .B(n2268), .Z(n2266) );
  XOR U6114 ( .A(n2269), .B(n2270), .Z(n2268) );
  XOR U6115 ( .A(DB[1492]), .B(DB[1461]), .Z(n2270) );
  AND U6116 ( .A(n324), .B(n2271), .Z(n2269) );
  XOR U6117 ( .A(n2272), .B(n2273), .Z(n2271) );
  XOR U6118 ( .A(DB[1461]), .B(DB[1430]), .Z(n2273) );
  AND U6119 ( .A(n328), .B(n2274), .Z(n2272) );
  XOR U6120 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U6121 ( .A(DB[1430]), .B(DB[1399]), .Z(n2276) );
  AND U6122 ( .A(n332), .B(n2277), .Z(n2275) );
  XOR U6123 ( .A(n2278), .B(n2279), .Z(n2277) );
  XOR U6124 ( .A(DB[1399]), .B(DB[1368]), .Z(n2279) );
  AND U6125 ( .A(n336), .B(n2280), .Z(n2278) );
  XOR U6126 ( .A(n2281), .B(n2282), .Z(n2280) );
  XOR U6127 ( .A(DB[1368]), .B(DB[1337]), .Z(n2282) );
  AND U6128 ( .A(n340), .B(n2283), .Z(n2281) );
  XOR U6129 ( .A(n2284), .B(n2285), .Z(n2283) );
  XOR U6130 ( .A(DB[1337]), .B(DB[1306]), .Z(n2285) );
  AND U6131 ( .A(n344), .B(n2286), .Z(n2284) );
  XOR U6132 ( .A(n2287), .B(n2288), .Z(n2286) );
  XOR U6133 ( .A(DB[1306]), .B(DB[1275]), .Z(n2288) );
  AND U6134 ( .A(n348), .B(n2289), .Z(n2287) );
  XOR U6135 ( .A(n2290), .B(n2291), .Z(n2289) );
  XOR U6136 ( .A(DB[1275]), .B(DB[1244]), .Z(n2291) );
  AND U6137 ( .A(n352), .B(n2292), .Z(n2290) );
  XOR U6138 ( .A(n2293), .B(n2294), .Z(n2292) );
  XOR U6139 ( .A(DB[1244]), .B(DB[1213]), .Z(n2294) );
  AND U6140 ( .A(n356), .B(n2295), .Z(n2293) );
  XOR U6141 ( .A(n2296), .B(n2297), .Z(n2295) );
  XOR U6142 ( .A(DB[1213]), .B(DB[1182]), .Z(n2297) );
  AND U6143 ( .A(n360), .B(n2298), .Z(n2296) );
  XOR U6144 ( .A(n2299), .B(n2300), .Z(n2298) );
  XOR U6145 ( .A(DB[1182]), .B(DB[1151]), .Z(n2300) );
  AND U6146 ( .A(n364), .B(n2301), .Z(n2299) );
  XOR U6147 ( .A(n2302), .B(n2303), .Z(n2301) );
  XOR U6148 ( .A(DB[1151]), .B(DB[1120]), .Z(n2303) );
  AND U6149 ( .A(n368), .B(n2304), .Z(n2302) );
  XOR U6150 ( .A(n2305), .B(n2306), .Z(n2304) );
  XOR U6151 ( .A(DB[1120]), .B(DB[1089]), .Z(n2306) );
  AND U6152 ( .A(n372), .B(n2307), .Z(n2305) );
  XOR U6153 ( .A(n2308), .B(n2309), .Z(n2307) );
  XOR U6154 ( .A(DB[1089]), .B(DB[1058]), .Z(n2309) );
  AND U6155 ( .A(n376), .B(n2310), .Z(n2308) );
  XOR U6156 ( .A(n2311), .B(n2312), .Z(n2310) );
  XOR U6157 ( .A(DB[1058]), .B(DB[1027]), .Z(n2312) );
  AND U6158 ( .A(n380), .B(n2313), .Z(n2311) );
  XOR U6159 ( .A(n2314), .B(n2315), .Z(n2313) );
  XOR U6160 ( .A(DB[996]), .B(DB[1027]), .Z(n2315) );
  AND U6161 ( .A(n384), .B(n2316), .Z(n2314) );
  XOR U6162 ( .A(n2317), .B(n2318), .Z(n2316) );
  XOR U6163 ( .A(DB[996]), .B(DB[965]), .Z(n2318) );
  AND U6164 ( .A(n388), .B(n2319), .Z(n2317) );
  XOR U6165 ( .A(n2320), .B(n2321), .Z(n2319) );
  XOR U6166 ( .A(DB[965]), .B(DB[934]), .Z(n2321) );
  AND U6167 ( .A(n392), .B(n2322), .Z(n2320) );
  XOR U6168 ( .A(n2323), .B(n2324), .Z(n2322) );
  XOR U6169 ( .A(DB[934]), .B(DB[903]), .Z(n2324) );
  AND U6170 ( .A(n396), .B(n2325), .Z(n2323) );
  XOR U6171 ( .A(n2326), .B(n2327), .Z(n2325) );
  XOR U6172 ( .A(DB[903]), .B(DB[872]), .Z(n2327) );
  AND U6173 ( .A(n400), .B(n2328), .Z(n2326) );
  XOR U6174 ( .A(n2329), .B(n2330), .Z(n2328) );
  XOR U6175 ( .A(DB[872]), .B(DB[841]), .Z(n2330) );
  AND U6176 ( .A(n404), .B(n2331), .Z(n2329) );
  XOR U6177 ( .A(n2332), .B(n2333), .Z(n2331) );
  XOR U6178 ( .A(DB[841]), .B(DB[810]), .Z(n2333) );
  AND U6179 ( .A(n408), .B(n2334), .Z(n2332) );
  XOR U6180 ( .A(n2335), .B(n2336), .Z(n2334) );
  XOR U6181 ( .A(DB[810]), .B(DB[779]), .Z(n2336) );
  AND U6182 ( .A(n412), .B(n2337), .Z(n2335) );
  XOR U6183 ( .A(n2338), .B(n2339), .Z(n2337) );
  XOR U6184 ( .A(DB[779]), .B(DB[748]), .Z(n2339) );
  AND U6185 ( .A(n416), .B(n2340), .Z(n2338) );
  XOR U6186 ( .A(n2341), .B(n2342), .Z(n2340) );
  XOR U6187 ( .A(DB[748]), .B(DB[717]), .Z(n2342) );
  AND U6188 ( .A(n420), .B(n2343), .Z(n2341) );
  XOR U6189 ( .A(n2344), .B(n2345), .Z(n2343) );
  XOR U6190 ( .A(DB[717]), .B(DB[686]), .Z(n2345) );
  AND U6191 ( .A(n424), .B(n2346), .Z(n2344) );
  XOR U6192 ( .A(n2347), .B(n2348), .Z(n2346) );
  XOR U6193 ( .A(DB[686]), .B(DB[655]), .Z(n2348) );
  AND U6194 ( .A(n428), .B(n2349), .Z(n2347) );
  XOR U6195 ( .A(n2350), .B(n2351), .Z(n2349) );
  XOR U6196 ( .A(DB[655]), .B(DB[624]), .Z(n2351) );
  AND U6197 ( .A(n432), .B(n2352), .Z(n2350) );
  XOR U6198 ( .A(n2353), .B(n2354), .Z(n2352) );
  XOR U6199 ( .A(DB[624]), .B(DB[593]), .Z(n2354) );
  AND U6200 ( .A(n436), .B(n2355), .Z(n2353) );
  XOR U6201 ( .A(n2356), .B(n2357), .Z(n2355) );
  XOR U6202 ( .A(DB[593]), .B(DB[562]), .Z(n2357) );
  AND U6203 ( .A(n440), .B(n2358), .Z(n2356) );
  XOR U6204 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U6205 ( .A(DB[562]), .B(DB[531]), .Z(n2360) );
  AND U6206 ( .A(n444), .B(n2361), .Z(n2359) );
  XOR U6207 ( .A(n2362), .B(n2363), .Z(n2361) );
  XOR U6208 ( .A(DB[531]), .B(DB[500]), .Z(n2363) );
  AND U6209 ( .A(n448), .B(n2364), .Z(n2362) );
  XOR U6210 ( .A(n2365), .B(n2366), .Z(n2364) );
  XOR U6211 ( .A(DB[500]), .B(DB[469]), .Z(n2366) );
  AND U6212 ( .A(n452), .B(n2367), .Z(n2365) );
  XOR U6213 ( .A(n2368), .B(n2369), .Z(n2367) );
  XOR U6214 ( .A(DB[469]), .B(DB[438]), .Z(n2369) );
  AND U6215 ( .A(n456), .B(n2370), .Z(n2368) );
  XOR U6216 ( .A(n2371), .B(n2372), .Z(n2370) );
  XOR U6217 ( .A(DB[438]), .B(DB[407]), .Z(n2372) );
  AND U6218 ( .A(n460), .B(n2373), .Z(n2371) );
  XOR U6219 ( .A(n2374), .B(n2375), .Z(n2373) );
  XOR U6220 ( .A(DB[407]), .B(DB[376]), .Z(n2375) );
  AND U6221 ( .A(n464), .B(n2376), .Z(n2374) );
  XOR U6222 ( .A(n2377), .B(n2378), .Z(n2376) );
  XOR U6223 ( .A(DB[376]), .B(DB[345]), .Z(n2378) );
  AND U6224 ( .A(n468), .B(n2379), .Z(n2377) );
  XOR U6225 ( .A(n2380), .B(n2381), .Z(n2379) );
  XOR U6226 ( .A(DB[345]), .B(DB[314]), .Z(n2381) );
  AND U6227 ( .A(n472), .B(n2382), .Z(n2380) );
  XOR U6228 ( .A(n2383), .B(n2384), .Z(n2382) );
  XOR U6229 ( .A(DB[314]), .B(DB[283]), .Z(n2384) );
  AND U6230 ( .A(n476), .B(n2385), .Z(n2383) );
  XOR U6231 ( .A(n2386), .B(n2387), .Z(n2385) );
  XOR U6232 ( .A(DB[283]), .B(DB[252]), .Z(n2387) );
  AND U6233 ( .A(n480), .B(n2388), .Z(n2386) );
  XOR U6234 ( .A(n2389), .B(n2390), .Z(n2388) );
  XOR U6235 ( .A(DB[252]), .B(DB[221]), .Z(n2390) );
  AND U6236 ( .A(n484), .B(n2391), .Z(n2389) );
  XOR U6237 ( .A(n2392), .B(n2393), .Z(n2391) );
  XOR U6238 ( .A(DB[221]), .B(DB[190]), .Z(n2393) );
  AND U6239 ( .A(n488), .B(n2394), .Z(n2392) );
  XOR U6240 ( .A(n2395), .B(n2396), .Z(n2394) );
  XOR U6241 ( .A(DB[190]), .B(DB[159]), .Z(n2396) );
  AND U6242 ( .A(n492), .B(n2397), .Z(n2395) );
  XOR U6243 ( .A(n2398), .B(n2399), .Z(n2397) );
  XOR U6244 ( .A(DB[159]), .B(DB[128]), .Z(n2399) );
  AND U6245 ( .A(n496), .B(n2400), .Z(n2398) );
  XOR U6246 ( .A(n2401), .B(n2402), .Z(n2400) );
  XOR U6247 ( .A(DB[97]), .B(DB[128]), .Z(n2402) );
  AND U6248 ( .A(n500), .B(n2403), .Z(n2401) );
  XOR U6249 ( .A(n2404), .B(n2405), .Z(n2403) );
  XOR U6250 ( .A(DB[97]), .B(DB[66]), .Z(n2405) );
  AND U6251 ( .A(n504), .B(n2406), .Z(n2404) );
  XOR U6252 ( .A(n2407), .B(n2408), .Z(n2406) );
  XOR U6253 ( .A(DB[66]), .B(DB[35]), .Z(n2408) );
  AND U6254 ( .A(n508), .B(n2409), .Z(n2407) );
  XOR U6255 ( .A(DB[4]), .B(DB[35]), .Z(n2409) );
  XOR U6256 ( .A(DB[3940]), .B(n2410), .Z(min_val_out[3]) );
  AND U6257 ( .A(n2), .B(n2411), .Z(n2410) );
  XOR U6258 ( .A(n2412), .B(n2413), .Z(n2411) );
  XOR U6259 ( .A(DB[3940]), .B(DB[3909]), .Z(n2413) );
  AND U6260 ( .A(n8), .B(n2414), .Z(n2412) );
  XOR U6261 ( .A(n2415), .B(n2416), .Z(n2414) );
  XOR U6262 ( .A(DB[3909]), .B(DB[3878]), .Z(n2416) );
  AND U6263 ( .A(n12), .B(n2417), .Z(n2415) );
  XOR U6264 ( .A(n2418), .B(n2419), .Z(n2417) );
  XOR U6265 ( .A(DB[3878]), .B(DB[3847]), .Z(n2419) );
  AND U6266 ( .A(n16), .B(n2420), .Z(n2418) );
  XOR U6267 ( .A(n2421), .B(n2422), .Z(n2420) );
  XOR U6268 ( .A(DB[3847]), .B(DB[3816]), .Z(n2422) );
  AND U6269 ( .A(n20), .B(n2423), .Z(n2421) );
  XOR U6270 ( .A(n2424), .B(n2425), .Z(n2423) );
  XOR U6271 ( .A(DB[3816]), .B(DB[3785]), .Z(n2425) );
  AND U6272 ( .A(n24), .B(n2426), .Z(n2424) );
  XOR U6273 ( .A(n2427), .B(n2428), .Z(n2426) );
  XOR U6274 ( .A(DB[3785]), .B(DB[3754]), .Z(n2428) );
  AND U6275 ( .A(n28), .B(n2429), .Z(n2427) );
  XOR U6276 ( .A(n2430), .B(n2431), .Z(n2429) );
  XOR U6277 ( .A(DB[3754]), .B(DB[3723]), .Z(n2431) );
  AND U6278 ( .A(n32), .B(n2432), .Z(n2430) );
  XOR U6279 ( .A(n2433), .B(n2434), .Z(n2432) );
  XOR U6280 ( .A(DB[3723]), .B(DB[3692]), .Z(n2434) );
  AND U6281 ( .A(n36), .B(n2435), .Z(n2433) );
  XOR U6282 ( .A(n2436), .B(n2437), .Z(n2435) );
  XOR U6283 ( .A(DB[3692]), .B(DB[3661]), .Z(n2437) );
  AND U6284 ( .A(n40), .B(n2438), .Z(n2436) );
  XOR U6285 ( .A(n2439), .B(n2440), .Z(n2438) );
  XOR U6286 ( .A(DB[3661]), .B(DB[3630]), .Z(n2440) );
  AND U6287 ( .A(n44), .B(n2441), .Z(n2439) );
  XOR U6288 ( .A(n2442), .B(n2443), .Z(n2441) );
  XOR U6289 ( .A(DB[3630]), .B(DB[3599]), .Z(n2443) );
  AND U6290 ( .A(n48), .B(n2444), .Z(n2442) );
  XOR U6291 ( .A(n2445), .B(n2446), .Z(n2444) );
  XOR U6292 ( .A(DB[3599]), .B(DB[3568]), .Z(n2446) );
  AND U6293 ( .A(n52), .B(n2447), .Z(n2445) );
  XOR U6294 ( .A(n2448), .B(n2449), .Z(n2447) );
  XOR U6295 ( .A(DB[3568]), .B(DB[3537]), .Z(n2449) );
  AND U6296 ( .A(n56), .B(n2450), .Z(n2448) );
  XOR U6297 ( .A(n2451), .B(n2452), .Z(n2450) );
  XOR U6298 ( .A(DB[3537]), .B(DB[3506]), .Z(n2452) );
  AND U6299 ( .A(n60), .B(n2453), .Z(n2451) );
  XOR U6300 ( .A(n2454), .B(n2455), .Z(n2453) );
  XOR U6301 ( .A(DB[3506]), .B(DB[3475]), .Z(n2455) );
  AND U6302 ( .A(n64), .B(n2456), .Z(n2454) );
  XOR U6303 ( .A(n2457), .B(n2458), .Z(n2456) );
  XOR U6304 ( .A(DB[3475]), .B(DB[3444]), .Z(n2458) );
  AND U6305 ( .A(n68), .B(n2459), .Z(n2457) );
  XOR U6306 ( .A(n2460), .B(n2461), .Z(n2459) );
  XOR U6307 ( .A(DB[3444]), .B(DB[3413]), .Z(n2461) );
  AND U6308 ( .A(n72), .B(n2462), .Z(n2460) );
  XOR U6309 ( .A(n2463), .B(n2464), .Z(n2462) );
  XOR U6310 ( .A(DB[3413]), .B(DB[3382]), .Z(n2464) );
  AND U6311 ( .A(n76), .B(n2465), .Z(n2463) );
  XOR U6312 ( .A(n2466), .B(n2467), .Z(n2465) );
  XOR U6313 ( .A(DB[3382]), .B(DB[3351]), .Z(n2467) );
  AND U6314 ( .A(n80), .B(n2468), .Z(n2466) );
  XOR U6315 ( .A(n2469), .B(n2470), .Z(n2468) );
  XOR U6316 ( .A(DB[3351]), .B(DB[3320]), .Z(n2470) );
  AND U6317 ( .A(n84), .B(n2471), .Z(n2469) );
  XOR U6318 ( .A(n2472), .B(n2473), .Z(n2471) );
  XOR U6319 ( .A(DB[3320]), .B(DB[3289]), .Z(n2473) );
  AND U6320 ( .A(n88), .B(n2474), .Z(n2472) );
  XOR U6321 ( .A(n2475), .B(n2476), .Z(n2474) );
  XOR U6322 ( .A(DB[3289]), .B(DB[3258]), .Z(n2476) );
  AND U6323 ( .A(n92), .B(n2477), .Z(n2475) );
  XOR U6324 ( .A(n2478), .B(n2479), .Z(n2477) );
  XOR U6325 ( .A(DB[3258]), .B(DB[3227]), .Z(n2479) );
  AND U6326 ( .A(n96), .B(n2480), .Z(n2478) );
  XOR U6327 ( .A(n2481), .B(n2482), .Z(n2480) );
  XOR U6328 ( .A(DB[3227]), .B(DB[3196]), .Z(n2482) );
  AND U6329 ( .A(n100), .B(n2483), .Z(n2481) );
  XOR U6330 ( .A(n2484), .B(n2485), .Z(n2483) );
  XOR U6331 ( .A(DB[3196]), .B(DB[3165]), .Z(n2485) );
  AND U6332 ( .A(n104), .B(n2486), .Z(n2484) );
  XOR U6333 ( .A(n2487), .B(n2488), .Z(n2486) );
  XOR U6334 ( .A(DB[3165]), .B(DB[3134]), .Z(n2488) );
  AND U6335 ( .A(n108), .B(n2489), .Z(n2487) );
  XOR U6336 ( .A(n2490), .B(n2491), .Z(n2489) );
  XOR U6337 ( .A(DB[3134]), .B(DB[3103]), .Z(n2491) );
  AND U6338 ( .A(n112), .B(n2492), .Z(n2490) );
  XOR U6339 ( .A(n2493), .B(n2494), .Z(n2492) );
  XOR U6340 ( .A(DB[3103]), .B(DB[3072]), .Z(n2494) );
  AND U6341 ( .A(n116), .B(n2495), .Z(n2493) );
  XOR U6342 ( .A(n2496), .B(n2497), .Z(n2495) );
  XOR U6343 ( .A(DB[3072]), .B(DB[3041]), .Z(n2497) );
  AND U6344 ( .A(n120), .B(n2498), .Z(n2496) );
  XOR U6345 ( .A(n2499), .B(n2500), .Z(n2498) );
  XOR U6346 ( .A(DB[3041]), .B(DB[3010]), .Z(n2500) );
  AND U6347 ( .A(n124), .B(n2501), .Z(n2499) );
  XOR U6348 ( .A(n2502), .B(n2503), .Z(n2501) );
  XOR U6349 ( .A(DB[3010]), .B(DB[2979]), .Z(n2503) );
  AND U6350 ( .A(n128), .B(n2504), .Z(n2502) );
  XOR U6351 ( .A(n2505), .B(n2506), .Z(n2504) );
  XOR U6352 ( .A(DB[2979]), .B(DB[2948]), .Z(n2506) );
  AND U6353 ( .A(n132), .B(n2507), .Z(n2505) );
  XOR U6354 ( .A(n2508), .B(n2509), .Z(n2507) );
  XOR U6355 ( .A(DB[2948]), .B(DB[2917]), .Z(n2509) );
  AND U6356 ( .A(n136), .B(n2510), .Z(n2508) );
  XOR U6357 ( .A(n2511), .B(n2512), .Z(n2510) );
  XOR U6358 ( .A(DB[2917]), .B(DB[2886]), .Z(n2512) );
  AND U6359 ( .A(n140), .B(n2513), .Z(n2511) );
  XOR U6360 ( .A(n2514), .B(n2515), .Z(n2513) );
  XOR U6361 ( .A(DB[2886]), .B(DB[2855]), .Z(n2515) );
  AND U6362 ( .A(n144), .B(n2516), .Z(n2514) );
  XOR U6363 ( .A(n2517), .B(n2518), .Z(n2516) );
  XOR U6364 ( .A(DB[2855]), .B(DB[2824]), .Z(n2518) );
  AND U6365 ( .A(n148), .B(n2519), .Z(n2517) );
  XOR U6366 ( .A(n2520), .B(n2521), .Z(n2519) );
  XOR U6367 ( .A(DB[2824]), .B(DB[2793]), .Z(n2521) );
  AND U6368 ( .A(n152), .B(n2522), .Z(n2520) );
  XOR U6369 ( .A(n2523), .B(n2524), .Z(n2522) );
  XOR U6370 ( .A(DB[2793]), .B(DB[2762]), .Z(n2524) );
  AND U6371 ( .A(n156), .B(n2525), .Z(n2523) );
  XOR U6372 ( .A(n2526), .B(n2527), .Z(n2525) );
  XOR U6373 ( .A(DB[2762]), .B(DB[2731]), .Z(n2527) );
  AND U6374 ( .A(n160), .B(n2528), .Z(n2526) );
  XOR U6375 ( .A(n2529), .B(n2530), .Z(n2528) );
  XOR U6376 ( .A(DB[2731]), .B(DB[2700]), .Z(n2530) );
  AND U6377 ( .A(n164), .B(n2531), .Z(n2529) );
  XOR U6378 ( .A(n2532), .B(n2533), .Z(n2531) );
  XOR U6379 ( .A(DB[2700]), .B(DB[2669]), .Z(n2533) );
  AND U6380 ( .A(n168), .B(n2534), .Z(n2532) );
  XOR U6381 ( .A(n2535), .B(n2536), .Z(n2534) );
  XOR U6382 ( .A(DB[2669]), .B(DB[2638]), .Z(n2536) );
  AND U6383 ( .A(n172), .B(n2537), .Z(n2535) );
  XOR U6384 ( .A(n2538), .B(n2539), .Z(n2537) );
  XOR U6385 ( .A(DB[2638]), .B(DB[2607]), .Z(n2539) );
  AND U6386 ( .A(n176), .B(n2540), .Z(n2538) );
  XOR U6387 ( .A(n2541), .B(n2542), .Z(n2540) );
  XOR U6388 ( .A(DB[2607]), .B(DB[2576]), .Z(n2542) );
  AND U6389 ( .A(n180), .B(n2543), .Z(n2541) );
  XOR U6390 ( .A(n2544), .B(n2545), .Z(n2543) );
  XOR U6391 ( .A(DB[2576]), .B(DB[2545]), .Z(n2545) );
  AND U6392 ( .A(n184), .B(n2546), .Z(n2544) );
  XOR U6393 ( .A(n2547), .B(n2548), .Z(n2546) );
  XOR U6394 ( .A(DB[2545]), .B(DB[2514]), .Z(n2548) );
  AND U6395 ( .A(n188), .B(n2549), .Z(n2547) );
  XOR U6396 ( .A(n2550), .B(n2551), .Z(n2549) );
  XOR U6397 ( .A(DB[2514]), .B(DB[2483]), .Z(n2551) );
  AND U6398 ( .A(n192), .B(n2552), .Z(n2550) );
  XOR U6399 ( .A(n2553), .B(n2554), .Z(n2552) );
  XOR U6400 ( .A(DB[2483]), .B(DB[2452]), .Z(n2554) );
  AND U6401 ( .A(n196), .B(n2555), .Z(n2553) );
  XOR U6402 ( .A(n2556), .B(n2557), .Z(n2555) );
  XOR U6403 ( .A(DB[2452]), .B(DB[2421]), .Z(n2557) );
  AND U6404 ( .A(n200), .B(n2558), .Z(n2556) );
  XOR U6405 ( .A(n2559), .B(n2560), .Z(n2558) );
  XOR U6406 ( .A(DB[2421]), .B(DB[2390]), .Z(n2560) );
  AND U6407 ( .A(n204), .B(n2561), .Z(n2559) );
  XOR U6408 ( .A(n2562), .B(n2563), .Z(n2561) );
  XOR U6409 ( .A(DB[2390]), .B(DB[2359]), .Z(n2563) );
  AND U6410 ( .A(n208), .B(n2564), .Z(n2562) );
  XOR U6411 ( .A(n2565), .B(n2566), .Z(n2564) );
  XOR U6412 ( .A(DB[2359]), .B(DB[2328]), .Z(n2566) );
  AND U6413 ( .A(n212), .B(n2567), .Z(n2565) );
  XOR U6414 ( .A(n2568), .B(n2569), .Z(n2567) );
  XOR U6415 ( .A(DB[2328]), .B(DB[2297]), .Z(n2569) );
  AND U6416 ( .A(n216), .B(n2570), .Z(n2568) );
  XOR U6417 ( .A(n2571), .B(n2572), .Z(n2570) );
  XOR U6418 ( .A(DB[2297]), .B(DB[2266]), .Z(n2572) );
  AND U6419 ( .A(n220), .B(n2573), .Z(n2571) );
  XOR U6420 ( .A(n2574), .B(n2575), .Z(n2573) );
  XOR U6421 ( .A(DB[2266]), .B(DB[2235]), .Z(n2575) );
  AND U6422 ( .A(n224), .B(n2576), .Z(n2574) );
  XOR U6423 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR U6424 ( .A(DB[2235]), .B(DB[2204]), .Z(n2578) );
  AND U6425 ( .A(n228), .B(n2579), .Z(n2577) );
  XOR U6426 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U6427 ( .A(DB[2204]), .B(DB[2173]), .Z(n2581) );
  AND U6428 ( .A(n232), .B(n2582), .Z(n2580) );
  XOR U6429 ( .A(n2583), .B(n2584), .Z(n2582) );
  XOR U6430 ( .A(DB[2173]), .B(DB[2142]), .Z(n2584) );
  AND U6431 ( .A(n236), .B(n2585), .Z(n2583) );
  XOR U6432 ( .A(n2586), .B(n2587), .Z(n2585) );
  XOR U6433 ( .A(DB[2142]), .B(DB[2111]), .Z(n2587) );
  AND U6434 ( .A(n240), .B(n2588), .Z(n2586) );
  XOR U6435 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR U6436 ( .A(DB[2111]), .B(DB[2080]), .Z(n2590) );
  AND U6437 ( .A(n244), .B(n2591), .Z(n2589) );
  XOR U6438 ( .A(n2592), .B(n2593), .Z(n2591) );
  XOR U6439 ( .A(DB[2080]), .B(DB[2049]), .Z(n2593) );
  AND U6440 ( .A(n248), .B(n2594), .Z(n2592) );
  XOR U6441 ( .A(n2595), .B(n2596), .Z(n2594) );
  XOR U6442 ( .A(DB[2049]), .B(DB[2018]), .Z(n2596) );
  AND U6443 ( .A(n252), .B(n2597), .Z(n2595) );
  XOR U6444 ( .A(n2598), .B(n2599), .Z(n2597) );
  XOR U6445 ( .A(DB[2018]), .B(DB[1987]), .Z(n2599) );
  AND U6446 ( .A(n256), .B(n2600), .Z(n2598) );
  XOR U6447 ( .A(n2601), .B(n2602), .Z(n2600) );
  XOR U6448 ( .A(DB[1987]), .B(DB[1956]), .Z(n2602) );
  AND U6449 ( .A(n260), .B(n2603), .Z(n2601) );
  XOR U6450 ( .A(n2604), .B(n2605), .Z(n2603) );
  XOR U6451 ( .A(DB[1956]), .B(DB[1925]), .Z(n2605) );
  AND U6452 ( .A(n264), .B(n2606), .Z(n2604) );
  XOR U6453 ( .A(n2607), .B(n2608), .Z(n2606) );
  XOR U6454 ( .A(DB[1925]), .B(DB[1894]), .Z(n2608) );
  AND U6455 ( .A(n268), .B(n2609), .Z(n2607) );
  XOR U6456 ( .A(n2610), .B(n2611), .Z(n2609) );
  XOR U6457 ( .A(DB[1894]), .B(DB[1863]), .Z(n2611) );
  AND U6458 ( .A(n272), .B(n2612), .Z(n2610) );
  XOR U6459 ( .A(n2613), .B(n2614), .Z(n2612) );
  XOR U6460 ( .A(DB[1863]), .B(DB[1832]), .Z(n2614) );
  AND U6461 ( .A(n276), .B(n2615), .Z(n2613) );
  XOR U6462 ( .A(n2616), .B(n2617), .Z(n2615) );
  XOR U6463 ( .A(DB[1832]), .B(DB[1801]), .Z(n2617) );
  AND U6464 ( .A(n280), .B(n2618), .Z(n2616) );
  XOR U6465 ( .A(n2619), .B(n2620), .Z(n2618) );
  XOR U6466 ( .A(DB[1801]), .B(DB[1770]), .Z(n2620) );
  AND U6467 ( .A(n284), .B(n2621), .Z(n2619) );
  XOR U6468 ( .A(n2622), .B(n2623), .Z(n2621) );
  XOR U6469 ( .A(DB[1770]), .B(DB[1739]), .Z(n2623) );
  AND U6470 ( .A(n288), .B(n2624), .Z(n2622) );
  XOR U6471 ( .A(n2625), .B(n2626), .Z(n2624) );
  XOR U6472 ( .A(DB[1739]), .B(DB[1708]), .Z(n2626) );
  AND U6473 ( .A(n292), .B(n2627), .Z(n2625) );
  XOR U6474 ( .A(n2628), .B(n2629), .Z(n2627) );
  XOR U6475 ( .A(DB[1708]), .B(DB[1677]), .Z(n2629) );
  AND U6476 ( .A(n296), .B(n2630), .Z(n2628) );
  XOR U6477 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U6478 ( .A(DB[1677]), .B(DB[1646]), .Z(n2632) );
  AND U6479 ( .A(n300), .B(n2633), .Z(n2631) );
  XOR U6480 ( .A(n2634), .B(n2635), .Z(n2633) );
  XOR U6481 ( .A(DB[1646]), .B(DB[1615]), .Z(n2635) );
  AND U6482 ( .A(n304), .B(n2636), .Z(n2634) );
  XOR U6483 ( .A(n2637), .B(n2638), .Z(n2636) );
  XOR U6484 ( .A(DB[1615]), .B(DB[1584]), .Z(n2638) );
  AND U6485 ( .A(n308), .B(n2639), .Z(n2637) );
  XOR U6486 ( .A(n2640), .B(n2641), .Z(n2639) );
  XOR U6487 ( .A(DB[1584]), .B(DB[1553]), .Z(n2641) );
  AND U6488 ( .A(n312), .B(n2642), .Z(n2640) );
  XOR U6489 ( .A(n2643), .B(n2644), .Z(n2642) );
  XOR U6490 ( .A(DB[1553]), .B(DB[1522]), .Z(n2644) );
  AND U6491 ( .A(n316), .B(n2645), .Z(n2643) );
  XOR U6492 ( .A(n2646), .B(n2647), .Z(n2645) );
  XOR U6493 ( .A(DB[1522]), .B(DB[1491]), .Z(n2647) );
  AND U6494 ( .A(n320), .B(n2648), .Z(n2646) );
  XOR U6495 ( .A(n2649), .B(n2650), .Z(n2648) );
  XOR U6496 ( .A(DB[1491]), .B(DB[1460]), .Z(n2650) );
  AND U6497 ( .A(n324), .B(n2651), .Z(n2649) );
  XOR U6498 ( .A(n2652), .B(n2653), .Z(n2651) );
  XOR U6499 ( .A(DB[1460]), .B(DB[1429]), .Z(n2653) );
  AND U6500 ( .A(n328), .B(n2654), .Z(n2652) );
  XOR U6501 ( .A(n2655), .B(n2656), .Z(n2654) );
  XOR U6502 ( .A(DB[1429]), .B(DB[1398]), .Z(n2656) );
  AND U6503 ( .A(n332), .B(n2657), .Z(n2655) );
  XOR U6504 ( .A(n2658), .B(n2659), .Z(n2657) );
  XOR U6505 ( .A(DB[1398]), .B(DB[1367]), .Z(n2659) );
  AND U6506 ( .A(n336), .B(n2660), .Z(n2658) );
  XOR U6507 ( .A(n2661), .B(n2662), .Z(n2660) );
  XOR U6508 ( .A(DB[1367]), .B(DB[1336]), .Z(n2662) );
  AND U6509 ( .A(n340), .B(n2663), .Z(n2661) );
  XOR U6510 ( .A(n2664), .B(n2665), .Z(n2663) );
  XOR U6511 ( .A(DB[1336]), .B(DB[1305]), .Z(n2665) );
  AND U6512 ( .A(n344), .B(n2666), .Z(n2664) );
  XOR U6513 ( .A(n2667), .B(n2668), .Z(n2666) );
  XOR U6514 ( .A(DB[1305]), .B(DB[1274]), .Z(n2668) );
  AND U6515 ( .A(n348), .B(n2669), .Z(n2667) );
  XOR U6516 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR U6517 ( .A(DB[1274]), .B(DB[1243]), .Z(n2671) );
  AND U6518 ( .A(n352), .B(n2672), .Z(n2670) );
  XOR U6519 ( .A(n2673), .B(n2674), .Z(n2672) );
  XOR U6520 ( .A(DB[1243]), .B(DB[1212]), .Z(n2674) );
  AND U6521 ( .A(n356), .B(n2675), .Z(n2673) );
  XOR U6522 ( .A(n2676), .B(n2677), .Z(n2675) );
  XOR U6523 ( .A(DB[1212]), .B(DB[1181]), .Z(n2677) );
  AND U6524 ( .A(n360), .B(n2678), .Z(n2676) );
  XOR U6525 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR U6526 ( .A(DB[1181]), .B(DB[1150]), .Z(n2680) );
  AND U6527 ( .A(n364), .B(n2681), .Z(n2679) );
  XOR U6528 ( .A(n2682), .B(n2683), .Z(n2681) );
  XOR U6529 ( .A(DB[1150]), .B(DB[1119]), .Z(n2683) );
  AND U6530 ( .A(n368), .B(n2684), .Z(n2682) );
  XOR U6531 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR U6532 ( .A(DB[1119]), .B(DB[1088]), .Z(n2686) );
  AND U6533 ( .A(n372), .B(n2687), .Z(n2685) );
  XOR U6534 ( .A(n2688), .B(n2689), .Z(n2687) );
  XOR U6535 ( .A(DB[1088]), .B(DB[1057]), .Z(n2689) );
  AND U6536 ( .A(n376), .B(n2690), .Z(n2688) );
  XOR U6537 ( .A(n2691), .B(n2692), .Z(n2690) );
  XOR U6538 ( .A(DB[1057]), .B(DB[1026]), .Z(n2692) );
  AND U6539 ( .A(n380), .B(n2693), .Z(n2691) );
  XOR U6540 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR U6541 ( .A(DB[995]), .B(DB[1026]), .Z(n2695) );
  AND U6542 ( .A(n384), .B(n2696), .Z(n2694) );
  XOR U6543 ( .A(n2697), .B(n2698), .Z(n2696) );
  XOR U6544 ( .A(DB[995]), .B(DB[964]), .Z(n2698) );
  AND U6545 ( .A(n388), .B(n2699), .Z(n2697) );
  XOR U6546 ( .A(n2700), .B(n2701), .Z(n2699) );
  XOR U6547 ( .A(DB[964]), .B(DB[933]), .Z(n2701) );
  AND U6548 ( .A(n392), .B(n2702), .Z(n2700) );
  XOR U6549 ( .A(n2703), .B(n2704), .Z(n2702) );
  XOR U6550 ( .A(DB[933]), .B(DB[902]), .Z(n2704) );
  AND U6551 ( .A(n396), .B(n2705), .Z(n2703) );
  XOR U6552 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U6553 ( .A(DB[902]), .B(DB[871]), .Z(n2707) );
  AND U6554 ( .A(n400), .B(n2708), .Z(n2706) );
  XOR U6555 ( .A(n2709), .B(n2710), .Z(n2708) );
  XOR U6556 ( .A(DB[871]), .B(DB[840]), .Z(n2710) );
  AND U6557 ( .A(n404), .B(n2711), .Z(n2709) );
  XOR U6558 ( .A(n2712), .B(n2713), .Z(n2711) );
  XOR U6559 ( .A(DB[840]), .B(DB[809]), .Z(n2713) );
  AND U6560 ( .A(n408), .B(n2714), .Z(n2712) );
  XOR U6561 ( .A(n2715), .B(n2716), .Z(n2714) );
  XOR U6562 ( .A(DB[809]), .B(DB[778]), .Z(n2716) );
  AND U6563 ( .A(n412), .B(n2717), .Z(n2715) );
  XOR U6564 ( .A(n2718), .B(n2719), .Z(n2717) );
  XOR U6565 ( .A(DB[778]), .B(DB[747]), .Z(n2719) );
  AND U6566 ( .A(n416), .B(n2720), .Z(n2718) );
  XOR U6567 ( .A(n2721), .B(n2722), .Z(n2720) );
  XOR U6568 ( .A(DB[747]), .B(DB[716]), .Z(n2722) );
  AND U6569 ( .A(n420), .B(n2723), .Z(n2721) );
  XOR U6570 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR U6571 ( .A(DB[716]), .B(DB[685]), .Z(n2725) );
  AND U6572 ( .A(n424), .B(n2726), .Z(n2724) );
  XOR U6573 ( .A(n2727), .B(n2728), .Z(n2726) );
  XOR U6574 ( .A(DB[685]), .B(DB[654]), .Z(n2728) );
  AND U6575 ( .A(n428), .B(n2729), .Z(n2727) );
  XOR U6576 ( .A(n2730), .B(n2731), .Z(n2729) );
  XOR U6577 ( .A(DB[654]), .B(DB[623]), .Z(n2731) );
  AND U6578 ( .A(n432), .B(n2732), .Z(n2730) );
  XOR U6579 ( .A(n2733), .B(n2734), .Z(n2732) );
  XOR U6580 ( .A(DB[623]), .B(DB[592]), .Z(n2734) );
  AND U6581 ( .A(n436), .B(n2735), .Z(n2733) );
  XOR U6582 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR U6583 ( .A(DB[592]), .B(DB[561]), .Z(n2737) );
  AND U6584 ( .A(n440), .B(n2738), .Z(n2736) );
  XOR U6585 ( .A(n2739), .B(n2740), .Z(n2738) );
  XOR U6586 ( .A(DB[561]), .B(DB[530]), .Z(n2740) );
  AND U6587 ( .A(n444), .B(n2741), .Z(n2739) );
  XOR U6588 ( .A(n2742), .B(n2743), .Z(n2741) );
  XOR U6589 ( .A(DB[530]), .B(DB[499]), .Z(n2743) );
  AND U6590 ( .A(n448), .B(n2744), .Z(n2742) );
  XOR U6591 ( .A(n2745), .B(n2746), .Z(n2744) );
  XOR U6592 ( .A(DB[499]), .B(DB[468]), .Z(n2746) );
  AND U6593 ( .A(n452), .B(n2747), .Z(n2745) );
  XOR U6594 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR U6595 ( .A(DB[468]), .B(DB[437]), .Z(n2749) );
  AND U6596 ( .A(n456), .B(n2750), .Z(n2748) );
  XOR U6597 ( .A(n2751), .B(n2752), .Z(n2750) );
  XOR U6598 ( .A(DB[437]), .B(DB[406]), .Z(n2752) );
  AND U6599 ( .A(n460), .B(n2753), .Z(n2751) );
  XOR U6600 ( .A(n2754), .B(n2755), .Z(n2753) );
  XOR U6601 ( .A(DB[406]), .B(DB[375]), .Z(n2755) );
  AND U6602 ( .A(n464), .B(n2756), .Z(n2754) );
  XOR U6603 ( .A(n2757), .B(n2758), .Z(n2756) );
  XOR U6604 ( .A(DB[375]), .B(DB[344]), .Z(n2758) );
  AND U6605 ( .A(n468), .B(n2759), .Z(n2757) );
  XOR U6606 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U6607 ( .A(DB[344]), .B(DB[313]), .Z(n2761) );
  AND U6608 ( .A(n472), .B(n2762), .Z(n2760) );
  XOR U6609 ( .A(n2763), .B(n2764), .Z(n2762) );
  XOR U6610 ( .A(DB[313]), .B(DB[282]), .Z(n2764) );
  AND U6611 ( .A(n476), .B(n2765), .Z(n2763) );
  XOR U6612 ( .A(n2766), .B(n2767), .Z(n2765) );
  XOR U6613 ( .A(DB[282]), .B(DB[251]), .Z(n2767) );
  AND U6614 ( .A(n480), .B(n2768), .Z(n2766) );
  XOR U6615 ( .A(n2769), .B(n2770), .Z(n2768) );
  XOR U6616 ( .A(DB[251]), .B(DB[220]), .Z(n2770) );
  AND U6617 ( .A(n484), .B(n2771), .Z(n2769) );
  XOR U6618 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U6619 ( .A(DB[220]), .B(DB[189]), .Z(n2773) );
  AND U6620 ( .A(n488), .B(n2774), .Z(n2772) );
  XOR U6621 ( .A(n2775), .B(n2776), .Z(n2774) );
  XOR U6622 ( .A(DB[189]), .B(DB[158]), .Z(n2776) );
  AND U6623 ( .A(n492), .B(n2777), .Z(n2775) );
  XOR U6624 ( .A(n2778), .B(n2779), .Z(n2777) );
  XOR U6625 ( .A(DB[158]), .B(DB[127]), .Z(n2779) );
  AND U6626 ( .A(n496), .B(n2780), .Z(n2778) );
  XOR U6627 ( .A(n2781), .B(n2782), .Z(n2780) );
  XOR U6628 ( .A(DB[96]), .B(DB[127]), .Z(n2782) );
  AND U6629 ( .A(n500), .B(n2783), .Z(n2781) );
  XOR U6630 ( .A(n2784), .B(n2785), .Z(n2783) );
  XOR U6631 ( .A(DB[96]), .B(DB[65]), .Z(n2785) );
  AND U6632 ( .A(n504), .B(n2786), .Z(n2784) );
  XOR U6633 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U6634 ( .A(DB[65]), .B(DB[34]), .Z(n2788) );
  AND U6635 ( .A(n508), .B(n2789), .Z(n2787) );
  XOR U6636 ( .A(DB[3]), .B(DB[34]), .Z(n2789) );
  XOR U6637 ( .A(DB[3967]), .B(n2790), .Z(min_val_out[30]) );
  AND U6638 ( .A(n2), .B(n2791), .Z(n2790) );
  XOR U6639 ( .A(n2792), .B(n2793), .Z(n2791) );
  XOR U6640 ( .A(DB[3967]), .B(DB[3936]), .Z(n2793) );
  AND U6641 ( .A(n8), .B(n2794), .Z(n2792) );
  XOR U6642 ( .A(n2795), .B(n2796), .Z(n2794) );
  XOR U6643 ( .A(DB[3936]), .B(DB[3905]), .Z(n2796) );
  AND U6644 ( .A(n12), .B(n2797), .Z(n2795) );
  XOR U6645 ( .A(n2798), .B(n2799), .Z(n2797) );
  XOR U6646 ( .A(DB[3905]), .B(DB[3874]), .Z(n2799) );
  AND U6647 ( .A(n16), .B(n2800), .Z(n2798) );
  XOR U6648 ( .A(n2801), .B(n2802), .Z(n2800) );
  XOR U6649 ( .A(DB[3874]), .B(DB[3843]), .Z(n2802) );
  AND U6650 ( .A(n20), .B(n2803), .Z(n2801) );
  XOR U6651 ( .A(n2804), .B(n2805), .Z(n2803) );
  XOR U6652 ( .A(DB[3843]), .B(DB[3812]), .Z(n2805) );
  AND U6653 ( .A(n24), .B(n2806), .Z(n2804) );
  XOR U6654 ( .A(n2807), .B(n2808), .Z(n2806) );
  XOR U6655 ( .A(DB[3812]), .B(DB[3781]), .Z(n2808) );
  AND U6656 ( .A(n28), .B(n2809), .Z(n2807) );
  XOR U6657 ( .A(n2810), .B(n2811), .Z(n2809) );
  XOR U6658 ( .A(DB[3781]), .B(DB[3750]), .Z(n2811) );
  AND U6659 ( .A(n32), .B(n2812), .Z(n2810) );
  XOR U6660 ( .A(n2813), .B(n2814), .Z(n2812) );
  XOR U6661 ( .A(DB[3750]), .B(DB[3719]), .Z(n2814) );
  AND U6662 ( .A(n36), .B(n2815), .Z(n2813) );
  XOR U6663 ( .A(n2816), .B(n2817), .Z(n2815) );
  XOR U6664 ( .A(DB[3719]), .B(DB[3688]), .Z(n2817) );
  AND U6665 ( .A(n40), .B(n2818), .Z(n2816) );
  XOR U6666 ( .A(n2819), .B(n2820), .Z(n2818) );
  XOR U6667 ( .A(DB[3688]), .B(DB[3657]), .Z(n2820) );
  AND U6668 ( .A(n44), .B(n2821), .Z(n2819) );
  XOR U6669 ( .A(n2822), .B(n2823), .Z(n2821) );
  XOR U6670 ( .A(DB[3657]), .B(DB[3626]), .Z(n2823) );
  AND U6671 ( .A(n48), .B(n2824), .Z(n2822) );
  XOR U6672 ( .A(n2825), .B(n2826), .Z(n2824) );
  XOR U6673 ( .A(DB[3626]), .B(DB[3595]), .Z(n2826) );
  AND U6674 ( .A(n52), .B(n2827), .Z(n2825) );
  XOR U6675 ( .A(n2828), .B(n2829), .Z(n2827) );
  XOR U6676 ( .A(DB[3595]), .B(DB[3564]), .Z(n2829) );
  AND U6677 ( .A(n56), .B(n2830), .Z(n2828) );
  XOR U6678 ( .A(n2831), .B(n2832), .Z(n2830) );
  XOR U6679 ( .A(DB[3564]), .B(DB[3533]), .Z(n2832) );
  AND U6680 ( .A(n60), .B(n2833), .Z(n2831) );
  XOR U6681 ( .A(n2834), .B(n2835), .Z(n2833) );
  XOR U6682 ( .A(DB[3533]), .B(DB[3502]), .Z(n2835) );
  AND U6683 ( .A(n64), .B(n2836), .Z(n2834) );
  XOR U6684 ( .A(n2837), .B(n2838), .Z(n2836) );
  XOR U6685 ( .A(DB[3502]), .B(DB[3471]), .Z(n2838) );
  AND U6686 ( .A(n68), .B(n2839), .Z(n2837) );
  XOR U6687 ( .A(n2840), .B(n2841), .Z(n2839) );
  XOR U6688 ( .A(DB[3471]), .B(DB[3440]), .Z(n2841) );
  AND U6689 ( .A(n72), .B(n2842), .Z(n2840) );
  XOR U6690 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR U6691 ( .A(DB[3440]), .B(DB[3409]), .Z(n2844) );
  AND U6692 ( .A(n76), .B(n2845), .Z(n2843) );
  XOR U6693 ( .A(n2846), .B(n2847), .Z(n2845) );
  XOR U6694 ( .A(DB[3409]), .B(DB[3378]), .Z(n2847) );
  AND U6695 ( .A(n80), .B(n2848), .Z(n2846) );
  XOR U6696 ( .A(n2849), .B(n2850), .Z(n2848) );
  XOR U6697 ( .A(DB[3378]), .B(DB[3347]), .Z(n2850) );
  AND U6698 ( .A(n84), .B(n2851), .Z(n2849) );
  XOR U6699 ( .A(n2852), .B(n2853), .Z(n2851) );
  XOR U6700 ( .A(DB[3347]), .B(DB[3316]), .Z(n2853) );
  AND U6701 ( .A(n88), .B(n2854), .Z(n2852) );
  XOR U6702 ( .A(n2855), .B(n2856), .Z(n2854) );
  XOR U6703 ( .A(DB[3316]), .B(DB[3285]), .Z(n2856) );
  AND U6704 ( .A(n92), .B(n2857), .Z(n2855) );
  XOR U6705 ( .A(n2858), .B(n2859), .Z(n2857) );
  XOR U6706 ( .A(DB[3285]), .B(DB[3254]), .Z(n2859) );
  AND U6707 ( .A(n96), .B(n2860), .Z(n2858) );
  XOR U6708 ( .A(n2861), .B(n2862), .Z(n2860) );
  XOR U6709 ( .A(DB[3254]), .B(DB[3223]), .Z(n2862) );
  AND U6710 ( .A(n100), .B(n2863), .Z(n2861) );
  XOR U6711 ( .A(n2864), .B(n2865), .Z(n2863) );
  XOR U6712 ( .A(DB[3223]), .B(DB[3192]), .Z(n2865) );
  AND U6713 ( .A(n104), .B(n2866), .Z(n2864) );
  XOR U6714 ( .A(n2867), .B(n2868), .Z(n2866) );
  XOR U6715 ( .A(DB[3192]), .B(DB[3161]), .Z(n2868) );
  AND U6716 ( .A(n108), .B(n2869), .Z(n2867) );
  XOR U6717 ( .A(n2870), .B(n2871), .Z(n2869) );
  XOR U6718 ( .A(DB[3161]), .B(DB[3130]), .Z(n2871) );
  AND U6719 ( .A(n112), .B(n2872), .Z(n2870) );
  XOR U6720 ( .A(n2873), .B(n2874), .Z(n2872) );
  XOR U6721 ( .A(DB[3130]), .B(DB[3099]), .Z(n2874) );
  AND U6722 ( .A(n116), .B(n2875), .Z(n2873) );
  XOR U6723 ( .A(n2876), .B(n2877), .Z(n2875) );
  XOR U6724 ( .A(DB[3099]), .B(DB[3068]), .Z(n2877) );
  AND U6725 ( .A(n120), .B(n2878), .Z(n2876) );
  XOR U6726 ( .A(n2879), .B(n2880), .Z(n2878) );
  XOR U6727 ( .A(DB[3068]), .B(DB[3037]), .Z(n2880) );
  AND U6728 ( .A(n124), .B(n2881), .Z(n2879) );
  XOR U6729 ( .A(n2882), .B(n2883), .Z(n2881) );
  XOR U6730 ( .A(DB[3037]), .B(DB[3006]), .Z(n2883) );
  AND U6731 ( .A(n128), .B(n2884), .Z(n2882) );
  XOR U6732 ( .A(n2885), .B(n2886), .Z(n2884) );
  XOR U6733 ( .A(DB[3006]), .B(DB[2975]), .Z(n2886) );
  AND U6734 ( .A(n132), .B(n2887), .Z(n2885) );
  XOR U6735 ( .A(n2888), .B(n2889), .Z(n2887) );
  XOR U6736 ( .A(DB[2975]), .B(DB[2944]), .Z(n2889) );
  AND U6737 ( .A(n136), .B(n2890), .Z(n2888) );
  XOR U6738 ( .A(n2891), .B(n2892), .Z(n2890) );
  XOR U6739 ( .A(DB[2944]), .B(DB[2913]), .Z(n2892) );
  AND U6740 ( .A(n140), .B(n2893), .Z(n2891) );
  XOR U6741 ( .A(n2894), .B(n2895), .Z(n2893) );
  XOR U6742 ( .A(DB[2913]), .B(DB[2882]), .Z(n2895) );
  AND U6743 ( .A(n144), .B(n2896), .Z(n2894) );
  XOR U6744 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR U6745 ( .A(DB[2882]), .B(DB[2851]), .Z(n2898) );
  AND U6746 ( .A(n148), .B(n2899), .Z(n2897) );
  XOR U6747 ( .A(n2900), .B(n2901), .Z(n2899) );
  XOR U6748 ( .A(DB[2851]), .B(DB[2820]), .Z(n2901) );
  AND U6749 ( .A(n152), .B(n2902), .Z(n2900) );
  XOR U6750 ( .A(n2903), .B(n2904), .Z(n2902) );
  XOR U6751 ( .A(DB[2820]), .B(DB[2789]), .Z(n2904) );
  AND U6752 ( .A(n156), .B(n2905), .Z(n2903) );
  XOR U6753 ( .A(n2906), .B(n2907), .Z(n2905) );
  XOR U6754 ( .A(DB[2789]), .B(DB[2758]), .Z(n2907) );
  AND U6755 ( .A(n160), .B(n2908), .Z(n2906) );
  XOR U6756 ( .A(n2909), .B(n2910), .Z(n2908) );
  XOR U6757 ( .A(DB[2758]), .B(DB[2727]), .Z(n2910) );
  AND U6758 ( .A(n164), .B(n2911), .Z(n2909) );
  XOR U6759 ( .A(n2912), .B(n2913), .Z(n2911) );
  XOR U6760 ( .A(DB[2727]), .B(DB[2696]), .Z(n2913) );
  AND U6761 ( .A(n168), .B(n2914), .Z(n2912) );
  XOR U6762 ( .A(n2915), .B(n2916), .Z(n2914) );
  XOR U6763 ( .A(DB[2696]), .B(DB[2665]), .Z(n2916) );
  AND U6764 ( .A(n172), .B(n2917), .Z(n2915) );
  XOR U6765 ( .A(n2918), .B(n2919), .Z(n2917) );
  XOR U6766 ( .A(DB[2665]), .B(DB[2634]), .Z(n2919) );
  AND U6767 ( .A(n176), .B(n2920), .Z(n2918) );
  XOR U6768 ( .A(n2921), .B(n2922), .Z(n2920) );
  XOR U6769 ( .A(DB[2634]), .B(DB[2603]), .Z(n2922) );
  AND U6770 ( .A(n180), .B(n2923), .Z(n2921) );
  XOR U6771 ( .A(n2924), .B(n2925), .Z(n2923) );
  XOR U6772 ( .A(DB[2603]), .B(DB[2572]), .Z(n2925) );
  AND U6773 ( .A(n184), .B(n2926), .Z(n2924) );
  XOR U6774 ( .A(n2927), .B(n2928), .Z(n2926) );
  XOR U6775 ( .A(DB[2572]), .B(DB[2541]), .Z(n2928) );
  AND U6776 ( .A(n188), .B(n2929), .Z(n2927) );
  XOR U6777 ( .A(n2930), .B(n2931), .Z(n2929) );
  XOR U6778 ( .A(DB[2541]), .B(DB[2510]), .Z(n2931) );
  AND U6779 ( .A(n192), .B(n2932), .Z(n2930) );
  XOR U6780 ( .A(n2933), .B(n2934), .Z(n2932) );
  XOR U6781 ( .A(DB[2510]), .B(DB[2479]), .Z(n2934) );
  AND U6782 ( .A(n196), .B(n2935), .Z(n2933) );
  XOR U6783 ( .A(n2936), .B(n2937), .Z(n2935) );
  XOR U6784 ( .A(DB[2479]), .B(DB[2448]), .Z(n2937) );
  AND U6785 ( .A(n200), .B(n2938), .Z(n2936) );
  XOR U6786 ( .A(n2939), .B(n2940), .Z(n2938) );
  XOR U6787 ( .A(DB[2448]), .B(DB[2417]), .Z(n2940) );
  AND U6788 ( .A(n204), .B(n2941), .Z(n2939) );
  XOR U6789 ( .A(n2942), .B(n2943), .Z(n2941) );
  XOR U6790 ( .A(DB[2417]), .B(DB[2386]), .Z(n2943) );
  AND U6791 ( .A(n208), .B(n2944), .Z(n2942) );
  XOR U6792 ( .A(n2945), .B(n2946), .Z(n2944) );
  XOR U6793 ( .A(DB[2386]), .B(DB[2355]), .Z(n2946) );
  AND U6794 ( .A(n212), .B(n2947), .Z(n2945) );
  XOR U6795 ( .A(n2948), .B(n2949), .Z(n2947) );
  XOR U6796 ( .A(DB[2355]), .B(DB[2324]), .Z(n2949) );
  AND U6797 ( .A(n216), .B(n2950), .Z(n2948) );
  XOR U6798 ( .A(n2951), .B(n2952), .Z(n2950) );
  XOR U6799 ( .A(DB[2324]), .B(DB[2293]), .Z(n2952) );
  AND U6800 ( .A(n220), .B(n2953), .Z(n2951) );
  XOR U6801 ( .A(n2954), .B(n2955), .Z(n2953) );
  XOR U6802 ( .A(DB[2293]), .B(DB[2262]), .Z(n2955) );
  AND U6803 ( .A(n224), .B(n2956), .Z(n2954) );
  XOR U6804 ( .A(n2957), .B(n2958), .Z(n2956) );
  XOR U6805 ( .A(DB[2262]), .B(DB[2231]), .Z(n2958) );
  AND U6806 ( .A(n228), .B(n2959), .Z(n2957) );
  XOR U6807 ( .A(n2960), .B(n2961), .Z(n2959) );
  XOR U6808 ( .A(DB[2231]), .B(DB[2200]), .Z(n2961) );
  AND U6809 ( .A(n232), .B(n2962), .Z(n2960) );
  XOR U6810 ( .A(n2963), .B(n2964), .Z(n2962) );
  XOR U6811 ( .A(DB[2200]), .B(DB[2169]), .Z(n2964) );
  AND U6812 ( .A(n236), .B(n2965), .Z(n2963) );
  XOR U6813 ( .A(n2966), .B(n2967), .Z(n2965) );
  XOR U6814 ( .A(DB[2169]), .B(DB[2138]), .Z(n2967) );
  AND U6815 ( .A(n240), .B(n2968), .Z(n2966) );
  XOR U6816 ( .A(n2969), .B(n2970), .Z(n2968) );
  XOR U6817 ( .A(DB[2138]), .B(DB[2107]), .Z(n2970) );
  AND U6818 ( .A(n244), .B(n2971), .Z(n2969) );
  XOR U6819 ( .A(n2972), .B(n2973), .Z(n2971) );
  XOR U6820 ( .A(DB[2107]), .B(DB[2076]), .Z(n2973) );
  AND U6821 ( .A(n248), .B(n2974), .Z(n2972) );
  XOR U6822 ( .A(n2975), .B(n2976), .Z(n2974) );
  XOR U6823 ( .A(DB[2076]), .B(DB[2045]), .Z(n2976) );
  AND U6824 ( .A(n252), .B(n2977), .Z(n2975) );
  XOR U6825 ( .A(n2978), .B(n2979), .Z(n2977) );
  XOR U6826 ( .A(DB[2045]), .B(DB[2014]), .Z(n2979) );
  AND U6827 ( .A(n256), .B(n2980), .Z(n2978) );
  XOR U6828 ( .A(n2981), .B(n2982), .Z(n2980) );
  XOR U6829 ( .A(DB[2014]), .B(DB[1983]), .Z(n2982) );
  AND U6830 ( .A(n260), .B(n2983), .Z(n2981) );
  XOR U6831 ( .A(n2984), .B(n2985), .Z(n2983) );
  XOR U6832 ( .A(DB[1983]), .B(DB[1952]), .Z(n2985) );
  AND U6833 ( .A(n264), .B(n2986), .Z(n2984) );
  XOR U6834 ( .A(n2987), .B(n2988), .Z(n2986) );
  XOR U6835 ( .A(DB[1952]), .B(DB[1921]), .Z(n2988) );
  AND U6836 ( .A(n268), .B(n2989), .Z(n2987) );
  XOR U6837 ( .A(n2990), .B(n2991), .Z(n2989) );
  XOR U6838 ( .A(DB[1921]), .B(DB[1890]), .Z(n2991) );
  AND U6839 ( .A(n272), .B(n2992), .Z(n2990) );
  XOR U6840 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U6841 ( .A(DB[1890]), .B(DB[1859]), .Z(n2994) );
  AND U6842 ( .A(n276), .B(n2995), .Z(n2993) );
  XOR U6843 ( .A(n2996), .B(n2997), .Z(n2995) );
  XOR U6844 ( .A(DB[1859]), .B(DB[1828]), .Z(n2997) );
  AND U6845 ( .A(n280), .B(n2998), .Z(n2996) );
  XOR U6846 ( .A(n2999), .B(n3000), .Z(n2998) );
  XOR U6847 ( .A(DB[1828]), .B(DB[1797]), .Z(n3000) );
  AND U6848 ( .A(n284), .B(n3001), .Z(n2999) );
  XOR U6849 ( .A(n3002), .B(n3003), .Z(n3001) );
  XOR U6850 ( .A(DB[1797]), .B(DB[1766]), .Z(n3003) );
  AND U6851 ( .A(n288), .B(n3004), .Z(n3002) );
  XOR U6852 ( .A(n3005), .B(n3006), .Z(n3004) );
  XOR U6853 ( .A(DB[1766]), .B(DB[1735]), .Z(n3006) );
  AND U6854 ( .A(n292), .B(n3007), .Z(n3005) );
  XOR U6855 ( .A(n3008), .B(n3009), .Z(n3007) );
  XOR U6856 ( .A(DB[1735]), .B(DB[1704]), .Z(n3009) );
  AND U6857 ( .A(n296), .B(n3010), .Z(n3008) );
  XOR U6858 ( .A(n3011), .B(n3012), .Z(n3010) );
  XOR U6859 ( .A(DB[1704]), .B(DB[1673]), .Z(n3012) );
  AND U6860 ( .A(n300), .B(n3013), .Z(n3011) );
  XOR U6861 ( .A(n3014), .B(n3015), .Z(n3013) );
  XOR U6862 ( .A(DB[1673]), .B(DB[1642]), .Z(n3015) );
  AND U6863 ( .A(n304), .B(n3016), .Z(n3014) );
  XOR U6864 ( .A(n3017), .B(n3018), .Z(n3016) );
  XOR U6865 ( .A(DB[1642]), .B(DB[1611]), .Z(n3018) );
  AND U6866 ( .A(n308), .B(n3019), .Z(n3017) );
  XOR U6867 ( .A(n3020), .B(n3021), .Z(n3019) );
  XOR U6868 ( .A(DB[1611]), .B(DB[1580]), .Z(n3021) );
  AND U6869 ( .A(n312), .B(n3022), .Z(n3020) );
  XOR U6870 ( .A(n3023), .B(n3024), .Z(n3022) );
  XOR U6871 ( .A(DB[1580]), .B(DB[1549]), .Z(n3024) );
  AND U6872 ( .A(n316), .B(n3025), .Z(n3023) );
  XOR U6873 ( .A(n3026), .B(n3027), .Z(n3025) );
  XOR U6874 ( .A(DB[1549]), .B(DB[1518]), .Z(n3027) );
  AND U6875 ( .A(n320), .B(n3028), .Z(n3026) );
  XOR U6876 ( .A(n3029), .B(n3030), .Z(n3028) );
  XOR U6877 ( .A(DB[1518]), .B(DB[1487]), .Z(n3030) );
  AND U6878 ( .A(n324), .B(n3031), .Z(n3029) );
  XOR U6879 ( .A(n3032), .B(n3033), .Z(n3031) );
  XOR U6880 ( .A(DB[1487]), .B(DB[1456]), .Z(n3033) );
  AND U6881 ( .A(n328), .B(n3034), .Z(n3032) );
  XOR U6882 ( .A(n3035), .B(n3036), .Z(n3034) );
  XOR U6883 ( .A(DB[1456]), .B(DB[1425]), .Z(n3036) );
  AND U6884 ( .A(n332), .B(n3037), .Z(n3035) );
  XOR U6885 ( .A(n3038), .B(n3039), .Z(n3037) );
  XOR U6886 ( .A(DB[1425]), .B(DB[1394]), .Z(n3039) );
  AND U6887 ( .A(n336), .B(n3040), .Z(n3038) );
  XOR U6888 ( .A(n3041), .B(n3042), .Z(n3040) );
  XOR U6889 ( .A(DB[1394]), .B(DB[1363]), .Z(n3042) );
  AND U6890 ( .A(n340), .B(n3043), .Z(n3041) );
  XOR U6891 ( .A(n3044), .B(n3045), .Z(n3043) );
  XOR U6892 ( .A(DB[1363]), .B(DB[1332]), .Z(n3045) );
  AND U6893 ( .A(n344), .B(n3046), .Z(n3044) );
  XOR U6894 ( .A(n3047), .B(n3048), .Z(n3046) );
  XOR U6895 ( .A(DB[1332]), .B(DB[1301]), .Z(n3048) );
  AND U6896 ( .A(n348), .B(n3049), .Z(n3047) );
  XOR U6897 ( .A(n3050), .B(n3051), .Z(n3049) );
  XOR U6898 ( .A(DB[1301]), .B(DB[1270]), .Z(n3051) );
  AND U6899 ( .A(n352), .B(n3052), .Z(n3050) );
  XOR U6900 ( .A(n3053), .B(n3054), .Z(n3052) );
  XOR U6901 ( .A(DB[1270]), .B(DB[1239]), .Z(n3054) );
  AND U6902 ( .A(n356), .B(n3055), .Z(n3053) );
  XOR U6903 ( .A(n3056), .B(n3057), .Z(n3055) );
  XOR U6904 ( .A(DB[1239]), .B(DB[1208]), .Z(n3057) );
  AND U6905 ( .A(n360), .B(n3058), .Z(n3056) );
  XOR U6906 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR U6907 ( .A(DB[1208]), .B(DB[1177]), .Z(n3060) );
  AND U6908 ( .A(n364), .B(n3061), .Z(n3059) );
  XOR U6909 ( .A(n3062), .B(n3063), .Z(n3061) );
  XOR U6910 ( .A(DB[1177]), .B(DB[1146]), .Z(n3063) );
  AND U6911 ( .A(n368), .B(n3064), .Z(n3062) );
  XOR U6912 ( .A(n3065), .B(n3066), .Z(n3064) );
  XOR U6913 ( .A(DB[1146]), .B(DB[1115]), .Z(n3066) );
  AND U6914 ( .A(n372), .B(n3067), .Z(n3065) );
  XOR U6915 ( .A(n3068), .B(n3069), .Z(n3067) );
  XOR U6916 ( .A(DB[1115]), .B(DB[1084]), .Z(n3069) );
  AND U6917 ( .A(n376), .B(n3070), .Z(n3068) );
  XOR U6918 ( .A(n3071), .B(n3072), .Z(n3070) );
  XOR U6919 ( .A(DB[1084]), .B(DB[1053]), .Z(n3072) );
  AND U6920 ( .A(n380), .B(n3073), .Z(n3071) );
  XOR U6921 ( .A(n3074), .B(n3075), .Z(n3073) );
  XOR U6922 ( .A(DB[1053]), .B(DB[1022]), .Z(n3075) );
  AND U6923 ( .A(n384), .B(n3076), .Z(n3074) );
  XOR U6924 ( .A(n3077), .B(n3078), .Z(n3076) );
  XOR U6925 ( .A(DB[991]), .B(DB[1022]), .Z(n3078) );
  AND U6926 ( .A(n388), .B(n3079), .Z(n3077) );
  XOR U6927 ( .A(n3080), .B(n3081), .Z(n3079) );
  XOR U6928 ( .A(DB[991]), .B(DB[960]), .Z(n3081) );
  AND U6929 ( .A(n392), .B(n3082), .Z(n3080) );
  XOR U6930 ( .A(n3083), .B(n3084), .Z(n3082) );
  XOR U6931 ( .A(DB[960]), .B(DB[929]), .Z(n3084) );
  AND U6932 ( .A(n396), .B(n3085), .Z(n3083) );
  XOR U6933 ( .A(n3086), .B(n3087), .Z(n3085) );
  XOR U6934 ( .A(DB[929]), .B(DB[898]), .Z(n3087) );
  AND U6935 ( .A(n400), .B(n3088), .Z(n3086) );
  XOR U6936 ( .A(n3089), .B(n3090), .Z(n3088) );
  XOR U6937 ( .A(DB[898]), .B(DB[867]), .Z(n3090) );
  AND U6938 ( .A(n404), .B(n3091), .Z(n3089) );
  XOR U6939 ( .A(n3092), .B(n3093), .Z(n3091) );
  XOR U6940 ( .A(DB[867]), .B(DB[836]), .Z(n3093) );
  AND U6941 ( .A(n408), .B(n3094), .Z(n3092) );
  XOR U6942 ( .A(n3095), .B(n3096), .Z(n3094) );
  XOR U6943 ( .A(DB[836]), .B(DB[805]), .Z(n3096) );
  AND U6944 ( .A(n412), .B(n3097), .Z(n3095) );
  XOR U6945 ( .A(n3098), .B(n3099), .Z(n3097) );
  XOR U6946 ( .A(DB[805]), .B(DB[774]), .Z(n3099) );
  AND U6947 ( .A(n416), .B(n3100), .Z(n3098) );
  XOR U6948 ( .A(n3101), .B(n3102), .Z(n3100) );
  XOR U6949 ( .A(DB[774]), .B(DB[743]), .Z(n3102) );
  AND U6950 ( .A(n420), .B(n3103), .Z(n3101) );
  XOR U6951 ( .A(n3104), .B(n3105), .Z(n3103) );
  XOR U6952 ( .A(DB[743]), .B(DB[712]), .Z(n3105) );
  AND U6953 ( .A(n424), .B(n3106), .Z(n3104) );
  XOR U6954 ( .A(n3107), .B(n3108), .Z(n3106) );
  XOR U6955 ( .A(DB[712]), .B(DB[681]), .Z(n3108) );
  AND U6956 ( .A(n428), .B(n3109), .Z(n3107) );
  XOR U6957 ( .A(n3110), .B(n3111), .Z(n3109) );
  XOR U6958 ( .A(DB[681]), .B(DB[650]), .Z(n3111) );
  AND U6959 ( .A(n432), .B(n3112), .Z(n3110) );
  XOR U6960 ( .A(n3113), .B(n3114), .Z(n3112) );
  XOR U6961 ( .A(DB[650]), .B(DB[619]), .Z(n3114) );
  AND U6962 ( .A(n436), .B(n3115), .Z(n3113) );
  XOR U6963 ( .A(n3116), .B(n3117), .Z(n3115) );
  XOR U6964 ( .A(DB[619]), .B(DB[588]), .Z(n3117) );
  AND U6965 ( .A(n440), .B(n3118), .Z(n3116) );
  XOR U6966 ( .A(n3119), .B(n3120), .Z(n3118) );
  XOR U6967 ( .A(DB[588]), .B(DB[557]), .Z(n3120) );
  AND U6968 ( .A(n444), .B(n3121), .Z(n3119) );
  XOR U6969 ( .A(n3122), .B(n3123), .Z(n3121) );
  XOR U6970 ( .A(DB[557]), .B(DB[526]), .Z(n3123) );
  AND U6971 ( .A(n448), .B(n3124), .Z(n3122) );
  XOR U6972 ( .A(n3125), .B(n3126), .Z(n3124) );
  XOR U6973 ( .A(DB[526]), .B(DB[495]), .Z(n3126) );
  AND U6974 ( .A(n452), .B(n3127), .Z(n3125) );
  XOR U6975 ( .A(n3128), .B(n3129), .Z(n3127) );
  XOR U6976 ( .A(DB[495]), .B(DB[464]), .Z(n3129) );
  AND U6977 ( .A(n456), .B(n3130), .Z(n3128) );
  XOR U6978 ( .A(n3131), .B(n3132), .Z(n3130) );
  XOR U6979 ( .A(DB[464]), .B(DB[433]), .Z(n3132) );
  AND U6980 ( .A(n460), .B(n3133), .Z(n3131) );
  XOR U6981 ( .A(n3134), .B(n3135), .Z(n3133) );
  XOR U6982 ( .A(DB[433]), .B(DB[402]), .Z(n3135) );
  AND U6983 ( .A(n464), .B(n3136), .Z(n3134) );
  XOR U6984 ( .A(n3137), .B(n3138), .Z(n3136) );
  XOR U6985 ( .A(DB[402]), .B(DB[371]), .Z(n3138) );
  AND U6986 ( .A(n468), .B(n3139), .Z(n3137) );
  XOR U6987 ( .A(n3140), .B(n3141), .Z(n3139) );
  XOR U6988 ( .A(DB[371]), .B(DB[340]), .Z(n3141) );
  AND U6989 ( .A(n472), .B(n3142), .Z(n3140) );
  XOR U6990 ( .A(n3143), .B(n3144), .Z(n3142) );
  XOR U6991 ( .A(DB[340]), .B(DB[309]), .Z(n3144) );
  AND U6992 ( .A(n476), .B(n3145), .Z(n3143) );
  XOR U6993 ( .A(n3146), .B(n3147), .Z(n3145) );
  XOR U6994 ( .A(DB[309]), .B(DB[278]), .Z(n3147) );
  AND U6995 ( .A(n480), .B(n3148), .Z(n3146) );
  XOR U6996 ( .A(n3149), .B(n3150), .Z(n3148) );
  XOR U6997 ( .A(DB[278]), .B(DB[247]), .Z(n3150) );
  AND U6998 ( .A(n484), .B(n3151), .Z(n3149) );
  XOR U6999 ( .A(n3152), .B(n3153), .Z(n3151) );
  XOR U7000 ( .A(DB[247]), .B(DB[216]), .Z(n3153) );
  AND U7001 ( .A(n488), .B(n3154), .Z(n3152) );
  XOR U7002 ( .A(n3155), .B(n3156), .Z(n3154) );
  XOR U7003 ( .A(DB[216]), .B(DB[185]), .Z(n3156) );
  AND U7004 ( .A(n492), .B(n3157), .Z(n3155) );
  XOR U7005 ( .A(n3158), .B(n3159), .Z(n3157) );
  XOR U7006 ( .A(DB[185]), .B(DB[154]), .Z(n3159) );
  AND U7007 ( .A(n496), .B(n3160), .Z(n3158) );
  XOR U7008 ( .A(n3161), .B(n3162), .Z(n3160) );
  XOR U7009 ( .A(DB[154]), .B(DB[123]), .Z(n3162) );
  AND U7010 ( .A(n500), .B(n3163), .Z(n3161) );
  XOR U7011 ( .A(n3164), .B(n3165), .Z(n3163) );
  XOR U7012 ( .A(DB[92]), .B(DB[123]), .Z(n3165) );
  AND U7013 ( .A(n504), .B(n3166), .Z(n3164) );
  XOR U7014 ( .A(n3167), .B(n3168), .Z(n3166) );
  XOR U7015 ( .A(DB[92]), .B(DB[61]), .Z(n3168) );
  AND U7016 ( .A(n508), .B(n3169), .Z(n3167) );
  XOR U7017 ( .A(DB[61]), .B(DB[30]), .Z(n3169) );
  XOR U7018 ( .A(DB[3939]), .B(n3170), .Z(min_val_out[2]) );
  AND U7019 ( .A(n2), .B(n3171), .Z(n3170) );
  XOR U7020 ( .A(n3172), .B(n3173), .Z(n3171) );
  XOR U7021 ( .A(DB[3939]), .B(DB[3908]), .Z(n3173) );
  AND U7022 ( .A(n8), .B(n3174), .Z(n3172) );
  XOR U7023 ( .A(n3175), .B(n3176), .Z(n3174) );
  XOR U7024 ( .A(DB[3908]), .B(DB[3877]), .Z(n3176) );
  AND U7025 ( .A(n12), .B(n3177), .Z(n3175) );
  XOR U7026 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U7027 ( .A(DB[3877]), .B(DB[3846]), .Z(n3179) );
  AND U7028 ( .A(n16), .B(n3180), .Z(n3178) );
  XOR U7029 ( .A(n3181), .B(n3182), .Z(n3180) );
  XOR U7030 ( .A(DB[3846]), .B(DB[3815]), .Z(n3182) );
  AND U7031 ( .A(n20), .B(n3183), .Z(n3181) );
  XOR U7032 ( .A(n3184), .B(n3185), .Z(n3183) );
  XOR U7033 ( .A(DB[3815]), .B(DB[3784]), .Z(n3185) );
  AND U7034 ( .A(n24), .B(n3186), .Z(n3184) );
  XOR U7035 ( .A(n3187), .B(n3188), .Z(n3186) );
  XOR U7036 ( .A(DB[3784]), .B(DB[3753]), .Z(n3188) );
  AND U7037 ( .A(n28), .B(n3189), .Z(n3187) );
  XOR U7038 ( .A(n3190), .B(n3191), .Z(n3189) );
  XOR U7039 ( .A(DB[3753]), .B(DB[3722]), .Z(n3191) );
  AND U7040 ( .A(n32), .B(n3192), .Z(n3190) );
  XOR U7041 ( .A(n3193), .B(n3194), .Z(n3192) );
  XOR U7042 ( .A(DB[3722]), .B(DB[3691]), .Z(n3194) );
  AND U7043 ( .A(n36), .B(n3195), .Z(n3193) );
  XOR U7044 ( .A(n3196), .B(n3197), .Z(n3195) );
  XOR U7045 ( .A(DB[3691]), .B(DB[3660]), .Z(n3197) );
  AND U7046 ( .A(n40), .B(n3198), .Z(n3196) );
  XOR U7047 ( .A(n3199), .B(n3200), .Z(n3198) );
  XOR U7048 ( .A(DB[3660]), .B(DB[3629]), .Z(n3200) );
  AND U7049 ( .A(n44), .B(n3201), .Z(n3199) );
  XOR U7050 ( .A(n3202), .B(n3203), .Z(n3201) );
  XOR U7051 ( .A(DB[3629]), .B(DB[3598]), .Z(n3203) );
  AND U7052 ( .A(n48), .B(n3204), .Z(n3202) );
  XOR U7053 ( .A(n3205), .B(n3206), .Z(n3204) );
  XOR U7054 ( .A(DB[3598]), .B(DB[3567]), .Z(n3206) );
  AND U7055 ( .A(n52), .B(n3207), .Z(n3205) );
  XOR U7056 ( .A(n3208), .B(n3209), .Z(n3207) );
  XOR U7057 ( .A(DB[3567]), .B(DB[3536]), .Z(n3209) );
  AND U7058 ( .A(n56), .B(n3210), .Z(n3208) );
  XOR U7059 ( .A(n3211), .B(n3212), .Z(n3210) );
  XOR U7060 ( .A(DB[3536]), .B(DB[3505]), .Z(n3212) );
  AND U7061 ( .A(n60), .B(n3213), .Z(n3211) );
  XOR U7062 ( .A(n3214), .B(n3215), .Z(n3213) );
  XOR U7063 ( .A(DB[3505]), .B(DB[3474]), .Z(n3215) );
  AND U7064 ( .A(n64), .B(n3216), .Z(n3214) );
  XOR U7065 ( .A(n3217), .B(n3218), .Z(n3216) );
  XOR U7066 ( .A(DB[3474]), .B(DB[3443]), .Z(n3218) );
  AND U7067 ( .A(n68), .B(n3219), .Z(n3217) );
  XOR U7068 ( .A(n3220), .B(n3221), .Z(n3219) );
  XOR U7069 ( .A(DB[3443]), .B(DB[3412]), .Z(n3221) );
  AND U7070 ( .A(n72), .B(n3222), .Z(n3220) );
  XOR U7071 ( .A(n3223), .B(n3224), .Z(n3222) );
  XOR U7072 ( .A(DB[3412]), .B(DB[3381]), .Z(n3224) );
  AND U7073 ( .A(n76), .B(n3225), .Z(n3223) );
  XOR U7074 ( .A(n3226), .B(n3227), .Z(n3225) );
  XOR U7075 ( .A(DB[3381]), .B(DB[3350]), .Z(n3227) );
  AND U7076 ( .A(n80), .B(n3228), .Z(n3226) );
  XOR U7077 ( .A(n3229), .B(n3230), .Z(n3228) );
  XOR U7078 ( .A(DB[3350]), .B(DB[3319]), .Z(n3230) );
  AND U7079 ( .A(n84), .B(n3231), .Z(n3229) );
  XOR U7080 ( .A(n3232), .B(n3233), .Z(n3231) );
  XOR U7081 ( .A(DB[3319]), .B(DB[3288]), .Z(n3233) );
  AND U7082 ( .A(n88), .B(n3234), .Z(n3232) );
  XOR U7083 ( .A(n3235), .B(n3236), .Z(n3234) );
  XOR U7084 ( .A(DB[3288]), .B(DB[3257]), .Z(n3236) );
  AND U7085 ( .A(n92), .B(n3237), .Z(n3235) );
  XOR U7086 ( .A(n3238), .B(n3239), .Z(n3237) );
  XOR U7087 ( .A(DB[3257]), .B(DB[3226]), .Z(n3239) );
  AND U7088 ( .A(n96), .B(n3240), .Z(n3238) );
  XOR U7089 ( .A(n3241), .B(n3242), .Z(n3240) );
  XOR U7090 ( .A(DB[3226]), .B(DB[3195]), .Z(n3242) );
  AND U7091 ( .A(n100), .B(n3243), .Z(n3241) );
  XOR U7092 ( .A(n3244), .B(n3245), .Z(n3243) );
  XOR U7093 ( .A(DB[3195]), .B(DB[3164]), .Z(n3245) );
  AND U7094 ( .A(n104), .B(n3246), .Z(n3244) );
  XOR U7095 ( .A(n3247), .B(n3248), .Z(n3246) );
  XOR U7096 ( .A(DB[3164]), .B(DB[3133]), .Z(n3248) );
  AND U7097 ( .A(n108), .B(n3249), .Z(n3247) );
  XOR U7098 ( .A(n3250), .B(n3251), .Z(n3249) );
  XOR U7099 ( .A(DB[3133]), .B(DB[3102]), .Z(n3251) );
  AND U7100 ( .A(n112), .B(n3252), .Z(n3250) );
  XOR U7101 ( .A(n3253), .B(n3254), .Z(n3252) );
  XOR U7102 ( .A(DB[3102]), .B(DB[3071]), .Z(n3254) );
  AND U7103 ( .A(n116), .B(n3255), .Z(n3253) );
  XOR U7104 ( .A(n3256), .B(n3257), .Z(n3255) );
  XOR U7105 ( .A(DB[3071]), .B(DB[3040]), .Z(n3257) );
  AND U7106 ( .A(n120), .B(n3258), .Z(n3256) );
  XOR U7107 ( .A(n3259), .B(n3260), .Z(n3258) );
  XOR U7108 ( .A(DB[3040]), .B(DB[3009]), .Z(n3260) );
  AND U7109 ( .A(n124), .B(n3261), .Z(n3259) );
  XOR U7110 ( .A(n3262), .B(n3263), .Z(n3261) );
  XOR U7111 ( .A(DB[3009]), .B(DB[2978]), .Z(n3263) );
  AND U7112 ( .A(n128), .B(n3264), .Z(n3262) );
  XOR U7113 ( .A(n3265), .B(n3266), .Z(n3264) );
  XOR U7114 ( .A(DB[2978]), .B(DB[2947]), .Z(n3266) );
  AND U7115 ( .A(n132), .B(n3267), .Z(n3265) );
  XOR U7116 ( .A(n3268), .B(n3269), .Z(n3267) );
  XOR U7117 ( .A(DB[2947]), .B(DB[2916]), .Z(n3269) );
  AND U7118 ( .A(n136), .B(n3270), .Z(n3268) );
  XOR U7119 ( .A(n3271), .B(n3272), .Z(n3270) );
  XOR U7120 ( .A(DB[2916]), .B(DB[2885]), .Z(n3272) );
  AND U7121 ( .A(n140), .B(n3273), .Z(n3271) );
  XOR U7122 ( .A(n3274), .B(n3275), .Z(n3273) );
  XOR U7123 ( .A(DB[2885]), .B(DB[2854]), .Z(n3275) );
  AND U7124 ( .A(n144), .B(n3276), .Z(n3274) );
  XOR U7125 ( .A(n3277), .B(n3278), .Z(n3276) );
  XOR U7126 ( .A(DB[2854]), .B(DB[2823]), .Z(n3278) );
  AND U7127 ( .A(n148), .B(n3279), .Z(n3277) );
  XOR U7128 ( .A(n3280), .B(n3281), .Z(n3279) );
  XOR U7129 ( .A(DB[2823]), .B(DB[2792]), .Z(n3281) );
  AND U7130 ( .A(n152), .B(n3282), .Z(n3280) );
  XOR U7131 ( .A(n3283), .B(n3284), .Z(n3282) );
  XOR U7132 ( .A(DB[2792]), .B(DB[2761]), .Z(n3284) );
  AND U7133 ( .A(n156), .B(n3285), .Z(n3283) );
  XOR U7134 ( .A(n3286), .B(n3287), .Z(n3285) );
  XOR U7135 ( .A(DB[2761]), .B(DB[2730]), .Z(n3287) );
  AND U7136 ( .A(n160), .B(n3288), .Z(n3286) );
  XOR U7137 ( .A(n3289), .B(n3290), .Z(n3288) );
  XOR U7138 ( .A(DB[2730]), .B(DB[2699]), .Z(n3290) );
  AND U7139 ( .A(n164), .B(n3291), .Z(n3289) );
  XOR U7140 ( .A(n3292), .B(n3293), .Z(n3291) );
  XOR U7141 ( .A(DB[2699]), .B(DB[2668]), .Z(n3293) );
  AND U7142 ( .A(n168), .B(n3294), .Z(n3292) );
  XOR U7143 ( .A(n3295), .B(n3296), .Z(n3294) );
  XOR U7144 ( .A(DB[2668]), .B(DB[2637]), .Z(n3296) );
  AND U7145 ( .A(n172), .B(n3297), .Z(n3295) );
  XOR U7146 ( .A(n3298), .B(n3299), .Z(n3297) );
  XOR U7147 ( .A(DB[2637]), .B(DB[2606]), .Z(n3299) );
  AND U7148 ( .A(n176), .B(n3300), .Z(n3298) );
  XOR U7149 ( .A(n3301), .B(n3302), .Z(n3300) );
  XOR U7150 ( .A(DB[2606]), .B(DB[2575]), .Z(n3302) );
  AND U7151 ( .A(n180), .B(n3303), .Z(n3301) );
  XOR U7152 ( .A(n3304), .B(n3305), .Z(n3303) );
  XOR U7153 ( .A(DB[2575]), .B(DB[2544]), .Z(n3305) );
  AND U7154 ( .A(n184), .B(n3306), .Z(n3304) );
  XOR U7155 ( .A(n3307), .B(n3308), .Z(n3306) );
  XOR U7156 ( .A(DB[2544]), .B(DB[2513]), .Z(n3308) );
  AND U7157 ( .A(n188), .B(n3309), .Z(n3307) );
  XOR U7158 ( .A(n3310), .B(n3311), .Z(n3309) );
  XOR U7159 ( .A(DB[2513]), .B(DB[2482]), .Z(n3311) );
  AND U7160 ( .A(n192), .B(n3312), .Z(n3310) );
  XOR U7161 ( .A(n3313), .B(n3314), .Z(n3312) );
  XOR U7162 ( .A(DB[2482]), .B(DB[2451]), .Z(n3314) );
  AND U7163 ( .A(n196), .B(n3315), .Z(n3313) );
  XOR U7164 ( .A(n3316), .B(n3317), .Z(n3315) );
  XOR U7165 ( .A(DB[2451]), .B(DB[2420]), .Z(n3317) );
  AND U7166 ( .A(n200), .B(n3318), .Z(n3316) );
  XOR U7167 ( .A(n3319), .B(n3320), .Z(n3318) );
  XOR U7168 ( .A(DB[2420]), .B(DB[2389]), .Z(n3320) );
  AND U7169 ( .A(n204), .B(n3321), .Z(n3319) );
  XOR U7170 ( .A(n3322), .B(n3323), .Z(n3321) );
  XOR U7171 ( .A(DB[2389]), .B(DB[2358]), .Z(n3323) );
  AND U7172 ( .A(n208), .B(n3324), .Z(n3322) );
  XOR U7173 ( .A(n3325), .B(n3326), .Z(n3324) );
  XOR U7174 ( .A(DB[2358]), .B(DB[2327]), .Z(n3326) );
  AND U7175 ( .A(n212), .B(n3327), .Z(n3325) );
  XOR U7176 ( .A(n3328), .B(n3329), .Z(n3327) );
  XOR U7177 ( .A(DB[2327]), .B(DB[2296]), .Z(n3329) );
  AND U7178 ( .A(n216), .B(n3330), .Z(n3328) );
  XOR U7179 ( .A(n3331), .B(n3332), .Z(n3330) );
  XOR U7180 ( .A(DB[2296]), .B(DB[2265]), .Z(n3332) );
  AND U7181 ( .A(n220), .B(n3333), .Z(n3331) );
  XOR U7182 ( .A(n3334), .B(n3335), .Z(n3333) );
  XOR U7183 ( .A(DB[2265]), .B(DB[2234]), .Z(n3335) );
  AND U7184 ( .A(n224), .B(n3336), .Z(n3334) );
  XOR U7185 ( .A(n3337), .B(n3338), .Z(n3336) );
  XOR U7186 ( .A(DB[2234]), .B(DB[2203]), .Z(n3338) );
  AND U7187 ( .A(n228), .B(n3339), .Z(n3337) );
  XOR U7188 ( .A(n3340), .B(n3341), .Z(n3339) );
  XOR U7189 ( .A(DB[2203]), .B(DB[2172]), .Z(n3341) );
  AND U7190 ( .A(n232), .B(n3342), .Z(n3340) );
  XOR U7191 ( .A(n3343), .B(n3344), .Z(n3342) );
  XOR U7192 ( .A(DB[2172]), .B(DB[2141]), .Z(n3344) );
  AND U7193 ( .A(n236), .B(n3345), .Z(n3343) );
  XOR U7194 ( .A(n3346), .B(n3347), .Z(n3345) );
  XOR U7195 ( .A(DB[2141]), .B(DB[2110]), .Z(n3347) );
  AND U7196 ( .A(n240), .B(n3348), .Z(n3346) );
  XOR U7197 ( .A(n3349), .B(n3350), .Z(n3348) );
  XOR U7198 ( .A(DB[2110]), .B(DB[2079]), .Z(n3350) );
  AND U7199 ( .A(n244), .B(n3351), .Z(n3349) );
  XOR U7200 ( .A(n3352), .B(n3353), .Z(n3351) );
  XOR U7201 ( .A(DB[2079]), .B(DB[2048]), .Z(n3353) );
  AND U7202 ( .A(n248), .B(n3354), .Z(n3352) );
  XOR U7203 ( .A(n3355), .B(n3356), .Z(n3354) );
  XOR U7204 ( .A(DB[2048]), .B(DB[2017]), .Z(n3356) );
  AND U7205 ( .A(n252), .B(n3357), .Z(n3355) );
  XOR U7206 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR U7207 ( .A(DB[2017]), .B(DB[1986]), .Z(n3359) );
  AND U7208 ( .A(n256), .B(n3360), .Z(n3358) );
  XOR U7209 ( .A(n3361), .B(n3362), .Z(n3360) );
  XOR U7210 ( .A(DB[1986]), .B(DB[1955]), .Z(n3362) );
  AND U7211 ( .A(n260), .B(n3363), .Z(n3361) );
  XOR U7212 ( .A(n3364), .B(n3365), .Z(n3363) );
  XOR U7213 ( .A(DB[1955]), .B(DB[1924]), .Z(n3365) );
  AND U7214 ( .A(n264), .B(n3366), .Z(n3364) );
  XOR U7215 ( .A(n3367), .B(n3368), .Z(n3366) );
  XOR U7216 ( .A(DB[1924]), .B(DB[1893]), .Z(n3368) );
  AND U7217 ( .A(n268), .B(n3369), .Z(n3367) );
  XOR U7218 ( .A(n3370), .B(n3371), .Z(n3369) );
  XOR U7219 ( .A(DB[1893]), .B(DB[1862]), .Z(n3371) );
  AND U7220 ( .A(n272), .B(n3372), .Z(n3370) );
  XOR U7221 ( .A(n3373), .B(n3374), .Z(n3372) );
  XOR U7222 ( .A(DB[1862]), .B(DB[1831]), .Z(n3374) );
  AND U7223 ( .A(n276), .B(n3375), .Z(n3373) );
  XOR U7224 ( .A(n3376), .B(n3377), .Z(n3375) );
  XOR U7225 ( .A(DB[1831]), .B(DB[1800]), .Z(n3377) );
  AND U7226 ( .A(n280), .B(n3378), .Z(n3376) );
  XOR U7227 ( .A(n3379), .B(n3380), .Z(n3378) );
  XOR U7228 ( .A(DB[1800]), .B(DB[1769]), .Z(n3380) );
  AND U7229 ( .A(n284), .B(n3381), .Z(n3379) );
  XOR U7230 ( .A(n3382), .B(n3383), .Z(n3381) );
  XOR U7231 ( .A(DB[1769]), .B(DB[1738]), .Z(n3383) );
  AND U7232 ( .A(n288), .B(n3384), .Z(n3382) );
  XOR U7233 ( .A(n3385), .B(n3386), .Z(n3384) );
  XOR U7234 ( .A(DB[1738]), .B(DB[1707]), .Z(n3386) );
  AND U7235 ( .A(n292), .B(n3387), .Z(n3385) );
  XOR U7236 ( .A(n3388), .B(n3389), .Z(n3387) );
  XOR U7237 ( .A(DB[1707]), .B(DB[1676]), .Z(n3389) );
  AND U7238 ( .A(n296), .B(n3390), .Z(n3388) );
  XOR U7239 ( .A(n3391), .B(n3392), .Z(n3390) );
  XOR U7240 ( .A(DB[1676]), .B(DB[1645]), .Z(n3392) );
  AND U7241 ( .A(n300), .B(n3393), .Z(n3391) );
  XOR U7242 ( .A(n3394), .B(n3395), .Z(n3393) );
  XOR U7243 ( .A(DB[1645]), .B(DB[1614]), .Z(n3395) );
  AND U7244 ( .A(n304), .B(n3396), .Z(n3394) );
  XOR U7245 ( .A(n3397), .B(n3398), .Z(n3396) );
  XOR U7246 ( .A(DB[1614]), .B(DB[1583]), .Z(n3398) );
  AND U7247 ( .A(n308), .B(n3399), .Z(n3397) );
  XOR U7248 ( .A(n3400), .B(n3401), .Z(n3399) );
  XOR U7249 ( .A(DB[1583]), .B(DB[1552]), .Z(n3401) );
  AND U7250 ( .A(n312), .B(n3402), .Z(n3400) );
  XOR U7251 ( .A(n3403), .B(n3404), .Z(n3402) );
  XOR U7252 ( .A(DB[1552]), .B(DB[1521]), .Z(n3404) );
  AND U7253 ( .A(n316), .B(n3405), .Z(n3403) );
  XOR U7254 ( .A(n3406), .B(n3407), .Z(n3405) );
  XOR U7255 ( .A(DB[1521]), .B(DB[1490]), .Z(n3407) );
  AND U7256 ( .A(n320), .B(n3408), .Z(n3406) );
  XOR U7257 ( .A(n3409), .B(n3410), .Z(n3408) );
  XOR U7258 ( .A(DB[1490]), .B(DB[1459]), .Z(n3410) );
  AND U7259 ( .A(n324), .B(n3411), .Z(n3409) );
  XOR U7260 ( .A(n3412), .B(n3413), .Z(n3411) );
  XOR U7261 ( .A(DB[1459]), .B(DB[1428]), .Z(n3413) );
  AND U7262 ( .A(n328), .B(n3414), .Z(n3412) );
  XOR U7263 ( .A(n3415), .B(n3416), .Z(n3414) );
  XOR U7264 ( .A(DB[1428]), .B(DB[1397]), .Z(n3416) );
  AND U7265 ( .A(n332), .B(n3417), .Z(n3415) );
  XOR U7266 ( .A(n3418), .B(n3419), .Z(n3417) );
  XOR U7267 ( .A(DB[1397]), .B(DB[1366]), .Z(n3419) );
  AND U7268 ( .A(n336), .B(n3420), .Z(n3418) );
  XOR U7269 ( .A(n3421), .B(n3422), .Z(n3420) );
  XOR U7270 ( .A(DB[1366]), .B(DB[1335]), .Z(n3422) );
  AND U7271 ( .A(n340), .B(n3423), .Z(n3421) );
  XOR U7272 ( .A(n3424), .B(n3425), .Z(n3423) );
  XOR U7273 ( .A(DB[1335]), .B(DB[1304]), .Z(n3425) );
  AND U7274 ( .A(n344), .B(n3426), .Z(n3424) );
  XOR U7275 ( .A(n3427), .B(n3428), .Z(n3426) );
  XOR U7276 ( .A(DB[1304]), .B(DB[1273]), .Z(n3428) );
  AND U7277 ( .A(n348), .B(n3429), .Z(n3427) );
  XOR U7278 ( .A(n3430), .B(n3431), .Z(n3429) );
  XOR U7279 ( .A(DB[1273]), .B(DB[1242]), .Z(n3431) );
  AND U7280 ( .A(n352), .B(n3432), .Z(n3430) );
  XOR U7281 ( .A(n3433), .B(n3434), .Z(n3432) );
  XOR U7282 ( .A(DB[1242]), .B(DB[1211]), .Z(n3434) );
  AND U7283 ( .A(n356), .B(n3435), .Z(n3433) );
  XOR U7284 ( .A(n3436), .B(n3437), .Z(n3435) );
  XOR U7285 ( .A(DB[1211]), .B(DB[1180]), .Z(n3437) );
  AND U7286 ( .A(n360), .B(n3438), .Z(n3436) );
  XOR U7287 ( .A(n3439), .B(n3440), .Z(n3438) );
  XOR U7288 ( .A(DB[1180]), .B(DB[1149]), .Z(n3440) );
  AND U7289 ( .A(n364), .B(n3441), .Z(n3439) );
  XOR U7290 ( .A(n3442), .B(n3443), .Z(n3441) );
  XOR U7291 ( .A(DB[1149]), .B(DB[1118]), .Z(n3443) );
  AND U7292 ( .A(n368), .B(n3444), .Z(n3442) );
  XOR U7293 ( .A(n3445), .B(n3446), .Z(n3444) );
  XOR U7294 ( .A(DB[1118]), .B(DB[1087]), .Z(n3446) );
  AND U7295 ( .A(n372), .B(n3447), .Z(n3445) );
  XOR U7296 ( .A(n3448), .B(n3449), .Z(n3447) );
  XOR U7297 ( .A(DB[1087]), .B(DB[1056]), .Z(n3449) );
  AND U7298 ( .A(n376), .B(n3450), .Z(n3448) );
  XOR U7299 ( .A(n3451), .B(n3452), .Z(n3450) );
  XOR U7300 ( .A(DB[1056]), .B(DB[1025]), .Z(n3452) );
  AND U7301 ( .A(n380), .B(n3453), .Z(n3451) );
  XOR U7302 ( .A(n3454), .B(n3455), .Z(n3453) );
  XOR U7303 ( .A(DB[994]), .B(DB[1025]), .Z(n3455) );
  AND U7304 ( .A(n384), .B(n3456), .Z(n3454) );
  XOR U7305 ( .A(n3457), .B(n3458), .Z(n3456) );
  XOR U7306 ( .A(DB[994]), .B(DB[963]), .Z(n3458) );
  AND U7307 ( .A(n388), .B(n3459), .Z(n3457) );
  XOR U7308 ( .A(n3460), .B(n3461), .Z(n3459) );
  XOR U7309 ( .A(DB[963]), .B(DB[932]), .Z(n3461) );
  AND U7310 ( .A(n392), .B(n3462), .Z(n3460) );
  XOR U7311 ( .A(n3463), .B(n3464), .Z(n3462) );
  XOR U7312 ( .A(DB[932]), .B(DB[901]), .Z(n3464) );
  AND U7313 ( .A(n396), .B(n3465), .Z(n3463) );
  XOR U7314 ( .A(n3466), .B(n3467), .Z(n3465) );
  XOR U7315 ( .A(DB[901]), .B(DB[870]), .Z(n3467) );
  AND U7316 ( .A(n400), .B(n3468), .Z(n3466) );
  XOR U7317 ( .A(n3469), .B(n3470), .Z(n3468) );
  XOR U7318 ( .A(DB[870]), .B(DB[839]), .Z(n3470) );
  AND U7319 ( .A(n404), .B(n3471), .Z(n3469) );
  XOR U7320 ( .A(n3472), .B(n3473), .Z(n3471) );
  XOR U7321 ( .A(DB[839]), .B(DB[808]), .Z(n3473) );
  AND U7322 ( .A(n408), .B(n3474), .Z(n3472) );
  XOR U7323 ( .A(n3475), .B(n3476), .Z(n3474) );
  XOR U7324 ( .A(DB[808]), .B(DB[777]), .Z(n3476) );
  AND U7325 ( .A(n412), .B(n3477), .Z(n3475) );
  XOR U7326 ( .A(n3478), .B(n3479), .Z(n3477) );
  XOR U7327 ( .A(DB[777]), .B(DB[746]), .Z(n3479) );
  AND U7328 ( .A(n416), .B(n3480), .Z(n3478) );
  XOR U7329 ( .A(n3481), .B(n3482), .Z(n3480) );
  XOR U7330 ( .A(DB[746]), .B(DB[715]), .Z(n3482) );
  AND U7331 ( .A(n420), .B(n3483), .Z(n3481) );
  XOR U7332 ( .A(n3484), .B(n3485), .Z(n3483) );
  XOR U7333 ( .A(DB[715]), .B(DB[684]), .Z(n3485) );
  AND U7334 ( .A(n424), .B(n3486), .Z(n3484) );
  XOR U7335 ( .A(n3487), .B(n3488), .Z(n3486) );
  XOR U7336 ( .A(DB[684]), .B(DB[653]), .Z(n3488) );
  AND U7337 ( .A(n428), .B(n3489), .Z(n3487) );
  XOR U7338 ( .A(n3490), .B(n3491), .Z(n3489) );
  XOR U7339 ( .A(DB[653]), .B(DB[622]), .Z(n3491) );
  AND U7340 ( .A(n432), .B(n3492), .Z(n3490) );
  XOR U7341 ( .A(n3493), .B(n3494), .Z(n3492) );
  XOR U7342 ( .A(DB[622]), .B(DB[591]), .Z(n3494) );
  AND U7343 ( .A(n436), .B(n3495), .Z(n3493) );
  XOR U7344 ( .A(n3496), .B(n3497), .Z(n3495) );
  XOR U7345 ( .A(DB[591]), .B(DB[560]), .Z(n3497) );
  AND U7346 ( .A(n440), .B(n3498), .Z(n3496) );
  XOR U7347 ( .A(n3499), .B(n3500), .Z(n3498) );
  XOR U7348 ( .A(DB[560]), .B(DB[529]), .Z(n3500) );
  AND U7349 ( .A(n444), .B(n3501), .Z(n3499) );
  XOR U7350 ( .A(n3502), .B(n3503), .Z(n3501) );
  XOR U7351 ( .A(DB[529]), .B(DB[498]), .Z(n3503) );
  AND U7352 ( .A(n448), .B(n3504), .Z(n3502) );
  XOR U7353 ( .A(n3505), .B(n3506), .Z(n3504) );
  XOR U7354 ( .A(DB[498]), .B(DB[467]), .Z(n3506) );
  AND U7355 ( .A(n452), .B(n3507), .Z(n3505) );
  XOR U7356 ( .A(n3508), .B(n3509), .Z(n3507) );
  XOR U7357 ( .A(DB[467]), .B(DB[436]), .Z(n3509) );
  AND U7358 ( .A(n456), .B(n3510), .Z(n3508) );
  XOR U7359 ( .A(n3511), .B(n3512), .Z(n3510) );
  XOR U7360 ( .A(DB[436]), .B(DB[405]), .Z(n3512) );
  AND U7361 ( .A(n460), .B(n3513), .Z(n3511) );
  XOR U7362 ( .A(n3514), .B(n3515), .Z(n3513) );
  XOR U7363 ( .A(DB[405]), .B(DB[374]), .Z(n3515) );
  AND U7364 ( .A(n464), .B(n3516), .Z(n3514) );
  XOR U7365 ( .A(n3517), .B(n3518), .Z(n3516) );
  XOR U7366 ( .A(DB[374]), .B(DB[343]), .Z(n3518) );
  AND U7367 ( .A(n468), .B(n3519), .Z(n3517) );
  XOR U7368 ( .A(n3520), .B(n3521), .Z(n3519) );
  XOR U7369 ( .A(DB[343]), .B(DB[312]), .Z(n3521) );
  AND U7370 ( .A(n472), .B(n3522), .Z(n3520) );
  XOR U7371 ( .A(n3523), .B(n3524), .Z(n3522) );
  XOR U7372 ( .A(DB[312]), .B(DB[281]), .Z(n3524) );
  AND U7373 ( .A(n476), .B(n3525), .Z(n3523) );
  XOR U7374 ( .A(n3526), .B(n3527), .Z(n3525) );
  XOR U7375 ( .A(DB[281]), .B(DB[250]), .Z(n3527) );
  AND U7376 ( .A(n480), .B(n3528), .Z(n3526) );
  XOR U7377 ( .A(n3529), .B(n3530), .Z(n3528) );
  XOR U7378 ( .A(DB[250]), .B(DB[219]), .Z(n3530) );
  AND U7379 ( .A(n484), .B(n3531), .Z(n3529) );
  XOR U7380 ( .A(n3532), .B(n3533), .Z(n3531) );
  XOR U7381 ( .A(DB[219]), .B(DB[188]), .Z(n3533) );
  AND U7382 ( .A(n488), .B(n3534), .Z(n3532) );
  XOR U7383 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U7384 ( .A(DB[188]), .B(DB[157]), .Z(n3536) );
  AND U7385 ( .A(n492), .B(n3537), .Z(n3535) );
  XOR U7386 ( .A(n3538), .B(n3539), .Z(n3537) );
  XOR U7387 ( .A(DB[157]), .B(DB[126]), .Z(n3539) );
  AND U7388 ( .A(n496), .B(n3540), .Z(n3538) );
  XOR U7389 ( .A(n3541), .B(n3542), .Z(n3540) );
  XOR U7390 ( .A(DB[95]), .B(DB[126]), .Z(n3542) );
  AND U7391 ( .A(n500), .B(n3543), .Z(n3541) );
  XOR U7392 ( .A(n3544), .B(n3545), .Z(n3543) );
  XOR U7393 ( .A(DB[95]), .B(DB[64]), .Z(n3545) );
  AND U7394 ( .A(n504), .B(n3546), .Z(n3544) );
  XOR U7395 ( .A(n3547), .B(n3548), .Z(n3546) );
  XOR U7396 ( .A(DB[64]), .B(DB[33]), .Z(n3548) );
  AND U7397 ( .A(n508), .B(n3549), .Z(n3547) );
  XOR U7398 ( .A(DB[33]), .B(DB[2]), .Z(n3549) );
  XOR U7399 ( .A(DB[3966]), .B(n3550), .Z(min_val_out[29]) );
  AND U7400 ( .A(n2), .B(n3551), .Z(n3550) );
  XOR U7401 ( .A(n3552), .B(n3553), .Z(n3551) );
  XOR U7402 ( .A(DB[3966]), .B(DB[3935]), .Z(n3553) );
  AND U7403 ( .A(n8), .B(n3554), .Z(n3552) );
  XOR U7404 ( .A(n3555), .B(n3556), .Z(n3554) );
  XOR U7405 ( .A(DB[3935]), .B(DB[3904]), .Z(n3556) );
  AND U7406 ( .A(n12), .B(n3557), .Z(n3555) );
  XOR U7407 ( .A(n3558), .B(n3559), .Z(n3557) );
  XOR U7408 ( .A(DB[3904]), .B(DB[3873]), .Z(n3559) );
  AND U7409 ( .A(n16), .B(n3560), .Z(n3558) );
  XOR U7410 ( .A(n3561), .B(n3562), .Z(n3560) );
  XOR U7411 ( .A(DB[3873]), .B(DB[3842]), .Z(n3562) );
  AND U7412 ( .A(n20), .B(n3563), .Z(n3561) );
  XOR U7413 ( .A(n3564), .B(n3565), .Z(n3563) );
  XOR U7414 ( .A(DB[3842]), .B(DB[3811]), .Z(n3565) );
  AND U7415 ( .A(n24), .B(n3566), .Z(n3564) );
  XOR U7416 ( .A(n3567), .B(n3568), .Z(n3566) );
  XOR U7417 ( .A(DB[3811]), .B(DB[3780]), .Z(n3568) );
  AND U7418 ( .A(n28), .B(n3569), .Z(n3567) );
  XOR U7419 ( .A(n3570), .B(n3571), .Z(n3569) );
  XOR U7420 ( .A(DB[3780]), .B(DB[3749]), .Z(n3571) );
  AND U7421 ( .A(n32), .B(n3572), .Z(n3570) );
  XOR U7422 ( .A(n3573), .B(n3574), .Z(n3572) );
  XOR U7423 ( .A(DB[3749]), .B(DB[3718]), .Z(n3574) );
  AND U7424 ( .A(n36), .B(n3575), .Z(n3573) );
  XOR U7425 ( .A(n3576), .B(n3577), .Z(n3575) );
  XOR U7426 ( .A(DB[3718]), .B(DB[3687]), .Z(n3577) );
  AND U7427 ( .A(n40), .B(n3578), .Z(n3576) );
  XOR U7428 ( .A(n3579), .B(n3580), .Z(n3578) );
  XOR U7429 ( .A(DB[3687]), .B(DB[3656]), .Z(n3580) );
  AND U7430 ( .A(n44), .B(n3581), .Z(n3579) );
  XOR U7431 ( .A(n3582), .B(n3583), .Z(n3581) );
  XOR U7432 ( .A(DB[3656]), .B(DB[3625]), .Z(n3583) );
  AND U7433 ( .A(n48), .B(n3584), .Z(n3582) );
  XOR U7434 ( .A(n3585), .B(n3586), .Z(n3584) );
  XOR U7435 ( .A(DB[3625]), .B(DB[3594]), .Z(n3586) );
  AND U7436 ( .A(n52), .B(n3587), .Z(n3585) );
  XOR U7437 ( .A(n3588), .B(n3589), .Z(n3587) );
  XOR U7438 ( .A(DB[3594]), .B(DB[3563]), .Z(n3589) );
  AND U7439 ( .A(n56), .B(n3590), .Z(n3588) );
  XOR U7440 ( .A(n3591), .B(n3592), .Z(n3590) );
  XOR U7441 ( .A(DB[3563]), .B(DB[3532]), .Z(n3592) );
  AND U7442 ( .A(n60), .B(n3593), .Z(n3591) );
  XOR U7443 ( .A(n3594), .B(n3595), .Z(n3593) );
  XOR U7444 ( .A(DB[3532]), .B(DB[3501]), .Z(n3595) );
  AND U7445 ( .A(n64), .B(n3596), .Z(n3594) );
  XOR U7446 ( .A(n3597), .B(n3598), .Z(n3596) );
  XOR U7447 ( .A(DB[3501]), .B(DB[3470]), .Z(n3598) );
  AND U7448 ( .A(n68), .B(n3599), .Z(n3597) );
  XOR U7449 ( .A(n3600), .B(n3601), .Z(n3599) );
  XOR U7450 ( .A(DB[3470]), .B(DB[3439]), .Z(n3601) );
  AND U7451 ( .A(n72), .B(n3602), .Z(n3600) );
  XOR U7452 ( .A(n3603), .B(n3604), .Z(n3602) );
  XOR U7453 ( .A(DB[3439]), .B(DB[3408]), .Z(n3604) );
  AND U7454 ( .A(n76), .B(n3605), .Z(n3603) );
  XOR U7455 ( .A(n3606), .B(n3607), .Z(n3605) );
  XOR U7456 ( .A(DB[3408]), .B(DB[3377]), .Z(n3607) );
  AND U7457 ( .A(n80), .B(n3608), .Z(n3606) );
  XOR U7458 ( .A(n3609), .B(n3610), .Z(n3608) );
  XOR U7459 ( .A(DB[3377]), .B(DB[3346]), .Z(n3610) );
  AND U7460 ( .A(n84), .B(n3611), .Z(n3609) );
  XOR U7461 ( .A(n3612), .B(n3613), .Z(n3611) );
  XOR U7462 ( .A(DB[3346]), .B(DB[3315]), .Z(n3613) );
  AND U7463 ( .A(n88), .B(n3614), .Z(n3612) );
  XOR U7464 ( .A(n3615), .B(n3616), .Z(n3614) );
  XOR U7465 ( .A(DB[3315]), .B(DB[3284]), .Z(n3616) );
  AND U7466 ( .A(n92), .B(n3617), .Z(n3615) );
  XOR U7467 ( .A(n3618), .B(n3619), .Z(n3617) );
  XOR U7468 ( .A(DB[3284]), .B(DB[3253]), .Z(n3619) );
  AND U7469 ( .A(n96), .B(n3620), .Z(n3618) );
  XOR U7470 ( .A(n3621), .B(n3622), .Z(n3620) );
  XOR U7471 ( .A(DB[3253]), .B(DB[3222]), .Z(n3622) );
  AND U7472 ( .A(n100), .B(n3623), .Z(n3621) );
  XOR U7473 ( .A(n3624), .B(n3625), .Z(n3623) );
  XOR U7474 ( .A(DB[3222]), .B(DB[3191]), .Z(n3625) );
  AND U7475 ( .A(n104), .B(n3626), .Z(n3624) );
  XOR U7476 ( .A(n3627), .B(n3628), .Z(n3626) );
  XOR U7477 ( .A(DB[3191]), .B(DB[3160]), .Z(n3628) );
  AND U7478 ( .A(n108), .B(n3629), .Z(n3627) );
  XOR U7479 ( .A(n3630), .B(n3631), .Z(n3629) );
  XOR U7480 ( .A(DB[3160]), .B(DB[3129]), .Z(n3631) );
  AND U7481 ( .A(n112), .B(n3632), .Z(n3630) );
  XOR U7482 ( .A(n3633), .B(n3634), .Z(n3632) );
  XOR U7483 ( .A(DB[3129]), .B(DB[3098]), .Z(n3634) );
  AND U7484 ( .A(n116), .B(n3635), .Z(n3633) );
  XOR U7485 ( .A(n3636), .B(n3637), .Z(n3635) );
  XOR U7486 ( .A(DB[3098]), .B(DB[3067]), .Z(n3637) );
  AND U7487 ( .A(n120), .B(n3638), .Z(n3636) );
  XOR U7488 ( .A(n3639), .B(n3640), .Z(n3638) );
  XOR U7489 ( .A(DB[3067]), .B(DB[3036]), .Z(n3640) );
  AND U7490 ( .A(n124), .B(n3641), .Z(n3639) );
  XOR U7491 ( .A(n3642), .B(n3643), .Z(n3641) );
  XOR U7492 ( .A(DB[3036]), .B(DB[3005]), .Z(n3643) );
  AND U7493 ( .A(n128), .B(n3644), .Z(n3642) );
  XOR U7494 ( .A(n3645), .B(n3646), .Z(n3644) );
  XOR U7495 ( .A(DB[3005]), .B(DB[2974]), .Z(n3646) );
  AND U7496 ( .A(n132), .B(n3647), .Z(n3645) );
  XOR U7497 ( .A(n3648), .B(n3649), .Z(n3647) );
  XOR U7498 ( .A(DB[2974]), .B(DB[2943]), .Z(n3649) );
  AND U7499 ( .A(n136), .B(n3650), .Z(n3648) );
  XOR U7500 ( .A(n3651), .B(n3652), .Z(n3650) );
  XOR U7501 ( .A(DB[2943]), .B(DB[2912]), .Z(n3652) );
  AND U7502 ( .A(n140), .B(n3653), .Z(n3651) );
  XOR U7503 ( .A(n3654), .B(n3655), .Z(n3653) );
  XOR U7504 ( .A(DB[2912]), .B(DB[2881]), .Z(n3655) );
  AND U7505 ( .A(n144), .B(n3656), .Z(n3654) );
  XOR U7506 ( .A(n3657), .B(n3658), .Z(n3656) );
  XOR U7507 ( .A(DB[2881]), .B(DB[2850]), .Z(n3658) );
  AND U7508 ( .A(n148), .B(n3659), .Z(n3657) );
  XOR U7509 ( .A(n3660), .B(n3661), .Z(n3659) );
  XOR U7510 ( .A(DB[2850]), .B(DB[2819]), .Z(n3661) );
  AND U7511 ( .A(n152), .B(n3662), .Z(n3660) );
  XOR U7512 ( .A(n3663), .B(n3664), .Z(n3662) );
  XOR U7513 ( .A(DB[2819]), .B(DB[2788]), .Z(n3664) );
  AND U7514 ( .A(n156), .B(n3665), .Z(n3663) );
  XOR U7515 ( .A(n3666), .B(n3667), .Z(n3665) );
  XOR U7516 ( .A(DB[2788]), .B(DB[2757]), .Z(n3667) );
  AND U7517 ( .A(n160), .B(n3668), .Z(n3666) );
  XOR U7518 ( .A(n3669), .B(n3670), .Z(n3668) );
  XOR U7519 ( .A(DB[2757]), .B(DB[2726]), .Z(n3670) );
  AND U7520 ( .A(n164), .B(n3671), .Z(n3669) );
  XOR U7521 ( .A(n3672), .B(n3673), .Z(n3671) );
  XOR U7522 ( .A(DB[2726]), .B(DB[2695]), .Z(n3673) );
  AND U7523 ( .A(n168), .B(n3674), .Z(n3672) );
  XOR U7524 ( .A(n3675), .B(n3676), .Z(n3674) );
  XOR U7525 ( .A(DB[2695]), .B(DB[2664]), .Z(n3676) );
  AND U7526 ( .A(n172), .B(n3677), .Z(n3675) );
  XOR U7527 ( .A(n3678), .B(n3679), .Z(n3677) );
  XOR U7528 ( .A(DB[2664]), .B(DB[2633]), .Z(n3679) );
  AND U7529 ( .A(n176), .B(n3680), .Z(n3678) );
  XOR U7530 ( .A(n3681), .B(n3682), .Z(n3680) );
  XOR U7531 ( .A(DB[2633]), .B(DB[2602]), .Z(n3682) );
  AND U7532 ( .A(n180), .B(n3683), .Z(n3681) );
  XOR U7533 ( .A(n3684), .B(n3685), .Z(n3683) );
  XOR U7534 ( .A(DB[2602]), .B(DB[2571]), .Z(n3685) );
  AND U7535 ( .A(n184), .B(n3686), .Z(n3684) );
  XOR U7536 ( .A(n3687), .B(n3688), .Z(n3686) );
  XOR U7537 ( .A(DB[2571]), .B(DB[2540]), .Z(n3688) );
  AND U7538 ( .A(n188), .B(n3689), .Z(n3687) );
  XOR U7539 ( .A(n3690), .B(n3691), .Z(n3689) );
  XOR U7540 ( .A(DB[2540]), .B(DB[2509]), .Z(n3691) );
  AND U7541 ( .A(n192), .B(n3692), .Z(n3690) );
  XOR U7542 ( .A(n3693), .B(n3694), .Z(n3692) );
  XOR U7543 ( .A(DB[2509]), .B(DB[2478]), .Z(n3694) );
  AND U7544 ( .A(n196), .B(n3695), .Z(n3693) );
  XOR U7545 ( .A(n3696), .B(n3697), .Z(n3695) );
  XOR U7546 ( .A(DB[2478]), .B(DB[2447]), .Z(n3697) );
  AND U7547 ( .A(n200), .B(n3698), .Z(n3696) );
  XOR U7548 ( .A(n3699), .B(n3700), .Z(n3698) );
  XOR U7549 ( .A(DB[2447]), .B(DB[2416]), .Z(n3700) );
  AND U7550 ( .A(n204), .B(n3701), .Z(n3699) );
  XOR U7551 ( .A(n3702), .B(n3703), .Z(n3701) );
  XOR U7552 ( .A(DB[2416]), .B(DB[2385]), .Z(n3703) );
  AND U7553 ( .A(n208), .B(n3704), .Z(n3702) );
  XOR U7554 ( .A(n3705), .B(n3706), .Z(n3704) );
  XOR U7555 ( .A(DB[2385]), .B(DB[2354]), .Z(n3706) );
  AND U7556 ( .A(n212), .B(n3707), .Z(n3705) );
  XOR U7557 ( .A(n3708), .B(n3709), .Z(n3707) );
  XOR U7558 ( .A(DB[2354]), .B(DB[2323]), .Z(n3709) );
  AND U7559 ( .A(n216), .B(n3710), .Z(n3708) );
  XOR U7560 ( .A(n3711), .B(n3712), .Z(n3710) );
  XOR U7561 ( .A(DB[2323]), .B(DB[2292]), .Z(n3712) );
  AND U7562 ( .A(n220), .B(n3713), .Z(n3711) );
  XOR U7563 ( .A(n3714), .B(n3715), .Z(n3713) );
  XOR U7564 ( .A(DB[2292]), .B(DB[2261]), .Z(n3715) );
  AND U7565 ( .A(n224), .B(n3716), .Z(n3714) );
  XOR U7566 ( .A(n3717), .B(n3718), .Z(n3716) );
  XOR U7567 ( .A(DB[2261]), .B(DB[2230]), .Z(n3718) );
  AND U7568 ( .A(n228), .B(n3719), .Z(n3717) );
  XOR U7569 ( .A(n3720), .B(n3721), .Z(n3719) );
  XOR U7570 ( .A(DB[2230]), .B(DB[2199]), .Z(n3721) );
  AND U7571 ( .A(n232), .B(n3722), .Z(n3720) );
  XOR U7572 ( .A(n3723), .B(n3724), .Z(n3722) );
  XOR U7573 ( .A(DB[2199]), .B(DB[2168]), .Z(n3724) );
  AND U7574 ( .A(n236), .B(n3725), .Z(n3723) );
  XOR U7575 ( .A(n3726), .B(n3727), .Z(n3725) );
  XOR U7576 ( .A(DB[2168]), .B(DB[2137]), .Z(n3727) );
  AND U7577 ( .A(n240), .B(n3728), .Z(n3726) );
  XOR U7578 ( .A(n3729), .B(n3730), .Z(n3728) );
  XOR U7579 ( .A(DB[2137]), .B(DB[2106]), .Z(n3730) );
  AND U7580 ( .A(n244), .B(n3731), .Z(n3729) );
  XOR U7581 ( .A(n3732), .B(n3733), .Z(n3731) );
  XOR U7582 ( .A(DB[2106]), .B(DB[2075]), .Z(n3733) );
  AND U7583 ( .A(n248), .B(n3734), .Z(n3732) );
  XOR U7584 ( .A(n3735), .B(n3736), .Z(n3734) );
  XOR U7585 ( .A(DB[2075]), .B(DB[2044]), .Z(n3736) );
  AND U7586 ( .A(n252), .B(n3737), .Z(n3735) );
  XOR U7587 ( .A(n3738), .B(n3739), .Z(n3737) );
  XOR U7588 ( .A(DB[2044]), .B(DB[2013]), .Z(n3739) );
  AND U7589 ( .A(n256), .B(n3740), .Z(n3738) );
  XOR U7590 ( .A(n3741), .B(n3742), .Z(n3740) );
  XOR U7591 ( .A(DB[2013]), .B(DB[1982]), .Z(n3742) );
  AND U7592 ( .A(n260), .B(n3743), .Z(n3741) );
  XOR U7593 ( .A(n3744), .B(n3745), .Z(n3743) );
  XOR U7594 ( .A(DB[1982]), .B(DB[1951]), .Z(n3745) );
  AND U7595 ( .A(n264), .B(n3746), .Z(n3744) );
  XOR U7596 ( .A(n3747), .B(n3748), .Z(n3746) );
  XOR U7597 ( .A(DB[1951]), .B(DB[1920]), .Z(n3748) );
  AND U7598 ( .A(n268), .B(n3749), .Z(n3747) );
  XOR U7599 ( .A(n3750), .B(n3751), .Z(n3749) );
  XOR U7600 ( .A(DB[1920]), .B(DB[1889]), .Z(n3751) );
  AND U7601 ( .A(n272), .B(n3752), .Z(n3750) );
  XOR U7602 ( .A(n3753), .B(n3754), .Z(n3752) );
  XOR U7603 ( .A(DB[1889]), .B(DB[1858]), .Z(n3754) );
  AND U7604 ( .A(n276), .B(n3755), .Z(n3753) );
  XOR U7605 ( .A(n3756), .B(n3757), .Z(n3755) );
  XOR U7606 ( .A(DB[1858]), .B(DB[1827]), .Z(n3757) );
  AND U7607 ( .A(n280), .B(n3758), .Z(n3756) );
  XOR U7608 ( .A(n3759), .B(n3760), .Z(n3758) );
  XOR U7609 ( .A(DB[1827]), .B(DB[1796]), .Z(n3760) );
  AND U7610 ( .A(n284), .B(n3761), .Z(n3759) );
  XOR U7611 ( .A(n3762), .B(n3763), .Z(n3761) );
  XOR U7612 ( .A(DB[1796]), .B(DB[1765]), .Z(n3763) );
  AND U7613 ( .A(n288), .B(n3764), .Z(n3762) );
  XOR U7614 ( .A(n3765), .B(n3766), .Z(n3764) );
  XOR U7615 ( .A(DB[1765]), .B(DB[1734]), .Z(n3766) );
  AND U7616 ( .A(n292), .B(n3767), .Z(n3765) );
  XOR U7617 ( .A(n3768), .B(n3769), .Z(n3767) );
  XOR U7618 ( .A(DB[1734]), .B(DB[1703]), .Z(n3769) );
  AND U7619 ( .A(n296), .B(n3770), .Z(n3768) );
  XOR U7620 ( .A(n3771), .B(n3772), .Z(n3770) );
  XOR U7621 ( .A(DB[1703]), .B(DB[1672]), .Z(n3772) );
  AND U7622 ( .A(n300), .B(n3773), .Z(n3771) );
  XOR U7623 ( .A(n3774), .B(n3775), .Z(n3773) );
  XOR U7624 ( .A(DB[1672]), .B(DB[1641]), .Z(n3775) );
  AND U7625 ( .A(n304), .B(n3776), .Z(n3774) );
  XOR U7626 ( .A(n3777), .B(n3778), .Z(n3776) );
  XOR U7627 ( .A(DB[1641]), .B(DB[1610]), .Z(n3778) );
  AND U7628 ( .A(n308), .B(n3779), .Z(n3777) );
  XOR U7629 ( .A(n3780), .B(n3781), .Z(n3779) );
  XOR U7630 ( .A(DB[1610]), .B(DB[1579]), .Z(n3781) );
  AND U7631 ( .A(n312), .B(n3782), .Z(n3780) );
  XOR U7632 ( .A(n3783), .B(n3784), .Z(n3782) );
  XOR U7633 ( .A(DB[1579]), .B(DB[1548]), .Z(n3784) );
  AND U7634 ( .A(n316), .B(n3785), .Z(n3783) );
  XOR U7635 ( .A(n3786), .B(n3787), .Z(n3785) );
  XOR U7636 ( .A(DB[1548]), .B(DB[1517]), .Z(n3787) );
  AND U7637 ( .A(n320), .B(n3788), .Z(n3786) );
  XOR U7638 ( .A(n3789), .B(n3790), .Z(n3788) );
  XOR U7639 ( .A(DB[1517]), .B(DB[1486]), .Z(n3790) );
  AND U7640 ( .A(n324), .B(n3791), .Z(n3789) );
  XOR U7641 ( .A(n3792), .B(n3793), .Z(n3791) );
  XOR U7642 ( .A(DB[1486]), .B(DB[1455]), .Z(n3793) );
  AND U7643 ( .A(n328), .B(n3794), .Z(n3792) );
  XOR U7644 ( .A(n3795), .B(n3796), .Z(n3794) );
  XOR U7645 ( .A(DB[1455]), .B(DB[1424]), .Z(n3796) );
  AND U7646 ( .A(n332), .B(n3797), .Z(n3795) );
  XOR U7647 ( .A(n3798), .B(n3799), .Z(n3797) );
  XOR U7648 ( .A(DB[1424]), .B(DB[1393]), .Z(n3799) );
  AND U7649 ( .A(n336), .B(n3800), .Z(n3798) );
  XOR U7650 ( .A(n3801), .B(n3802), .Z(n3800) );
  XOR U7651 ( .A(DB[1393]), .B(DB[1362]), .Z(n3802) );
  AND U7652 ( .A(n340), .B(n3803), .Z(n3801) );
  XOR U7653 ( .A(n3804), .B(n3805), .Z(n3803) );
  XOR U7654 ( .A(DB[1362]), .B(DB[1331]), .Z(n3805) );
  AND U7655 ( .A(n344), .B(n3806), .Z(n3804) );
  XOR U7656 ( .A(n3807), .B(n3808), .Z(n3806) );
  XOR U7657 ( .A(DB[1331]), .B(DB[1300]), .Z(n3808) );
  AND U7658 ( .A(n348), .B(n3809), .Z(n3807) );
  XOR U7659 ( .A(n3810), .B(n3811), .Z(n3809) );
  XOR U7660 ( .A(DB[1300]), .B(DB[1269]), .Z(n3811) );
  AND U7661 ( .A(n352), .B(n3812), .Z(n3810) );
  XOR U7662 ( .A(n3813), .B(n3814), .Z(n3812) );
  XOR U7663 ( .A(DB[1269]), .B(DB[1238]), .Z(n3814) );
  AND U7664 ( .A(n356), .B(n3815), .Z(n3813) );
  XOR U7665 ( .A(n3816), .B(n3817), .Z(n3815) );
  XOR U7666 ( .A(DB[1238]), .B(DB[1207]), .Z(n3817) );
  AND U7667 ( .A(n360), .B(n3818), .Z(n3816) );
  XOR U7668 ( .A(n3819), .B(n3820), .Z(n3818) );
  XOR U7669 ( .A(DB[1207]), .B(DB[1176]), .Z(n3820) );
  AND U7670 ( .A(n364), .B(n3821), .Z(n3819) );
  XOR U7671 ( .A(n3822), .B(n3823), .Z(n3821) );
  XOR U7672 ( .A(DB[1176]), .B(DB[1145]), .Z(n3823) );
  AND U7673 ( .A(n368), .B(n3824), .Z(n3822) );
  XOR U7674 ( .A(n3825), .B(n3826), .Z(n3824) );
  XOR U7675 ( .A(DB[1145]), .B(DB[1114]), .Z(n3826) );
  AND U7676 ( .A(n372), .B(n3827), .Z(n3825) );
  XOR U7677 ( .A(n3828), .B(n3829), .Z(n3827) );
  XOR U7678 ( .A(DB[1114]), .B(DB[1083]), .Z(n3829) );
  AND U7679 ( .A(n376), .B(n3830), .Z(n3828) );
  XOR U7680 ( .A(n3831), .B(n3832), .Z(n3830) );
  XOR U7681 ( .A(DB[1083]), .B(DB[1052]), .Z(n3832) );
  AND U7682 ( .A(n380), .B(n3833), .Z(n3831) );
  XOR U7683 ( .A(n3834), .B(n3835), .Z(n3833) );
  XOR U7684 ( .A(DB[1052]), .B(DB[1021]), .Z(n3835) );
  AND U7685 ( .A(n384), .B(n3836), .Z(n3834) );
  XOR U7686 ( .A(n3837), .B(n3838), .Z(n3836) );
  XOR U7687 ( .A(DB[990]), .B(DB[1021]), .Z(n3838) );
  AND U7688 ( .A(n388), .B(n3839), .Z(n3837) );
  XOR U7689 ( .A(n3840), .B(n3841), .Z(n3839) );
  XOR U7690 ( .A(DB[990]), .B(DB[959]), .Z(n3841) );
  AND U7691 ( .A(n392), .B(n3842), .Z(n3840) );
  XOR U7692 ( .A(n3843), .B(n3844), .Z(n3842) );
  XOR U7693 ( .A(DB[959]), .B(DB[928]), .Z(n3844) );
  AND U7694 ( .A(n396), .B(n3845), .Z(n3843) );
  XOR U7695 ( .A(n3846), .B(n3847), .Z(n3845) );
  XOR U7696 ( .A(DB[928]), .B(DB[897]), .Z(n3847) );
  AND U7697 ( .A(n400), .B(n3848), .Z(n3846) );
  XOR U7698 ( .A(n3849), .B(n3850), .Z(n3848) );
  XOR U7699 ( .A(DB[897]), .B(DB[866]), .Z(n3850) );
  AND U7700 ( .A(n404), .B(n3851), .Z(n3849) );
  XOR U7701 ( .A(n3852), .B(n3853), .Z(n3851) );
  XOR U7702 ( .A(DB[866]), .B(DB[835]), .Z(n3853) );
  AND U7703 ( .A(n408), .B(n3854), .Z(n3852) );
  XOR U7704 ( .A(n3855), .B(n3856), .Z(n3854) );
  XOR U7705 ( .A(DB[835]), .B(DB[804]), .Z(n3856) );
  AND U7706 ( .A(n412), .B(n3857), .Z(n3855) );
  XOR U7707 ( .A(n3858), .B(n3859), .Z(n3857) );
  XOR U7708 ( .A(DB[804]), .B(DB[773]), .Z(n3859) );
  AND U7709 ( .A(n416), .B(n3860), .Z(n3858) );
  XOR U7710 ( .A(n3861), .B(n3862), .Z(n3860) );
  XOR U7711 ( .A(DB[773]), .B(DB[742]), .Z(n3862) );
  AND U7712 ( .A(n420), .B(n3863), .Z(n3861) );
  XOR U7713 ( .A(n3864), .B(n3865), .Z(n3863) );
  XOR U7714 ( .A(DB[742]), .B(DB[711]), .Z(n3865) );
  AND U7715 ( .A(n424), .B(n3866), .Z(n3864) );
  XOR U7716 ( .A(n3867), .B(n3868), .Z(n3866) );
  XOR U7717 ( .A(DB[711]), .B(DB[680]), .Z(n3868) );
  AND U7718 ( .A(n428), .B(n3869), .Z(n3867) );
  XOR U7719 ( .A(n3870), .B(n3871), .Z(n3869) );
  XOR U7720 ( .A(DB[680]), .B(DB[649]), .Z(n3871) );
  AND U7721 ( .A(n432), .B(n3872), .Z(n3870) );
  XOR U7722 ( .A(n3873), .B(n3874), .Z(n3872) );
  XOR U7723 ( .A(DB[649]), .B(DB[618]), .Z(n3874) );
  AND U7724 ( .A(n436), .B(n3875), .Z(n3873) );
  XOR U7725 ( .A(n3876), .B(n3877), .Z(n3875) );
  XOR U7726 ( .A(DB[618]), .B(DB[587]), .Z(n3877) );
  AND U7727 ( .A(n440), .B(n3878), .Z(n3876) );
  XOR U7728 ( .A(n3879), .B(n3880), .Z(n3878) );
  XOR U7729 ( .A(DB[587]), .B(DB[556]), .Z(n3880) );
  AND U7730 ( .A(n444), .B(n3881), .Z(n3879) );
  XOR U7731 ( .A(n3882), .B(n3883), .Z(n3881) );
  XOR U7732 ( .A(DB[556]), .B(DB[525]), .Z(n3883) );
  AND U7733 ( .A(n448), .B(n3884), .Z(n3882) );
  XOR U7734 ( .A(n3885), .B(n3886), .Z(n3884) );
  XOR U7735 ( .A(DB[525]), .B(DB[494]), .Z(n3886) );
  AND U7736 ( .A(n452), .B(n3887), .Z(n3885) );
  XOR U7737 ( .A(n3888), .B(n3889), .Z(n3887) );
  XOR U7738 ( .A(DB[494]), .B(DB[463]), .Z(n3889) );
  AND U7739 ( .A(n456), .B(n3890), .Z(n3888) );
  XOR U7740 ( .A(n3891), .B(n3892), .Z(n3890) );
  XOR U7741 ( .A(DB[463]), .B(DB[432]), .Z(n3892) );
  AND U7742 ( .A(n460), .B(n3893), .Z(n3891) );
  XOR U7743 ( .A(n3894), .B(n3895), .Z(n3893) );
  XOR U7744 ( .A(DB[432]), .B(DB[401]), .Z(n3895) );
  AND U7745 ( .A(n464), .B(n3896), .Z(n3894) );
  XOR U7746 ( .A(n3897), .B(n3898), .Z(n3896) );
  XOR U7747 ( .A(DB[401]), .B(DB[370]), .Z(n3898) );
  AND U7748 ( .A(n468), .B(n3899), .Z(n3897) );
  XOR U7749 ( .A(n3900), .B(n3901), .Z(n3899) );
  XOR U7750 ( .A(DB[370]), .B(DB[339]), .Z(n3901) );
  AND U7751 ( .A(n472), .B(n3902), .Z(n3900) );
  XOR U7752 ( .A(n3903), .B(n3904), .Z(n3902) );
  XOR U7753 ( .A(DB[339]), .B(DB[308]), .Z(n3904) );
  AND U7754 ( .A(n476), .B(n3905), .Z(n3903) );
  XOR U7755 ( .A(n3906), .B(n3907), .Z(n3905) );
  XOR U7756 ( .A(DB[308]), .B(DB[277]), .Z(n3907) );
  AND U7757 ( .A(n480), .B(n3908), .Z(n3906) );
  XOR U7758 ( .A(n3909), .B(n3910), .Z(n3908) );
  XOR U7759 ( .A(DB[277]), .B(DB[246]), .Z(n3910) );
  AND U7760 ( .A(n484), .B(n3911), .Z(n3909) );
  XOR U7761 ( .A(n3912), .B(n3913), .Z(n3911) );
  XOR U7762 ( .A(DB[246]), .B(DB[215]), .Z(n3913) );
  AND U7763 ( .A(n488), .B(n3914), .Z(n3912) );
  XOR U7764 ( .A(n3915), .B(n3916), .Z(n3914) );
  XOR U7765 ( .A(DB[215]), .B(DB[184]), .Z(n3916) );
  AND U7766 ( .A(n492), .B(n3917), .Z(n3915) );
  XOR U7767 ( .A(n3918), .B(n3919), .Z(n3917) );
  XOR U7768 ( .A(DB[184]), .B(DB[153]), .Z(n3919) );
  AND U7769 ( .A(n496), .B(n3920), .Z(n3918) );
  XOR U7770 ( .A(n3921), .B(n3922), .Z(n3920) );
  XOR U7771 ( .A(DB[153]), .B(DB[122]), .Z(n3922) );
  AND U7772 ( .A(n500), .B(n3923), .Z(n3921) );
  XOR U7773 ( .A(n3924), .B(n3925), .Z(n3923) );
  XOR U7774 ( .A(DB[91]), .B(DB[122]), .Z(n3925) );
  AND U7775 ( .A(n504), .B(n3926), .Z(n3924) );
  XOR U7776 ( .A(n3927), .B(n3928), .Z(n3926) );
  XOR U7777 ( .A(DB[91]), .B(DB[60]), .Z(n3928) );
  AND U7778 ( .A(n508), .B(n3929), .Z(n3927) );
  XOR U7779 ( .A(DB[60]), .B(DB[29]), .Z(n3929) );
  XOR U7780 ( .A(DB[3965]), .B(n3930), .Z(min_val_out[28]) );
  AND U7781 ( .A(n2), .B(n3931), .Z(n3930) );
  XOR U7782 ( .A(n3932), .B(n3933), .Z(n3931) );
  XOR U7783 ( .A(n3934), .B(n3935), .Z(n3933) );
  IV U7784 ( .A(DB[3965]), .Z(n3934) );
  AND U7785 ( .A(n8), .B(n3936), .Z(n3932) );
  XOR U7786 ( .A(n3937), .B(n3938), .Z(n3936) );
  XOR U7787 ( .A(DB[3934]), .B(DB[3903]), .Z(n3938) );
  AND U7788 ( .A(n12), .B(n3939), .Z(n3937) );
  XOR U7789 ( .A(n3940), .B(n3941), .Z(n3939) );
  XOR U7790 ( .A(DB[3903]), .B(DB[3872]), .Z(n3941) );
  AND U7791 ( .A(n16), .B(n3942), .Z(n3940) );
  XOR U7792 ( .A(n3943), .B(n3944), .Z(n3942) );
  XOR U7793 ( .A(DB[3872]), .B(DB[3841]), .Z(n3944) );
  AND U7794 ( .A(n20), .B(n3945), .Z(n3943) );
  XOR U7795 ( .A(n3946), .B(n3947), .Z(n3945) );
  XOR U7796 ( .A(DB[3841]), .B(DB[3810]), .Z(n3947) );
  AND U7797 ( .A(n24), .B(n3948), .Z(n3946) );
  XOR U7798 ( .A(n3949), .B(n3950), .Z(n3948) );
  XOR U7799 ( .A(DB[3810]), .B(DB[3779]), .Z(n3950) );
  AND U7800 ( .A(n28), .B(n3951), .Z(n3949) );
  XOR U7801 ( .A(n3952), .B(n3953), .Z(n3951) );
  XOR U7802 ( .A(DB[3779]), .B(DB[3748]), .Z(n3953) );
  AND U7803 ( .A(n32), .B(n3954), .Z(n3952) );
  XOR U7804 ( .A(n3955), .B(n3956), .Z(n3954) );
  XOR U7805 ( .A(DB[3748]), .B(DB[3717]), .Z(n3956) );
  AND U7806 ( .A(n36), .B(n3957), .Z(n3955) );
  XOR U7807 ( .A(n3958), .B(n3959), .Z(n3957) );
  XOR U7808 ( .A(DB[3717]), .B(DB[3686]), .Z(n3959) );
  AND U7809 ( .A(n40), .B(n3960), .Z(n3958) );
  XOR U7810 ( .A(n3961), .B(n3962), .Z(n3960) );
  XOR U7811 ( .A(DB[3686]), .B(DB[3655]), .Z(n3962) );
  AND U7812 ( .A(n44), .B(n3963), .Z(n3961) );
  XOR U7813 ( .A(n3964), .B(n3965), .Z(n3963) );
  XOR U7814 ( .A(DB[3655]), .B(DB[3624]), .Z(n3965) );
  AND U7815 ( .A(n48), .B(n3966), .Z(n3964) );
  XOR U7816 ( .A(n3967), .B(n3968), .Z(n3966) );
  XOR U7817 ( .A(DB[3624]), .B(DB[3593]), .Z(n3968) );
  AND U7818 ( .A(n52), .B(n3969), .Z(n3967) );
  XOR U7819 ( .A(n3970), .B(n3971), .Z(n3969) );
  XOR U7820 ( .A(DB[3593]), .B(DB[3562]), .Z(n3971) );
  AND U7821 ( .A(n56), .B(n3972), .Z(n3970) );
  XOR U7822 ( .A(n3973), .B(n3974), .Z(n3972) );
  XOR U7823 ( .A(DB[3562]), .B(DB[3531]), .Z(n3974) );
  AND U7824 ( .A(n60), .B(n3975), .Z(n3973) );
  XOR U7825 ( .A(n3976), .B(n3977), .Z(n3975) );
  XOR U7826 ( .A(DB[3531]), .B(DB[3500]), .Z(n3977) );
  AND U7827 ( .A(n64), .B(n3978), .Z(n3976) );
  XOR U7828 ( .A(n3979), .B(n3980), .Z(n3978) );
  XOR U7829 ( .A(DB[3500]), .B(DB[3469]), .Z(n3980) );
  AND U7830 ( .A(n68), .B(n3981), .Z(n3979) );
  XOR U7831 ( .A(n3982), .B(n3983), .Z(n3981) );
  XOR U7832 ( .A(DB[3469]), .B(DB[3438]), .Z(n3983) );
  AND U7833 ( .A(n72), .B(n3984), .Z(n3982) );
  XOR U7834 ( .A(n3985), .B(n3986), .Z(n3984) );
  XOR U7835 ( .A(DB[3438]), .B(DB[3407]), .Z(n3986) );
  AND U7836 ( .A(n76), .B(n3987), .Z(n3985) );
  XOR U7837 ( .A(n3988), .B(n3989), .Z(n3987) );
  XOR U7838 ( .A(DB[3407]), .B(DB[3376]), .Z(n3989) );
  AND U7839 ( .A(n80), .B(n3990), .Z(n3988) );
  XOR U7840 ( .A(n3991), .B(n3992), .Z(n3990) );
  XOR U7841 ( .A(DB[3376]), .B(DB[3345]), .Z(n3992) );
  AND U7842 ( .A(n84), .B(n3993), .Z(n3991) );
  XOR U7843 ( .A(n3994), .B(n3995), .Z(n3993) );
  XOR U7844 ( .A(DB[3345]), .B(DB[3314]), .Z(n3995) );
  AND U7845 ( .A(n88), .B(n3996), .Z(n3994) );
  XOR U7846 ( .A(n3997), .B(n3998), .Z(n3996) );
  XOR U7847 ( .A(DB[3314]), .B(DB[3283]), .Z(n3998) );
  AND U7848 ( .A(n92), .B(n3999), .Z(n3997) );
  XOR U7849 ( .A(n4000), .B(n4001), .Z(n3999) );
  XOR U7850 ( .A(DB[3283]), .B(DB[3252]), .Z(n4001) );
  AND U7851 ( .A(n96), .B(n4002), .Z(n4000) );
  XOR U7852 ( .A(n4003), .B(n4004), .Z(n4002) );
  XOR U7853 ( .A(DB[3252]), .B(DB[3221]), .Z(n4004) );
  AND U7854 ( .A(n100), .B(n4005), .Z(n4003) );
  XOR U7855 ( .A(n4006), .B(n4007), .Z(n4005) );
  XOR U7856 ( .A(DB[3221]), .B(DB[3190]), .Z(n4007) );
  AND U7857 ( .A(n104), .B(n4008), .Z(n4006) );
  XOR U7858 ( .A(n4009), .B(n4010), .Z(n4008) );
  XOR U7859 ( .A(DB[3190]), .B(DB[3159]), .Z(n4010) );
  AND U7860 ( .A(n108), .B(n4011), .Z(n4009) );
  XOR U7861 ( .A(n4012), .B(n4013), .Z(n4011) );
  XOR U7862 ( .A(DB[3159]), .B(DB[3128]), .Z(n4013) );
  AND U7863 ( .A(n112), .B(n4014), .Z(n4012) );
  XOR U7864 ( .A(n4015), .B(n4016), .Z(n4014) );
  XOR U7865 ( .A(DB[3128]), .B(DB[3097]), .Z(n4016) );
  AND U7866 ( .A(n116), .B(n4017), .Z(n4015) );
  XOR U7867 ( .A(n4018), .B(n4019), .Z(n4017) );
  XOR U7868 ( .A(DB[3097]), .B(DB[3066]), .Z(n4019) );
  AND U7869 ( .A(n120), .B(n4020), .Z(n4018) );
  XOR U7870 ( .A(n4021), .B(n4022), .Z(n4020) );
  XOR U7871 ( .A(DB[3066]), .B(DB[3035]), .Z(n4022) );
  AND U7872 ( .A(n124), .B(n4023), .Z(n4021) );
  XOR U7873 ( .A(n4024), .B(n4025), .Z(n4023) );
  XOR U7874 ( .A(DB[3035]), .B(DB[3004]), .Z(n4025) );
  AND U7875 ( .A(n128), .B(n4026), .Z(n4024) );
  XOR U7876 ( .A(n4027), .B(n4028), .Z(n4026) );
  XOR U7877 ( .A(DB[3004]), .B(DB[2973]), .Z(n4028) );
  AND U7878 ( .A(n132), .B(n4029), .Z(n4027) );
  XOR U7879 ( .A(n4030), .B(n4031), .Z(n4029) );
  XOR U7880 ( .A(DB[2973]), .B(DB[2942]), .Z(n4031) );
  AND U7881 ( .A(n136), .B(n4032), .Z(n4030) );
  XOR U7882 ( .A(n4033), .B(n4034), .Z(n4032) );
  XOR U7883 ( .A(DB[2942]), .B(DB[2911]), .Z(n4034) );
  AND U7884 ( .A(n140), .B(n4035), .Z(n4033) );
  XOR U7885 ( .A(n4036), .B(n4037), .Z(n4035) );
  XOR U7886 ( .A(DB[2911]), .B(DB[2880]), .Z(n4037) );
  AND U7887 ( .A(n144), .B(n4038), .Z(n4036) );
  XOR U7888 ( .A(n4039), .B(n4040), .Z(n4038) );
  XOR U7889 ( .A(DB[2880]), .B(DB[2849]), .Z(n4040) );
  AND U7890 ( .A(n148), .B(n4041), .Z(n4039) );
  XOR U7891 ( .A(n4042), .B(n4043), .Z(n4041) );
  XOR U7892 ( .A(DB[2849]), .B(DB[2818]), .Z(n4043) );
  AND U7893 ( .A(n152), .B(n4044), .Z(n4042) );
  XOR U7894 ( .A(n4045), .B(n4046), .Z(n4044) );
  XOR U7895 ( .A(DB[2818]), .B(DB[2787]), .Z(n4046) );
  AND U7896 ( .A(n156), .B(n4047), .Z(n4045) );
  XOR U7897 ( .A(n4048), .B(n4049), .Z(n4047) );
  XOR U7898 ( .A(DB[2787]), .B(DB[2756]), .Z(n4049) );
  AND U7899 ( .A(n160), .B(n4050), .Z(n4048) );
  XOR U7900 ( .A(n4051), .B(n4052), .Z(n4050) );
  XOR U7901 ( .A(DB[2756]), .B(DB[2725]), .Z(n4052) );
  AND U7902 ( .A(n164), .B(n4053), .Z(n4051) );
  XOR U7903 ( .A(n4054), .B(n4055), .Z(n4053) );
  XOR U7904 ( .A(DB[2725]), .B(DB[2694]), .Z(n4055) );
  AND U7905 ( .A(n168), .B(n4056), .Z(n4054) );
  XOR U7906 ( .A(n4057), .B(n4058), .Z(n4056) );
  XOR U7907 ( .A(DB[2694]), .B(DB[2663]), .Z(n4058) );
  AND U7908 ( .A(n172), .B(n4059), .Z(n4057) );
  XOR U7909 ( .A(n4060), .B(n4061), .Z(n4059) );
  XOR U7910 ( .A(DB[2663]), .B(DB[2632]), .Z(n4061) );
  AND U7911 ( .A(n176), .B(n4062), .Z(n4060) );
  XOR U7912 ( .A(n4063), .B(n4064), .Z(n4062) );
  XOR U7913 ( .A(DB[2632]), .B(DB[2601]), .Z(n4064) );
  AND U7914 ( .A(n180), .B(n4065), .Z(n4063) );
  XOR U7915 ( .A(n4066), .B(n4067), .Z(n4065) );
  XOR U7916 ( .A(DB[2601]), .B(DB[2570]), .Z(n4067) );
  AND U7917 ( .A(n184), .B(n4068), .Z(n4066) );
  XOR U7918 ( .A(n4069), .B(n4070), .Z(n4068) );
  XOR U7919 ( .A(DB[2570]), .B(DB[2539]), .Z(n4070) );
  AND U7920 ( .A(n188), .B(n4071), .Z(n4069) );
  XOR U7921 ( .A(n4072), .B(n4073), .Z(n4071) );
  XOR U7922 ( .A(DB[2539]), .B(DB[2508]), .Z(n4073) );
  AND U7923 ( .A(n192), .B(n4074), .Z(n4072) );
  XOR U7924 ( .A(n4075), .B(n4076), .Z(n4074) );
  XOR U7925 ( .A(DB[2508]), .B(DB[2477]), .Z(n4076) );
  AND U7926 ( .A(n196), .B(n4077), .Z(n4075) );
  XOR U7927 ( .A(n4078), .B(n4079), .Z(n4077) );
  XOR U7928 ( .A(DB[2477]), .B(DB[2446]), .Z(n4079) );
  AND U7929 ( .A(n200), .B(n4080), .Z(n4078) );
  XOR U7930 ( .A(n4081), .B(n4082), .Z(n4080) );
  XOR U7931 ( .A(DB[2446]), .B(DB[2415]), .Z(n4082) );
  AND U7932 ( .A(n204), .B(n4083), .Z(n4081) );
  XOR U7933 ( .A(n4084), .B(n4085), .Z(n4083) );
  XOR U7934 ( .A(DB[2415]), .B(DB[2384]), .Z(n4085) );
  AND U7935 ( .A(n208), .B(n4086), .Z(n4084) );
  XOR U7936 ( .A(n4087), .B(n4088), .Z(n4086) );
  XOR U7937 ( .A(DB[2384]), .B(DB[2353]), .Z(n4088) );
  AND U7938 ( .A(n212), .B(n4089), .Z(n4087) );
  XOR U7939 ( .A(n4090), .B(n4091), .Z(n4089) );
  XOR U7940 ( .A(DB[2353]), .B(DB[2322]), .Z(n4091) );
  AND U7941 ( .A(n216), .B(n4092), .Z(n4090) );
  XOR U7942 ( .A(n4093), .B(n4094), .Z(n4092) );
  XOR U7943 ( .A(DB[2322]), .B(DB[2291]), .Z(n4094) );
  AND U7944 ( .A(n220), .B(n4095), .Z(n4093) );
  XOR U7945 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U7946 ( .A(DB[2291]), .B(DB[2260]), .Z(n4097) );
  AND U7947 ( .A(n224), .B(n4098), .Z(n4096) );
  XOR U7948 ( .A(n4099), .B(n4100), .Z(n4098) );
  XOR U7949 ( .A(DB[2260]), .B(DB[2229]), .Z(n4100) );
  AND U7950 ( .A(n228), .B(n4101), .Z(n4099) );
  XOR U7951 ( .A(n4102), .B(n4103), .Z(n4101) );
  XOR U7952 ( .A(DB[2229]), .B(DB[2198]), .Z(n4103) );
  AND U7953 ( .A(n232), .B(n4104), .Z(n4102) );
  XOR U7954 ( .A(n4105), .B(n4106), .Z(n4104) );
  XOR U7955 ( .A(DB[2198]), .B(DB[2167]), .Z(n4106) );
  AND U7956 ( .A(n236), .B(n4107), .Z(n4105) );
  XOR U7957 ( .A(n4108), .B(n4109), .Z(n4107) );
  XOR U7958 ( .A(DB[2167]), .B(DB[2136]), .Z(n4109) );
  AND U7959 ( .A(n240), .B(n4110), .Z(n4108) );
  XOR U7960 ( .A(n4111), .B(n4112), .Z(n4110) );
  XOR U7961 ( .A(DB[2136]), .B(DB[2105]), .Z(n4112) );
  AND U7962 ( .A(n244), .B(n4113), .Z(n4111) );
  XOR U7963 ( .A(n4114), .B(n4115), .Z(n4113) );
  XOR U7964 ( .A(DB[2105]), .B(DB[2074]), .Z(n4115) );
  AND U7965 ( .A(n248), .B(n4116), .Z(n4114) );
  XOR U7966 ( .A(n4117), .B(n4118), .Z(n4116) );
  XOR U7967 ( .A(DB[2074]), .B(DB[2043]), .Z(n4118) );
  AND U7968 ( .A(n252), .B(n4119), .Z(n4117) );
  XOR U7969 ( .A(n4120), .B(n4121), .Z(n4119) );
  XOR U7970 ( .A(DB[2043]), .B(DB[2012]), .Z(n4121) );
  AND U7971 ( .A(n256), .B(n4122), .Z(n4120) );
  XOR U7972 ( .A(n4123), .B(n4124), .Z(n4122) );
  XOR U7973 ( .A(DB[2012]), .B(DB[1981]), .Z(n4124) );
  AND U7974 ( .A(n260), .B(n4125), .Z(n4123) );
  XOR U7975 ( .A(n4126), .B(n4127), .Z(n4125) );
  XOR U7976 ( .A(DB[1981]), .B(DB[1950]), .Z(n4127) );
  AND U7977 ( .A(n264), .B(n4128), .Z(n4126) );
  XOR U7978 ( .A(n4129), .B(n4130), .Z(n4128) );
  XOR U7979 ( .A(DB[1950]), .B(DB[1919]), .Z(n4130) );
  AND U7980 ( .A(n268), .B(n4131), .Z(n4129) );
  XOR U7981 ( .A(n4132), .B(n4133), .Z(n4131) );
  XOR U7982 ( .A(DB[1919]), .B(DB[1888]), .Z(n4133) );
  AND U7983 ( .A(n272), .B(n4134), .Z(n4132) );
  XOR U7984 ( .A(n4135), .B(n4136), .Z(n4134) );
  XOR U7985 ( .A(DB[1888]), .B(DB[1857]), .Z(n4136) );
  AND U7986 ( .A(n276), .B(n4137), .Z(n4135) );
  XOR U7987 ( .A(n4138), .B(n4139), .Z(n4137) );
  XOR U7988 ( .A(DB[1857]), .B(DB[1826]), .Z(n4139) );
  AND U7989 ( .A(n280), .B(n4140), .Z(n4138) );
  XOR U7990 ( .A(n4141), .B(n4142), .Z(n4140) );
  XOR U7991 ( .A(DB[1826]), .B(DB[1795]), .Z(n4142) );
  AND U7992 ( .A(n284), .B(n4143), .Z(n4141) );
  XOR U7993 ( .A(n4144), .B(n4145), .Z(n4143) );
  XOR U7994 ( .A(DB[1795]), .B(DB[1764]), .Z(n4145) );
  AND U7995 ( .A(n288), .B(n4146), .Z(n4144) );
  XOR U7996 ( .A(n4147), .B(n4148), .Z(n4146) );
  XOR U7997 ( .A(DB[1764]), .B(DB[1733]), .Z(n4148) );
  AND U7998 ( .A(n292), .B(n4149), .Z(n4147) );
  XOR U7999 ( .A(n4150), .B(n4151), .Z(n4149) );
  XOR U8000 ( .A(DB[1733]), .B(DB[1702]), .Z(n4151) );
  AND U8001 ( .A(n296), .B(n4152), .Z(n4150) );
  XOR U8002 ( .A(n4153), .B(n4154), .Z(n4152) );
  XOR U8003 ( .A(DB[1702]), .B(DB[1671]), .Z(n4154) );
  AND U8004 ( .A(n300), .B(n4155), .Z(n4153) );
  XOR U8005 ( .A(n4156), .B(n4157), .Z(n4155) );
  XOR U8006 ( .A(DB[1671]), .B(DB[1640]), .Z(n4157) );
  AND U8007 ( .A(n304), .B(n4158), .Z(n4156) );
  XOR U8008 ( .A(n4159), .B(n4160), .Z(n4158) );
  XOR U8009 ( .A(DB[1640]), .B(DB[1609]), .Z(n4160) );
  AND U8010 ( .A(n308), .B(n4161), .Z(n4159) );
  XOR U8011 ( .A(n4162), .B(n4163), .Z(n4161) );
  XOR U8012 ( .A(DB[1609]), .B(DB[1578]), .Z(n4163) );
  AND U8013 ( .A(n312), .B(n4164), .Z(n4162) );
  XOR U8014 ( .A(n4165), .B(n4166), .Z(n4164) );
  XOR U8015 ( .A(DB[1578]), .B(DB[1547]), .Z(n4166) );
  AND U8016 ( .A(n316), .B(n4167), .Z(n4165) );
  XOR U8017 ( .A(n4168), .B(n4169), .Z(n4167) );
  XOR U8018 ( .A(DB[1547]), .B(DB[1516]), .Z(n4169) );
  AND U8019 ( .A(n320), .B(n4170), .Z(n4168) );
  XOR U8020 ( .A(n4171), .B(n4172), .Z(n4170) );
  XOR U8021 ( .A(DB[1516]), .B(DB[1485]), .Z(n4172) );
  AND U8022 ( .A(n324), .B(n4173), .Z(n4171) );
  XOR U8023 ( .A(n4174), .B(n4175), .Z(n4173) );
  XOR U8024 ( .A(DB[1485]), .B(DB[1454]), .Z(n4175) );
  AND U8025 ( .A(n328), .B(n4176), .Z(n4174) );
  XOR U8026 ( .A(n4177), .B(n4178), .Z(n4176) );
  XOR U8027 ( .A(DB[1454]), .B(DB[1423]), .Z(n4178) );
  AND U8028 ( .A(n332), .B(n4179), .Z(n4177) );
  XOR U8029 ( .A(n4180), .B(n4181), .Z(n4179) );
  XOR U8030 ( .A(DB[1423]), .B(DB[1392]), .Z(n4181) );
  AND U8031 ( .A(n336), .B(n4182), .Z(n4180) );
  XOR U8032 ( .A(n4183), .B(n4184), .Z(n4182) );
  XOR U8033 ( .A(DB[1392]), .B(DB[1361]), .Z(n4184) );
  AND U8034 ( .A(n340), .B(n4185), .Z(n4183) );
  XOR U8035 ( .A(n4186), .B(n4187), .Z(n4185) );
  XOR U8036 ( .A(DB[1361]), .B(DB[1330]), .Z(n4187) );
  AND U8037 ( .A(n344), .B(n4188), .Z(n4186) );
  XOR U8038 ( .A(n4189), .B(n4190), .Z(n4188) );
  XOR U8039 ( .A(DB[1330]), .B(DB[1299]), .Z(n4190) );
  AND U8040 ( .A(n348), .B(n4191), .Z(n4189) );
  XOR U8041 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR U8042 ( .A(DB[1299]), .B(DB[1268]), .Z(n4193) );
  AND U8043 ( .A(n352), .B(n4194), .Z(n4192) );
  XOR U8044 ( .A(n4195), .B(n4196), .Z(n4194) );
  XOR U8045 ( .A(DB[1268]), .B(DB[1237]), .Z(n4196) );
  AND U8046 ( .A(n356), .B(n4197), .Z(n4195) );
  XOR U8047 ( .A(n4198), .B(n4199), .Z(n4197) );
  XOR U8048 ( .A(DB[1237]), .B(DB[1206]), .Z(n4199) );
  AND U8049 ( .A(n360), .B(n4200), .Z(n4198) );
  XOR U8050 ( .A(n4201), .B(n4202), .Z(n4200) );
  XOR U8051 ( .A(DB[1206]), .B(DB[1175]), .Z(n4202) );
  AND U8052 ( .A(n364), .B(n4203), .Z(n4201) );
  XOR U8053 ( .A(n4204), .B(n4205), .Z(n4203) );
  XOR U8054 ( .A(DB[1175]), .B(DB[1144]), .Z(n4205) );
  AND U8055 ( .A(n368), .B(n4206), .Z(n4204) );
  XOR U8056 ( .A(n4207), .B(n4208), .Z(n4206) );
  XOR U8057 ( .A(DB[1144]), .B(DB[1113]), .Z(n4208) );
  AND U8058 ( .A(n372), .B(n4209), .Z(n4207) );
  XOR U8059 ( .A(n4210), .B(n4211), .Z(n4209) );
  XOR U8060 ( .A(DB[1113]), .B(DB[1082]), .Z(n4211) );
  AND U8061 ( .A(n376), .B(n4212), .Z(n4210) );
  XOR U8062 ( .A(n4213), .B(n4214), .Z(n4212) );
  XOR U8063 ( .A(DB[1082]), .B(DB[1051]), .Z(n4214) );
  AND U8064 ( .A(n380), .B(n4215), .Z(n4213) );
  XOR U8065 ( .A(n4216), .B(n4217), .Z(n4215) );
  XOR U8066 ( .A(DB[1051]), .B(DB[1020]), .Z(n4217) );
  AND U8067 ( .A(n384), .B(n4218), .Z(n4216) );
  XOR U8068 ( .A(n4219), .B(n4220), .Z(n4218) );
  XOR U8069 ( .A(DB[989]), .B(DB[1020]), .Z(n4220) );
  AND U8070 ( .A(n388), .B(n4221), .Z(n4219) );
  XOR U8071 ( .A(n4222), .B(n4223), .Z(n4221) );
  XOR U8072 ( .A(DB[989]), .B(DB[958]), .Z(n4223) );
  AND U8073 ( .A(n392), .B(n4224), .Z(n4222) );
  XOR U8074 ( .A(n4225), .B(n4226), .Z(n4224) );
  XOR U8075 ( .A(DB[958]), .B(DB[927]), .Z(n4226) );
  AND U8076 ( .A(n396), .B(n4227), .Z(n4225) );
  XOR U8077 ( .A(n4228), .B(n4229), .Z(n4227) );
  XOR U8078 ( .A(DB[927]), .B(DB[896]), .Z(n4229) );
  AND U8079 ( .A(n400), .B(n4230), .Z(n4228) );
  XOR U8080 ( .A(n4231), .B(n4232), .Z(n4230) );
  XOR U8081 ( .A(DB[896]), .B(DB[865]), .Z(n4232) );
  AND U8082 ( .A(n404), .B(n4233), .Z(n4231) );
  XOR U8083 ( .A(n4234), .B(n4235), .Z(n4233) );
  XOR U8084 ( .A(DB[865]), .B(DB[834]), .Z(n4235) );
  AND U8085 ( .A(n408), .B(n4236), .Z(n4234) );
  XOR U8086 ( .A(n4237), .B(n4238), .Z(n4236) );
  XOR U8087 ( .A(DB[834]), .B(DB[803]), .Z(n4238) );
  AND U8088 ( .A(n412), .B(n4239), .Z(n4237) );
  XOR U8089 ( .A(n4240), .B(n4241), .Z(n4239) );
  XOR U8090 ( .A(DB[803]), .B(DB[772]), .Z(n4241) );
  AND U8091 ( .A(n416), .B(n4242), .Z(n4240) );
  XOR U8092 ( .A(n4243), .B(n4244), .Z(n4242) );
  XOR U8093 ( .A(DB[772]), .B(DB[741]), .Z(n4244) );
  AND U8094 ( .A(n420), .B(n4245), .Z(n4243) );
  XOR U8095 ( .A(n4246), .B(n4247), .Z(n4245) );
  XOR U8096 ( .A(DB[741]), .B(DB[710]), .Z(n4247) );
  AND U8097 ( .A(n424), .B(n4248), .Z(n4246) );
  XOR U8098 ( .A(n4249), .B(n4250), .Z(n4248) );
  XOR U8099 ( .A(DB[710]), .B(DB[679]), .Z(n4250) );
  AND U8100 ( .A(n428), .B(n4251), .Z(n4249) );
  XOR U8101 ( .A(n4252), .B(n4253), .Z(n4251) );
  XOR U8102 ( .A(DB[679]), .B(DB[648]), .Z(n4253) );
  AND U8103 ( .A(n432), .B(n4254), .Z(n4252) );
  XOR U8104 ( .A(n4255), .B(n4256), .Z(n4254) );
  XOR U8105 ( .A(DB[648]), .B(DB[617]), .Z(n4256) );
  AND U8106 ( .A(n436), .B(n4257), .Z(n4255) );
  XOR U8107 ( .A(n4258), .B(n4259), .Z(n4257) );
  XOR U8108 ( .A(DB[617]), .B(DB[586]), .Z(n4259) );
  AND U8109 ( .A(n440), .B(n4260), .Z(n4258) );
  XOR U8110 ( .A(n4261), .B(n4262), .Z(n4260) );
  XOR U8111 ( .A(DB[586]), .B(DB[555]), .Z(n4262) );
  AND U8112 ( .A(n444), .B(n4263), .Z(n4261) );
  XOR U8113 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U8114 ( .A(DB[555]), .B(DB[524]), .Z(n4265) );
  AND U8115 ( .A(n448), .B(n4266), .Z(n4264) );
  XOR U8116 ( .A(n4267), .B(n4268), .Z(n4266) );
  XOR U8117 ( .A(DB[524]), .B(DB[493]), .Z(n4268) );
  AND U8118 ( .A(n452), .B(n4269), .Z(n4267) );
  XOR U8119 ( .A(n4270), .B(n4271), .Z(n4269) );
  XOR U8120 ( .A(DB[493]), .B(DB[462]), .Z(n4271) );
  AND U8121 ( .A(n456), .B(n4272), .Z(n4270) );
  XOR U8122 ( .A(n4273), .B(n4274), .Z(n4272) );
  XOR U8123 ( .A(DB[462]), .B(DB[431]), .Z(n4274) );
  AND U8124 ( .A(n460), .B(n4275), .Z(n4273) );
  XOR U8125 ( .A(n4276), .B(n4277), .Z(n4275) );
  XOR U8126 ( .A(DB[431]), .B(DB[400]), .Z(n4277) );
  AND U8127 ( .A(n464), .B(n4278), .Z(n4276) );
  XOR U8128 ( .A(n4279), .B(n4280), .Z(n4278) );
  XOR U8129 ( .A(DB[400]), .B(DB[369]), .Z(n4280) );
  AND U8130 ( .A(n468), .B(n4281), .Z(n4279) );
  XOR U8131 ( .A(n4282), .B(n4283), .Z(n4281) );
  XOR U8132 ( .A(DB[369]), .B(DB[338]), .Z(n4283) );
  AND U8133 ( .A(n472), .B(n4284), .Z(n4282) );
  XOR U8134 ( .A(n4285), .B(n4286), .Z(n4284) );
  XOR U8135 ( .A(DB[338]), .B(DB[307]), .Z(n4286) );
  AND U8136 ( .A(n476), .B(n4287), .Z(n4285) );
  XOR U8137 ( .A(n4288), .B(n4289), .Z(n4287) );
  XOR U8138 ( .A(DB[307]), .B(DB[276]), .Z(n4289) );
  AND U8139 ( .A(n480), .B(n4290), .Z(n4288) );
  XOR U8140 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR U8141 ( .A(DB[276]), .B(DB[245]), .Z(n4292) );
  AND U8142 ( .A(n484), .B(n4293), .Z(n4291) );
  XOR U8143 ( .A(n4294), .B(n4295), .Z(n4293) );
  XOR U8144 ( .A(DB[245]), .B(DB[214]), .Z(n4295) );
  AND U8145 ( .A(n488), .B(n4296), .Z(n4294) );
  XOR U8146 ( .A(n4297), .B(n4298), .Z(n4296) );
  XOR U8147 ( .A(DB[214]), .B(DB[183]), .Z(n4298) );
  AND U8148 ( .A(n492), .B(n4299), .Z(n4297) );
  XOR U8149 ( .A(n4300), .B(n4301), .Z(n4299) );
  XOR U8150 ( .A(DB[183]), .B(DB[152]), .Z(n4301) );
  AND U8151 ( .A(n496), .B(n4302), .Z(n4300) );
  XOR U8152 ( .A(n4303), .B(n4304), .Z(n4302) );
  XOR U8153 ( .A(DB[152]), .B(DB[121]), .Z(n4304) );
  AND U8154 ( .A(n500), .B(n4305), .Z(n4303) );
  XOR U8155 ( .A(n4306), .B(n4307), .Z(n4305) );
  XOR U8156 ( .A(DB[90]), .B(DB[121]), .Z(n4307) );
  AND U8157 ( .A(n504), .B(n4308), .Z(n4306) );
  XOR U8158 ( .A(n4309), .B(n4310), .Z(n4308) );
  XOR U8159 ( .A(DB[90]), .B(DB[59]), .Z(n4310) );
  AND U8160 ( .A(n508), .B(n4311), .Z(n4309) );
  XOR U8161 ( .A(DB[59]), .B(DB[28]), .Z(n4311) );
  XOR U8162 ( .A(DB[3964]), .B(n4312), .Z(min_val_out[27]) );
  AND U8163 ( .A(n2), .B(n4313), .Z(n4312) );
  XOR U8164 ( .A(n4314), .B(n4315), .Z(n4313) );
  XOR U8165 ( .A(n4316), .B(n4317), .Z(n4315) );
  IV U8166 ( .A(DB[3964]), .Z(n4316) );
  AND U8167 ( .A(n8), .B(n4318), .Z(n4314) );
  XOR U8168 ( .A(n4319), .B(n4320), .Z(n4318) );
  XOR U8169 ( .A(DB[3933]), .B(DB[3902]), .Z(n4320) );
  AND U8170 ( .A(n12), .B(n4321), .Z(n4319) );
  XOR U8171 ( .A(n4322), .B(n4323), .Z(n4321) );
  XOR U8172 ( .A(DB[3902]), .B(DB[3871]), .Z(n4323) );
  AND U8173 ( .A(n16), .B(n4324), .Z(n4322) );
  XOR U8174 ( .A(n4325), .B(n4326), .Z(n4324) );
  XOR U8175 ( .A(DB[3871]), .B(DB[3840]), .Z(n4326) );
  AND U8176 ( .A(n20), .B(n4327), .Z(n4325) );
  XOR U8177 ( .A(n4328), .B(n4329), .Z(n4327) );
  XOR U8178 ( .A(DB[3840]), .B(DB[3809]), .Z(n4329) );
  AND U8179 ( .A(n24), .B(n4330), .Z(n4328) );
  XOR U8180 ( .A(n4331), .B(n4332), .Z(n4330) );
  XOR U8181 ( .A(DB[3809]), .B(DB[3778]), .Z(n4332) );
  AND U8182 ( .A(n28), .B(n4333), .Z(n4331) );
  XOR U8183 ( .A(n4334), .B(n4335), .Z(n4333) );
  XOR U8184 ( .A(DB[3778]), .B(DB[3747]), .Z(n4335) );
  AND U8185 ( .A(n32), .B(n4336), .Z(n4334) );
  XOR U8186 ( .A(n4337), .B(n4338), .Z(n4336) );
  XOR U8187 ( .A(DB[3747]), .B(DB[3716]), .Z(n4338) );
  AND U8188 ( .A(n36), .B(n4339), .Z(n4337) );
  XOR U8189 ( .A(n4340), .B(n4341), .Z(n4339) );
  XOR U8190 ( .A(DB[3716]), .B(DB[3685]), .Z(n4341) );
  AND U8191 ( .A(n40), .B(n4342), .Z(n4340) );
  XOR U8192 ( .A(n4343), .B(n4344), .Z(n4342) );
  XOR U8193 ( .A(DB[3685]), .B(DB[3654]), .Z(n4344) );
  AND U8194 ( .A(n44), .B(n4345), .Z(n4343) );
  XOR U8195 ( .A(n4346), .B(n4347), .Z(n4345) );
  XOR U8196 ( .A(DB[3654]), .B(DB[3623]), .Z(n4347) );
  AND U8197 ( .A(n48), .B(n4348), .Z(n4346) );
  XOR U8198 ( .A(n4349), .B(n4350), .Z(n4348) );
  XOR U8199 ( .A(DB[3623]), .B(DB[3592]), .Z(n4350) );
  AND U8200 ( .A(n52), .B(n4351), .Z(n4349) );
  XOR U8201 ( .A(n4352), .B(n4353), .Z(n4351) );
  XOR U8202 ( .A(DB[3592]), .B(DB[3561]), .Z(n4353) );
  AND U8203 ( .A(n56), .B(n4354), .Z(n4352) );
  XOR U8204 ( .A(n4355), .B(n4356), .Z(n4354) );
  XOR U8205 ( .A(DB[3561]), .B(DB[3530]), .Z(n4356) );
  AND U8206 ( .A(n60), .B(n4357), .Z(n4355) );
  XOR U8207 ( .A(n4358), .B(n4359), .Z(n4357) );
  XOR U8208 ( .A(DB[3530]), .B(DB[3499]), .Z(n4359) );
  AND U8209 ( .A(n64), .B(n4360), .Z(n4358) );
  XOR U8210 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U8211 ( .A(DB[3499]), .B(DB[3468]), .Z(n4362) );
  AND U8212 ( .A(n68), .B(n4363), .Z(n4361) );
  XOR U8213 ( .A(n4364), .B(n4365), .Z(n4363) );
  XOR U8214 ( .A(DB[3468]), .B(DB[3437]), .Z(n4365) );
  AND U8215 ( .A(n72), .B(n4366), .Z(n4364) );
  XOR U8216 ( .A(n4367), .B(n4368), .Z(n4366) );
  XOR U8217 ( .A(DB[3437]), .B(DB[3406]), .Z(n4368) );
  AND U8218 ( .A(n76), .B(n4369), .Z(n4367) );
  XOR U8219 ( .A(n4370), .B(n4371), .Z(n4369) );
  XOR U8220 ( .A(DB[3406]), .B(DB[3375]), .Z(n4371) );
  AND U8221 ( .A(n80), .B(n4372), .Z(n4370) );
  XOR U8222 ( .A(n4373), .B(n4374), .Z(n4372) );
  XOR U8223 ( .A(DB[3375]), .B(DB[3344]), .Z(n4374) );
  AND U8224 ( .A(n84), .B(n4375), .Z(n4373) );
  XOR U8225 ( .A(n4376), .B(n4377), .Z(n4375) );
  XOR U8226 ( .A(DB[3344]), .B(DB[3313]), .Z(n4377) );
  AND U8227 ( .A(n88), .B(n4378), .Z(n4376) );
  XOR U8228 ( .A(n4379), .B(n4380), .Z(n4378) );
  XOR U8229 ( .A(DB[3313]), .B(DB[3282]), .Z(n4380) );
  AND U8230 ( .A(n92), .B(n4381), .Z(n4379) );
  XOR U8231 ( .A(n4382), .B(n4383), .Z(n4381) );
  XOR U8232 ( .A(DB[3282]), .B(DB[3251]), .Z(n4383) );
  AND U8233 ( .A(n96), .B(n4384), .Z(n4382) );
  XOR U8234 ( .A(n4385), .B(n4386), .Z(n4384) );
  XOR U8235 ( .A(DB[3251]), .B(DB[3220]), .Z(n4386) );
  AND U8236 ( .A(n100), .B(n4387), .Z(n4385) );
  XOR U8237 ( .A(n4388), .B(n4389), .Z(n4387) );
  XOR U8238 ( .A(DB[3220]), .B(DB[3189]), .Z(n4389) );
  AND U8239 ( .A(n104), .B(n4390), .Z(n4388) );
  XOR U8240 ( .A(n4391), .B(n4392), .Z(n4390) );
  XOR U8241 ( .A(DB[3189]), .B(DB[3158]), .Z(n4392) );
  AND U8242 ( .A(n108), .B(n4393), .Z(n4391) );
  XOR U8243 ( .A(n4394), .B(n4395), .Z(n4393) );
  XOR U8244 ( .A(DB[3158]), .B(DB[3127]), .Z(n4395) );
  AND U8245 ( .A(n112), .B(n4396), .Z(n4394) );
  XOR U8246 ( .A(n4397), .B(n4398), .Z(n4396) );
  XOR U8247 ( .A(DB[3127]), .B(DB[3096]), .Z(n4398) );
  AND U8248 ( .A(n116), .B(n4399), .Z(n4397) );
  XOR U8249 ( .A(n4400), .B(n4401), .Z(n4399) );
  XOR U8250 ( .A(DB[3096]), .B(DB[3065]), .Z(n4401) );
  AND U8251 ( .A(n120), .B(n4402), .Z(n4400) );
  XOR U8252 ( .A(n4403), .B(n4404), .Z(n4402) );
  XOR U8253 ( .A(DB[3065]), .B(DB[3034]), .Z(n4404) );
  AND U8254 ( .A(n124), .B(n4405), .Z(n4403) );
  XOR U8255 ( .A(n4406), .B(n4407), .Z(n4405) );
  XOR U8256 ( .A(DB[3034]), .B(DB[3003]), .Z(n4407) );
  AND U8257 ( .A(n128), .B(n4408), .Z(n4406) );
  XOR U8258 ( .A(n4409), .B(n4410), .Z(n4408) );
  XOR U8259 ( .A(DB[3003]), .B(DB[2972]), .Z(n4410) );
  AND U8260 ( .A(n132), .B(n4411), .Z(n4409) );
  XOR U8261 ( .A(n4412), .B(n4413), .Z(n4411) );
  XOR U8262 ( .A(DB[2972]), .B(DB[2941]), .Z(n4413) );
  AND U8263 ( .A(n136), .B(n4414), .Z(n4412) );
  XOR U8264 ( .A(n4415), .B(n4416), .Z(n4414) );
  XOR U8265 ( .A(DB[2941]), .B(DB[2910]), .Z(n4416) );
  AND U8266 ( .A(n140), .B(n4417), .Z(n4415) );
  XOR U8267 ( .A(n4418), .B(n4419), .Z(n4417) );
  XOR U8268 ( .A(DB[2910]), .B(DB[2879]), .Z(n4419) );
  AND U8269 ( .A(n144), .B(n4420), .Z(n4418) );
  XOR U8270 ( .A(n4421), .B(n4422), .Z(n4420) );
  XOR U8271 ( .A(DB[2879]), .B(DB[2848]), .Z(n4422) );
  AND U8272 ( .A(n148), .B(n4423), .Z(n4421) );
  XOR U8273 ( .A(n4424), .B(n4425), .Z(n4423) );
  XOR U8274 ( .A(DB[2848]), .B(DB[2817]), .Z(n4425) );
  AND U8275 ( .A(n152), .B(n4426), .Z(n4424) );
  XOR U8276 ( .A(n4427), .B(n4428), .Z(n4426) );
  XOR U8277 ( .A(DB[2817]), .B(DB[2786]), .Z(n4428) );
  AND U8278 ( .A(n156), .B(n4429), .Z(n4427) );
  XOR U8279 ( .A(n4430), .B(n4431), .Z(n4429) );
  XOR U8280 ( .A(DB[2786]), .B(DB[2755]), .Z(n4431) );
  AND U8281 ( .A(n160), .B(n4432), .Z(n4430) );
  XOR U8282 ( .A(n4433), .B(n4434), .Z(n4432) );
  XOR U8283 ( .A(DB[2755]), .B(DB[2724]), .Z(n4434) );
  AND U8284 ( .A(n164), .B(n4435), .Z(n4433) );
  XOR U8285 ( .A(n4436), .B(n4437), .Z(n4435) );
  XOR U8286 ( .A(DB[2724]), .B(DB[2693]), .Z(n4437) );
  AND U8287 ( .A(n168), .B(n4438), .Z(n4436) );
  XOR U8288 ( .A(n4439), .B(n4440), .Z(n4438) );
  XOR U8289 ( .A(DB[2693]), .B(DB[2662]), .Z(n4440) );
  AND U8290 ( .A(n172), .B(n4441), .Z(n4439) );
  XOR U8291 ( .A(n4442), .B(n4443), .Z(n4441) );
  XOR U8292 ( .A(DB[2662]), .B(DB[2631]), .Z(n4443) );
  AND U8293 ( .A(n176), .B(n4444), .Z(n4442) );
  XOR U8294 ( .A(n4445), .B(n4446), .Z(n4444) );
  XOR U8295 ( .A(DB[2631]), .B(DB[2600]), .Z(n4446) );
  AND U8296 ( .A(n180), .B(n4447), .Z(n4445) );
  XOR U8297 ( .A(n4448), .B(n4449), .Z(n4447) );
  XOR U8298 ( .A(DB[2600]), .B(DB[2569]), .Z(n4449) );
  AND U8299 ( .A(n184), .B(n4450), .Z(n4448) );
  XOR U8300 ( .A(n4451), .B(n4452), .Z(n4450) );
  XOR U8301 ( .A(DB[2569]), .B(DB[2538]), .Z(n4452) );
  AND U8302 ( .A(n188), .B(n4453), .Z(n4451) );
  XOR U8303 ( .A(n4454), .B(n4455), .Z(n4453) );
  XOR U8304 ( .A(DB[2538]), .B(DB[2507]), .Z(n4455) );
  AND U8305 ( .A(n192), .B(n4456), .Z(n4454) );
  XOR U8306 ( .A(n4457), .B(n4458), .Z(n4456) );
  XOR U8307 ( .A(DB[2507]), .B(DB[2476]), .Z(n4458) );
  AND U8308 ( .A(n196), .B(n4459), .Z(n4457) );
  XOR U8309 ( .A(n4460), .B(n4461), .Z(n4459) );
  XOR U8310 ( .A(DB[2476]), .B(DB[2445]), .Z(n4461) );
  AND U8311 ( .A(n200), .B(n4462), .Z(n4460) );
  XOR U8312 ( .A(n4463), .B(n4464), .Z(n4462) );
  XOR U8313 ( .A(DB[2445]), .B(DB[2414]), .Z(n4464) );
  AND U8314 ( .A(n204), .B(n4465), .Z(n4463) );
  XOR U8315 ( .A(n4466), .B(n4467), .Z(n4465) );
  XOR U8316 ( .A(DB[2414]), .B(DB[2383]), .Z(n4467) );
  AND U8317 ( .A(n208), .B(n4468), .Z(n4466) );
  XOR U8318 ( .A(n4469), .B(n4470), .Z(n4468) );
  XOR U8319 ( .A(DB[2383]), .B(DB[2352]), .Z(n4470) );
  AND U8320 ( .A(n212), .B(n4471), .Z(n4469) );
  XOR U8321 ( .A(n4472), .B(n4473), .Z(n4471) );
  XOR U8322 ( .A(DB[2352]), .B(DB[2321]), .Z(n4473) );
  AND U8323 ( .A(n216), .B(n4474), .Z(n4472) );
  XOR U8324 ( .A(n4475), .B(n4476), .Z(n4474) );
  XOR U8325 ( .A(DB[2321]), .B(DB[2290]), .Z(n4476) );
  AND U8326 ( .A(n220), .B(n4477), .Z(n4475) );
  XOR U8327 ( .A(n4478), .B(n4479), .Z(n4477) );
  XOR U8328 ( .A(DB[2290]), .B(DB[2259]), .Z(n4479) );
  AND U8329 ( .A(n224), .B(n4480), .Z(n4478) );
  XOR U8330 ( .A(n4481), .B(n4482), .Z(n4480) );
  XOR U8331 ( .A(DB[2259]), .B(DB[2228]), .Z(n4482) );
  AND U8332 ( .A(n228), .B(n4483), .Z(n4481) );
  XOR U8333 ( .A(n4484), .B(n4485), .Z(n4483) );
  XOR U8334 ( .A(DB[2228]), .B(DB[2197]), .Z(n4485) );
  AND U8335 ( .A(n232), .B(n4486), .Z(n4484) );
  XOR U8336 ( .A(n4487), .B(n4488), .Z(n4486) );
  XOR U8337 ( .A(DB[2197]), .B(DB[2166]), .Z(n4488) );
  AND U8338 ( .A(n236), .B(n4489), .Z(n4487) );
  XOR U8339 ( .A(n4490), .B(n4491), .Z(n4489) );
  XOR U8340 ( .A(DB[2166]), .B(DB[2135]), .Z(n4491) );
  AND U8341 ( .A(n240), .B(n4492), .Z(n4490) );
  XOR U8342 ( .A(n4493), .B(n4494), .Z(n4492) );
  XOR U8343 ( .A(DB[2135]), .B(DB[2104]), .Z(n4494) );
  AND U8344 ( .A(n244), .B(n4495), .Z(n4493) );
  XOR U8345 ( .A(n4496), .B(n4497), .Z(n4495) );
  XOR U8346 ( .A(DB[2104]), .B(DB[2073]), .Z(n4497) );
  AND U8347 ( .A(n248), .B(n4498), .Z(n4496) );
  XOR U8348 ( .A(n4499), .B(n4500), .Z(n4498) );
  XOR U8349 ( .A(DB[2073]), .B(DB[2042]), .Z(n4500) );
  AND U8350 ( .A(n252), .B(n4501), .Z(n4499) );
  XOR U8351 ( .A(n4502), .B(n4503), .Z(n4501) );
  XOR U8352 ( .A(DB[2042]), .B(DB[2011]), .Z(n4503) );
  AND U8353 ( .A(n256), .B(n4504), .Z(n4502) );
  XOR U8354 ( .A(n4505), .B(n4506), .Z(n4504) );
  XOR U8355 ( .A(DB[2011]), .B(DB[1980]), .Z(n4506) );
  AND U8356 ( .A(n260), .B(n4507), .Z(n4505) );
  XOR U8357 ( .A(n4508), .B(n4509), .Z(n4507) );
  XOR U8358 ( .A(DB[1980]), .B(DB[1949]), .Z(n4509) );
  AND U8359 ( .A(n264), .B(n4510), .Z(n4508) );
  XOR U8360 ( .A(n4511), .B(n4512), .Z(n4510) );
  XOR U8361 ( .A(DB[1949]), .B(DB[1918]), .Z(n4512) );
  AND U8362 ( .A(n268), .B(n4513), .Z(n4511) );
  XOR U8363 ( .A(n4514), .B(n4515), .Z(n4513) );
  XOR U8364 ( .A(DB[1918]), .B(DB[1887]), .Z(n4515) );
  AND U8365 ( .A(n272), .B(n4516), .Z(n4514) );
  XOR U8366 ( .A(n4517), .B(n4518), .Z(n4516) );
  XOR U8367 ( .A(DB[1887]), .B(DB[1856]), .Z(n4518) );
  AND U8368 ( .A(n276), .B(n4519), .Z(n4517) );
  XOR U8369 ( .A(n4520), .B(n4521), .Z(n4519) );
  XOR U8370 ( .A(DB[1856]), .B(DB[1825]), .Z(n4521) );
  AND U8371 ( .A(n280), .B(n4522), .Z(n4520) );
  XOR U8372 ( .A(n4523), .B(n4524), .Z(n4522) );
  XOR U8373 ( .A(DB[1825]), .B(DB[1794]), .Z(n4524) );
  AND U8374 ( .A(n284), .B(n4525), .Z(n4523) );
  XOR U8375 ( .A(n4526), .B(n4527), .Z(n4525) );
  XOR U8376 ( .A(DB[1794]), .B(DB[1763]), .Z(n4527) );
  AND U8377 ( .A(n288), .B(n4528), .Z(n4526) );
  XOR U8378 ( .A(n4529), .B(n4530), .Z(n4528) );
  XOR U8379 ( .A(DB[1763]), .B(DB[1732]), .Z(n4530) );
  AND U8380 ( .A(n292), .B(n4531), .Z(n4529) );
  XOR U8381 ( .A(n4532), .B(n4533), .Z(n4531) );
  XOR U8382 ( .A(DB[1732]), .B(DB[1701]), .Z(n4533) );
  AND U8383 ( .A(n296), .B(n4534), .Z(n4532) );
  XOR U8384 ( .A(n4535), .B(n4536), .Z(n4534) );
  XOR U8385 ( .A(DB[1701]), .B(DB[1670]), .Z(n4536) );
  AND U8386 ( .A(n300), .B(n4537), .Z(n4535) );
  XOR U8387 ( .A(n4538), .B(n4539), .Z(n4537) );
  XOR U8388 ( .A(DB[1670]), .B(DB[1639]), .Z(n4539) );
  AND U8389 ( .A(n304), .B(n4540), .Z(n4538) );
  XOR U8390 ( .A(n4541), .B(n4542), .Z(n4540) );
  XOR U8391 ( .A(DB[1639]), .B(DB[1608]), .Z(n4542) );
  AND U8392 ( .A(n308), .B(n4543), .Z(n4541) );
  XOR U8393 ( .A(n4544), .B(n4545), .Z(n4543) );
  XOR U8394 ( .A(DB[1608]), .B(DB[1577]), .Z(n4545) );
  AND U8395 ( .A(n312), .B(n4546), .Z(n4544) );
  XOR U8396 ( .A(n4547), .B(n4548), .Z(n4546) );
  XOR U8397 ( .A(DB[1577]), .B(DB[1546]), .Z(n4548) );
  AND U8398 ( .A(n316), .B(n4549), .Z(n4547) );
  XOR U8399 ( .A(n4550), .B(n4551), .Z(n4549) );
  XOR U8400 ( .A(DB[1546]), .B(DB[1515]), .Z(n4551) );
  AND U8401 ( .A(n320), .B(n4552), .Z(n4550) );
  XOR U8402 ( .A(n4553), .B(n4554), .Z(n4552) );
  XOR U8403 ( .A(DB[1515]), .B(DB[1484]), .Z(n4554) );
  AND U8404 ( .A(n324), .B(n4555), .Z(n4553) );
  XOR U8405 ( .A(n4556), .B(n4557), .Z(n4555) );
  XOR U8406 ( .A(DB[1484]), .B(DB[1453]), .Z(n4557) );
  AND U8407 ( .A(n328), .B(n4558), .Z(n4556) );
  XOR U8408 ( .A(n4559), .B(n4560), .Z(n4558) );
  XOR U8409 ( .A(DB[1453]), .B(DB[1422]), .Z(n4560) );
  AND U8410 ( .A(n332), .B(n4561), .Z(n4559) );
  XOR U8411 ( .A(n4562), .B(n4563), .Z(n4561) );
  XOR U8412 ( .A(DB[1422]), .B(DB[1391]), .Z(n4563) );
  AND U8413 ( .A(n336), .B(n4564), .Z(n4562) );
  XOR U8414 ( .A(n4565), .B(n4566), .Z(n4564) );
  XOR U8415 ( .A(DB[1391]), .B(DB[1360]), .Z(n4566) );
  AND U8416 ( .A(n340), .B(n4567), .Z(n4565) );
  XOR U8417 ( .A(n4568), .B(n4569), .Z(n4567) );
  XOR U8418 ( .A(DB[1360]), .B(DB[1329]), .Z(n4569) );
  AND U8419 ( .A(n344), .B(n4570), .Z(n4568) );
  XOR U8420 ( .A(n4571), .B(n4572), .Z(n4570) );
  XOR U8421 ( .A(DB[1329]), .B(DB[1298]), .Z(n4572) );
  AND U8422 ( .A(n348), .B(n4573), .Z(n4571) );
  XOR U8423 ( .A(n4574), .B(n4575), .Z(n4573) );
  XOR U8424 ( .A(DB[1298]), .B(DB[1267]), .Z(n4575) );
  AND U8425 ( .A(n352), .B(n4576), .Z(n4574) );
  XOR U8426 ( .A(n4577), .B(n4578), .Z(n4576) );
  XOR U8427 ( .A(DB[1267]), .B(DB[1236]), .Z(n4578) );
  AND U8428 ( .A(n356), .B(n4579), .Z(n4577) );
  XOR U8429 ( .A(n4580), .B(n4581), .Z(n4579) );
  XOR U8430 ( .A(DB[1236]), .B(DB[1205]), .Z(n4581) );
  AND U8431 ( .A(n360), .B(n4582), .Z(n4580) );
  XOR U8432 ( .A(n4583), .B(n4584), .Z(n4582) );
  XOR U8433 ( .A(DB[1205]), .B(DB[1174]), .Z(n4584) );
  AND U8434 ( .A(n364), .B(n4585), .Z(n4583) );
  XOR U8435 ( .A(n4586), .B(n4587), .Z(n4585) );
  XOR U8436 ( .A(DB[1174]), .B(DB[1143]), .Z(n4587) );
  AND U8437 ( .A(n368), .B(n4588), .Z(n4586) );
  XOR U8438 ( .A(n4589), .B(n4590), .Z(n4588) );
  XOR U8439 ( .A(DB[1143]), .B(DB[1112]), .Z(n4590) );
  AND U8440 ( .A(n372), .B(n4591), .Z(n4589) );
  XOR U8441 ( .A(n4592), .B(n4593), .Z(n4591) );
  XOR U8442 ( .A(DB[1112]), .B(DB[1081]), .Z(n4593) );
  AND U8443 ( .A(n376), .B(n4594), .Z(n4592) );
  XOR U8444 ( .A(n4595), .B(n4596), .Z(n4594) );
  XOR U8445 ( .A(DB[1081]), .B(DB[1050]), .Z(n4596) );
  AND U8446 ( .A(n380), .B(n4597), .Z(n4595) );
  XOR U8447 ( .A(n4598), .B(n4599), .Z(n4597) );
  XOR U8448 ( .A(DB[1050]), .B(DB[1019]), .Z(n4599) );
  AND U8449 ( .A(n384), .B(n4600), .Z(n4598) );
  XOR U8450 ( .A(n4601), .B(n4602), .Z(n4600) );
  XOR U8451 ( .A(DB[988]), .B(DB[1019]), .Z(n4602) );
  AND U8452 ( .A(n388), .B(n4603), .Z(n4601) );
  XOR U8453 ( .A(n4604), .B(n4605), .Z(n4603) );
  XOR U8454 ( .A(DB[988]), .B(DB[957]), .Z(n4605) );
  AND U8455 ( .A(n392), .B(n4606), .Z(n4604) );
  XOR U8456 ( .A(n4607), .B(n4608), .Z(n4606) );
  XOR U8457 ( .A(DB[957]), .B(DB[926]), .Z(n4608) );
  AND U8458 ( .A(n396), .B(n4609), .Z(n4607) );
  XOR U8459 ( .A(n4610), .B(n4611), .Z(n4609) );
  XOR U8460 ( .A(DB[926]), .B(DB[895]), .Z(n4611) );
  AND U8461 ( .A(n400), .B(n4612), .Z(n4610) );
  XOR U8462 ( .A(n4613), .B(n4614), .Z(n4612) );
  XOR U8463 ( .A(DB[895]), .B(DB[864]), .Z(n4614) );
  AND U8464 ( .A(n404), .B(n4615), .Z(n4613) );
  XOR U8465 ( .A(n4616), .B(n4617), .Z(n4615) );
  XOR U8466 ( .A(DB[864]), .B(DB[833]), .Z(n4617) );
  AND U8467 ( .A(n408), .B(n4618), .Z(n4616) );
  XOR U8468 ( .A(n4619), .B(n4620), .Z(n4618) );
  XOR U8469 ( .A(DB[833]), .B(DB[802]), .Z(n4620) );
  AND U8470 ( .A(n412), .B(n4621), .Z(n4619) );
  XOR U8471 ( .A(n4622), .B(n4623), .Z(n4621) );
  XOR U8472 ( .A(DB[802]), .B(DB[771]), .Z(n4623) );
  AND U8473 ( .A(n416), .B(n4624), .Z(n4622) );
  XOR U8474 ( .A(n4625), .B(n4626), .Z(n4624) );
  XOR U8475 ( .A(DB[771]), .B(DB[740]), .Z(n4626) );
  AND U8476 ( .A(n420), .B(n4627), .Z(n4625) );
  XOR U8477 ( .A(n4628), .B(n4629), .Z(n4627) );
  XOR U8478 ( .A(DB[740]), .B(DB[709]), .Z(n4629) );
  AND U8479 ( .A(n424), .B(n4630), .Z(n4628) );
  XOR U8480 ( .A(n4631), .B(n4632), .Z(n4630) );
  XOR U8481 ( .A(DB[709]), .B(DB[678]), .Z(n4632) );
  AND U8482 ( .A(n428), .B(n4633), .Z(n4631) );
  XOR U8483 ( .A(n4634), .B(n4635), .Z(n4633) );
  XOR U8484 ( .A(DB[678]), .B(DB[647]), .Z(n4635) );
  AND U8485 ( .A(n432), .B(n4636), .Z(n4634) );
  XOR U8486 ( .A(n4637), .B(n4638), .Z(n4636) );
  XOR U8487 ( .A(DB[647]), .B(DB[616]), .Z(n4638) );
  AND U8488 ( .A(n436), .B(n4639), .Z(n4637) );
  XOR U8489 ( .A(n4640), .B(n4641), .Z(n4639) );
  XOR U8490 ( .A(DB[616]), .B(DB[585]), .Z(n4641) );
  AND U8491 ( .A(n440), .B(n4642), .Z(n4640) );
  XOR U8492 ( .A(n4643), .B(n4644), .Z(n4642) );
  XOR U8493 ( .A(DB[585]), .B(DB[554]), .Z(n4644) );
  AND U8494 ( .A(n444), .B(n4645), .Z(n4643) );
  XOR U8495 ( .A(n4646), .B(n4647), .Z(n4645) );
  XOR U8496 ( .A(DB[554]), .B(DB[523]), .Z(n4647) );
  AND U8497 ( .A(n448), .B(n4648), .Z(n4646) );
  XOR U8498 ( .A(n4649), .B(n4650), .Z(n4648) );
  XOR U8499 ( .A(DB[523]), .B(DB[492]), .Z(n4650) );
  AND U8500 ( .A(n452), .B(n4651), .Z(n4649) );
  XOR U8501 ( .A(n4652), .B(n4653), .Z(n4651) );
  XOR U8502 ( .A(DB[492]), .B(DB[461]), .Z(n4653) );
  AND U8503 ( .A(n456), .B(n4654), .Z(n4652) );
  XOR U8504 ( .A(n4655), .B(n4656), .Z(n4654) );
  XOR U8505 ( .A(DB[461]), .B(DB[430]), .Z(n4656) );
  AND U8506 ( .A(n460), .B(n4657), .Z(n4655) );
  XOR U8507 ( .A(n4658), .B(n4659), .Z(n4657) );
  XOR U8508 ( .A(DB[430]), .B(DB[399]), .Z(n4659) );
  AND U8509 ( .A(n464), .B(n4660), .Z(n4658) );
  XOR U8510 ( .A(n4661), .B(n4662), .Z(n4660) );
  XOR U8511 ( .A(DB[399]), .B(DB[368]), .Z(n4662) );
  AND U8512 ( .A(n468), .B(n4663), .Z(n4661) );
  XOR U8513 ( .A(n4664), .B(n4665), .Z(n4663) );
  XOR U8514 ( .A(DB[368]), .B(DB[337]), .Z(n4665) );
  AND U8515 ( .A(n472), .B(n4666), .Z(n4664) );
  XOR U8516 ( .A(n4667), .B(n4668), .Z(n4666) );
  XOR U8517 ( .A(DB[337]), .B(DB[306]), .Z(n4668) );
  AND U8518 ( .A(n476), .B(n4669), .Z(n4667) );
  XOR U8519 ( .A(n4670), .B(n4671), .Z(n4669) );
  XOR U8520 ( .A(DB[306]), .B(DB[275]), .Z(n4671) );
  AND U8521 ( .A(n480), .B(n4672), .Z(n4670) );
  XOR U8522 ( .A(n4673), .B(n4674), .Z(n4672) );
  XOR U8523 ( .A(DB[275]), .B(DB[244]), .Z(n4674) );
  AND U8524 ( .A(n484), .B(n4675), .Z(n4673) );
  XOR U8525 ( .A(n4676), .B(n4677), .Z(n4675) );
  XOR U8526 ( .A(DB[244]), .B(DB[213]), .Z(n4677) );
  AND U8527 ( .A(n488), .B(n4678), .Z(n4676) );
  XOR U8528 ( .A(n4679), .B(n4680), .Z(n4678) );
  XOR U8529 ( .A(DB[213]), .B(DB[182]), .Z(n4680) );
  AND U8530 ( .A(n492), .B(n4681), .Z(n4679) );
  XOR U8531 ( .A(n4682), .B(n4683), .Z(n4681) );
  XOR U8532 ( .A(DB[182]), .B(DB[151]), .Z(n4683) );
  AND U8533 ( .A(n496), .B(n4684), .Z(n4682) );
  XOR U8534 ( .A(n4685), .B(n4686), .Z(n4684) );
  XOR U8535 ( .A(DB[151]), .B(DB[120]), .Z(n4686) );
  AND U8536 ( .A(n500), .B(n4687), .Z(n4685) );
  XOR U8537 ( .A(n4688), .B(n4689), .Z(n4687) );
  XOR U8538 ( .A(DB[89]), .B(DB[120]), .Z(n4689) );
  AND U8539 ( .A(n504), .B(n4690), .Z(n4688) );
  XOR U8540 ( .A(n4691), .B(n4692), .Z(n4690) );
  XOR U8541 ( .A(DB[89]), .B(DB[58]), .Z(n4692) );
  AND U8542 ( .A(n508), .B(n4693), .Z(n4691) );
  XOR U8543 ( .A(DB[58]), .B(DB[27]), .Z(n4693) );
  XOR U8544 ( .A(DB[3963]), .B(n4694), .Z(min_val_out[26]) );
  AND U8545 ( .A(n2), .B(n4695), .Z(n4694) );
  XOR U8546 ( .A(n4696), .B(n4697), .Z(n4695) );
  XOR U8547 ( .A(DB[3963]), .B(DB[3932]), .Z(n4697) );
  AND U8548 ( .A(n8), .B(n4698), .Z(n4696) );
  XOR U8549 ( .A(n4699), .B(n4700), .Z(n4698) );
  XOR U8550 ( .A(DB[3932]), .B(DB[3901]), .Z(n4700) );
  AND U8551 ( .A(n12), .B(n4701), .Z(n4699) );
  XOR U8552 ( .A(n4702), .B(n4703), .Z(n4701) );
  XOR U8553 ( .A(DB[3901]), .B(DB[3870]), .Z(n4703) );
  AND U8554 ( .A(n16), .B(n4704), .Z(n4702) );
  XOR U8555 ( .A(n4705), .B(n4706), .Z(n4704) );
  XOR U8556 ( .A(DB[3870]), .B(DB[3839]), .Z(n4706) );
  AND U8557 ( .A(n20), .B(n4707), .Z(n4705) );
  XOR U8558 ( .A(n4708), .B(n4709), .Z(n4707) );
  XOR U8559 ( .A(DB[3839]), .B(DB[3808]), .Z(n4709) );
  AND U8560 ( .A(n24), .B(n4710), .Z(n4708) );
  XOR U8561 ( .A(n4711), .B(n4712), .Z(n4710) );
  XOR U8562 ( .A(DB[3808]), .B(DB[3777]), .Z(n4712) );
  AND U8563 ( .A(n28), .B(n4713), .Z(n4711) );
  XOR U8564 ( .A(n4714), .B(n4715), .Z(n4713) );
  XOR U8565 ( .A(DB[3777]), .B(DB[3746]), .Z(n4715) );
  AND U8566 ( .A(n32), .B(n4716), .Z(n4714) );
  XOR U8567 ( .A(n4717), .B(n4718), .Z(n4716) );
  XOR U8568 ( .A(DB[3746]), .B(DB[3715]), .Z(n4718) );
  AND U8569 ( .A(n36), .B(n4719), .Z(n4717) );
  XOR U8570 ( .A(n4720), .B(n4721), .Z(n4719) );
  XOR U8571 ( .A(DB[3715]), .B(DB[3684]), .Z(n4721) );
  AND U8572 ( .A(n40), .B(n4722), .Z(n4720) );
  XOR U8573 ( .A(n4723), .B(n4724), .Z(n4722) );
  XOR U8574 ( .A(DB[3684]), .B(DB[3653]), .Z(n4724) );
  AND U8575 ( .A(n44), .B(n4725), .Z(n4723) );
  XOR U8576 ( .A(n4726), .B(n4727), .Z(n4725) );
  XOR U8577 ( .A(DB[3653]), .B(DB[3622]), .Z(n4727) );
  AND U8578 ( .A(n48), .B(n4728), .Z(n4726) );
  XOR U8579 ( .A(n4729), .B(n4730), .Z(n4728) );
  XOR U8580 ( .A(DB[3622]), .B(DB[3591]), .Z(n4730) );
  AND U8581 ( .A(n52), .B(n4731), .Z(n4729) );
  XOR U8582 ( .A(n4732), .B(n4733), .Z(n4731) );
  XOR U8583 ( .A(DB[3591]), .B(DB[3560]), .Z(n4733) );
  AND U8584 ( .A(n56), .B(n4734), .Z(n4732) );
  XOR U8585 ( .A(n4735), .B(n4736), .Z(n4734) );
  XOR U8586 ( .A(DB[3560]), .B(DB[3529]), .Z(n4736) );
  AND U8587 ( .A(n60), .B(n4737), .Z(n4735) );
  XOR U8588 ( .A(n4738), .B(n4739), .Z(n4737) );
  XOR U8589 ( .A(DB[3529]), .B(DB[3498]), .Z(n4739) );
  AND U8590 ( .A(n64), .B(n4740), .Z(n4738) );
  XOR U8591 ( .A(n4741), .B(n4742), .Z(n4740) );
  XOR U8592 ( .A(DB[3498]), .B(DB[3467]), .Z(n4742) );
  AND U8593 ( .A(n68), .B(n4743), .Z(n4741) );
  XOR U8594 ( .A(n4744), .B(n4745), .Z(n4743) );
  XOR U8595 ( .A(DB[3467]), .B(DB[3436]), .Z(n4745) );
  AND U8596 ( .A(n72), .B(n4746), .Z(n4744) );
  XOR U8597 ( .A(n4747), .B(n4748), .Z(n4746) );
  XOR U8598 ( .A(DB[3436]), .B(DB[3405]), .Z(n4748) );
  AND U8599 ( .A(n76), .B(n4749), .Z(n4747) );
  XOR U8600 ( .A(n4750), .B(n4751), .Z(n4749) );
  XOR U8601 ( .A(DB[3405]), .B(DB[3374]), .Z(n4751) );
  AND U8602 ( .A(n80), .B(n4752), .Z(n4750) );
  XOR U8603 ( .A(n4753), .B(n4754), .Z(n4752) );
  XOR U8604 ( .A(DB[3374]), .B(DB[3343]), .Z(n4754) );
  AND U8605 ( .A(n84), .B(n4755), .Z(n4753) );
  XOR U8606 ( .A(n4756), .B(n4757), .Z(n4755) );
  XOR U8607 ( .A(DB[3343]), .B(DB[3312]), .Z(n4757) );
  AND U8608 ( .A(n88), .B(n4758), .Z(n4756) );
  XOR U8609 ( .A(n4759), .B(n4760), .Z(n4758) );
  XOR U8610 ( .A(DB[3312]), .B(DB[3281]), .Z(n4760) );
  AND U8611 ( .A(n92), .B(n4761), .Z(n4759) );
  XOR U8612 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U8613 ( .A(DB[3281]), .B(DB[3250]), .Z(n4763) );
  AND U8614 ( .A(n96), .B(n4764), .Z(n4762) );
  XOR U8615 ( .A(n4765), .B(n4766), .Z(n4764) );
  XOR U8616 ( .A(DB[3250]), .B(DB[3219]), .Z(n4766) );
  AND U8617 ( .A(n100), .B(n4767), .Z(n4765) );
  XOR U8618 ( .A(n4768), .B(n4769), .Z(n4767) );
  XOR U8619 ( .A(DB[3219]), .B(DB[3188]), .Z(n4769) );
  AND U8620 ( .A(n104), .B(n4770), .Z(n4768) );
  XOR U8621 ( .A(n4771), .B(n4772), .Z(n4770) );
  XOR U8622 ( .A(DB[3188]), .B(DB[3157]), .Z(n4772) );
  AND U8623 ( .A(n108), .B(n4773), .Z(n4771) );
  XOR U8624 ( .A(n4774), .B(n4775), .Z(n4773) );
  XOR U8625 ( .A(DB[3157]), .B(DB[3126]), .Z(n4775) );
  AND U8626 ( .A(n112), .B(n4776), .Z(n4774) );
  XOR U8627 ( .A(n4777), .B(n4778), .Z(n4776) );
  XOR U8628 ( .A(DB[3126]), .B(DB[3095]), .Z(n4778) );
  AND U8629 ( .A(n116), .B(n4779), .Z(n4777) );
  XOR U8630 ( .A(n4780), .B(n4781), .Z(n4779) );
  XOR U8631 ( .A(DB[3095]), .B(DB[3064]), .Z(n4781) );
  AND U8632 ( .A(n120), .B(n4782), .Z(n4780) );
  XOR U8633 ( .A(n4783), .B(n4784), .Z(n4782) );
  XOR U8634 ( .A(DB[3064]), .B(DB[3033]), .Z(n4784) );
  AND U8635 ( .A(n124), .B(n4785), .Z(n4783) );
  XOR U8636 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U8637 ( .A(DB[3033]), .B(DB[3002]), .Z(n4787) );
  AND U8638 ( .A(n128), .B(n4788), .Z(n4786) );
  XOR U8639 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U8640 ( .A(DB[3002]), .B(DB[2971]), .Z(n4790) );
  AND U8641 ( .A(n132), .B(n4791), .Z(n4789) );
  XOR U8642 ( .A(n4792), .B(n4793), .Z(n4791) );
  XOR U8643 ( .A(DB[2971]), .B(DB[2940]), .Z(n4793) );
  AND U8644 ( .A(n136), .B(n4794), .Z(n4792) );
  XOR U8645 ( .A(n4795), .B(n4796), .Z(n4794) );
  XOR U8646 ( .A(DB[2940]), .B(DB[2909]), .Z(n4796) );
  AND U8647 ( .A(n140), .B(n4797), .Z(n4795) );
  XOR U8648 ( .A(n4798), .B(n4799), .Z(n4797) );
  XOR U8649 ( .A(DB[2909]), .B(DB[2878]), .Z(n4799) );
  AND U8650 ( .A(n144), .B(n4800), .Z(n4798) );
  XOR U8651 ( .A(n4801), .B(n4802), .Z(n4800) );
  XOR U8652 ( .A(DB[2878]), .B(DB[2847]), .Z(n4802) );
  AND U8653 ( .A(n148), .B(n4803), .Z(n4801) );
  XOR U8654 ( .A(n4804), .B(n4805), .Z(n4803) );
  XOR U8655 ( .A(DB[2847]), .B(DB[2816]), .Z(n4805) );
  AND U8656 ( .A(n152), .B(n4806), .Z(n4804) );
  XOR U8657 ( .A(n4807), .B(n4808), .Z(n4806) );
  XOR U8658 ( .A(DB[2816]), .B(DB[2785]), .Z(n4808) );
  AND U8659 ( .A(n156), .B(n4809), .Z(n4807) );
  XOR U8660 ( .A(n4810), .B(n4811), .Z(n4809) );
  XOR U8661 ( .A(DB[2785]), .B(DB[2754]), .Z(n4811) );
  AND U8662 ( .A(n160), .B(n4812), .Z(n4810) );
  XOR U8663 ( .A(n4813), .B(n4814), .Z(n4812) );
  XOR U8664 ( .A(DB[2754]), .B(DB[2723]), .Z(n4814) );
  AND U8665 ( .A(n164), .B(n4815), .Z(n4813) );
  XOR U8666 ( .A(n4816), .B(n4817), .Z(n4815) );
  XOR U8667 ( .A(DB[2723]), .B(DB[2692]), .Z(n4817) );
  AND U8668 ( .A(n168), .B(n4818), .Z(n4816) );
  XOR U8669 ( .A(n4819), .B(n4820), .Z(n4818) );
  XOR U8670 ( .A(DB[2692]), .B(DB[2661]), .Z(n4820) );
  AND U8671 ( .A(n172), .B(n4821), .Z(n4819) );
  XOR U8672 ( .A(n4822), .B(n4823), .Z(n4821) );
  XOR U8673 ( .A(DB[2661]), .B(DB[2630]), .Z(n4823) );
  AND U8674 ( .A(n176), .B(n4824), .Z(n4822) );
  XOR U8675 ( .A(n4825), .B(n4826), .Z(n4824) );
  XOR U8676 ( .A(DB[2630]), .B(DB[2599]), .Z(n4826) );
  AND U8677 ( .A(n180), .B(n4827), .Z(n4825) );
  XOR U8678 ( .A(n4828), .B(n4829), .Z(n4827) );
  XOR U8679 ( .A(DB[2599]), .B(DB[2568]), .Z(n4829) );
  AND U8680 ( .A(n184), .B(n4830), .Z(n4828) );
  XOR U8681 ( .A(n4831), .B(n4832), .Z(n4830) );
  XOR U8682 ( .A(DB[2568]), .B(DB[2537]), .Z(n4832) );
  AND U8683 ( .A(n188), .B(n4833), .Z(n4831) );
  XOR U8684 ( .A(n4834), .B(n4835), .Z(n4833) );
  XOR U8685 ( .A(DB[2537]), .B(DB[2506]), .Z(n4835) );
  AND U8686 ( .A(n192), .B(n4836), .Z(n4834) );
  XOR U8687 ( .A(n4837), .B(n4838), .Z(n4836) );
  XOR U8688 ( .A(DB[2506]), .B(DB[2475]), .Z(n4838) );
  AND U8689 ( .A(n196), .B(n4839), .Z(n4837) );
  XOR U8690 ( .A(n4840), .B(n4841), .Z(n4839) );
  XOR U8691 ( .A(DB[2475]), .B(DB[2444]), .Z(n4841) );
  AND U8692 ( .A(n200), .B(n4842), .Z(n4840) );
  XOR U8693 ( .A(n4843), .B(n4844), .Z(n4842) );
  XOR U8694 ( .A(DB[2444]), .B(DB[2413]), .Z(n4844) );
  AND U8695 ( .A(n204), .B(n4845), .Z(n4843) );
  XOR U8696 ( .A(n4846), .B(n4847), .Z(n4845) );
  XOR U8697 ( .A(DB[2413]), .B(DB[2382]), .Z(n4847) );
  AND U8698 ( .A(n208), .B(n4848), .Z(n4846) );
  XOR U8699 ( .A(n4849), .B(n4850), .Z(n4848) );
  XOR U8700 ( .A(DB[2382]), .B(DB[2351]), .Z(n4850) );
  AND U8701 ( .A(n212), .B(n4851), .Z(n4849) );
  XOR U8702 ( .A(n4852), .B(n4853), .Z(n4851) );
  XOR U8703 ( .A(DB[2351]), .B(DB[2320]), .Z(n4853) );
  AND U8704 ( .A(n216), .B(n4854), .Z(n4852) );
  XOR U8705 ( .A(n4855), .B(n4856), .Z(n4854) );
  XOR U8706 ( .A(DB[2320]), .B(DB[2289]), .Z(n4856) );
  AND U8707 ( .A(n220), .B(n4857), .Z(n4855) );
  XOR U8708 ( .A(n4858), .B(n4859), .Z(n4857) );
  XOR U8709 ( .A(DB[2289]), .B(DB[2258]), .Z(n4859) );
  AND U8710 ( .A(n224), .B(n4860), .Z(n4858) );
  XOR U8711 ( .A(n4861), .B(n4862), .Z(n4860) );
  XOR U8712 ( .A(DB[2258]), .B(DB[2227]), .Z(n4862) );
  AND U8713 ( .A(n228), .B(n4863), .Z(n4861) );
  XOR U8714 ( .A(n4864), .B(n4865), .Z(n4863) );
  XOR U8715 ( .A(DB[2227]), .B(DB[2196]), .Z(n4865) );
  AND U8716 ( .A(n232), .B(n4866), .Z(n4864) );
  XOR U8717 ( .A(n4867), .B(n4868), .Z(n4866) );
  XOR U8718 ( .A(DB[2196]), .B(DB[2165]), .Z(n4868) );
  AND U8719 ( .A(n236), .B(n4869), .Z(n4867) );
  XOR U8720 ( .A(n4870), .B(n4871), .Z(n4869) );
  XOR U8721 ( .A(DB[2165]), .B(DB[2134]), .Z(n4871) );
  AND U8722 ( .A(n240), .B(n4872), .Z(n4870) );
  XOR U8723 ( .A(n4873), .B(n4874), .Z(n4872) );
  XOR U8724 ( .A(DB[2134]), .B(DB[2103]), .Z(n4874) );
  AND U8725 ( .A(n244), .B(n4875), .Z(n4873) );
  XOR U8726 ( .A(n4876), .B(n4877), .Z(n4875) );
  XOR U8727 ( .A(DB[2103]), .B(DB[2072]), .Z(n4877) );
  AND U8728 ( .A(n248), .B(n4878), .Z(n4876) );
  XOR U8729 ( .A(n4879), .B(n4880), .Z(n4878) );
  XOR U8730 ( .A(DB[2072]), .B(DB[2041]), .Z(n4880) );
  AND U8731 ( .A(n252), .B(n4881), .Z(n4879) );
  XOR U8732 ( .A(n4882), .B(n4883), .Z(n4881) );
  XOR U8733 ( .A(DB[2041]), .B(DB[2010]), .Z(n4883) );
  AND U8734 ( .A(n256), .B(n4884), .Z(n4882) );
  XOR U8735 ( .A(n4885), .B(n4886), .Z(n4884) );
  XOR U8736 ( .A(DB[2010]), .B(DB[1979]), .Z(n4886) );
  AND U8737 ( .A(n260), .B(n4887), .Z(n4885) );
  XOR U8738 ( .A(n4888), .B(n4889), .Z(n4887) );
  XOR U8739 ( .A(DB[1979]), .B(DB[1948]), .Z(n4889) );
  AND U8740 ( .A(n264), .B(n4890), .Z(n4888) );
  XOR U8741 ( .A(n4891), .B(n4892), .Z(n4890) );
  XOR U8742 ( .A(DB[1948]), .B(DB[1917]), .Z(n4892) );
  AND U8743 ( .A(n268), .B(n4893), .Z(n4891) );
  XOR U8744 ( .A(n4894), .B(n4895), .Z(n4893) );
  XOR U8745 ( .A(DB[1917]), .B(DB[1886]), .Z(n4895) );
  AND U8746 ( .A(n272), .B(n4896), .Z(n4894) );
  XOR U8747 ( .A(n4897), .B(n4898), .Z(n4896) );
  XOR U8748 ( .A(DB[1886]), .B(DB[1855]), .Z(n4898) );
  AND U8749 ( .A(n276), .B(n4899), .Z(n4897) );
  XOR U8750 ( .A(n4900), .B(n4901), .Z(n4899) );
  XOR U8751 ( .A(DB[1855]), .B(DB[1824]), .Z(n4901) );
  AND U8752 ( .A(n280), .B(n4902), .Z(n4900) );
  XOR U8753 ( .A(n4903), .B(n4904), .Z(n4902) );
  XOR U8754 ( .A(DB[1824]), .B(DB[1793]), .Z(n4904) );
  AND U8755 ( .A(n284), .B(n4905), .Z(n4903) );
  XOR U8756 ( .A(n4906), .B(n4907), .Z(n4905) );
  XOR U8757 ( .A(DB[1793]), .B(DB[1762]), .Z(n4907) );
  AND U8758 ( .A(n288), .B(n4908), .Z(n4906) );
  XOR U8759 ( .A(n4909), .B(n4910), .Z(n4908) );
  XOR U8760 ( .A(DB[1762]), .B(DB[1731]), .Z(n4910) );
  AND U8761 ( .A(n292), .B(n4911), .Z(n4909) );
  XOR U8762 ( .A(n4912), .B(n4913), .Z(n4911) );
  XOR U8763 ( .A(DB[1731]), .B(DB[1700]), .Z(n4913) );
  AND U8764 ( .A(n296), .B(n4914), .Z(n4912) );
  XOR U8765 ( .A(n4915), .B(n4916), .Z(n4914) );
  XOR U8766 ( .A(DB[1700]), .B(DB[1669]), .Z(n4916) );
  AND U8767 ( .A(n300), .B(n4917), .Z(n4915) );
  XOR U8768 ( .A(n4918), .B(n4919), .Z(n4917) );
  XOR U8769 ( .A(DB[1669]), .B(DB[1638]), .Z(n4919) );
  AND U8770 ( .A(n304), .B(n4920), .Z(n4918) );
  XOR U8771 ( .A(n4921), .B(n4922), .Z(n4920) );
  XOR U8772 ( .A(DB[1638]), .B(DB[1607]), .Z(n4922) );
  AND U8773 ( .A(n308), .B(n4923), .Z(n4921) );
  XOR U8774 ( .A(n4924), .B(n4925), .Z(n4923) );
  XOR U8775 ( .A(DB[1607]), .B(DB[1576]), .Z(n4925) );
  AND U8776 ( .A(n312), .B(n4926), .Z(n4924) );
  XOR U8777 ( .A(n4927), .B(n4928), .Z(n4926) );
  XOR U8778 ( .A(DB[1576]), .B(DB[1545]), .Z(n4928) );
  AND U8779 ( .A(n316), .B(n4929), .Z(n4927) );
  XOR U8780 ( .A(n4930), .B(n4931), .Z(n4929) );
  XOR U8781 ( .A(DB[1545]), .B(DB[1514]), .Z(n4931) );
  AND U8782 ( .A(n320), .B(n4932), .Z(n4930) );
  XOR U8783 ( .A(n4933), .B(n4934), .Z(n4932) );
  XOR U8784 ( .A(DB[1514]), .B(DB[1483]), .Z(n4934) );
  AND U8785 ( .A(n324), .B(n4935), .Z(n4933) );
  XOR U8786 ( .A(n4936), .B(n4937), .Z(n4935) );
  XOR U8787 ( .A(DB[1483]), .B(DB[1452]), .Z(n4937) );
  AND U8788 ( .A(n328), .B(n4938), .Z(n4936) );
  XOR U8789 ( .A(n4939), .B(n4940), .Z(n4938) );
  XOR U8790 ( .A(DB[1452]), .B(DB[1421]), .Z(n4940) );
  AND U8791 ( .A(n332), .B(n4941), .Z(n4939) );
  XOR U8792 ( .A(n4942), .B(n4943), .Z(n4941) );
  XOR U8793 ( .A(DB[1421]), .B(DB[1390]), .Z(n4943) );
  AND U8794 ( .A(n336), .B(n4944), .Z(n4942) );
  XOR U8795 ( .A(n4945), .B(n4946), .Z(n4944) );
  XOR U8796 ( .A(DB[1390]), .B(DB[1359]), .Z(n4946) );
  AND U8797 ( .A(n340), .B(n4947), .Z(n4945) );
  XOR U8798 ( .A(n4948), .B(n4949), .Z(n4947) );
  XOR U8799 ( .A(DB[1359]), .B(DB[1328]), .Z(n4949) );
  AND U8800 ( .A(n344), .B(n4950), .Z(n4948) );
  XOR U8801 ( .A(n4951), .B(n4952), .Z(n4950) );
  XOR U8802 ( .A(DB[1328]), .B(DB[1297]), .Z(n4952) );
  AND U8803 ( .A(n348), .B(n4953), .Z(n4951) );
  XOR U8804 ( .A(n4954), .B(n4955), .Z(n4953) );
  XOR U8805 ( .A(DB[1297]), .B(DB[1266]), .Z(n4955) );
  AND U8806 ( .A(n352), .B(n4956), .Z(n4954) );
  XOR U8807 ( .A(n4957), .B(n4958), .Z(n4956) );
  XOR U8808 ( .A(DB[1266]), .B(DB[1235]), .Z(n4958) );
  AND U8809 ( .A(n356), .B(n4959), .Z(n4957) );
  XOR U8810 ( .A(n4960), .B(n4961), .Z(n4959) );
  XOR U8811 ( .A(DB[1235]), .B(DB[1204]), .Z(n4961) );
  AND U8812 ( .A(n360), .B(n4962), .Z(n4960) );
  XOR U8813 ( .A(n4963), .B(n4964), .Z(n4962) );
  XOR U8814 ( .A(DB[1204]), .B(DB[1173]), .Z(n4964) );
  AND U8815 ( .A(n364), .B(n4965), .Z(n4963) );
  XOR U8816 ( .A(n4966), .B(n4967), .Z(n4965) );
  XOR U8817 ( .A(DB[1173]), .B(DB[1142]), .Z(n4967) );
  AND U8818 ( .A(n368), .B(n4968), .Z(n4966) );
  XOR U8819 ( .A(n4969), .B(n4970), .Z(n4968) );
  XOR U8820 ( .A(DB[1142]), .B(DB[1111]), .Z(n4970) );
  AND U8821 ( .A(n372), .B(n4971), .Z(n4969) );
  XOR U8822 ( .A(n4972), .B(n4973), .Z(n4971) );
  XOR U8823 ( .A(DB[1111]), .B(DB[1080]), .Z(n4973) );
  AND U8824 ( .A(n376), .B(n4974), .Z(n4972) );
  XOR U8825 ( .A(n4975), .B(n4976), .Z(n4974) );
  XOR U8826 ( .A(DB[1080]), .B(DB[1049]), .Z(n4976) );
  AND U8827 ( .A(n380), .B(n4977), .Z(n4975) );
  XOR U8828 ( .A(n4978), .B(n4979), .Z(n4977) );
  XOR U8829 ( .A(DB[1049]), .B(DB[1018]), .Z(n4979) );
  AND U8830 ( .A(n384), .B(n4980), .Z(n4978) );
  XOR U8831 ( .A(n4981), .B(n4982), .Z(n4980) );
  XOR U8832 ( .A(DB[987]), .B(DB[1018]), .Z(n4982) );
  AND U8833 ( .A(n388), .B(n4983), .Z(n4981) );
  XOR U8834 ( .A(n4984), .B(n4985), .Z(n4983) );
  XOR U8835 ( .A(DB[987]), .B(DB[956]), .Z(n4985) );
  AND U8836 ( .A(n392), .B(n4986), .Z(n4984) );
  XOR U8837 ( .A(n4987), .B(n4988), .Z(n4986) );
  XOR U8838 ( .A(DB[956]), .B(DB[925]), .Z(n4988) );
  AND U8839 ( .A(n396), .B(n4989), .Z(n4987) );
  XOR U8840 ( .A(n4990), .B(n4991), .Z(n4989) );
  XOR U8841 ( .A(DB[925]), .B(DB[894]), .Z(n4991) );
  AND U8842 ( .A(n400), .B(n4992), .Z(n4990) );
  XOR U8843 ( .A(n4993), .B(n4994), .Z(n4992) );
  XOR U8844 ( .A(DB[894]), .B(DB[863]), .Z(n4994) );
  AND U8845 ( .A(n404), .B(n4995), .Z(n4993) );
  XOR U8846 ( .A(n4996), .B(n4997), .Z(n4995) );
  XOR U8847 ( .A(DB[863]), .B(DB[832]), .Z(n4997) );
  AND U8848 ( .A(n408), .B(n4998), .Z(n4996) );
  XOR U8849 ( .A(n4999), .B(n5000), .Z(n4998) );
  XOR U8850 ( .A(DB[832]), .B(DB[801]), .Z(n5000) );
  AND U8851 ( .A(n412), .B(n5001), .Z(n4999) );
  XOR U8852 ( .A(n5002), .B(n5003), .Z(n5001) );
  XOR U8853 ( .A(DB[801]), .B(DB[770]), .Z(n5003) );
  AND U8854 ( .A(n416), .B(n5004), .Z(n5002) );
  XOR U8855 ( .A(n5005), .B(n5006), .Z(n5004) );
  XOR U8856 ( .A(DB[770]), .B(DB[739]), .Z(n5006) );
  AND U8857 ( .A(n420), .B(n5007), .Z(n5005) );
  XOR U8858 ( .A(n5008), .B(n5009), .Z(n5007) );
  XOR U8859 ( .A(DB[739]), .B(DB[708]), .Z(n5009) );
  AND U8860 ( .A(n424), .B(n5010), .Z(n5008) );
  XOR U8861 ( .A(n5011), .B(n5012), .Z(n5010) );
  XOR U8862 ( .A(DB[708]), .B(DB[677]), .Z(n5012) );
  AND U8863 ( .A(n428), .B(n5013), .Z(n5011) );
  XOR U8864 ( .A(n5014), .B(n5015), .Z(n5013) );
  XOR U8865 ( .A(DB[677]), .B(DB[646]), .Z(n5015) );
  AND U8866 ( .A(n432), .B(n5016), .Z(n5014) );
  XOR U8867 ( .A(n5017), .B(n5018), .Z(n5016) );
  XOR U8868 ( .A(DB[646]), .B(DB[615]), .Z(n5018) );
  AND U8869 ( .A(n436), .B(n5019), .Z(n5017) );
  XOR U8870 ( .A(n5020), .B(n5021), .Z(n5019) );
  XOR U8871 ( .A(DB[615]), .B(DB[584]), .Z(n5021) );
  AND U8872 ( .A(n440), .B(n5022), .Z(n5020) );
  XOR U8873 ( .A(n5023), .B(n5024), .Z(n5022) );
  XOR U8874 ( .A(DB[584]), .B(DB[553]), .Z(n5024) );
  AND U8875 ( .A(n444), .B(n5025), .Z(n5023) );
  XOR U8876 ( .A(n5026), .B(n5027), .Z(n5025) );
  XOR U8877 ( .A(DB[553]), .B(DB[522]), .Z(n5027) );
  AND U8878 ( .A(n448), .B(n5028), .Z(n5026) );
  XOR U8879 ( .A(n5029), .B(n5030), .Z(n5028) );
  XOR U8880 ( .A(DB[522]), .B(DB[491]), .Z(n5030) );
  AND U8881 ( .A(n452), .B(n5031), .Z(n5029) );
  XOR U8882 ( .A(n5032), .B(n5033), .Z(n5031) );
  XOR U8883 ( .A(DB[491]), .B(DB[460]), .Z(n5033) );
  AND U8884 ( .A(n456), .B(n5034), .Z(n5032) );
  XOR U8885 ( .A(n5035), .B(n5036), .Z(n5034) );
  XOR U8886 ( .A(DB[460]), .B(DB[429]), .Z(n5036) );
  AND U8887 ( .A(n460), .B(n5037), .Z(n5035) );
  XOR U8888 ( .A(n5038), .B(n5039), .Z(n5037) );
  XOR U8889 ( .A(DB[429]), .B(DB[398]), .Z(n5039) );
  AND U8890 ( .A(n464), .B(n5040), .Z(n5038) );
  XOR U8891 ( .A(n5041), .B(n5042), .Z(n5040) );
  XOR U8892 ( .A(DB[398]), .B(DB[367]), .Z(n5042) );
  AND U8893 ( .A(n468), .B(n5043), .Z(n5041) );
  XOR U8894 ( .A(n5044), .B(n5045), .Z(n5043) );
  XOR U8895 ( .A(DB[367]), .B(DB[336]), .Z(n5045) );
  AND U8896 ( .A(n472), .B(n5046), .Z(n5044) );
  XOR U8897 ( .A(n5047), .B(n5048), .Z(n5046) );
  XOR U8898 ( .A(DB[336]), .B(DB[305]), .Z(n5048) );
  AND U8899 ( .A(n476), .B(n5049), .Z(n5047) );
  XOR U8900 ( .A(n5050), .B(n5051), .Z(n5049) );
  XOR U8901 ( .A(DB[305]), .B(DB[274]), .Z(n5051) );
  AND U8902 ( .A(n480), .B(n5052), .Z(n5050) );
  XOR U8903 ( .A(n5053), .B(n5054), .Z(n5052) );
  XOR U8904 ( .A(DB[274]), .B(DB[243]), .Z(n5054) );
  AND U8905 ( .A(n484), .B(n5055), .Z(n5053) );
  XOR U8906 ( .A(n5056), .B(n5057), .Z(n5055) );
  XOR U8907 ( .A(DB[243]), .B(DB[212]), .Z(n5057) );
  AND U8908 ( .A(n488), .B(n5058), .Z(n5056) );
  XOR U8909 ( .A(n5059), .B(n5060), .Z(n5058) );
  XOR U8910 ( .A(DB[212]), .B(DB[181]), .Z(n5060) );
  AND U8911 ( .A(n492), .B(n5061), .Z(n5059) );
  XOR U8912 ( .A(n5062), .B(n5063), .Z(n5061) );
  XOR U8913 ( .A(DB[181]), .B(DB[150]), .Z(n5063) );
  AND U8914 ( .A(n496), .B(n5064), .Z(n5062) );
  XOR U8915 ( .A(n5065), .B(n5066), .Z(n5064) );
  XOR U8916 ( .A(DB[150]), .B(DB[119]), .Z(n5066) );
  AND U8917 ( .A(n500), .B(n5067), .Z(n5065) );
  XOR U8918 ( .A(n5068), .B(n5069), .Z(n5067) );
  XOR U8919 ( .A(DB[88]), .B(DB[119]), .Z(n5069) );
  AND U8920 ( .A(n504), .B(n5070), .Z(n5068) );
  XOR U8921 ( .A(n5071), .B(n5072), .Z(n5070) );
  XOR U8922 ( .A(DB[88]), .B(DB[57]), .Z(n5072) );
  AND U8923 ( .A(n508), .B(n5073), .Z(n5071) );
  XOR U8924 ( .A(DB[57]), .B(DB[26]), .Z(n5073) );
  XOR U8925 ( .A(DB[3962]), .B(n5074), .Z(min_val_out[25]) );
  AND U8926 ( .A(n2), .B(n5075), .Z(n5074) );
  XOR U8927 ( .A(n5076), .B(n5077), .Z(n5075) );
  XOR U8928 ( .A(n5078), .B(n5079), .Z(n5077) );
  IV U8929 ( .A(DB[3962]), .Z(n5078) );
  AND U8930 ( .A(n8), .B(n5080), .Z(n5076) );
  XOR U8931 ( .A(n5081), .B(n5082), .Z(n5080) );
  XOR U8932 ( .A(DB[3931]), .B(DB[3900]), .Z(n5082) );
  AND U8933 ( .A(n12), .B(n5083), .Z(n5081) );
  XOR U8934 ( .A(n5084), .B(n5085), .Z(n5083) );
  XOR U8935 ( .A(DB[3900]), .B(DB[3869]), .Z(n5085) );
  AND U8936 ( .A(n16), .B(n5086), .Z(n5084) );
  XOR U8937 ( .A(n5087), .B(n5088), .Z(n5086) );
  XOR U8938 ( .A(DB[3869]), .B(DB[3838]), .Z(n5088) );
  AND U8939 ( .A(n20), .B(n5089), .Z(n5087) );
  XOR U8940 ( .A(n5090), .B(n5091), .Z(n5089) );
  XOR U8941 ( .A(DB[3838]), .B(DB[3807]), .Z(n5091) );
  AND U8942 ( .A(n24), .B(n5092), .Z(n5090) );
  XOR U8943 ( .A(n5093), .B(n5094), .Z(n5092) );
  XOR U8944 ( .A(DB[3807]), .B(DB[3776]), .Z(n5094) );
  AND U8945 ( .A(n28), .B(n5095), .Z(n5093) );
  XOR U8946 ( .A(n5096), .B(n5097), .Z(n5095) );
  XOR U8947 ( .A(DB[3776]), .B(DB[3745]), .Z(n5097) );
  AND U8948 ( .A(n32), .B(n5098), .Z(n5096) );
  XOR U8949 ( .A(n5099), .B(n5100), .Z(n5098) );
  XOR U8950 ( .A(DB[3745]), .B(DB[3714]), .Z(n5100) );
  AND U8951 ( .A(n36), .B(n5101), .Z(n5099) );
  XOR U8952 ( .A(n5102), .B(n5103), .Z(n5101) );
  XOR U8953 ( .A(DB[3714]), .B(DB[3683]), .Z(n5103) );
  AND U8954 ( .A(n40), .B(n5104), .Z(n5102) );
  XOR U8955 ( .A(n5105), .B(n5106), .Z(n5104) );
  XOR U8956 ( .A(DB[3683]), .B(DB[3652]), .Z(n5106) );
  AND U8957 ( .A(n44), .B(n5107), .Z(n5105) );
  XOR U8958 ( .A(n5108), .B(n5109), .Z(n5107) );
  XOR U8959 ( .A(DB[3652]), .B(DB[3621]), .Z(n5109) );
  AND U8960 ( .A(n48), .B(n5110), .Z(n5108) );
  XOR U8961 ( .A(n5111), .B(n5112), .Z(n5110) );
  XOR U8962 ( .A(DB[3621]), .B(DB[3590]), .Z(n5112) );
  AND U8963 ( .A(n52), .B(n5113), .Z(n5111) );
  XOR U8964 ( .A(n5114), .B(n5115), .Z(n5113) );
  XOR U8965 ( .A(DB[3590]), .B(DB[3559]), .Z(n5115) );
  AND U8966 ( .A(n56), .B(n5116), .Z(n5114) );
  XOR U8967 ( .A(n5117), .B(n5118), .Z(n5116) );
  XOR U8968 ( .A(DB[3559]), .B(DB[3528]), .Z(n5118) );
  AND U8969 ( .A(n60), .B(n5119), .Z(n5117) );
  XOR U8970 ( .A(n5120), .B(n5121), .Z(n5119) );
  XOR U8971 ( .A(DB[3528]), .B(DB[3497]), .Z(n5121) );
  AND U8972 ( .A(n64), .B(n5122), .Z(n5120) );
  XOR U8973 ( .A(n5123), .B(n5124), .Z(n5122) );
  XOR U8974 ( .A(DB[3497]), .B(DB[3466]), .Z(n5124) );
  AND U8975 ( .A(n68), .B(n5125), .Z(n5123) );
  XOR U8976 ( .A(n5126), .B(n5127), .Z(n5125) );
  XOR U8977 ( .A(DB[3466]), .B(DB[3435]), .Z(n5127) );
  AND U8978 ( .A(n72), .B(n5128), .Z(n5126) );
  XOR U8979 ( .A(n5129), .B(n5130), .Z(n5128) );
  XOR U8980 ( .A(DB[3435]), .B(DB[3404]), .Z(n5130) );
  AND U8981 ( .A(n76), .B(n5131), .Z(n5129) );
  XOR U8982 ( .A(n5132), .B(n5133), .Z(n5131) );
  XOR U8983 ( .A(DB[3404]), .B(DB[3373]), .Z(n5133) );
  AND U8984 ( .A(n80), .B(n5134), .Z(n5132) );
  XOR U8985 ( .A(n5135), .B(n5136), .Z(n5134) );
  XOR U8986 ( .A(DB[3373]), .B(DB[3342]), .Z(n5136) );
  AND U8987 ( .A(n84), .B(n5137), .Z(n5135) );
  XOR U8988 ( .A(n5138), .B(n5139), .Z(n5137) );
  XOR U8989 ( .A(DB[3342]), .B(DB[3311]), .Z(n5139) );
  AND U8990 ( .A(n88), .B(n5140), .Z(n5138) );
  XOR U8991 ( .A(n5141), .B(n5142), .Z(n5140) );
  XOR U8992 ( .A(DB[3311]), .B(DB[3280]), .Z(n5142) );
  AND U8993 ( .A(n92), .B(n5143), .Z(n5141) );
  XOR U8994 ( .A(n5144), .B(n5145), .Z(n5143) );
  XOR U8995 ( .A(DB[3280]), .B(DB[3249]), .Z(n5145) );
  AND U8996 ( .A(n96), .B(n5146), .Z(n5144) );
  XOR U8997 ( .A(n5147), .B(n5148), .Z(n5146) );
  XOR U8998 ( .A(DB[3249]), .B(DB[3218]), .Z(n5148) );
  AND U8999 ( .A(n100), .B(n5149), .Z(n5147) );
  XOR U9000 ( .A(n5150), .B(n5151), .Z(n5149) );
  XOR U9001 ( .A(DB[3218]), .B(DB[3187]), .Z(n5151) );
  AND U9002 ( .A(n104), .B(n5152), .Z(n5150) );
  XOR U9003 ( .A(n5153), .B(n5154), .Z(n5152) );
  XOR U9004 ( .A(DB[3187]), .B(DB[3156]), .Z(n5154) );
  AND U9005 ( .A(n108), .B(n5155), .Z(n5153) );
  XOR U9006 ( .A(n5156), .B(n5157), .Z(n5155) );
  XOR U9007 ( .A(DB[3156]), .B(DB[3125]), .Z(n5157) );
  AND U9008 ( .A(n112), .B(n5158), .Z(n5156) );
  XOR U9009 ( .A(n5159), .B(n5160), .Z(n5158) );
  XOR U9010 ( .A(DB[3125]), .B(DB[3094]), .Z(n5160) );
  AND U9011 ( .A(n116), .B(n5161), .Z(n5159) );
  XOR U9012 ( .A(n5162), .B(n5163), .Z(n5161) );
  XOR U9013 ( .A(DB[3094]), .B(DB[3063]), .Z(n5163) );
  AND U9014 ( .A(n120), .B(n5164), .Z(n5162) );
  XOR U9015 ( .A(n5165), .B(n5166), .Z(n5164) );
  XOR U9016 ( .A(DB[3063]), .B(DB[3032]), .Z(n5166) );
  AND U9017 ( .A(n124), .B(n5167), .Z(n5165) );
  XOR U9018 ( .A(n5168), .B(n5169), .Z(n5167) );
  XOR U9019 ( .A(DB[3032]), .B(DB[3001]), .Z(n5169) );
  AND U9020 ( .A(n128), .B(n5170), .Z(n5168) );
  XOR U9021 ( .A(n5171), .B(n5172), .Z(n5170) );
  XOR U9022 ( .A(DB[3001]), .B(DB[2970]), .Z(n5172) );
  AND U9023 ( .A(n132), .B(n5173), .Z(n5171) );
  XOR U9024 ( .A(n5174), .B(n5175), .Z(n5173) );
  XOR U9025 ( .A(DB[2970]), .B(DB[2939]), .Z(n5175) );
  AND U9026 ( .A(n136), .B(n5176), .Z(n5174) );
  XOR U9027 ( .A(n5177), .B(n5178), .Z(n5176) );
  XOR U9028 ( .A(DB[2939]), .B(DB[2908]), .Z(n5178) );
  AND U9029 ( .A(n140), .B(n5179), .Z(n5177) );
  XOR U9030 ( .A(n5180), .B(n5181), .Z(n5179) );
  XOR U9031 ( .A(DB[2908]), .B(DB[2877]), .Z(n5181) );
  AND U9032 ( .A(n144), .B(n5182), .Z(n5180) );
  XOR U9033 ( .A(n5183), .B(n5184), .Z(n5182) );
  XOR U9034 ( .A(DB[2877]), .B(DB[2846]), .Z(n5184) );
  AND U9035 ( .A(n148), .B(n5185), .Z(n5183) );
  XOR U9036 ( .A(n5186), .B(n5187), .Z(n5185) );
  XOR U9037 ( .A(DB[2846]), .B(DB[2815]), .Z(n5187) );
  AND U9038 ( .A(n152), .B(n5188), .Z(n5186) );
  XOR U9039 ( .A(n5189), .B(n5190), .Z(n5188) );
  XOR U9040 ( .A(DB[2815]), .B(DB[2784]), .Z(n5190) );
  AND U9041 ( .A(n156), .B(n5191), .Z(n5189) );
  XOR U9042 ( .A(n5192), .B(n5193), .Z(n5191) );
  XOR U9043 ( .A(DB[2784]), .B(DB[2753]), .Z(n5193) );
  AND U9044 ( .A(n160), .B(n5194), .Z(n5192) );
  XOR U9045 ( .A(n5195), .B(n5196), .Z(n5194) );
  XOR U9046 ( .A(DB[2753]), .B(DB[2722]), .Z(n5196) );
  AND U9047 ( .A(n164), .B(n5197), .Z(n5195) );
  XOR U9048 ( .A(n5198), .B(n5199), .Z(n5197) );
  XOR U9049 ( .A(DB[2722]), .B(DB[2691]), .Z(n5199) );
  AND U9050 ( .A(n168), .B(n5200), .Z(n5198) );
  XOR U9051 ( .A(n5201), .B(n5202), .Z(n5200) );
  XOR U9052 ( .A(DB[2691]), .B(DB[2660]), .Z(n5202) );
  AND U9053 ( .A(n172), .B(n5203), .Z(n5201) );
  XOR U9054 ( .A(n5204), .B(n5205), .Z(n5203) );
  XOR U9055 ( .A(DB[2660]), .B(DB[2629]), .Z(n5205) );
  AND U9056 ( .A(n176), .B(n5206), .Z(n5204) );
  XOR U9057 ( .A(n5207), .B(n5208), .Z(n5206) );
  XOR U9058 ( .A(DB[2629]), .B(DB[2598]), .Z(n5208) );
  AND U9059 ( .A(n180), .B(n5209), .Z(n5207) );
  XOR U9060 ( .A(n5210), .B(n5211), .Z(n5209) );
  XOR U9061 ( .A(DB[2598]), .B(DB[2567]), .Z(n5211) );
  AND U9062 ( .A(n184), .B(n5212), .Z(n5210) );
  XOR U9063 ( .A(n5213), .B(n5214), .Z(n5212) );
  XOR U9064 ( .A(DB[2567]), .B(DB[2536]), .Z(n5214) );
  AND U9065 ( .A(n188), .B(n5215), .Z(n5213) );
  XOR U9066 ( .A(n5216), .B(n5217), .Z(n5215) );
  XOR U9067 ( .A(DB[2536]), .B(DB[2505]), .Z(n5217) );
  AND U9068 ( .A(n192), .B(n5218), .Z(n5216) );
  XOR U9069 ( .A(n5219), .B(n5220), .Z(n5218) );
  XOR U9070 ( .A(DB[2505]), .B(DB[2474]), .Z(n5220) );
  AND U9071 ( .A(n196), .B(n5221), .Z(n5219) );
  XOR U9072 ( .A(n5222), .B(n5223), .Z(n5221) );
  XOR U9073 ( .A(DB[2474]), .B(DB[2443]), .Z(n5223) );
  AND U9074 ( .A(n200), .B(n5224), .Z(n5222) );
  XOR U9075 ( .A(n5225), .B(n5226), .Z(n5224) );
  XOR U9076 ( .A(DB[2443]), .B(DB[2412]), .Z(n5226) );
  AND U9077 ( .A(n204), .B(n5227), .Z(n5225) );
  XOR U9078 ( .A(n5228), .B(n5229), .Z(n5227) );
  XOR U9079 ( .A(DB[2412]), .B(DB[2381]), .Z(n5229) );
  AND U9080 ( .A(n208), .B(n5230), .Z(n5228) );
  XOR U9081 ( .A(n5231), .B(n5232), .Z(n5230) );
  XOR U9082 ( .A(DB[2381]), .B(DB[2350]), .Z(n5232) );
  AND U9083 ( .A(n212), .B(n5233), .Z(n5231) );
  XOR U9084 ( .A(n5234), .B(n5235), .Z(n5233) );
  XOR U9085 ( .A(DB[2350]), .B(DB[2319]), .Z(n5235) );
  AND U9086 ( .A(n216), .B(n5236), .Z(n5234) );
  XOR U9087 ( .A(n5237), .B(n5238), .Z(n5236) );
  XOR U9088 ( .A(DB[2319]), .B(DB[2288]), .Z(n5238) );
  AND U9089 ( .A(n220), .B(n5239), .Z(n5237) );
  XOR U9090 ( .A(n5240), .B(n5241), .Z(n5239) );
  XOR U9091 ( .A(DB[2288]), .B(DB[2257]), .Z(n5241) );
  AND U9092 ( .A(n224), .B(n5242), .Z(n5240) );
  XOR U9093 ( .A(n5243), .B(n5244), .Z(n5242) );
  XOR U9094 ( .A(DB[2257]), .B(DB[2226]), .Z(n5244) );
  AND U9095 ( .A(n228), .B(n5245), .Z(n5243) );
  XOR U9096 ( .A(n5246), .B(n5247), .Z(n5245) );
  XOR U9097 ( .A(DB[2226]), .B(DB[2195]), .Z(n5247) );
  AND U9098 ( .A(n232), .B(n5248), .Z(n5246) );
  XOR U9099 ( .A(n5249), .B(n5250), .Z(n5248) );
  XOR U9100 ( .A(DB[2195]), .B(DB[2164]), .Z(n5250) );
  AND U9101 ( .A(n236), .B(n5251), .Z(n5249) );
  XOR U9102 ( .A(n5252), .B(n5253), .Z(n5251) );
  XOR U9103 ( .A(DB[2164]), .B(DB[2133]), .Z(n5253) );
  AND U9104 ( .A(n240), .B(n5254), .Z(n5252) );
  XOR U9105 ( .A(n5255), .B(n5256), .Z(n5254) );
  XOR U9106 ( .A(DB[2133]), .B(DB[2102]), .Z(n5256) );
  AND U9107 ( .A(n244), .B(n5257), .Z(n5255) );
  XOR U9108 ( .A(n5258), .B(n5259), .Z(n5257) );
  XOR U9109 ( .A(DB[2102]), .B(DB[2071]), .Z(n5259) );
  AND U9110 ( .A(n248), .B(n5260), .Z(n5258) );
  XOR U9111 ( .A(n5261), .B(n5262), .Z(n5260) );
  XOR U9112 ( .A(DB[2071]), .B(DB[2040]), .Z(n5262) );
  AND U9113 ( .A(n252), .B(n5263), .Z(n5261) );
  XOR U9114 ( .A(n5264), .B(n5265), .Z(n5263) );
  XOR U9115 ( .A(DB[2040]), .B(DB[2009]), .Z(n5265) );
  AND U9116 ( .A(n256), .B(n5266), .Z(n5264) );
  XOR U9117 ( .A(n5267), .B(n5268), .Z(n5266) );
  XOR U9118 ( .A(DB[2009]), .B(DB[1978]), .Z(n5268) );
  AND U9119 ( .A(n260), .B(n5269), .Z(n5267) );
  XOR U9120 ( .A(n5270), .B(n5271), .Z(n5269) );
  XOR U9121 ( .A(DB[1978]), .B(DB[1947]), .Z(n5271) );
  AND U9122 ( .A(n264), .B(n5272), .Z(n5270) );
  XOR U9123 ( .A(n5273), .B(n5274), .Z(n5272) );
  XOR U9124 ( .A(DB[1947]), .B(DB[1916]), .Z(n5274) );
  AND U9125 ( .A(n268), .B(n5275), .Z(n5273) );
  XOR U9126 ( .A(n5276), .B(n5277), .Z(n5275) );
  XOR U9127 ( .A(DB[1916]), .B(DB[1885]), .Z(n5277) );
  AND U9128 ( .A(n272), .B(n5278), .Z(n5276) );
  XOR U9129 ( .A(n5279), .B(n5280), .Z(n5278) );
  XOR U9130 ( .A(DB[1885]), .B(DB[1854]), .Z(n5280) );
  AND U9131 ( .A(n276), .B(n5281), .Z(n5279) );
  XOR U9132 ( .A(n5282), .B(n5283), .Z(n5281) );
  XOR U9133 ( .A(DB[1854]), .B(DB[1823]), .Z(n5283) );
  AND U9134 ( .A(n280), .B(n5284), .Z(n5282) );
  XOR U9135 ( .A(n5285), .B(n5286), .Z(n5284) );
  XOR U9136 ( .A(DB[1823]), .B(DB[1792]), .Z(n5286) );
  AND U9137 ( .A(n284), .B(n5287), .Z(n5285) );
  XOR U9138 ( .A(n5288), .B(n5289), .Z(n5287) );
  XOR U9139 ( .A(DB[1792]), .B(DB[1761]), .Z(n5289) );
  AND U9140 ( .A(n288), .B(n5290), .Z(n5288) );
  XOR U9141 ( .A(n5291), .B(n5292), .Z(n5290) );
  XOR U9142 ( .A(DB[1761]), .B(DB[1730]), .Z(n5292) );
  AND U9143 ( .A(n292), .B(n5293), .Z(n5291) );
  XOR U9144 ( .A(n5294), .B(n5295), .Z(n5293) );
  XOR U9145 ( .A(DB[1730]), .B(DB[1699]), .Z(n5295) );
  AND U9146 ( .A(n296), .B(n5296), .Z(n5294) );
  XOR U9147 ( .A(n5297), .B(n5298), .Z(n5296) );
  XOR U9148 ( .A(DB[1699]), .B(DB[1668]), .Z(n5298) );
  AND U9149 ( .A(n300), .B(n5299), .Z(n5297) );
  XOR U9150 ( .A(n5300), .B(n5301), .Z(n5299) );
  XOR U9151 ( .A(DB[1668]), .B(DB[1637]), .Z(n5301) );
  AND U9152 ( .A(n304), .B(n5302), .Z(n5300) );
  XOR U9153 ( .A(n5303), .B(n5304), .Z(n5302) );
  XOR U9154 ( .A(DB[1637]), .B(DB[1606]), .Z(n5304) );
  AND U9155 ( .A(n308), .B(n5305), .Z(n5303) );
  XOR U9156 ( .A(n5306), .B(n5307), .Z(n5305) );
  XOR U9157 ( .A(DB[1606]), .B(DB[1575]), .Z(n5307) );
  AND U9158 ( .A(n312), .B(n5308), .Z(n5306) );
  XOR U9159 ( .A(n5309), .B(n5310), .Z(n5308) );
  XOR U9160 ( .A(DB[1575]), .B(DB[1544]), .Z(n5310) );
  AND U9161 ( .A(n316), .B(n5311), .Z(n5309) );
  XOR U9162 ( .A(n5312), .B(n5313), .Z(n5311) );
  XOR U9163 ( .A(DB[1544]), .B(DB[1513]), .Z(n5313) );
  AND U9164 ( .A(n320), .B(n5314), .Z(n5312) );
  XOR U9165 ( .A(n5315), .B(n5316), .Z(n5314) );
  XOR U9166 ( .A(DB[1513]), .B(DB[1482]), .Z(n5316) );
  AND U9167 ( .A(n324), .B(n5317), .Z(n5315) );
  XOR U9168 ( .A(n5318), .B(n5319), .Z(n5317) );
  XOR U9169 ( .A(DB[1482]), .B(DB[1451]), .Z(n5319) );
  AND U9170 ( .A(n328), .B(n5320), .Z(n5318) );
  XOR U9171 ( .A(n5321), .B(n5322), .Z(n5320) );
  XOR U9172 ( .A(DB[1451]), .B(DB[1420]), .Z(n5322) );
  AND U9173 ( .A(n332), .B(n5323), .Z(n5321) );
  XOR U9174 ( .A(n5324), .B(n5325), .Z(n5323) );
  XOR U9175 ( .A(DB[1420]), .B(DB[1389]), .Z(n5325) );
  AND U9176 ( .A(n336), .B(n5326), .Z(n5324) );
  XOR U9177 ( .A(n5327), .B(n5328), .Z(n5326) );
  XOR U9178 ( .A(DB[1389]), .B(DB[1358]), .Z(n5328) );
  AND U9179 ( .A(n340), .B(n5329), .Z(n5327) );
  XOR U9180 ( .A(n5330), .B(n5331), .Z(n5329) );
  XOR U9181 ( .A(DB[1358]), .B(DB[1327]), .Z(n5331) );
  AND U9182 ( .A(n344), .B(n5332), .Z(n5330) );
  XOR U9183 ( .A(n5333), .B(n5334), .Z(n5332) );
  XOR U9184 ( .A(DB[1327]), .B(DB[1296]), .Z(n5334) );
  AND U9185 ( .A(n348), .B(n5335), .Z(n5333) );
  XOR U9186 ( .A(n5336), .B(n5337), .Z(n5335) );
  XOR U9187 ( .A(DB[1296]), .B(DB[1265]), .Z(n5337) );
  AND U9188 ( .A(n352), .B(n5338), .Z(n5336) );
  XOR U9189 ( .A(n5339), .B(n5340), .Z(n5338) );
  XOR U9190 ( .A(DB[1265]), .B(DB[1234]), .Z(n5340) );
  AND U9191 ( .A(n356), .B(n5341), .Z(n5339) );
  XOR U9192 ( .A(n5342), .B(n5343), .Z(n5341) );
  XOR U9193 ( .A(DB[1234]), .B(DB[1203]), .Z(n5343) );
  AND U9194 ( .A(n360), .B(n5344), .Z(n5342) );
  XOR U9195 ( .A(n5345), .B(n5346), .Z(n5344) );
  XOR U9196 ( .A(DB[1203]), .B(DB[1172]), .Z(n5346) );
  AND U9197 ( .A(n364), .B(n5347), .Z(n5345) );
  XOR U9198 ( .A(n5348), .B(n5349), .Z(n5347) );
  XOR U9199 ( .A(DB[1172]), .B(DB[1141]), .Z(n5349) );
  AND U9200 ( .A(n368), .B(n5350), .Z(n5348) );
  XOR U9201 ( .A(n5351), .B(n5352), .Z(n5350) );
  XOR U9202 ( .A(DB[1141]), .B(DB[1110]), .Z(n5352) );
  AND U9203 ( .A(n372), .B(n5353), .Z(n5351) );
  XOR U9204 ( .A(n5354), .B(n5355), .Z(n5353) );
  XOR U9205 ( .A(DB[1110]), .B(DB[1079]), .Z(n5355) );
  AND U9206 ( .A(n376), .B(n5356), .Z(n5354) );
  XOR U9207 ( .A(n5357), .B(n5358), .Z(n5356) );
  XOR U9208 ( .A(DB[1079]), .B(DB[1048]), .Z(n5358) );
  AND U9209 ( .A(n380), .B(n5359), .Z(n5357) );
  XOR U9210 ( .A(n5360), .B(n5361), .Z(n5359) );
  XOR U9211 ( .A(DB[1048]), .B(DB[1017]), .Z(n5361) );
  AND U9212 ( .A(n384), .B(n5362), .Z(n5360) );
  XOR U9213 ( .A(n5363), .B(n5364), .Z(n5362) );
  XOR U9214 ( .A(DB[986]), .B(DB[1017]), .Z(n5364) );
  AND U9215 ( .A(n388), .B(n5365), .Z(n5363) );
  XOR U9216 ( .A(n5366), .B(n5367), .Z(n5365) );
  XOR U9217 ( .A(DB[986]), .B(DB[955]), .Z(n5367) );
  AND U9218 ( .A(n392), .B(n5368), .Z(n5366) );
  XOR U9219 ( .A(n5369), .B(n5370), .Z(n5368) );
  XOR U9220 ( .A(DB[955]), .B(DB[924]), .Z(n5370) );
  AND U9221 ( .A(n396), .B(n5371), .Z(n5369) );
  XOR U9222 ( .A(n5372), .B(n5373), .Z(n5371) );
  XOR U9223 ( .A(DB[924]), .B(DB[893]), .Z(n5373) );
  AND U9224 ( .A(n400), .B(n5374), .Z(n5372) );
  XOR U9225 ( .A(n5375), .B(n5376), .Z(n5374) );
  XOR U9226 ( .A(DB[893]), .B(DB[862]), .Z(n5376) );
  AND U9227 ( .A(n404), .B(n5377), .Z(n5375) );
  XOR U9228 ( .A(n5378), .B(n5379), .Z(n5377) );
  XOR U9229 ( .A(DB[862]), .B(DB[831]), .Z(n5379) );
  AND U9230 ( .A(n408), .B(n5380), .Z(n5378) );
  XOR U9231 ( .A(n5381), .B(n5382), .Z(n5380) );
  XOR U9232 ( .A(DB[831]), .B(DB[800]), .Z(n5382) );
  AND U9233 ( .A(n412), .B(n5383), .Z(n5381) );
  XOR U9234 ( .A(n5384), .B(n5385), .Z(n5383) );
  XOR U9235 ( .A(DB[800]), .B(DB[769]), .Z(n5385) );
  AND U9236 ( .A(n416), .B(n5386), .Z(n5384) );
  XOR U9237 ( .A(n5387), .B(n5388), .Z(n5386) );
  XOR U9238 ( .A(DB[769]), .B(DB[738]), .Z(n5388) );
  AND U9239 ( .A(n420), .B(n5389), .Z(n5387) );
  XOR U9240 ( .A(n5390), .B(n5391), .Z(n5389) );
  XOR U9241 ( .A(DB[738]), .B(DB[707]), .Z(n5391) );
  AND U9242 ( .A(n424), .B(n5392), .Z(n5390) );
  XOR U9243 ( .A(n5393), .B(n5394), .Z(n5392) );
  XOR U9244 ( .A(DB[707]), .B(DB[676]), .Z(n5394) );
  AND U9245 ( .A(n428), .B(n5395), .Z(n5393) );
  XOR U9246 ( .A(n5396), .B(n5397), .Z(n5395) );
  XOR U9247 ( .A(DB[676]), .B(DB[645]), .Z(n5397) );
  AND U9248 ( .A(n432), .B(n5398), .Z(n5396) );
  XOR U9249 ( .A(n5399), .B(n5400), .Z(n5398) );
  XOR U9250 ( .A(DB[645]), .B(DB[614]), .Z(n5400) );
  AND U9251 ( .A(n436), .B(n5401), .Z(n5399) );
  XOR U9252 ( .A(n5402), .B(n5403), .Z(n5401) );
  XOR U9253 ( .A(DB[614]), .B(DB[583]), .Z(n5403) );
  AND U9254 ( .A(n440), .B(n5404), .Z(n5402) );
  XOR U9255 ( .A(n5405), .B(n5406), .Z(n5404) );
  XOR U9256 ( .A(DB[583]), .B(DB[552]), .Z(n5406) );
  AND U9257 ( .A(n444), .B(n5407), .Z(n5405) );
  XOR U9258 ( .A(n5408), .B(n5409), .Z(n5407) );
  XOR U9259 ( .A(DB[552]), .B(DB[521]), .Z(n5409) );
  AND U9260 ( .A(n448), .B(n5410), .Z(n5408) );
  XOR U9261 ( .A(n5411), .B(n5412), .Z(n5410) );
  XOR U9262 ( .A(DB[521]), .B(DB[490]), .Z(n5412) );
  AND U9263 ( .A(n452), .B(n5413), .Z(n5411) );
  XOR U9264 ( .A(n5414), .B(n5415), .Z(n5413) );
  XOR U9265 ( .A(DB[490]), .B(DB[459]), .Z(n5415) );
  AND U9266 ( .A(n456), .B(n5416), .Z(n5414) );
  XOR U9267 ( .A(n5417), .B(n5418), .Z(n5416) );
  XOR U9268 ( .A(DB[459]), .B(DB[428]), .Z(n5418) );
  AND U9269 ( .A(n460), .B(n5419), .Z(n5417) );
  XOR U9270 ( .A(n5420), .B(n5421), .Z(n5419) );
  XOR U9271 ( .A(DB[428]), .B(DB[397]), .Z(n5421) );
  AND U9272 ( .A(n464), .B(n5422), .Z(n5420) );
  XOR U9273 ( .A(n5423), .B(n5424), .Z(n5422) );
  XOR U9274 ( .A(DB[397]), .B(DB[366]), .Z(n5424) );
  AND U9275 ( .A(n468), .B(n5425), .Z(n5423) );
  XOR U9276 ( .A(n5426), .B(n5427), .Z(n5425) );
  XOR U9277 ( .A(DB[366]), .B(DB[335]), .Z(n5427) );
  AND U9278 ( .A(n472), .B(n5428), .Z(n5426) );
  XOR U9279 ( .A(n5429), .B(n5430), .Z(n5428) );
  XOR U9280 ( .A(DB[335]), .B(DB[304]), .Z(n5430) );
  AND U9281 ( .A(n476), .B(n5431), .Z(n5429) );
  XOR U9282 ( .A(n5432), .B(n5433), .Z(n5431) );
  XOR U9283 ( .A(DB[304]), .B(DB[273]), .Z(n5433) );
  AND U9284 ( .A(n480), .B(n5434), .Z(n5432) );
  XOR U9285 ( .A(n5435), .B(n5436), .Z(n5434) );
  XOR U9286 ( .A(DB[273]), .B(DB[242]), .Z(n5436) );
  AND U9287 ( .A(n484), .B(n5437), .Z(n5435) );
  XOR U9288 ( .A(n5438), .B(n5439), .Z(n5437) );
  XOR U9289 ( .A(DB[242]), .B(DB[211]), .Z(n5439) );
  AND U9290 ( .A(n488), .B(n5440), .Z(n5438) );
  XOR U9291 ( .A(n5441), .B(n5442), .Z(n5440) );
  XOR U9292 ( .A(DB[211]), .B(DB[180]), .Z(n5442) );
  AND U9293 ( .A(n492), .B(n5443), .Z(n5441) );
  XOR U9294 ( .A(n5444), .B(n5445), .Z(n5443) );
  XOR U9295 ( .A(DB[180]), .B(DB[149]), .Z(n5445) );
  AND U9296 ( .A(n496), .B(n5446), .Z(n5444) );
  XOR U9297 ( .A(n5447), .B(n5448), .Z(n5446) );
  XOR U9298 ( .A(DB[149]), .B(DB[118]), .Z(n5448) );
  AND U9299 ( .A(n500), .B(n5449), .Z(n5447) );
  XOR U9300 ( .A(n5450), .B(n5451), .Z(n5449) );
  XOR U9301 ( .A(DB[87]), .B(DB[118]), .Z(n5451) );
  AND U9302 ( .A(n504), .B(n5452), .Z(n5450) );
  XOR U9303 ( .A(n5453), .B(n5454), .Z(n5452) );
  XOR U9304 ( .A(DB[87]), .B(DB[56]), .Z(n5454) );
  AND U9305 ( .A(n508), .B(n5455), .Z(n5453) );
  XOR U9306 ( .A(DB[56]), .B(DB[25]), .Z(n5455) );
  XOR U9307 ( .A(DB[3961]), .B(n5456), .Z(min_val_out[24]) );
  AND U9308 ( .A(n2), .B(n5457), .Z(n5456) );
  XOR U9309 ( .A(n5458), .B(n5459), .Z(n5457) );
  XOR U9310 ( .A(n5460), .B(n5461), .Z(n5459) );
  IV U9311 ( .A(DB[3961]), .Z(n5460) );
  AND U9312 ( .A(n8), .B(n5462), .Z(n5458) );
  XOR U9313 ( .A(n5463), .B(n5464), .Z(n5462) );
  XOR U9314 ( .A(DB[3930]), .B(DB[3899]), .Z(n5464) );
  AND U9315 ( .A(n12), .B(n5465), .Z(n5463) );
  XOR U9316 ( .A(n5466), .B(n5467), .Z(n5465) );
  XOR U9317 ( .A(DB[3899]), .B(DB[3868]), .Z(n5467) );
  AND U9318 ( .A(n16), .B(n5468), .Z(n5466) );
  XOR U9319 ( .A(n5469), .B(n5470), .Z(n5468) );
  XOR U9320 ( .A(DB[3868]), .B(DB[3837]), .Z(n5470) );
  AND U9321 ( .A(n20), .B(n5471), .Z(n5469) );
  XOR U9322 ( .A(n5472), .B(n5473), .Z(n5471) );
  XOR U9323 ( .A(DB[3837]), .B(DB[3806]), .Z(n5473) );
  AND U9324 ( .A(n24), .B(n5474), .Z(n5472) );
  XOR U9325 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U9326 ( .A(DB[3806]), .B(DB[3775]), .Z(n5476) );
  AND U9327 ( .A(n28), .B(n5477), .Z(n5475) );
  XOR U9328 ( .A(n5478), .B(n5479), .Z(n5477) );
  XOR U9329 ( .A(DB[3775]), .B(DB[3744]), .Z(n5479) );
  AND U9330 ( .A(n32), .B(n5480), .Z(n5478) );
  XOR U9331 ( .A(n5481), .B(n5482), .Z(n5480) );
  XOR U9332 ( .A(DB[3744]), .B(DB[3713]), .Z(n5482) );
  AND U9333 ( .A(n36), .B(n5483), .Z(n5481) );
  XOR U9334 ( .A(n5484), .B(n5485), .Z(n5483) );
  XOR U9335 ( .A(DB[3713]), .B(DB[3682]), .Z(n5485) );
  AND U9336 ( .A(n40), .B(n5486), .Z(n5484) );
  XOR U9337 ( .A(n5487), .B(n5488), .Z(n5486) );
  XOR U9338 ( .A(DB[3682]), .B(DB[3651]), .Z(n5488) );
  AND U9339 ( .A(n44), .B(n5489), .Z(n5487) );
  XOR U9340 ( .A(n5490), .B(n5491), .Z(n5489) );
  XOR U9341 ( .A(DB[3651]), .B(DB[3620]), .Z(n5491) );
  AND U9342 ( .A(n48), .B(n5492), .Z(n5490) );
  XOR U9343 ( .A(n5493), .B(n5494), .Z(n5492) );
  XOR U9344 ( .A(DB[3620]), .B(DB[3589]), .Z(n5494) );
  AND U9345 ( .A(n52), .B(n5495), .Z(n5493) );
  XOR U9346 ( .A(n5496), .B(n5497), .Z(n5495) );
  XOR U9347 ( .A(DB[3589]), .B(DB[3558]), .Z(n5497) );
  AND U9348 ( .A(n56), .B(n5498), .Z(n5496) );
  XOR U9349 ( .A(n5499), .B(n5500), .Z(n5498) );
  XOR U9350 ( .A(DB[3558]), .B(DB[3527]), .Z(n5500) );
  AND U9351 ( .A(n60), .B(n5501), .Z(n5499) );
  XOR U9352 ( .A(n5502), .B(n5503), .Z(n5501) );
  XOR U9353 ( .A(DB[3527]), .B(DB[3496]), .Z(n5503) );
  AND U9354 ( .A(n64), .B(n5504), .Z(n5502) );
  XOR U9355 ( .A(n5505), .B(n5506), .Z(n5504) );
  XOR U9356 ( .A(DB[3496]), .B(DB[3465]), .Z(n5506) );
  AND U9357 ( .A(n68), .B(n5507), .Z(n5505) );
  XOR U9358 ( .A(n5508), .B(n5509), .Z(n5507) );
  XOR U9359 ( .A(DB[3465]), .B(DB[3434]), .Z(n5509) );
  AND U9360 ( .A(n72), .B(n5510), .Z(n5508) );
  XOR U9361 ( .A(n5511), .B(n5512), .Z(n5510) );
  XOR U9362 ( .A(DB[3434]), .B(DB[3403]), .Z(n5512) );
  AND U9363 ( .A(n76), .B(n5513), .Z(n5511) );
  XOR U9364 ( .A(n5514), .B(n5515), .Z(n5513) );
  XOR U9365 ( .A(DB[3403]), .B(DB[3372]), .Z(n5515) );
  AND U9366 ( .A(n80), .B(n5516), .Z(n5514) );
  XOR U9367 ( .A(n5517), .B(n5518), .Z(n5516) );
  XOR U9368 ( .A(DB[3372]), .B(DB[3341]), .Z(n5518) );
  AND U9369 ( .A(n84), .B(n5519), .Z(n5517) );
  XOR U9370 ( .A(n5520), .B(n5521), .Z(n5519) );
  XOR U9371 ( .A(DB[3341]), .B(DB[3310]), .Z(n5521) );
  AND U9372 ( .A(n88), .B(n5522), .Z(n5520) );
  XOR U9373 ( .A(n5523), .B(n5524), .Z(n5522) );
  XOR U9374 ( .A(DB[3310]), .B(DB[3279]), .Z(n5524) );
  AND U9375 ( .A(n92), .B(n5525), .Z(n5523) );
  XOR U9376 ( .A(n5526), .B(n5527), .Z(n5525) );
  XOR U9377 ( .A(DB[3279]), .B(DB[3248]), .Z(n5527) );
  AND U9378 ( .A(n96), .B(n5528), .Z(n5526) );
  XOR U9379 ( .A(n5529), .B(n5530), .Z(n5528) );
  XOR U9380 ( .A(DB[3248]), .B(DB[3217]), .Z(n5530) );
  AND U9381 ( .A(n100), .B(n5531), .Z(n5529) );
  XOR U9382 ( .A(n5532), .B(n5533), .Z(n5531) );
  XOR U9383 ( .A(DB[3217]), .B(DB[3186]), .Z(n5533) );
  AND U9384 ( .A(n104), .B(n5534), .Z(n5532) );
  XOR U9385 ( .A(n5535), .B(n5536), .Z(n5534) );
  XOR U9386 ( .A(DB[3186]), .B(DB[3155]), .Z(n5536) );
  AND U9387 ( .A(n108), .B(n5537), .Z(n5535) );
  XOR U9388 ( .A(n5538), .B(n5539), .Z(n5537) );
  XOR U9389 ( .A(DB[3155]), .B(DB[3124]), .Z(n5539) );
  AND U9390 ( .A(n112), .B(n5540), .Z(n5538) );
  XOR U9391 ( .A(n5541), .B(n5542), .Z(n5540) );
  XOR U9392 ( .A(DB[3124]), .B(DB[3093]), .Z(n5542) );
  AND U9393 ( .A(n116), .B(n5543), .Z(n5541) );
  XOR U9394 ( .A(n5544), .B(n5545), .Z(n5543) );
  XOR U9395 ( .A(DB[3093]), .B(DB[3062]), .Z(n5545) );
  AND U9396 ( .A(n120), .B(n5546), .Z(n5544) );
  XOR U9397 ( .A(n5547), .B(n5548), .Z(n5546) );
  XOR U9398 ( .A(DB[3062]), .B(DB[3031]), .Z(n5548) );
  AND U9399 ( .A(n124), .B(n5549), .Z(n5547) );
  XOR U9400 ( .A(n5550), .B(n5551), .Z(n5549) );
  XOR U9401 ( .A(DB[3031]), .B(DB[3000]), .Z(n5551) );
  AND U9402 ( .A(n128), .B(n5552), .Z(n5550) );
  XOR U9403 ( .A(n5553), .B(n5554), .Z(n5552) );
  XOR U9404 ( .A(DB[3000]), .B(DB[2969]), .Z(n5554) );
  AND U9405 ( .A(n132), .B(n5555), .Z(n5553) );
  XOR U9406 ( .A(n5556), .B(n5557), .Z(n5555) );
  XOR U9407 ( .A(DB[2969]), .B(DB[2938]), .Z(n5557) );
  AND U9408 ( .A(n136), .B(n5558), .Z(n5556) );
  XOR U9409 ( .A(n5559), .B(n5560), .Z(n5558) );
  XOR U9410 ( .A(DB[2938]), .B(DB[2907]), .Z(n5560) );
  AND U9411 ( .A(n140), .B(n5561), .Z(n5559) );
  XOR U9412 ( .A(n5562), .B(n5563), .Z(n5561) );
  XOR U9413 ( .A(DB[2907]), .B(DB[2876]), .Z(n5563) );
  AND U9414 ( .A(n144), .B(n5564), .Z(n5562) );
  XOR U9415 ( .A(n5565), .B(n5566), .Z(n5564) );
  XOR U9416 ( .A(DB[2876]), .B(DB[2845]), .Z(n5566) );
  AND U9417 ( .A(n148), .B(n5567), .Z(n5565) );
  XOR U9418 ( .A(n5568), .B(n5569), .Z(n5567) );
  XOR U9419 ( .A(DB[2845]), .B(DB[2814]), .Z(n5569) );
  AND U9420 ( .A(n152), .B(n5570), .Z(n5568) );
  XOR U9421 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U9422 ( .A(DB[2814]), .B(DB[2783]), .Z(n5572) );
  AND U9423 ( .A(n156), .B(n5573), .Z(n5571) );
  XOR U9424 ( .A(n5574), .B(n5575), .Z(n5573) );
  XOR U9425 ( .A(DB[2783]), .B(DB[2752]), .Z(n5575) );
  AND U9426 ( .A(n160), .B(n5576), .Z(n5574) );
  XOR U9427 ( .A(n5577), .B(n5578), .Z(n5576) );
  XOR U9428 ( .A(DB[2752]), .B(DB[2721]), .Z(n5578) );
  AND U9429 ( .A(n164), .B(n5579), .Z(n5577) );
  XOR U9430 ( .A(n5580), .B(n5581), .Z(n5579) );
  XOR U9431 ( .A(DB[2721]), .B(DB[2690]), .Z(n5581) );
  AND U9432 ( .A(n168), .B(n5582), .Z(n5580) );
  XOR U9433 ( .A(n5583), .B(n5584), .Z(n5582) );
  XOR U9434 ( .A(DB[2690]), .B(DB[2659]), .Z(n5584) );
  AND U9435 ( .A(n172), .B(n5585), .Z(n5583) );
  XOR U9436 ( .A(n5586), .B(n5587), .Z(n5585) );
  XOR U9437 ( .A(DB[2659]), .B(DB[2628]), .Z(n5587) );
  AND U9438 ( .A(n176), .B(n5588), .Z(n5586) );
  XOR U9439 ( .A(n5589), .B(n5590), .Z(n5588) );
  XOR U9440 ( .A(DB[2628]), .B(DB[2597]), .Z(n5590) );
  AND U9441 ( .A(n180), .B(n5591), .Z(n5589) );
  XOR U9442 ( .A(n5592), .B(n5593), .Z(n5591) );
  XOR U9443 ( .A(DB[2597]), .B(DB[2566]), .Z(n5593) );
  AND U9444 ( .A(n184), .B(n5594), .Z(n5592) );
  XOR U9445 ( .A(n5595), .B(n5596), .Z(n5594) );
  XOR U9446 ( .A(DB[2566]), .B(DB[2535]), .Z(n5596) );
  AND U9447 ( .A(n188), .B(n5597), .Z(n5595) );
  XOR U9448 ( .A(n5598), .B(n5599), .Z(n5597) );
  XOR U9449 ( .A(DB[2535]), .B(DB[2504]), .Z(n5599) );
  AND U9450 ( .A(n192), .B(n5600), .Z(n5598) );
  XOR U9451 ( .A(n5601), .B(n5602), .Z(n5600) );
  XOR U9452 ( .A(DB[2504]), .B(DB[2473]), .Z(n5602) );
  AND U9453 ( .A(n196), .B(n5603), .Z(n5601) );
  XOR U9454 ( .A(n5604), .B(n5605), .Z(n5603) );
  XOR U9455 ( .A(DB[2473]), .B(DB[2442]), .Z(n5605) );
  AND U9456 ( .A(n200), .B(n5606), .Z(n5604) );
  XOR U9457 ( .A(n5607), .B(n5608), .Z(n5606) );
  XOR U9458 ( .A(DB[2442]), .B(DB[2411]), .Z(n5608) );
  AND U9459 ( .A(n204), .B(n5609), .Z(n5607) );
  XOR U9460 ( .A(n5610), .B(n5611), .Z(n5609) );
  XOR U9461 ( .A(DB[2411]), .B(DB[2380]), .Z(n5611) );
  AND U9462 ( .A(n208), .B(n5612), .Z(n5610) );
  XOR U9463 ( .A(n5613), .B(n5614), .Z(n5612) );
  XOR U9464 ( .A(DB[2380]), .B(DB[2349]), .Z(n5614) );
  AND U9465 ( .A(n212), .B(n5615), .Z(n5613) );
  XOR U9466 ( .A(n5616), .B(n5617), .Z(n5615) );
  XOR U9467 ( .A(DB[2349]), .B(DB[2318]), .Z(n5617) );
  AND U9468 ( .A(n216), .B(n5618), .Z(n5616) );
  XOR U9469 ( .A(n5619), .B(n5620), .Z(n5618) );
  XOR U9470 ( .A(DB[2318]), .B(DB[2287]), .Z(n5620) );
  AND U9471 ( .A(n220), .B(n5621), .Z(n5619) );
  XOR U9472 ( .A(n5622), .B(n5623), .Z(n5621) );
  XOR U9473 ( .A(DB[2287]), .B(DB[2256]), .Z(n5623) );
  AND U9474 ( .A(n224), .B(n5624), .Z(n5622) );
  XOR U9475 ( .A(n5625), .B(n5626), .Z(n5624) );
  XOR U9476 ( .A(DB[2256]), .B(DB[2225]), .Z(n5626) );
  AND U9477 ( .A(n228), .B(n5627), .Z(n5625) );
  XOR U9478 ( .A(n5628), .B(n5629), .Z(n5627) );
  XOR U9479 ( .A(DB[2225]), .B(DB[2194]), .Z(n5629) );
  AND U9480 ( .A(n232), .B(n5630), .Z(n5628) );
  XOR U9481 ( .A(n5631), .B(n5632), .Z(n5630) );
  XOR U9482 ( .A(DB[2194]), .B(DB[2163]), .Z(n5632) );
  AND U9483 ( .A(n236), .B(n5633), .Z(n5631) );
  XOR U9484 ( .A(n5634), .B(n5635), .Z(n5633) );
  XOR U9485 ( .A(DB[2163]), .B(DB[2132]), .Z(n5635) );
  AND U9486 ( .A(n240), .B(n5636), .Z(n5634) );
  XOR U9487 ( .A(n5637), .B(n5638), .Z(n5636) );
  XOR U9488 ( .A(DB[2132]), .B(DB[2101]), .Z(n5638) );
  AND U9489 ( .A(n244), .B(n5639), .Z(n5637) );
  XOR U9490 ( .A(n5640), .B(n5641), .Z(n5639) );
  XOR U9491 ( .A(DB[2101]), .B(DB[2070]), .Z(n5641) );
  AND U9492 ( .A(n248), .B(n5642), .Z(n5640) );
  XOR U9493 ( .A(n5643), .B(n5644), .Z(n5642) );
  XOR U9494 ( .A(DB[2070]), .B(DB[2039]), .Z(n5644) );
  AND U9495 ( .A(n252), .B(n5645), .Z(n5643) );
  XOR U9496 ( .A(n5646), .B(n5647), .Z(n5645) );
  XOR U9497 ( .A(DB[2039]), .B(DB[2008]), .Z(n5647) );
  AND U9498 ( .A(n256), .B(n5648), .Z(n5646) );
  XOR U9499 ( .A(n5649), .B(n5650), .Z(n5648) );
  XOR U9500 ( .A(DB[2008]), .B(DB[1977]), .Z(n5650) );
  AND U9501 ( .A(n260), .B(n5651), .Z(n5649) );
  XOR U9502 ( .A(n5652), .B(n5653), .Z(n5651) );
  XOR U9503 ( .A(DB[1977]), .B(DB[1946]), .Z(n5653) );
  AND U9504 ( .A(n264), .B(n5654), .Z(n5652) );
  XOR U9505 ( .A(n5655), .B(n5656), .Z(n5654) );
  XOR U9506 ( .A(DB[1946]), .B(DB[1915]), .Z(n5656) );
  AND U9507 ( .A(n268), .B(n5657), .Z(n5655) );
  XOR U9508 ( .A(n5658), .B(n5659), .Z(n5657) );
  XOR U9509 ( .A(DB[1915]), .B(DB[1884]), .Z(n5659) );
  AND U9510 ( .A(n272), .B(n5660), .Z(n5658) );
  XOR U9511 ( .A(n5661), .B(n5662), .Z(n5660) );
  XOR U9512 ( .A(DB[1884]), .B(DB[1853]), .Z(n5662) );
  AND U9513 ( .A(n276), .B(n5663), .Z(n5661) );
  XOR U9514 ( .A(n5664), .B(n5665), .Z(n5663) );
  XOR U9515 ( .A(DB[1853]), .B(DB[1822]), .Z(n5665) );
  AND U9516 ( .A(n280), .B(n5666), .Z(n5664) );
  XOR U9517 ( .A(n5667), .B(n5668), .Z(n5666) );
  XOR U9518 ( .A(DB[1822]), .B(DB[1791]), .Z(n5668) );
  AND U9519 ( .A(n284), .B(n5669), .Z(n5667) );
  XOR U9520 ( .A(n5670), .B(n5671), .Z(n5669) );
  XOR U9521 ( .A(DB[1791]), .B(DB[1760]), .Z(n5671) );
  AND U9522 ( .A(n288), .B(n5672), .Z(n5670) );
  XOR U9523 ( .A(n5673), .B(n5674), .Z(n5672) );
  XOR U9524 ( .A(DB[1760]), .B(DB[1729]), .Z(n5674) );
  AND U9525 ( .A(n292), .B(n5675), .Z(n5673) );
  XOR U9526 ( .A(n5676), .B(n5677), .Z(n5675) );
  XOR U9527 ( .A(DB[1729]), .B(DB[1698]), .Z(n5677) );
  AND U9528 ( .A(n296), .B(n5678), .Z(n5676) );
  XOR U9529 ( .A(n5679), .B(n5680), .Z(n5678) );
  XOR U9530 ( .A(DB[1698]), .B(DB[1667]), .Z(n5680) );
  AND U9531 ( .A(n300), .B(n5681), .Z(n5679) );
  XOR U9532 ( .A(n5682), .B(n5683), .Z(n5681) );
  XOR U9533 ( .A(DB[1667]), .B(DB[1636]), .Z(n5683) );
  AND U9534 ( .A(n304), .B(n5684), .Z(n5682) );
  XOR U9535 ( .A(n5685), .B(n5686), .Z(n5684) );
  XOR U9536 ( .A(DB[1636]), .B(DB[1605]), .Z(n5686) );
  AND U9537 ( .A(n308), .B(n5687), .Z(n5685) );
  XOR U9538 ( .A(n5688), .B(n5689), .Z(n5687) );
  XOR U9539 ( .A(DB[1605]), .B(DB[1574]), .Z(n5689) );
  AND U9540 ( .A(n312), .B(n5690), .Z(n5688) );
  XOR U9541 ( .A(n5691), .B(n5692), .Z(n5690) );
  XOR U9542 ( .A(DB[1574]), .B(DB[1543]), .Z(n5692) );
  AND U9543 ( .A(n316), .B(n5693), .Z(n5691) );
  XOR U9544 ( .A(n5694), .B(n5695), .Z(n5693) );
  XOR U9545 ( .A(DB[1543]), .B(DB[1512]), .Z(n5695) );
  AND U9546 ( .A(n320), .B(n5696), .Z(n5694) );
  XOR U9547 ( .A(n5697), .B(n5698), .Z(n5696) );
  XOR U9548 ( .A(DB[1512]), .B(DB[1481]), .Z(n5698) );
  AND U9549 ( .A(n324), .B(n5699), .Z(n5697) );
  XOR U9550 ( .A(n5700), .B(n5701), .Z(n5699) );
  XOR U9551 ( .A(DB[1481]), .B(DB[1450]), .Z(n5701) );
  AND U9552 ( .A(n328), .B(n5702), .Z(n5700) );
  XOR U9553 ( .A(n5703), .B(n5704), .Z(n5702) );
  XOR U9554 ( .A(DB[1450]), .B(DB[1419]), .Z(n5704) );
  AND U9555 ( .A(n332), .B(n5705), .Z(n5703) );
  XOR U9556 ( .A(n5706), .B(n5707), .Z(n5705) );
  XOR U9557 ( .A(DB[1419]), .B(DB[1388]), .Z(n5707) );
  AND U9558 ( .A(n336), .B(n5708), .Z(n5706) );
  XOR U9559 ( .A(n5709), .B(n5710), .Z(n5708) );
  XOR U9560 ( .A(DB[1388]), .B(DB[1357]), .Z(n5710) );
  AND U9561 ( .A(n340), .B(n5711), .Z(n5709) );
  XOR U9562 ( .A(n5712), .B(n5713), .Z(n5711) );
  XOR U9563 ( .A(DB[1357]), .B(DB[1326]), .Z(n5713) );
  AND U9564 ( .A(n344), .B(n5714), .Z(n5712) );
  XOR U9565 ( .A(n5715), .B(n5716), .Z(n5714) );
  XOR U9566 ( .A(DB[1326]), .B(DB[1295]), .Z(n5716) );
  AND U9567 ( .A(n348), .B(n5717), .Z(n5715) );
  XOR U9568 ( .A(n5718), .B(n5719), .Z(n5717) );
  XOR U9569 ( .A(DB[1295]), .B(DB[1264]), .Z(n5719) );
  AND U9570 ( .A(n352), .B(n5720), .Z(n5718) );
  XOR U9571 ( .A(n5721), .B(n5722), .Z(n5720) );
  XOR U9572 ( .A(DB[1264]), .B(DB[1233]), .Z(n5722) );
  AND U9573 ( .A(n356), .B(n5723), .Z(n5721) );
  XOR U9574 ( .A(n5724), .B(n5725), .Z(n5723) );
  XOR U9575 ( .A(DB[1233]), .B(DB[1202]), .Z(n5725) );
  AND U9576 ( .A(n360), .B(n5726), .Z(n5724) );
  XOR U9577 ( .A(n5727), .B(n5728), .Z(n5726) );
  XOR U9578 ( .A(DB[1202]), .B(DB[1171]), .Z(n5728) );
  AND U9579 ( .A(n364), .B(n5729), .Z(n5727) );
  XOR U9580 ( .A(n5730), .B(n5731), .Z(n5729) );
  XOR U9581 ( .A(DB[1171]), .B(DB[1140]), .Z(n5731) );
  AND U9582 ( .A(n368), .B(n5732), .Z(n5730) );
  XOR U9583 ( .A(n5733), .B(n5734), .Z(n5732) );
  XOR U9584 ( .A(DB[1140]), .B(DB[1109]), .Z(n5734) );
  AND U9585 ( .A(n372), .B(n5735), .Z(n5733) );
  XOR U9586 ( .A(n5736), .B(n5737), .Z(n5735) );
  XOR U9587 ( .A(DB[1109]), .B(DB[1078]), .Z(n5737) );
  AND U9588 ( .A(n376), .B(n5738), .Z(n5736) );
  XOR U9589 ( .A(n5739), .B(n5740), .Z(n5738) );
  XOR U9590 ( .A(DB[1078]), .B(DB[1047]), .Z(n5740) );
  AND U9591 ( .A(n380), .B(n5741), .Z(n5739) );
  XOR U9592 ( .A(n5742), .B(n5743), .Z(n5741) );
  XOR U9593 ( .A(DB[1047]), .B(DB[1016]), .Z(n5743) );
  AND U9594 ( .A(n384), .B(n5744), .Z(n5742) );
  XOR U9595 ( .A(n5745), .B(n5746), .Z(n5744) );
  XOR U9596 ( .A(DB[985]), .B(DB[1016]), .Z(n5746) );
  AND U9597 ( .A(n388), .B(n5747), .Z(n5745) );
  XOR U9598 ( .A(n5748), .B(n5749), .Z(n5747) );
  XOR U9599 ( .A(DB[985]), .B(DB[954]), .Z(n5749) );
  AND U9600 ( .A(n392), .B(n5750), .Z(n5748) );
  XOR U9601 ( .A(n5751), .B(n5752), .Z(n5750) );
  XOR U9602 ( .A(DB[954]), .B(DB[923]), .Z(n5752) );
  AND U9603 ( .A(n396), .B(n5753), .Z(n5751) );
  XOR U9604 ( .A(n5754), .B(n5755), .Z(n5753) );
  XOR U9605 ( .A(DB[923]), .B(DB[892]), .Z(n5755) );
  AND U9606 ( .A(n400), .B(n5756), .Z(n5754) );
  XOR U9607 ( .A(n5757), .B(n5758), .Z(n5756) );
  XOR U9608 ( .A(DB[892]), .B(DB[861]), .Z(n5758) );
  AND U9609 ( .A(n404), .B(n5759), .Z(n5757) );
  XOR U9610 ( .A(n5760), .B(n5761), .Z(n5759) );
  XOR U9611 ( .A(DB[861]), .B(DB[830]), .Z(n5761) );
  AND U9612 ( .A(n408), .B(n5762), .Z(n5760) );
  XOR U9613 ( .A(n5763), .B(n5764), .Z(n5762) );
  XOR U9614 ( .A(DB[830]), .B(DB[799]), .Z(n5764) );
  AND U9615 ( .A(n412), .B(n5765), .Z(n5763) );
  XOR U9616 ( .A(n5766), .B(n5767), .Z(n5765) );
  XOR U9617 ( .A(DB[799]), .B(DB[768]), .Z(n5767) );
  AND U9618 ( .A(n416), .B(n5768), .Z(n5766) );
  XOR U9619 ( .A(n5769), .B(n5770), .Z(n5768) );
  XOR U9620 ( .A(DB[768]), .B(DB[737]), .Z(n5770) );
  AND U9621 ( .A(n420), .B(n5771), .Z(n5769) );
  XOR U9622 ( .A(n5772), .B(n5773), .Z(n5771) );
  XOR U9623 ( .A(DB[737]), .B(DB[706]), .Z(n5773) );
  AND U9624 ( .A(n424), .B(n5774), .Z(n5772) );
  XOR U9625 ( .A(n5775), .B(n5776), .Z(n5774) );
  XOR U9626 ( .A(DB[706]), .B(DB[675]), .Z(n5776) );
  AND U9627 ( .A(n428), .B(n5777), .Z(n5775) );
  XOR U9628 ( .A(n5778), .B(n5779), .Z(n5777) );
  XOR U9629 ( .A(DB[675]), .B(DB[644]), .Z(n5779) );
  AND U9630 ( .A(n432), .B(n5780), .Z(n5778) );
  XOR U9631 ( .A(n5781), .B(n5782), .Z(n5780) );
  XOR U9632 ( .A(DB[644]), .B(DB[613]), .Z(n5782) );
  AND U9633 ( .A(n436), .B(n5783), .Z(n5781) );
  XOR U9634 ( .A(n5784), .B(n5785), .Z(n5783) );
  XOR U9635 ( .A(DB[613]), .B(DB[582]), .Z(n5785) );
  AND U9636 ( .A(n440), .B(n5786), .Z(n5784) );
  XOR U9637 ( .A(n5787), .B(n5788), .Z(n5786) );
  XOR U9638 ( .A(DB[582]), .B(DB[551]), .Z(n5788) );
  AND U9639 ( .A(n444), .B(n5789), .Z(n5787) );
  XOR U9640 ( .A(n5790), .B(n5791), .Z(n5789) );
  XOR U9641 ( .A(DB[551]), .B(DB[520]), .Z(n5791) );
  AND U9642 ( .A(n448), .B(n5792), .Z(n5790) );
  XOR U9643 ( .A(n5793), .B(n5794), .Z(n5792) );
  XOR U9644 ( .A(DB[520]), .B(DB[489]), .Z(n5794) );
  AND U9645 ( .A(n452), .B(n5795), .Z(n5793) );
  XOR U9646 ( .A(n5796), .B(n5797), .Z(n5795) );
  XOR U9647 ( .A(DB[489]), .B(DB[458]), .Z(n5797) );
  AND U9648 ( .A(n456), .B(n5798), .Z(n5796) );
  XOR U9649 ( .A(n5799), .B(n5800), .Z(n5798) );
  XOR U9650 ( .A(DB[458]), .B(DB[427]), .Z(n5800) );
  AND U9651 ( .A(n460), .B(n5801), .Z(n5799) );
  XOR U9652 ( .A(n5802), .B(n5803), .Z(n5801) );
  XOR U9653 ( .A(DB[427]), .B(DB[396]), .Z(n5803) );
  AND U9654 ( .A(n464), .B(n5804), .Z(n5802) );
  XOR U9655 ( .A(n5805), .B(n5806), .Z(n5804) );
  XOR U9656 ( .A(DB[396]), .B(DB[365]), .Z(n5806) );
  AND U9657 ( .A(n468), .B(n5807), .Z(n5805) );
  XOR U9658 ( .A(n5808), .B(n5809), .Z(n5807) );
  XOR U9659 ( .A(DB[365]), .B(DB[334]), .Z(n5809) );
  AND U9660 ( .A(n472), .B(n5810), .Z(n5808) );
  XOR U9661 ( .A(n5811), .B(n5812), .Z(n5810) );
  XOR U9662 ( .A(DB[334]), .B(DB[303]), .Z(n5812) );
  AND U9663 ( .A(n476), .B(n5813), .Z(n5811) );
  XOR U9664 ( .A(n5814), .B(n5815), .Z(n5813) );
  XOR U9665 ( .A(DB[303]), .B(DB[272]), .Z(n5815) );
  AND U9666 ( .A(n480), .B(n5816), .Z(n5814) );
  XOR U9667 ( .A(n5817), .B(n5818), .Z(n5816) );
  XOR U9668 ( .A(DB[272]), .B(DB[241]), .Z(n5818) );
  AND U9669 ( .A(n484), .B(n5819), .Z(n5817) );
  XOR U9670 ( .A(n5820), .B(n5821), .Z(n5819) );
  XOR U9671 ( .A(DB[241]), .B(DB[210]), .Z(n5821) );
  AND U9672 ( .A(n488), .B(n5822), .Z(n5820) );
  XOR U9673 ( .A(n5823), .B(n5824), .Z(n5822) );
  XOR U9674 ( .A(DB[210]), .B(DB[179]), .Z(n5824) );
  AND U9675 ( .A(n492), .B(n5825), .Z(n5823) );
  XOR U9676 ( .A(n5826), .B(n5827), .Z(n5825) );
  XOR U9677 ( .A(DB[179]), .B(DB[148]), .Z(n5827) );
  AND U9678 ( .A(n496), .B(n5828), .Z(n5826) );
  XOR U9679 ( .A(n5829), .B(n5830), .Z(n5828) );
  XOR U9680 ( .A(DB[148]), .B(DB[117]), .Z(n5830) );
  AND U9681 ( .A(n500), .B(n5831), .Z(n5829) );
  XOR U9682 ( .A(n5832), .B(n5833), .Z(n5831) );
  XOR U9683 ( .A(DB[86]), .B(DB[117]), .Z(n5833) );
  AND U9684 ( .A(n504), .B(n5834), .Z(n5832) );
  XOR U9685 ( .A(n5835), .B(n5836), .Z(n5834) );
  XOR U9686 ( .A(DB[86]), .B(DB[55]), .Z(n5836) );
  AND U9687 ( .A(n508), .B(n5837), .Z(n5835) );
  XOR U9688 ( .A(DB[55]), .B(DB[24]), .Z(n5837) );
  XOR U9689 ( .A(DB[3960]), .B(n5838), .Z(min_val_out[23]) );
  AND U9690 ( .A(n2), .B(n5839), .Z(n5838) );
  XOR U9691 ( .A(n5840), .B(n5841), .Z(n5839) );
  XOR U9692 ( .A(DB[3960]), .B(DB[3929]), .Z(n5841) );
  AND U9693 ( .A(n8), .B(n5842), .Z(n5840) );
  XOR U9694 ( .A(n5843), .B(n5844), .Z(n5842) );
  XOR U9695 ( .A(DB[3929]), .B(DB[3898]), .Z(n5844) );
  AND U9696 ( .A(n12), .B(n5845), .Z(n5843) );
  XOR U9697 ( .A(n5846), .B(n5847), .Z(n5845) );
  XOR U9698 ( .A(DB[3898]), .B(DB[3867]), .Z(n5847) );
  AND U9699 ( .A(n16), .B(n5848), .Z(n5846) );
  XOR U9700 ( .A(n5849), .B(n5850), .Z(n5848) );
  XOR U9701 ( .A(DB[3867]), .B(DB[3836]), .Z(n5850) );
  AND U9702 ( .A(n20), .B(n5851), .Z(n5849) );
  XOR U9703 ( .A(n5852), .B(n5853), .Z(n5851) );
  XOR U9704 ( .A(DB[3836]), .B(DB[3805]), .Z(n5853) );
  AND U9705 ( .A(n24), .B(n5854), .Z(n5852) );
  XOR U9706 ( .A(n5855), .B(n5856), .Z(n5854) );
  XOR U9707 ( .A(DB[3805]), .B(DB[3774]), .Z(n5856) );
  AND U9708 ( .A(n28), .B(n5857), .Z(n5855) );
  XOR U9709 ( .A(n5858), .B(n5859), .Z(n5857) );
  XOR U9710 ( .A(DB[3774]), .B(DB[3743]), .Z(n5859) );
  AND U9711 ( .A(n32), .B(n5860), .Z(n5858) );
  XOR U9712 ( .A(n5861), .B(n5862), .Z(n5860) );
  XOR U9713 ( .A(DB[3743]), .B(DB[3712]), .Z(n5862) );
  AND U9714 ( .A(n36), .B(n5863), .Z(n5861) );
  XOR U9715 ( .A(n5864), .B(n5865), .Z(n5863) );
  XOR U9716 ( .A(DB[3712]), .B(DB[3681]), .Z(n5865) );
  AND U9717 ( .A(n40), .B(n5866), .Z(n5864) );
  XOR U9718 ( .A(n5867), .B(n5868), .Z(n5866) );
  XOR U9719 ( .A(DB[3681]), .B(DB[3650]), .Z(n5868) );
  AND U9720 ( .A(n44), .B(n5869), .Z(n5867) );
  XOR U9721 ( .A(n5870), .B(n5871), .Z(n5869) );
  XOR U9722 ( .A(DB[3650]), .B(DB[3619]), .Z(n5871) );
  AND U9723 ( .A(n48), .B(n5872), .Z(n5870) );
  XOR U9724 ( .A(n5873), .B(n5874), .Z(n5872) );
  XOR U9725 ( .A(DB[3619]), .B(DB[3588]), .Z(n5874) );
  AND U9726 ( .A(n52), .B(n5875), .Z(n5873) );
  XOR U9727 ( .A(n5876), .B(n5877), .Z(n5875) );
  XOR U9728 ( .A(DB[3588]), .B(DB[3557]), .Z(n5877) );
  AND U9729 ( .A(n56), .B(n5878), .Z(n5876) );
  XOR U9730 ( .A(n5879), .B(n5880), .Z(n5878) );
  XOR U9731 ( .A(DB[3557]), .B(DB[3526]), .Z(n5880) );
  AND U9732 ( .A(n60), .B(n5881), .Z(n5879) );
  XOR U9733 ( .A(n5882), .B(n5883), .Z(n5881) );
  XOR U9734 ( .A(DB[3526]), .B(DB[3495]), .Z(n5883) );
  AND U9735 ( .A(n64), .B(n5884), .Z(n5882) );
  XOR U9736 ( .A(n5885), .B(n5886), .Z(n5884) );
  XOR U9737 ( .A(DB[3495]), .B(DB[3464]), .Z(n5886) );
  AND U9738 ( .A(n68), .B(n5887), .Z(n5885) );
  XOR U9739 ( .A(n5888), .B(n5889), .Z(n5887) );
  XOR U9740 ( .A(DB[3464]), .B(DB[3433]), .Z(n5889) );
  AND U9741 ( .A(n72), .B(n5890), .Z(n5888) );
  XOR U9742 ( .A(n5891), .B(n5892), .Z(n5890) );
  XOR U9743 ( .A(DB[3433]), .B(DB[3402]), .Z(n5892) );
  AND U9744 ( .A(n76), .B(n5893), .Z(n5891) );
  XOR U9745 ( .A(n5894), .B(n5895), .Z(n5893) );
  XOR U9746 ( .A(DB[3402]), .B(DB[3371]), .Z(n5895) );
  AND U9747 ( .A(n80), .B(n5896), .Z(n5894) );
  XOR U9748 ( .A(n5897), .B(n5898), .Z(n5896) );
  XOR U9749 ( .A(DB[3371]), .B(DB[3340]), .Z(n5898) );
  AND U9750 ( .A(n84), .B(n5899), .Z(n5897) );
  XOR U9751 ( .A(n5900), .B(n5901), .Z(n5899) );
  XOR U9752 ( .A(DB[3340]), .B(DB[3309]), .Z(n5901) );
  AND U9753 ( .A(n88), .B(n5902), .Z(n5900) );
  XOR U9754 ( .A(n5903), .B(n5904), .Z(n5902) );
  XOR U9755 ( .A(DB[3309]), .B(DB[3278]), .Z(n5904) );
  AND U9756 ( .A(n92), .B(n5905), .Z(n5903) );
  XOR U9757 ( .A(n5906), .B(n5907), .Z(n5905) );
  XOR U9758 ( .A(DB[3278]), .B(DB[3247]), .Z(n5907) );
  AND U9759 ( .A(n96), .B(n5908), .Z(n5906) );
  XOR U9760 ( .A(n5909), .B(n5910), .Z(n5908) );
  XOR U9761 ( .A(DB[3247]), .B(DB[3216]), .Z(n5910) );
  AND U9762 ( .A(n100), .B(n5911), .Z(n5909) );
  XOR U9763 ( .A(n5912), .B(n5913), .Z(n5911) );
  XOR U9764 ( .A(DB[3216]), .B(DB[3185]), .Z(n5913) );
  AND U9765 ( .A(n104), .B(n5914), .Z(n5912) );
  XOR U9766 ( .A(n5915), .B(n5916), .Z(n5914) );
  XOR U9767 ( .A(DB[3185]), .B(DB[3154]), .Z(n5916) );
  AND U9768 ( .A(n108), .B(n5917), .Z(n5915) );
  XOR U9769 ( .A(n5918), .B(n5919), .Z(n5917) );
  XOR U9770 ( .A(DB[3154]), .B(DB[3123]), .Z(n5919) );
  AND U9771 ( .A(n112), .B(n5920), .Z(n5918) );
  XOR U9772 ( .A(n5921), .B(n5922), .Z(n5920) );
  XOR U9773 ( .A(DB[3123]), .B(DB[3092]), .Z(n5922) );
  AND U9774 ( .A(n116), .B(n5923), .Z(n5921) );
  XOR U9775 ( .A(n5924), .B(n5925), .Z(n5923) );
  XOR U9776 ( .A(DB[3092]), .B(DB[3061]), .Z(n5925) );
  AND U9777 ( .A(n120), .B(n5926), .Z(n5924) );
  XOR U9778 ( .A(n5927), .B(n5928), .Z(n5926) );
  XOR U9779 ( .A(DB[3061]), .B(DB[3030]), .Z(n5928) );
  AND U9780 ( .A(n124), .B(n5929), .Z(n5927) );
  XOR U9781 ( .A(n5930), .B(n5931), .Z(n5929) );
  XOR U9782 ( .A(DB[3030]), .B(DB[2999]), .Z(n5931) );
  AND U9783 ( .A(n128), .B(n5932), .Z(n5930) );
  XOR U9784 ( .A(n5933), .B(n5934), .Z(n5932) );
  XOR U9785 ( .A(DB[2999]), .B(DB[2968]), .Z(n5934) );
  AND U9786 ( .A(n132), .B(n5935), .Z(n5933) );
  XOR U9787 ( .A(n5936), .B(n5937), .Z(n5935) );
  XOR U9788 ( .A(DB[2968]), .B(DB[2937]), .Z(n5937) );
  AND U9789 ( .A(n136), .B(n5938), .Z(n5936) );
  XOR U9790 ( .A(n5939), .B(n5940), .Z(n5938) );
  XOR U9791 ( .A(DB[2937]), .B(DB[2906]), .Z(n5940) );
  AND U9792 ( .A(n140), .B(n5941), .Z(n5939) );
  XOR U9793 ( .A(n5942), .B(n5943), .Z(n5941) );
  XOR U9794 ( .A(DB[2906]), .B(DB[2875]), .Z(n5943) );
  AND U9795 ( .A(n144), .B(n5944), .Z(n5942) );
  XOR U9796 ( .A(n5945), .B(n5946), .Z(n5944) );
  XOR U9797 ( .A(DB[2875]), .B(DB[2844]), .Z(n5946) );
  AND U9798 ( .A(n148), .B(n5947), .Z(n5945) );
  XOR U9799 ( .A(n5948), .B(n5949), .Z(n5947) );
  XOR U9800 ( .A(DB[2844]), .B(DB[2813]), .Z(n5949) );
  AND U9801 ( .A(n152), .B(n5950), .Z(n5948) );
  XOR U9802 ( .A(n5951), .B(n5952), .Z(n5950) );
  XOR U9803 ( .A(DB[2813]), .B(DB[2782]), .Z(n5952) );
  AND U9804 ( .A(n156), .B(n5953), .Z(n5951) );
  XOR U9805 ( .A(n5954), .B(n5955), .Z(n5953) );
  XOR U9806 ( .A(DB[2782]), .B(DB[2751]), .Z(n5955) );
  AND U9807 ( .A(n160), .B(n5956), .Z(n5954) );
  XOR U9808 ( .A(n5957), .B(n5958), .Z(n5956) );
  XOR U9809 ( .A(DB[2751]), .B(DB[2720]), .Z(n5958) );
  AND U9810 ( .A(n164), .B(n5959), .Z(n5957) );
  XOR U9811 ( .A(n5960), .B(n5961), .Z(n5959) );
  XOR U9812 ( .A(DB[2720]), .B(DB[2689]), .Z(n5961) );
  AND U9813 ( .A(n168), .B(n5962), .Z(n5960) );
  XOR U9814 ( .A(n5963), .B(n5964), .Z(n5962) );
  XOR U9815 ( .A(DB[2689]), .B(DB[2658]), .Z(n5964) );
  AND U9816 ( .A(n172), .B(n5965), .Z(n5963) );
  XOR U9817 ( .A(n5966), .B(n5967), .Z(n5965) );
  XOR U9818 ( .A(DB[2658]), .B(DB[2627]), .Z(n5967) );
  AND U9819 ( .A(n176), .B(n5968), .Z(n5966) );
  XOR U9820 ( .A(n5969), .B(n5970), .Z(n5968) );
  XOR U9821 ( .A(DB[2627]), .B(DB[2596]), .Z(n5970) );
  AND U9822 ( .A(n180), .B(n5971), .Z(n5969) );
  XOR U9823 ( .A(n5972), .B(n5973), .Z(n5971) );
  XOR U9824 ( .A(DB[2596]), .B(DB[2565]), .Z(n5973) );
  AND U9825 ( .A(n184), .B(n5974), .Z(n5972) );
  XOR U9826 ( .A(n5975), .B(n5976), .Z(n5974) );
  XOR U9827 ( .A(DB[2565]), .B(DB[2534]), .Z(n5976) );
  AND U9828 ( .A(n188), .B(n5977), .Z(n5975) );
  XOR U9829 ( .A(n5978), .B(n5979), .Z(n5977) );
  XOR U9830 ( .A(DB[2534]), .B(DB[2503]), .Z(n5979) );
  AND U9831 ( .A(n192), .B(n5980), .Z(n5978) );
  XOR U9832 ( .A(n5981), .B(n5982), .Z(n5980) );
  XOR U9833 ( .A(DB[2503]), .B(DB[2472]), .Z(n5982) );
  AND U9834 ( .A(n196), .B(n5983), .Z(n5981) );
  XOR U9835 ( .A(n5984), .B(n5985), .Z(n5983) );
  XOR U9836 ( .A(DB[2472]), .B(DB[2441]), .Z(n5985) );
  AND U9837 ( .A(n200), .B(n5986), .Z(n5984) );
  XOR U9838 ( .A(n5987), .B(n5988), .Z(n5986) );
  XOR U9839 ( .A(DB[2441]), .B(DB[2410]), .Z(n5988) );
  AND U9840 ( .A(n204), .B(n5989), .Z(n5987) );
  XOR U9841 ( .A(n5990), .B(n5991), .Z(n5989) );
  XOR U9842 ( .A(DB[2410]), .B(DB[2379]), .Z(n5991) );
  AND U9843 ( .A(n208), .B(n5992), .Z(n5990) );
  XOR U9844 ( .A(n5993), .B(n5994), .Z(n5992) );
  XOR U9845 ( .A(DB[2379]), .B(DB[2348]), .Z(n5994) );
  AND U9846 ( .A(n212), .B(n5995), .Z(n5993) );
  XOR U9847 ( .A(n5996), .B(n5997), .Z(n5995) );
  XOR U9848 ( .A(DB[2348]), .B(DB[2317]), .Z(n5997) );
  AND U9849 ( .A(n216), .B(n5998), .Z(n5996) );
  XOR U9850 ( .A(n5999), .B(n6000), .Z(n5998) );
  XOR U9851 ( .A(DB[2317]), .B(DB[2286]), .Z(n6000) );
  AND U9852 ( .A(n220), .B(n6001), .Z(n5999) );
  XOR U9853 ( .A(n6002), .B(n6003), .Z(n6001) );
  XOR U9854 ( .A(DB[2286]), .B(DB[2255]), .Z(n6003) );
  AND U9855 ( .A(n224), .B(n6004), .Z(n6002) );
  XOR U9856 ( .A(n6005), .B(n6006), .Z(n6004) );
  XOR U9857 ( .A(DB[2255]), .B(DB[2224]), .Z(n6006) );
  AND U9858 ( .A(n228), .B(n6007), .Z(n6005) );
  XOR U9859 ( .A(n6008), .B(n6009), .Z(n6007) );
  XOR U9860 ( .A(DB[2224]), .B(DB[2193]), .Z(n6009) );
  AND U9861 ( .A(n232), .B(n6010), .Z(n6008) );
  XOR U9862 ( .A(n6011), .B(n6012), .Z(n6010) );
  XOR U9863 ( .A(DB[2193]), .B(DB[2162]), .Z(n6012) );
  AND U9864 ( .A(n236), .B(n6013), .Z(n6011) );
  XOR U9865 ( .A(n6014), .B(n6015), .Z(n6013) );
  XOR U9866 ( .A(DB[2162]), .B(DB[2131]), .Z(n6015) );
  AND U9867 ( .A(n240), .B(n6016), .Z(n6014) );
  XOR U9868 ( .A(n6017), .B(n6018), .Z(n6016) );
  XOR U9869 ( .A(DB[2131]), .B(DB[2100]), .Z(n6018) );
  AND U9870 ( .A(n244), .B(n6019), .Z(n6017) );
  XOR U9871 ( .A(n6020), .B(n6021), .Z(n6019) );
  XOR U9872 ( .A(DB[2100]), .B(DB[2069]), .Z(n6021) );
  AND U9873 ( .A(n248), .B(n6022), .Z(n6020) );
  XOR U9874 ( .A(n6023), .B(n6024), .Z(n6022) );
  XOR U9875 ( .A(DB[2069]), .B(DB[2038]), .Z(n6024) );
  AND U9876 ( .A(n252), .B(n6025), .Z(n6023) );
  XOR U9877 ( .A(n6026), .B(n6027), .Z(n6025) );
  XOR U9878 ( .A(DB[2038]), .B(DB[2007]), .Z(n6027) );
  AND U9879 ( .A(n256), .B(n6028), .Z(n6026) );
  XOR U9880 ( .A(n6029), .B(n6030), .Z(n6028) );
  XOR U9881 ( .A(DB[2007]), .B(DB[1976]), .Z(n6030) );
  AND U9882 ( .A(n260), .B(n6031), .Z(n6029) );
  XOR U9883 ( .A(n6032), .B(n6033), .Z(n6031) );
  XOR U9884 ( .A(DB[1976]), .B(DB[1945]), .Z(n6033) );
  AND U9885 ( .A(n264), .B(n6034), .Z(n6032) );
  XOR U9886 ( .A(n6035), .B(n6036), .Z(n6034) );
  XOR U9887 ( .A(DB[1945]), .B(DB[1914]), .Z(n6036) );
  AND U9888 ( .A(n268), .B(n6037), .Z(n6035) );
  XOR U9889 ( .A(n6038), .B(n6039), .Z(n6037) );
  XOR U9890 ( .A(DB[1914]), .B(DB[1883]), .Z(n6039) );
  AND U9891 ( .A(n272), .B(n6040), .Z(n6038) );
  XOR U9892 ( .A(n6041), .B(n6042), .Z(n6040) );
  XOR U9893 ( .A(DB[1883]), .B(DB[1852]), .Z(n6042) );
  AND U9894 ( .A(n276), .B(n6043), .Z(n6041) );
  XOR U9895 ( .A(n6044), .B(n6045), .Z(n6043) );
  XOR U9896 ( .A(DB[1852]), .B(DB[1821]), .Z(n6045) );
  AND U9897 ( .A(n280), .B(n6046), .Z(n6044) );
  XOR U9898 ( .A(n6047), .B(n6048), .Z(n6046) );
  XOR U9899 ( .A(DB[1821]), .B(DB[1790]), .Z(n6048) );
  AND U9900 ( .A(n284), .B(n6049), .Z(n6047) );
  XOR U9901 ( .A(n6050), .B(n6051), .Z(n6049) );
  XOR U9902 ( .A(DB[1790]), .B(DB[1759]), .Z(n6051) );
  AND U9903 ( .A(n288), .B(n6052), .Z(n6050) );
  XOR U9904 ( .A(n6053), .B(n6054), .Z(n6052) );
  XOR U9905 ( .A(DB[1759]), .B(DB[1728]), .Z(n6054) );
  AND U9906 ( .A(n292), .B(n6055), .Z(n6053) );
  XOR U9907 ( .A(n6056), .B(n6057), .Z(n6055) );
  XOR U9908 ( .A(DB[1728]), .B(DB[1697]), .Z(n6057) );
  AND U9909 ( .A(n296), .B(n6058), .Z(n6056) );
  XOR U9910 ( .A(n6059), .B(n6060), .Z(n6058) );
  XOR U9911 ( .A(DB[1697]), .B(DB[1666]), .Z(n6060) );
  AND U9912 ( .A(n300), .B(n6061), .Z(n6059) );
  XOR U9913 ( .A(n6062), .B(n6063), .Z(n6061) );
  XOR U9914 ( .A(DB[1666]), .B(DB[1635]), .Z(n6063) );
  AND U9915 ( .A(n304), .B(n6064), .Z(n6062) );
  XOR U9916 ( .A(n6065), .B(n6066), .Z(n6064) );
  XOR U9917 ( .A(DB[1635]), .B(DB[1604]), .Z(n6066) );
  AND U9918 ( .A(n308), .B(n6067), .Z(n6065) );
  XOR U9919 ( .A(n6068), .B(n6069), .Z(n6067) );
  XOR U9920 ( .A(DB[1604]), .B(DB[1573]), .Z(n6069) );
  AND U9921 ( .A(n312), .B(n6070), .Z(n6068) );
  XOR U9922 ( .A(n6071), .B(n6072), .Z(n6070) );
  XOR U9923 ( .A(DB[1573]), .B(DB[1542]), .Z(n6072) );
  AND U9924 ( .A(n316), .B(n6073), .Z(n6071) );
  XOR U9925 ( .A(n6074), .B(n6075), .Z(n6073) );
  XOR U9926 ( .A(DB[1542]), .B(DB[1511]), .Z(n6075) );
  AND U9927 ( .A(n320), .B(n6076), .Z(n6074) );
  XOR U9928 ( .A(n6077), .B(n6078), .Z(n6076) );
  XOR U9929 ( .A(DB[1511]), .B(DB[1480]), .Z(n6078) );
  AND U9930 ( .A(n324), .B(n6079), .Z(n6077) );
  XOR U9931 ( .A(n6080), .B(n6081), .Z(n6079) );
  XOR U9932 ( .A(DB[1480]), .B(DB[1449]), .Z(n6081) );
  AND U9933 ( .A(n328), .B(n6082), .Z(n6080) );
  XOR U9934 ( .A(n6083), .B(n6084), .Z(n6082) );
  XOR U9935 ( .A(DB[1449]), .B(DB[1418]), .Z(n6084) );
  AND U9936 ( .A(n332), .B(n6085), .Z(n6083) );
  XOR U9937 ( .A(n6086), .B(n6087), .Z(n6085) );
  XOR U9938 ( .A(DB[1418]), .B(DB[1387]), .Z(n6087) );
  AND U9939 ( .A(n336), .B(n6088), .Z(n6086) );
  XOR U9940 ( .A(n6089), .B(n6090), .Z(n6088) );
  XOR U9941 ( .A(DB[1387]), .B(DB[1356]), .Z(n6090) );
  AND U9942 ( .A(n340), .B(n6091), .Z(n6089) );
  XOR U9943 ( .A(n6092), .B(n6093), .Z(n6091) );
  XOR U9944 ( .A(DB[1356]), .B(DB[1325]), .Z(n6093) );
  AND U9945 ( .A(n344), .B(n6094), .Z(n6092) );
  XOR U9946 ( .A(n6095), .B(n6096), .Z(n6094) );
  XOR U9947 ( .A(DB[1325]), .B(DB[1294]), .Z(n6096) );
  AND U9948 ( .A(n348), .B(n6097), .Z(n6095) );
  XOR U9949 ( .A(n6098), .B(n6099), .Z(n6097) );
  XOR U9950 ( .A(DB[1294]), .B(DB[1263]), .Z(n6099) );
  AND U9951 ( .A(n352), .B(n6100), .Z(n6098) );
  XOR U9952 ( .A(n6101), .B(n6102), .Z(n6100) );
  XOR U9953 ( .A(DB[1263]), .B(DB[1232]), .Z(n6102) );
  AND U9954 ( .A(n356), .B(n6103), .Z(n6101) );
  XOR U9955 ( .A(n6104), .B(n6105), .Z(n6103) );
  XOR U9956 ( .A(DB[1232]), .B(DB[1201]), .Z(n6105) );
  AND U9957 ( .A(n360), .B(n6106), .Z(n6104) );
  XOR U9958 ( .A(n6107), .B(n6108), .Z(n6106) );
  XOR U9959 ( .A(DB[1201]), .B(DB[1170]), .Z(n6108) );
  AND U9960 ( .A(n364), .B(n6109), .Z(n6107) );
  XOR U9961 ( .A(n6110), .B(n6111), .Z(n6109) );
  XOR U9962 ( .A(DB[1170]), .B(DB[1139]), .Z(n6111) );
  AND U9963 ( .A(n368), .B(n6112), .Z(n6110) );
  XOR U9964 ( .A(n6113), .B(n6114), .Z(n6112) );
  XOR U9965 ( .A(DB[1139]), .B(DB[1108]), .Z(n6114) );
  AND U9966 ( .A(n372), .B(n6115), .Z(n6113) );
  XOR U9967 ( .A(n6116), .B(n6117), .Z(n6115) );
  XOR U9968 ( .A(DB[1108]), .B(DB[1077]), .Z(n6117) );
  AND U9969 ( .A(n376), .B(n6118), .Z(n6116) );
  XOR U9970 ( .A(n6119), .B(n6120), .Z(n6118) );
  XOR U9971 ( .A(DB[1077]), .B(DB[1046]), .Z(n6120) );
  AND U9972 ( .A(n380), .B(n6121), .Z(n6119) );
  XOR U9973 ( .A(n6122), .B(n6123), .Z(n6121) );
  XOR U9974 ( .A(DB[1046]), .B(DB[1015]), .Z(n6123) );
  AND U9975 ( .A(n384), .B(n6124), .Z(n6122) );
  XOR U9976 ( .A(n6125), .B(n6126), .Z(n6124) );
  XOR U9977 ( .A(DB[984]), .B(DB[1015]), .Z(n6126) );
  AND U9978 ( .A(n388), .B(n6127), .Z(n6125) );
  XOR U9979 ( .A(n6128), .B(n6129), .Z(n6127) );
  XOR U9980 ( .A(DB[984]), .B(DB[953]), .Z(n6129) );
  AND U9981 ( .A(n392), .B(n6130), .Z(n6128) );
  XOR U9982 ( .A(n6131), .B(n6132), .Z(n6130) );
  XOR U9983 ( .A(DB[953]), .B(DB[922]), .Z(n6132) );
  AND U9984 ( .A(n396), .B(n6133), .Z(n6131) );
  XOR U9985 ( .A(n6134), .B(n6135), .Z(n6133) );
  XOR U9986 ( .A(DB[922]), .B(DB[891]), .Z(n6135) );
  AND U9987 ( .A(n400), .B(n6136), .Z(n6134) );
  XOR U9988 ( .A(n6137), .B(n6138), .Z(n6136) );
  XOR U9989 ( .A(DB[891]), .B(DB[860]), .Z(n6138) );
  AND U9990 ( .A(n404), .B(n6139), .Z(n6137) );
  XOR U9991 ( .A(n6140), .B(n6141), .Z(n6139) );
  XOR U9992 ( .A(DB[860]), .B(DB[829]), .Z(n6141) );
  AND U9993 ( .A(n408), .B(n6142), .Z(n6140) );
  XOR U9994 ( .A(n6143), .B(n6144), .Z(n6142) );
  XOR U9995 ( .A(DB[829]), .B(DB[798]), .Z(n6144) );
  AND U9996 ( .A(n412), .B(n6145), .Z(n6143) );
  XOR U9997 ( .A(n6146), .B(n6147), .Z(n6145) );
  XOR U9998 ( .A(DB[798]), .B(DB[767]), .Z(n6147) );
  AND U9999 ( .A(n416), .B(n6148), .Z(n6146) );
  XOR U10000 ( .A(n6149), .B(n6150), .Z(n6148) );
  XOR U10001 ( .A(DB[767]), .B(DB[736]), .Z(n6150) );
  AND U10002 ( .A(n420), .B(n6151), .Z(n6149) );
  XOR U10003 ( .A(n6152), .B(n6153), .Z(n6151) );
  XOR U10004 ( .A(DB[736]), .B(DB[705]), .Z(n6153) );
  AND U10005 ( .A(n424), .B(n6154), .Z(n6152) );
  XOR U10006 ( .A(n6155), .B(n6156), .Z(n6154) );
  XOR U10007 ( .A(DB[705]), .B(DB[674]), .Z(n6156) );
  AND U10008 ( .A(n428), .B(n6157), .Z(n6155) );
  XOR U10009 ( .A(n6158), .B(n6159), .Z(n6157) );
  XOR U10010 ( .A(DB[674]), .B(DB[643]), .Z(n6159) );
  AND U10011 ( .A(n432), .B(n6160), .Z(n6158) );
  XOR U10012 ( .A(n6161), .B(n6162), .Z(n6160) );
  XOR U10013 ( .A(DB[643]), .B(DB[612]), .Z(n6162) );
  AND U10014 ( .A(n436), .B(n6163), .Z(n6161) );
  XOR U10015 ( .A(n6164), .B(n6165), .Z(n6163) );
  XOR U10016 ( .A(DB[612]), .B(DB[581]), .Z(n6165) );
  AND U10017 ( .A(n440), .B(n6166), .Z(n6164) );
  XOR U10018 ( .A(n6167), .B(n6168), .Z(n6166) );
  XOR U10019 ( .A(DB[581]), .B(DB[550]), .Z(n6168) );
  AND U10020 ( .A(n444), .B(n6169), .Z(n6167) );
  XOR U10021 ( .A(n6170), .B(n6171), .Z(n6169) );
  XOR U10022 ( .A(DB[550]), .B(DB[519]), .Z(n6171) );
  AND U10023 ( .A(n448), .B(n6172), .Z(n6170) );
  XOR U10024 ( .A(n6173), .B(n6174), .Z(n6172) );
  XOR U10025 ( .A(DB[519]), .B(DB[488]), .Z(n6174) );
  AND U10026 ( .A(n452), .B(n6175), .Z(n6173) );
  XOR U10027 ( .A(n6176), .B(n6177), .Z(n6175) );
  XOR U10028 ( .A(DB[488]), .B(DB[457]), .Z(n6177) );
  AND U10029 ( .A(n456), .B(n6178), .Z(n6176) );
  XOR U10030 ( .A(n6179), .B(n6180), .Z(n6178) );
  XOR U10031 ( .A(DB[457]), .B(DB[426]), .Z(n6180) );
  AND U10032 ( .A(n460), .B(n6181), .Z(n6179) );
  XOR U10033 ( .A(n6182), .B(n6183), .Z(n6181) );
  XOR U10034 ( .A(DB[426]), .B(DB[395]), .Z(n6183) );
  AND U10035 ( .A(n464), .B(n6184), .Z(n6182) );
  XOR U10036 ( .A(n6185), .B(n6186), .Z(n6184) );
  XOR U10037 ( .A(DB[395]), .B(DB[364]), .Z(n6186) );
  AND U10038 ( .A(n468), .B(n6187), .Z(n6185) );
  XOR U10039 ( .A(n6188), .B(n6189), .Z(n6187) );
  XOR U10040 ( .A(DB[364]), .B(DB[333]), .Z(n6189) );
  AND U10041 ( .A(n472), .B(n6190), .Z(n6188) );
  XOR U10042 ( .A(n6191), .B(n6192), .Z(n6190) );
  XOR U10043 ( .A(DB[333]), .B(DB[302]), .Z(n6192) );
  AND U10044 ( .A(n476), .B(n6193), .Z(n6191) );
  XOR U10045 ( .A(n6194), .B(n6195), .Z(n6193) );
  XOR U10046 ( .A(DB[302]), .B(DB[271]), .Z(n6195) );
  AND U10047 ( .A(n480), .B(n6196), .Z(n6194) );
  XOR U10048 ( .A(n6197), .B(n6198), .Z(n6196) );
  XOR U10049 ( .A(DB[271]), .B(DB[240]), .Z(n6198) );
  AND U10050 ( .A(n484), .B(n6199), .Z(n6197) );
  XOR U10051 ( .A(n6200), .B(n6201), .Z(n6199) );
  XOR U10052 ( .A(DB[240]), .B(DB[209]), .Z(n6201) );
  AND U10053 ( .A(n488), .B(n6202), .Z(n6200) );
  XOR U10054 ( .A(n6203), .B(n6204), .Z(n6202) );
  XOR U10055 ( .A(DB[209]), .B(DB[178]), .Z(n6204) );
  AND U10056 ( .A(n492), .B(n6205), .Z(n6203) );
  XOR U10057 ( .A(n6206), .B(n6207), .Z(n6205) );
  XOR U10058 ( .A(DB[178]), .B(DB[147]), .Z(n6207) );
  AND U10059 ( .A(n496), .B(n6208), .Z(n6206) );
  XOR U10060 ( .A(n6209), .B(n6210), .Z(n6208) );
  XOR U10061 ( .A(DB[147]), .B(DB[116]), .Z(n6210) );
  AND U10062 ( .A(n500), .B(n6211), .Z(n6209) );
  XOR U10063 ( .A(n6212), .B(n6213), .Z(n6211) );
  XOR U10064 ( .A(DB[85]), .B(DB[116]), .Z(n6213) );
  AND U10065 ( .A(n504), .B(n6214), .Z(n6212) );
  XOR U10066 ( .A(n6215), .B(n6216), .Z(n6214) );
  XOR U10067 ( .A(DB[85]), .B(DB[54]), .Z(n6216) );
  AND U10068 ( .A(n508), .B(n6217), .Z(n6215) );
  XOR U10069 ( .A(DB[54]), .B(DB[23]), .Z(n6217) );
  XOR U10070 ( .A(DB[3959]), .B(n6218), .Z(min_val_out[22]) );
  AND U10071 ( .A(n2), .B(n6219), .Z(n6218) );
  XOR U10072 ( .A(n6220), .B(n6221), .Z(n6219) );
  XOR U10073 ( .A(DB[3959]), .B(DB[3928]), .Z(n6221) );
  AND U10074 ( .A(n8), .B(n6222), .Z(n6220) );
  XOR U10075 ( .A(n6223), .B(n6224), .Z(n6222) );
  XOR U10076 ( .A(DB[3928]), .B(DB[3897]), .Z(n6224) );
  AND U10077 ( .A(n12), .B(n6225), .Z(n6223) );
  XOR U10078 ( .A(n6226), .B(n6227), .Z(n6225) );
  XOR U10079 ( .A(DB[3897]), .B(DB[3866]), .Z(n6227) );
  AND U10080 ( .A(n16), .B(n6228), .Z(n6226) );
  XOR U10081 ( .A(n6229), .B(n6230), .Z(n6228) );
  XOR U10082 ( .A(DB[3866]), .B(DB[3835]), .Z(n6230) );
  AND U10083 ( .A(n20), .B(n6231), .Z(n6229) );
  XOR U10084 ( .A(n6232), .B(n6233), .Z(n6231) );
  XOR U10085 ( .A(DB[3835]), .B(DB[3804]), .Z(n6233) );
  AND U10086 ( .A(n24), .B(n6234), .Z(n6232) );
  XOR U10087 ( .A(n6235), .B(n6236), .Z(n6234) );
  XOR U10088 ( .A(DB[3804]), .B(DB[3773]), .Z(n6236) );
  AND U10089 ( .A(n28), .B(n6237), .Z(n6235) );
  XOR U10090 ( .A(n6238), .B(n6239), .Z(n6237) );
  XOR U10091 ( .A(DB[3773]), .B(DB[3742]), .Z(n6239) );
  AND U10092 ( .A(n32), .B(n6240), .Z(n6238) );
  XOR U10093 ( .A(n6241), .B(n6242), .Z(n6240) );
  XOR U10094 ( .A(DB[3742]), .B(DB[3711]), .Z(n6242) );
  AND U10095 ( .A(n36), .B(n6243), .Z(n6241) );
  XOR U10096 ( .A(n6244), .B(n6245), .Z(n6243) );
  XOR U10097 ( .A(DB[3711]), .B(DB[3680]), .Z(n6245) );
  AND U10098 ( .A(n40), .B(n6246), .Z(n6244) );
  XOR U10099 ( .A(n6247), .B(n6248), .Z(n6246) );
  XOR U10100 ( .A(DB[3680]), .B(DB[3649]), .Z(n6248) );
  AND U10101 ( .A(n44), .B(n6249), .Z(n6247) );
  XOR U10102 ( .A(n6250), .B(n6251), .Z(n6249) );
  XOR U10103 ( .A(DB[3649]), .B(DB[3618]), .Z(n6251) );
  AND U10104 ( .A(n48), .B(n6252), .Z(n6250) );
  XOR U10105 ( .A(n6253), .B(n6254), .Z(n6252) );
  XOR U10106 ( .A(DB[3618]), .B(DB[3587]), .Z(n6254) );
  AND U10107 ( .A(n52), .B(n6255), .Z(n6253) );
  XOR U10108 ( .A(n6256), .B(n6257), .Z(n6255) );
  XOR U10109 ( .A(DB[3587]), .B(DB[3556]), .Z(n6257) );
  AND U10110 ( .A(n56), .B(n6258), .Z(n6256) );
  XOR U10111 ( .A(n6259), .B(n6260), .Z(n6258) );
  XOR U10112 ( .A(DB[3556]), .B(DB[3525]), .Z(n6260) );
  AND U10113 ( .A(n60), .B(n6261), .Z(n6259) );
  XOR U10114 ( .A(n6262), .B(n6263), .Z(n6261) );
  XOR U10115 ( .A(DB[3525]), .B(DB[3494]), .Z(n6263) );
  AND U10116 ( .A(n64), .B(n6264), .Z(n6262) );
  XOR U10117 ( .A(n6265), .B(n6266), .Z(n6264) );
  XOR U10118 ( .A(DB[3494]), .B(DB[3463]), .Z(n6266) );
  AND U10119 ( .A(n68), .B(n6267), .Z(n6265) );
  XOR U10120 ( .A(n6268), .B(n6269), .Z(n6267) );
  XOR U10121 ( .A(DB[3463]), .B(DB[3432]), .Z(n6269) );
  AND U10122 ( .A(n72), .B(n6270), .Z(n6268) );
  XOR U10123 ( .A(n6271), .B(n6272), .Z(n6270) );
  XOR U10124 ( .A(DB[3432]), .B(DB[3401]), .Z(n6272) );
  AND U10125 ( .A(n76), .B(n6273), .Z(n6271) );
  XOR U10126 ( .A(n6274), .B(n6275), .Z(n6273) );
  XOR U10127 ( .A(DB[3401]), .B(DB[3370]), .Z(n6275) );
  AND U10128 ( .A(n80), .B(n6276), .Z(n6274) );
  XOR U10129 ( .A(n6277), .B(n6278), .Z(n6276) );
  XOR U10130 ( .A(DB[3370]), .B(DB[3339]), .Z(n6278) );
  AND U10131 ( .A(n84), .B(n6279), .Z(n6277) );
  XOR U10132 ( .A(n6280), .B(n6281), .Z(n6279) );
  XOR U10133 ( .A(DB[3339]), .B(DB[3308]), .Z(n6281) );
  AND U10134 ( .A(n88), .B(n6282), .Z(n6280) );
  XOR U10135 ( .A(n6283), .B(n6284), .Z(n6282) );
  XOR U10136 ( .A(DB[3308]), .B(DB[3277]), .Z(n6284) );
  AND U10137 ( .A(n92), .B(n6285), .Z(n6283) );
  XOR U10138 ( .A(n6286), .B(n6287), .Z(n6285) );
  XOR U10139 ( .A(DB[3277]), .B(DB[3246]), .Z(n6287) );
  AND U10140 ( .A(n96), .B(n6288), .Z(n6286) );
  XOR U10141 ( .A(n6289), .B(n6290), .Z(n6288) );
  XOR U10142 ( .A(DB[3246]), .B(DB[3215]), .Z(n6290) );
  AND U10143 ( .A(n100), .B(n6291), .Z(n6289) );
  XOR U10144 ( .A(n6292), .B(n6293), .Z(n6291) );
  XOR U10145 ( .A(DB[3215]), .B(DB[3184]), .Z(n6293) );
  AND U10146 ( .A(n104), .B(n6294), .Z(n6292) );
  XOR U10147 ( .A(n6295), .B(n6296), .Z(n6294) );
  XOR U10148 ( .A(DB[3184]), .B(DB[3153]), .Z(n6296) );
  AND U10149 ( .A(n108), .B(n6297), .Z(n6295) );
  XOR U10150 ( .A(n6298), .B(n6299), .Z(n6297) );
  XOR U10151 ( .A(DB[3153]), .B(DB[3122]), .Z(n6299) );
  AND U10152 ( .A(n112), .B(n6300), .Z(n6298) );
  XOR U10153 ( .A(n6301), .B(n6302), .Z(n6300) );
  XOR U10154 ( .A(DB[3122]), .B(DB[3091]), .Z(n6302) );
  AND U10155 ( .A(n116), .B(n6303), .Z(n6301) );
  XOR U10156 ( .A(n6304), .B(n6305), .Z(n6303) );
  XOR U10157 ( .A(DB[3091]), .B(DB[3060]), .Z(n6305) );
  AND U10158 ( .A(n120), .B(n6306), .Z(n6304) );
  XOR U10159 ( .A(n6307), .B(n6308), .Z(n6306) );
  XOR U10160 ( .A(DB[3060]), .B(DB[3029]), .Z(n6308) );
  AND U10161 ( .A(n124), .B(n6309), .Z(n6307) );
  XOR U10162 ( .A(n6310), .B(n6311), .Z(n6309) );
  XOR U10163 ( .A(DB[3029]), .B(DB[2998]), .Z(n6311) );
  AND U10164 ( .A(n128), .B(n6312), .Z(n6310) );
  XOR U10165 ( .A(n6313), .B(n6314), .Z(n6312) );
  XOR U10166 ( .A(DB[2998]), .B(DB[2967]), .Z(n6314) );
  AND U10167 ( .A(n132), .B(n6315), .Z(n6313) );
  XOR U10168 ( .A(n6316), .B(n6317), .Z(n6315) );
  XOR U10169 ( .A(DB[2967]), .B(DB[2936]), .Z(n6317) );
  AND U10170 ( .A(n136), .B(n6318), .Z(n6316) );
  XOR U10171 ( .A(n6319), .B(n6320), .Z(n6318) );
  XOR U10172 ( .A(DB[2936]), .B(DB[2905]), .Z(n6320) );
  AND U10173 ( .A(n140), .B(n6321), .Z(n6319) );
  XOR U10174 ( .A(n6322), .B(n6323), .Z(n6321) );
  XOR U10175 ( .A(DB[2905]), .B(DB[2874]), .Z(n6323) );
  AND U10176 ( .A(n144), .B(n6324), .Z(n6322) );
  XOR U10177 ( .A(n6325), .B(n6326), .Z(n6324) );
  XOR U10178 ( .A(DB[2874]), .B(DB[2843]), .Z(n6326) );
  AND U10179 ( .A(n148), .B(n6327), .Z(n6325) );
  XOR U10180 ( .A(n6328), .B(n6329), .Z(n6327) );
  XOR U10181 ( .A(DB[2843]), .B(DB[2812]), .Z(n6329) );
  AND U10182 ( .A(n152), .B(n6330), .Z(n6328) );
  XOR U10183 ( .A(n6331), .B(n6332), .Z(n6330) );
  XOR U10184 ( .A(DB[2812]), .B(DB[2781]), .Z(n6332) );
  AND U10185 ( .A(n156), .B(n6333), .Z(n6331) );
  XOR U10186 ( .A(n6334), .B(n6335), .Z(n6333) );
  XOR U10187 ( .A(DB[2781]), .B(DB[2750]), .Z(n6335) );
  AND U10188 ( .A(n160), .B(n6336), .Z(n6334) );
  XOR U10189 ( .A(n6337), .B(n6338), .Z(n6336) );
  XOR U10190 ( .A(DB[2750]), .B(DB[2719]), .Z(n6338) );
  AND U10191 ( .A(n164), .B(n6339), .Z(n6337) );
  XOR U10192 ( .A(n6340), .B(n6341), .Z(n6339) );
  XOR U10193 ( .A(DB[2719]), .B(DB[2688]), .Z(n6341) );
  AND U10194 ( .A(n168), .B(n6342), .Z(n6340) );
  XOR U10195 ( .A(n6343), .B(n6344), .Z(n6342) );
  XOR U10196 ( .A(DB[2688]), .B(DB[2657]), .Z(n6344) );
  AND U10197 ( .A(n172), .B(n6345), .Z(n6343) );
  XOR U10198 ( .A(n6346), .B(n6347), .Z(n6345) );
  XOR U10199 ( .A(DB[2657]), .B(DB[2626]), .Z(n6347) );
  AND U10200 ( .A(n176), .B(n6348), .Z(n6346) );
  XOR U10201 ( .A(n6349), .B(n6350), .Z(n6348) );
  XOR U10202 ( .A(DB[2626]), .B(DB[2595]), .Z(n6350) );
  AND U10203 ( .A(n180), .B(n6351), .Z(n6349) );
  XOR U10204 ( .A(n6352), .B(n6353), .Z(n6351) );
  XOR U10205 ( .A(DB[2595]), .B(DB[2564]), .Z(n6353) );
  AND U10206 ( .A(n184), .B(n6354), .Z(n6352) );
  XOR U10207 ( .A(n6355), .B(n6356), .Z(n6354) );
  XOR U10208 ( .A(DB[2564]), .B(DB[2533]), .Z(n6356) );
  AND U10209 ( .A(n188), .B(n6357), .Z(n6355) );
  XOR U10210 ( .A(n6358), .B(n6359), .Z(n6357) );
  XOR U10211 ( .A(DB[2533]), .B(DB[2502]), .Z(n6359) );
  AND U10212 ( .A(n192), .B(n6360), .Z(n6358) );
  XOR U10213 ( .A(n6361), .B(n6362), .Z(n6360) );
  XOR U10214 ( .A(DB[2502]), .B(DB[2471]), .Z(n6362) );
  AND U10215 ( .A(n196), .B(n6363), .Z(n6361) );
  XOR U10216 ( .A(n6364), .B(n6365), .Z(n6363) );
  XOR U10217 ( .A(DB[2471]), .B(DB[2440]), .Z(n6365) );
  AND U10218 ( .A(n200), .B(n6366), .Z(n6364) );
  XOR U10219 ( .A(n6367), .B(n6368), .Z(n6366) );
  XOR U10220 ( .A(DB[2440]), .B(DB[2409]), .Z(n6368) );
  AND U10221 ( .A(n204), .B(n6369), .Z(n6367) );
  XOR U10222 ( .A(n6370), .B(n6371), .Z(n6369) );
  XOR U10223 ( .A(DB[2409]), .B(DB[2378]), .Z(n6371) );
  AND U10224 ( .A(n208), .B(n6372), .Z(n6370) );
  XOR U10225 ( .A(n6373), .B(n6374), .Z(n6372) );
  XOR U10226 ( .A(DB[2378]), .B(DB[2347]), .Z(n6374) );
  AND U10227 ( .A(n212), .B(n6375), .Z(n6373) );
  XOR U10228 ( .A(n6376), .B(n6377), .Z(n6375) );
  XOR U10229 ( .A(DB[2347]), .B(DB[2316]), .Z(n6377) );
  AND U10230 ( .A(n216), .B(n6378), .Z(n6376) );
  XOR U10231 ( .A(n6379), .B(n6380), .Z(n6378) );
  XOR U10232 ( .A(DB[2316]), .B(DB[2285]), .Z(n6380) );
  AND U10233 ( .A(n220), .B(n6381), .Z(n6379) );
  XOR U10234 ( .A(n6382), .B(n6383), .Z(n6381) );
  XOR U10235 ( .A(DB[2285]), .B(DB[2254]), .Z(n6383) );
  AND U10236 ( .A(n224), .B(n6384), .Z(n6382) );
  XOR U10237 ( .A(n6385), .B(n6386), .Z(n6384) );
  XOR U10238 ( .A(DB[2254]), .B(DB[2223]), .Z(n6386) );
  AND U10239 ( .A(n228), .B(n6387), .Z(n6385) );
  XOR U10240 ( .A(n6388), .B(n6389), .Z(n6387) );
  XOR U10241 ( .A(DB[2223]), .B(DB[2192]), .Z(n6389) );
  AND U10242 ( .A(n232), .B(n6390), .Z(n6388) );
  XOR U10243 ( .A(n6391), .B(n6392), .Z(n6390) );
  XOR U10244 ( .A(DB[2192]), .B(DB[2161]), .Z(n6392) );
  AND U10245 ( .A(n236), .B(n6393), .Z(n6391) );
  XOR U10246 ( .A(n6394), .B(n6395), .Z(n6393) );
  XOR U10247 ( .A(DB[2161]), .B(DB[2130]), .Z(n6395) );
  AND U10248 ( .A(n240), .B(n6396), .Z(n6394) );
  XOR U10249 ( .A(n6397), .B(n6398), .Z(n6396) );
  XOR U10250 ( .A(DB[2130]), .B(DB[2099]), .Z(n6398) );
  AND U10251 ( .A(n244), .B(n6399), .Z(n6397) );
  XOR U10252 ( .A(n6400), .B(n6401), .Z(n6399) );
  XOR U10253 ( .A(DB[2099]), .B(DB[2068]), .Z(n6401) );
  AND U10254 ( .A(n248), .B(n6402), .Z(n6400) );
  XOR U10255 ( .A(n6403), .B(n6404), .Z(n6402) );
  XOR U10256 ( .A(DB[2068]), .B(DB[2037]), .Z(n6404) );
  AND U10257 ( .A(n252), .B(n6405), .Z(n6403) );
  XOR U10258 ( .A(n6406), .B(n6407), .Z(n6405) );
  XOR U10259 ( .A(DB[2037]), .B(DB[2006]), .Z(n6407) );
  AND U10260 ( .A(n256), .B(n6408), .Z(n6406) );
  XOR U10261 ( .A(n6409), .B(n6410), .Z(n6408) );
  XOR U10262 ( .A(DB[2006]), .B(DB[1975]), .Z(n6410) );
  AND U10263 ( .A(n260), .B(n6411), .Z(n6409) );
  XOR U10264 ( .A(n6412), .B(n6413), .Z(n6411) );
  XOR U10265 ( .A(DB[1975]), .B(DB[1944]), .Z(n6413) );
  AND U10266 ( .A(n264), .B(n6414), .Z(n6412) );
  XOR U10267 ( .A(n6415), .B(n6416), .Z(n6414) );
  XOR U10268 ( .A(DB[1944]), .B(DB[1913]), .Z(n6416) );
  AND U10269 ( .A(n268), .B(n6417), .Z(n6415) );
  XOR U10270 ( .A(n6418), .B(n6419), .Z(n6417) );
  XOR U10271 ( .A(DB[1913]), .B(DB[1882]), .Z(n6419) );
  AND U10272 ( .A(n272), .B(n6420), .Z(n6418) );
  XOR U10273 ( .A(n6421), .B(n6422), .Z(n6420) );
  XOR U10274 ( .A(DB[1882]), .B(DB[1851]), .Z(n6422) );
  AND U10275 ( .A(n276), .B(n6423), .Z(n6421) );
  XOR U10276 ( .A(n6424), .B(n6425), .Z(n6423) );
  XOR U10277 ( .A(DB[1851]), .B(DB[1820]), .Z(n6425) );
  AND U10278 ( .A(n280), .B(n6426), .Z(n6424) );
  XOR U10279 ( .A(n6427), .B(n6428), .Z(n6426) );
  XOR U10280 ( .A(DB[1820]), .B(DB[1789]), .Z(n6428) );
  AND U10281 ( .A(n284), .B(n6429), .Z(n6427) );
  XOR U10282 ( .A(n6430), .B(n6431), .Z(n6429) );
  XOR U10283 ( .A(DB[1789]), .B(DB[1758]), .Z(n6431) );
  AND U10284 ( .A(n288), .B(n6432), .Z(n6430) );
  XOR U10285 ( .A(n6433), .B(n6434), .Z(n6432) );
  XOR U10286 ( .A(DB[1758]), .B(DB[1727]), .Z(n6434) );
  AND U10287 ( .A(n292), .B(n6435), .Z(n6433) );
  XOR U10288 ( .A(n6436), .B(n6437), .Z(n6435) );
  XOR U10289 ( .A(DB[1727]), .B(DB[1696]), .Z(n6437) );
  AND U10290 ( .A(n296), .B(n6438), .Z(n6436) );
  XOR U10291 ( .A(n6439), .B(n6440), .Z(n6438) );
  XOR U10292 ( .A(DB[1696]), .B(DB[1665]), .Z(n6440) );
  AND U10293 ( .A(n300), .B(n6441), .Z(n6439) );
  XOR U10294 ( .A(n6442), .B(n6443), .Z(n6441) );
  XOR U10295 ( .A(DB[1665]), .B(DB[1634]), .Z(n6443) );
  AND U10296 ( .A(n304), .B(n6444), .Z(n6442) );
  XOR U10297 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U10298 ( .A(DB[1634]), .B(DB[1603]), .Z(n6446) );
  AND U10299 ( .A(n308), .B(n6447), .Z(n6445) );
  XOR U10300 ( .A(n6448), .B(n6449), .Z(n6447) );
  XOR U10301 ( .A(DB[1603]), .B(DB[1572]), .Z(n6449) );
  AND U10302 ( .A(n312), .B(n6450), .Z(n6448) );
  XOR U10303 ( .A(n6451), .B(n6452), .Z(n6450) );
  XOR U10304 ( .A(DB[1572]), .B(DB[1541]), .Z(n6452) );
  AND U10305 ( .A(n316), .B(n6453), .Z(n6451) );
  XOR U10306 ( .A(n6454), .B(n6455), .Z(n6453) );
  XOR U10307 ( .A(DB[1541]), .B(DB[1510]), .Z(n6455) );
  AND U10308 ( .A(n320), .B(n6456), .Z(n6454) );
  XOR U10309 ( .A(n6457), .B(n6458), .Z(n6456) );
  XOR U10310 ( .A(DB[1510]), .B(DB[1479]), .Z(n6458) );
  AND U10311 ( .A(n324), .B(n6459), .Z(n6457) );
  XOR U10312 ( .A(n6460), .B(n6461), .Z(n6459) );
  XOR U10313 ( .A(DB[1479]), .B(DB[1448]), .Z(n6461) );
  AND U10314 ( .A(n328), .B(n6462), .Z(n6460) );
  XOR U10315 ( .A(n6463), .B(n6464), .Z(n6462) );
  XOR U10316 ( .A(DB[1448]), .B(DB[1417]), .Z(n6464) );
  AND U10317 ( .A(n332), .B(n6465), .Z(n6463) );
  XOR U10318 ( .A(n6466), .B(n6467), .Z(n6465) );
  XOR U10319 ( .A(DB[1417]), .B(DB[1386]), .Z(n6467) );
  AND U10320 ( .A(n336), .B(n6468), .Z(n6466) );
  XOR U10321 ( .A(n6469), .B(n6470), .Z(n6468) );
  XOR U10322 ( .A(DB[1386]), .B(DB[1355]), .Z(n6470) );
  AND U10323 ( .A(n340), .B(n6471), .Z(n6469) );
  XOR U10324 ( .A(n6472), .B(n6473), .Z(n6471) );
  XOR U10325 ( .A(DB[1355]), .B(DB[1324]), .Z(n6473) );
  AND U10326 ( .A(n344), .B(n6474), .Z(n6472) );
  XOR U10327 ( .A(n6475), .B(n6476), .Z(n6474) );
  XOR U10328 ( .A(DB[1324]), .B(DB[1293]), .Z(n6476) );
  AND U10329 ( .A(n348), .B(n6477), .Z(n6475) );
  XOR U10330 ( .A(n6478), .B(n6479), .Z(n6477) );
  XOR U10331 ( .A(DB[1293]), .B(DB[1262]), .Z(n6479) );
  AND U10332 ( .A(n352), .B(n6480), .Z(n6478) );
  XOR U10333 ( .A(n6481), .B(n6482), .Z(n6480) );
  XOR U10334 ( .A(DB[1262]), .B(DB[1231]), .Z(n6482) );
  AND U10335 ( .A(n356), .B(n6483), .Z(n6481) );
  XOR U10336 ( .A(n6484), .B(n6485), .Z(n6483) );
  XOR U10337 ( .A(DB[1231]), .B(DB[1200]), .Z(n6485) );
  AND U10338 ( .A(n360), .B(n6486), .Z(n6484) );
  XOR U10339 ( .A(n6487), .B(n6488), .Z(n6486) );
  XOR U10340 ( .A(DB[1200]), .B(DB[1169]), .Z(n6488) );
  AND U10341 ( .A(n364), .B(n6489), .Z(n6487) );
  XOR U10342 ( .A(n6490), .B(n6491), .Z(n6489) );
  XOR U10343 ( .A(DB[1169]), .B(DB[1138]), .Z(n6491) );
  AND U10344 ( .A(n368), .B(n6492), .Z(n6490) );
  XOR U10345 ( .A(n6493), .B(n6494), .Z(n6492) );
  XOR U10346 ( .A(DB[1138]), .B(DB[1107]), .Z(n6494) );
  AND U10347 ( .A(n372), .B(n6495), .Z(n6493) );
  XOR U10348 ( .A(n6496), .B(n6497), .Z(n6495) );
  XOR U10349 ( .A(DB[1107]), .B(DB[1076]), .Z(n6497) );
  AND U10350 ( .A(n376), .B(n6498), .Z(n6496) );
  XOR U10351 ( .A(n6499), .B(n6500), .Z(n6498) );
  XOR U10352 ( .A(DB[1076]), .B(DB[1045]), .Z(n6500) );
  AND U10353 ( .A(n380), .B(n6501), .Z(n6499) );
  XOR U10354 ( .A(n6502), .B(n6503), .Z(n6501) );
  XOR U10355 ( .A(DB[1045]), .B(DB[1014]), .Z(n6503) );
  AND U10356 ( .A(n384), .B(n6504), .Z(n6502) );
  XOR U10357 ( .A(n6505), .B(n6506), .Z(n6504) );
  XOR U10358 ( .A(DB[983]), .B(DB[1014]), .Z(n6506) );
  AND U10359 ( .A(n388), .B(n6507), .Z(n6505) );
  XOR U10360 ( .A(n6508), .B(n6509), .Z(n6507) );
  XOR U10361 ( .A(DB[983]), .B(DB[952]), .Z(n6509) );
  AND U10362 ( .A(n392), .B(n6510), .Z(n6508) );
  XOR U10363 ( .A(n6511), .B(n6512), .Z(n6510) );
  XOR U10364 ( .A(DB[952]), .B(DB[921]), .Z(n6512) );
  AND U10365 ( .A(n396), .B(n6513), .Z(n6511) );
  XOR U10366 ( .A(n6514), .B(n6515), .Z(n6513) );
  XOR U10367 ( .A(DB[921]), .B(DB[890]), .Z(n6515) );
  AND U10368 ( .A(n400), .B(n6516), .Z(n6514) );
  XOR U10369 ( .A(n6517), .B(n6518), .Z(n6516) );
  XOR U10370 ( .A(DB[890]), .B(DB[859]), .Z(n6518) );
  AND U10371 ( .A(n404), .B(n6519), .Z(n6517) );
  XOR U10372 ( .A(n6520), .B(n6521), .Z(n6519) );
  XOR U10373 ( .A(DB[859]), .B(DB[828]), .Z(n6521) );
  AND U10374 ( .A(n408), .B(n6522), .Z(n6520) );
  XOR U10375 ( .A(n6523), .B(n6524), .Z(n6522) );
  XOR U10376 ( .A(DB[828]), .B(DB[797]), .Z(n6524) );
  AND U10377 ( .A(n412), .B(n6525), .Z(n6523) );
  XOR U10378 ( .A(n6526), .B(n6527), .Z(n6525) );
  XOR U10379 ( .A(DB[797]), .B(DB[766]), .Z(n6527) );
  AND U10380 ( .A(n416), .B(n6528), .Z(n6526) );
  XOR U10381 ( .A(n6529), .B(n6530), .Z(n6528) );
  XOR U10382 ( .A(DB[766]), .B(DB[735]), .Z(n6530) );
  AND U10383 ( .A(n420), .B(n6531), .Z(n6529) );
  XOR U10384 ( .A(n6532), .B(n6533), .Z(n6531) );
  XOR U10385 ( .A(DB[735]), .B(DB[704]), .Z(n6533) );
  AND U10386 ( .A(n424), .B(n6534), .Z(n6532) );
  XOR U10387 ( .A(n6535), .B(n6536), .Z(n6534) );
  XOR U10388 ( .A(DB[704]), .B(DB[673]), .Z(n6536) );
  AND U10389 ( .A(n428), .B(n6537), .Z(n6535) );
  XOR U10390 ( .A(n6538), .B(n6539), .Z(n6537) );
  XOR U10391 ( .A(DB[673]), .B(DB[642]), .Z(n6539) );
  AND U10392 ( .A(n432), .B(n6540), .Z(n6538) );
  XOR U10393 ( .A(n6541), .B(n6542), .Z(n6540) );
  XOR U10394 ( .A(DB[642]), .B(DB[611]), .Z(n6542) );
  AND U10395 ( .A(n436), .B(n6543), .Z(n6541) );
  XOR U10396 ( .A(n6544), .B(n6545), .Z(n6543) );
  XOR U10397 ( .A(DB[611]), .B(DB[580]), .Z(n6545) );
  AND U10398 ( .A(n440), .B(n6546), .Z(n6544) );
  XOR U10399 ( .A(n6547), .B(n6548), .Z(n6546) );
  XOR U10400 ( .A(DB[580]), .B(DB[549]), .Z(n6548) );
  AND U10401 ( .A(n444), .B(n6549), .Z(n6547) );
  XOR U10402 ( .A(n6550), .B(n6551), .Z(n6549) );
  XOR U10403 ( .A(DB[549]), .B(DB[518]), .Z(n6551) );
  AND U10404 ( .A(n448), .B(n6552), .Z(n6550) );
  XOR U10405 ( .A(n6553), .B(n6554), .Z(n6552) );
  XOR U10406 ( .A(DB[518]), .B(DB[487]), .Z(n6554) );
  AND U10407 ( .A(n452), .B(n6555), .Z(n6553) );
  XOR U10408 ( .A(n6556), .B(n6557), .Z(n6555) );
  XOR U10409 ( .A(DB[487]), .B(DB[456]), .Z(n6557) );
  AND U10410 ( .A(n456), .B(n6558), .Z(n6556) );
  XOR U10411 ( .A(n6559), .B(n6560), .Z(n6558) );
  XOR U10412 ( .A(DB[456]), .B(DB[425]), .Z(n6560) );
  AND U10413 ( .A(n460), .B(n6561), .Z(n6559) );
  XOR U10414 ( .A(n6562), .B(n6563), .Z(n6561) );
  XOR U10415 ( .A(DB[425]), .B(DB[394]), .Z(n6563) );
  AND U10416 ( .A(n464), .B(n6564), .Z(n6562) );
  XOR U10417 ( .A(n6565), .B(n6566), .Z(n6564) );
  XOR U10418 ( .A(DB[394]), .B(DB[363]), .Z(n6566) );
  AND U10419 ( .A(n468), .B(n6567), .Z(n6565) );
  XOR U10420 ( .A(n6568), .B(n6569), .Z(n6567) );
  XOR U10421 ( .A(DB[363]), .B(DB[332]), .Z(n6569) );
  AND U10422 ( .A(n472), .B(n6570), .Z(n6568) );
  XOR U10423 ( .A(n6571), .B(n6572), .Z(n6570) );
  XOR U10424 ( .A(DB[332]), .B(DB[301]), .Z(n6572) );
  AND U10425 ( .A(n476), .B(n6573), .Z(n6571) );
  XOR U10426 ( .A(n6574), .B(n6575), .Z(n6573) );
  XOR U10427 ( .A(DB[301]), .B(DB[270]), .Z(n6575) );
  AND U10428 ( .A(n480), .B(n6576), .Z(n6574) );
  XOR U10429 ( .A(n6577), .B(n6578), .Z(n6576) );
  XOR U10430 ( .A(DB[270]), .B(DB[239]), .Z(n6578) );
  AND U10431 ( .A(n484), .B(n6579), .Z(n6577) );
  XOR U10432 ( .A(n6580), .B(n6581), .Z(n6579) );
  XOR U10433 ( .A(DB[239]), .B(DB[208]), .Z(n6581) );
  AND U10434 ( .A(n488), .B(n6582), .Z(n6580) );
  XOR U10435 ( .A(n6583), .B(n6584), .Z(n6582) );
  XOR U10436 ( .A(DB[208]), .B(DB[177]), .Z(n6584) );
  AND U10437 ( .A(n492), .B(n6585), .Z(n6583) );
  XOR U10438 ( .A(n6586), .B(n6587), .Z(n6585) );
  XOR U10439 ( .A(DB[177]), .B(DB[146]), .Z(n6587) );
  AND U10440 ( .A(n496), .B(n6588), .Z(n6586) );
  XOR U10441 ( .A(n6589), .B(n6590), .Z(n6588) );
  XOR U10442 ( .A(DB[146]), .B(DB[115]), .Z(n6590) );
  AND U10443 ( .A(n500), .B(n6591), .Z(n6589) );
  XOR U10444 ( .A(n6592), .B(n6593), .Z(n6591) );
  XOR U10445 ( .A(DB[84]), .B(DB[115]), .Z(n6593) );
  AND U10446 ( .A(n504), .B(n6594), .Z(n6592) );
  XOR U10447 ( .A(n6595), .B(n6596), .Z(n6594) );
  XOR U10448 ( .A(DB[84]), .B(DB[53]), .Z(n6596) );
  AND U10449 ( .A(n508), .B(n6597), .Z(n6595) );
  XOR U10450 ( .A(DB[53]), .B(DB[22]), .Z(n6597) );
  XOR U10451 ( .A(DB[3958]), .B(n6598), .Z(min_val_out[21]) );
  AND U10452 ( .A(n2), .B(n6599), .Z(n6598) );
  XOR U10453 ( .A(n6600), .B(n6601), .Z(n6599) );
  XOR U10454 ( .A(n6602), .B(n6603), .Z(n6601) );
  IV U10455 ( .A(DB[3958]), .Z(n6602) );
  AND U10456 ( .A(n8), .B(n6604), .Z(n6600) );
  XOR U10457 ( .A(n6605), .B(n6606), .Z(n6604) );
  XOR U10458 ( .A(DB[3927]), .B(DB[3896]), .Z(n6606) );
  AND U10459 ( .A(n12), .B(n6607), .Z(n6605) );
  XOR U10460 ( .A(n6608), .B(n6609), .Z(n6607) );
  XOR U10461 ( .A(DB[3896]), .B(DB[3865]), .Z(n6609) );
  AND U10462 ( .A(n16), .B(n6610), .Z(n6608) );
  XOR U10463 ( .A(n6611), .B(n6612), .Z(n6610) );
  XOR U10464 ( .A(DB[3865]), .B(DB[3834]), .Z(n6612) );
  AND U10465 ( .A(n20), .B(n6613), .Z(n6611) );
  XOR U10466 ( .A(n6614), .B(n6615), .Z(n6613) );
  XOR U10467 ( .A(DB[3834]), .B(DB[3803]), .Z(n6615) );
  AND U10468 ( .A(n24), .B(n6616), .Z(n6614) );
  XOR U10469 ( .A(n6617), .B(n6618), .Z(n6616) );
  XOR U10470 ( .A(DB[3803]), .B(DB[3772]), .Z(n6618) );
  AND U10471 ( .A(n28), .B(n6619), .Z(n6617) );
  XOR U10472 ( .A(n6620), .B(n6621), .Z(n6619) );
  XOR U10473 ( .A(DB[3772]), .B(DB[3741]), .Z(n6621) );
  AND U10474 ( .A(n32), .B(n6622), .Z(n6620) );
  XOR U10475 ( .A(n6623), .B(n6624), .Z(n6622) );
  XOR U10476 ( .A(DB[3741]), .B(DB[3710]), .Z(n6624) );
  AND U10477 ( .A(n36), .B(n6625), .Z(n6623) );
  XOR U10478 ( .A(n6626), .B(n6627), .Z(n6625) );
  XOR U10479 ( .A(DB[3710]), .B(DB[3679]), .Z(n6627) );
  AND U10480 ( .A(n40), .B(n6628), .Z(n6626) );
  XOR U10481 ( .A(n6629), .B(n6630), .Z(n6628) );
  XOR U10482 ( .A(DB[3679]), .B(DB[3648]), .Z(n6630) );
  AND U10483 ( .A(n44), .B(n6631), .Z(n6629) );
  XOR U10484 ( .A(n6632), .B(n6633), .Z(n6631) );
  XOR U10485 ( .A(DB[3648]), .B(DB[3617]), .Z(n6633) );
  AND U10486 ( .A(n48), .B(n6634), .Z(n6632) );
  XOR U10487 ( .A(n6635), .B(n6636), .Z(n6634) );
  XOR U10488 ( .A(DB[3617]), .B(DB[3586]), .Z(n6636) );
  AND U10489 ( .A(n52), .B(n6637), .Z(n6635) );
  XOR U10490 ( .A(n6638), .B(n6639), .Z(n6637) );
  XOR U10491 ( .A(DB[3586]), .B(DB[3555]), .Z(n6639) );
  AND U10492 ( .A(n56), .B(n6640), .Z(n6638) );
  XOR U10493 ( .A(n6641), .B(n6642), .Z(n6640) );
  XOR U10494 ( .A(DB[3555]), .B(DB[3524]), .Z(n6642) );
  AND U10495 ( .A(n60), .B(n6643), .Z(n6641) );
  XOR U10496 ( .A(n6644), .B(n6645), .Z(n6643) );
  XOR U10497 ( .A(DB[3524]), .B(DB[3493]), .Z(n6645) );
  AND U10498 ( .A(n64), .B(n6646), .Z(n6644) );
  XOR U10499 ( .A(n6647), .B(n6648), .Z(n6646) );
  XOR U10500 ( .A(DB[3493]), .B(DB[3462]), .Z(n6648) );
  AND U10501 ( .A(n68), .B(n6649), .Z(n6647) );
  XOR U10502 ( .A(n6650), .B(n6651), .Z(n6649) );
  XOR U10503 ( .A(DB[3462]), .B(DB[3431]), .Z(n6651) );
  AND U10504 ( .A(n72), .B(n6652), .Z(n6650) );
  XOR U10505 ( .A(n6653), .B(n6654), .Z(n6652) );
  XOR U10506 ( .A(DB[3431]), .B(DB[3400]), .Z(n6654) );
  AND U10507 ( .A(n76), .B(n6655), .Z(n6653) );
  XOR U10508 ( .A(n6656), .B(n6657), .Z(n6655) );
  XOR U10509 ( .A(DB[3400]), .B(DB[3369]), .Z(n6657) );
  AND U10510 ( .A(n80), .B(n6658), .Z(n6656) );
  XOR U10511 ( .A(n6659), .B(n6660), .Z(n6658) );
  XOR U10512 ( .A(DB[3369]), .B(DB[3338]), .Z(n6660) );
  AND U10513 ( .A(n84), .B(n6661), .Z(n6659) );
  XOR U10514 ( .A(n6662), .B(n6663), .Z(n6661) );
  XOR U10515 ( .A(DB[3338]), .B(DB[3307]), .Z(n6663) );
  AND U10516 ( .A(n88), .B(n6664), .Z(n6662) );
  XOR U10517 ( .A(n6665), .B(n6666), .Z(n6664) );
  XOR U10518 ( .A(DB[3307]), .B(DB[3276]), .Z(n6666) );
  AND U10519 ( .A(n92), .B(n6667), .Z(n6665) );
  XOR U10520 ( .A(n6668), .B(n6669), .Z(n6667) );
  XOR U10521 ( .A(DB[3276]), .B(DB[3245]), .Z(n6669) );
  AND U10522 ( .A(n96), .B(n6670), .Z(n6668) );
  XOR U10523 ( .A(n6671), .B(n6672), .Z(n6670) );
  XOR U10524 ( .A(DB[3245]), .B(DB[3214]), .Z(n6672) );
  AND U10525 ( .A(n100), .B(n6673), .Z(n6671) );
  XOR U10526 ( .A(n6674), .B(n6675), .Z(n6673) );
  XOR U10527 ( .A(DB[3214]), .B(DB[3183]), .Z(n6675) );
  AND U10528 ( .A(n104), .B(n6676), .Z(n6674) );
  XOR U10529 ( .A(n6677), .B(n6678), .Z(n6676) );
  XOR U10530 ( .A(DB[3183]), .B(DB[3152]), .Z(n6678) );
  AND U10531 ( .A(n108), .B(n6679), .Z(n6677) );
  XOR U10532 ( .A(n6680), .B(n6681), .Z(n6679) );
  XOR U10533 ( .A(DB[3152]), .B(DB[3121]), .Z(n6681) );
  AND U10534 ( .A(n112), .B(n6682), .Z(n6680) );
  XOR U10535 ( .A(n6683), .B(n6684), .Z(n6682) );
  XOR U10536 ( .A(DB[3121]), .B(DB[3090]), .Z(n6684) );
  AND U10537 ( .A(n116), .B(n6685), .Z(n6683) );
  XOR U10538 ( .A(n6686), .B(n6687), .Z(n6685) );
  XOR U10539 ( .A(DB[3090]), .B(DB[3059]), .Z(n6687) );
  AND U10540 ( .A(n120), .B(n6688), .Z(n6686) );
  XOR U10541 ( .A(n6689), .B(n6690), .Z(n6688) );
  XOR U10542 ( .A(DB[3059]), .B(DB[3028]), .Z(n6690) );
  AND U10543 ( .A(n124), .B(n6691), .Z(n6689) );
  XOR U10544 ( .A(n6692), .B(n6693), .Z(n6691) );
  XOR U10545 ( .A(DB[3028]), .B(DB[2997]), .Z(n6693) );
  AND U10546 ( .A(n128), .B(n6694), .Z(n6692) );
  XOR U10547 ( .A(n6695), .B(n6696), .Z(n6694) );
  XOR U10548 ( .A(DB[2997]), .B(DB[2966]), .Z(n6696) );
  AND U10549 ( .A(n132), .B(n6697), .Z(n6695) );
  XOR U10550 ( .A(n6698), .B(n6699), .Z(n6697) );
  XOR U10551 ( .A(DB[2966]), .B(DB[2935]), .Z(n6699) );
  AND U10552 ( .A(n136), .B(n6700), .Z(n6698) );
  XOR U10553 ( .A(n6701), .B(n6702), .Z(n6700) );
  XOR U10554 ( .A(DB[2935]), .B(DB[2904]), .Z(n6702) );
  AND U10555 ( .A(n140), .B(n6703), .Z(n6701) );
  XOR U10556 ( .A(n6704), .B(n6705), .Z(n6703) );
  XOR U10557 ( .A(DB[2904]), .B(DB[2873]), .Z(n6705) );
  AND U10558 ( .A(n144), .B(n6706), .Z(n6704) );
  XOR U10559 ( .A(n6707), .B(n6708), .Z(n6706) );
  XOR U10560 ( .A(DB[2873]), .B(DB[2842]), .Z(n6708) );
  AND U10561 ( .A(n148), .B(n6709), .Z(n6707) );
  XOR U10562 ( .A(n6710), .B(n6711), .Z(n6709) );
  XOR U10563 ( .A(DB[2842]), .B(DB[2811]), .Z(n6711) );
  AND U10564 ( .A(n152), .B(n6712), .Z(n6710) );
  XOR U10565 ( .A(n6713), .B(n6714), .Z(n6712) );
  XOR U10566 ( .A(DB[2811]), .B(DB[2780]), .Z(n6714) );
  AND U10567 ( .A(n156), .B(n6715), .Z(n6713) );
  XOR U10568 ( .A(n6716), .B(n6717), .Z(n6715) );
  XOR U10569 ( .A(DB[2780]), .B(DB[2749]), .Z(n6717) );
  AND U10570 ( .A(n160), .B(n6718), .Z(n6716) );
  XOR U10571 ( .A(n6719), .B(n6720), .Z(n6718) );
  XOR U10572 ( .A(DB[2749]), .B(DB[2718]), .Z(n6720) );
  AND U10573 ( .A(n164), .B(n6721), .Z(n6719) );
  XOR U10574 ( .A(n6722), .B(n6723), .Z(n6721) );
  XOR U10575 ( .A(DB[2718]), .B(DB[2687]), .Z(n6723) );
  AND U10576 ( .A(n168), .B(n6724), .Z(n6722) );
  XOR U10577 ( .A(n6725), .B(n6726), .Z(n6724) );
  XOR U10578 ( .A(DB[2687]), .B(DB[2656]), .Z(n6726) );
  AND U10579 ( .A(n172), .B(n6727), .Z(n6725) );
  XOR U10580 ( .A(n6728), .B(n6729), .Z(n6727) );
  XOR U10581 ( .A(DB[2656]), .B(DB[2625]), .Z(n6729) );
  AND U10582 ( .A(n176), .B(n6730), .Z(n6728) );
  XOR U10583 ( .A(n6731), .B(n6732), .Z(n6730) );
  XOR U10584 ( .A(DB[2625]), .B(DB[2594]), .Z(n6732) );
  AND U10585 ( .A(n180), .B(n6733), .Z(n6731) );
  XOR U10586 ( .A(n6734), .B(n6735), .Z(n6733) );
  XOR U10587 ( .A(DB[2594]), .B(DB[2563]), .Z(n6735) );
  AND U10588 ( .A(n184), .B(n6736), .Z(n6734) );
  XOR U10589 ( .A(n6737), .B(n6738), .Z(n6736) );
  XOR U10590 ( .A(DB[2563]), .B(DB[2532]), .Z(n6738) );
  AND U10591 ( .A(n188), .B(n6739), .Z(n6737) );
  XOR U10592 ( .A(n6740), .B(n6741), .Z(n6739) );
  XOR U10593 ( .A(DB[2532]), .B(DB[2501]), .Z(n6741) );
  AND U10594 ( .A(n192), .B(n6742), .Z(n6740) );
  XOR U10595 ( .A(n6743), .B(n6744), .Z(n6742) );
  XOR U10596 ( .A(DB[2501]), .B(DB[2470]), .Z(n6744) );
  AND U10597 ( .A(n196), .B(n6745), .Z(n6743) );
  XOR U10598 ( .A(n6746), .B(n6747), .Z(n6745) );
  XOR U10599 ( .A(DB[2470]), .B(DB[2439]), .Z(n6747) );
  AND U10600 ( .A(n200), .B(n6748), .Z(n6746) );
  XOR U10601 ( .A(n6749), .B(n6750), .Z(n6748) );
  XOR U10602 ( .A(DB[2439]), .B(DB[2408]), .Z(n6750) );
  AND U10603 ( .A(n204), .B(n6751), .Z(n6749) );
  XOR U10604 ( .A(n6752), .B(n6753), .Z(n6751) );
  XOR U10605 ( .A(DB[2408]), .B(DB[2377]), .Z(n6753) );
  AND U10606 ( .A(n208), .B(n6754), .Z(n6752) );
  XOR U10607 ( .A(n6755), .B(n6756), .Z(n6754) );
  XOR U10608 ( .A(DB[2377]), .B(DB[2346]), .Z(n6756) );
  AND U10609 ( .A(n212), .B(n6757), .Z(n6755) );
  XOR U10610 ( .A(n6758), .B(n6759), .Z(n6757) );
  XOR U10611 ( .A(DB[2346]), .B(DB[2315]), .Z(n6759) );
  AND U10612 ( .A(n216), .B(n6760), .Z(n6758) );
  XOR U10613 ( .A(n6761), .B(n6762), .Z(n6760) );
  XOR U10614 ( .A(DB[2315]), .B(DB[2284]), .Z(n6762) );
  AND U10615 ( .A(n220), .B(n6763), .Z(n6761) );
  XOR U10616 ( .A(n6764), .B(n6765), .Z(n6763) );
  XOR U10617 ( .A(DB[2284]), .B(DB[2253]), .Z(n6765) );
  AND U10618 ( .A(n224), .B(n6766), .Z(n6764) );
  XOR U10619 ( .A(n6767), .B(n6768), .Z(n6766) );
  XOR U10620 ( .A(DB[2253]), .B(DB[2222]), .Z(n6768) );
  AND U10621 ( .A(n228), .B(n6769), .Z(n6767) );
  XOR U10622 ( .A(n6770), .B(n6771), .Z(n6769) );
  XOR U10623 ( .A(DB[2222]), .B(DB[2191]), .Z(n6771) );
  AND U10624 ( .A(n232), .B(n6772), .Z(n6770) );
  XOR U10625 ( .A(n6773), .B(n6774), .Z(n6772) );
  XOR U10626 ( .A(DB[2191]), .B(DB[2160]), .Z(n6774) );
  AND U10627 ( .A(n236), .B(n6775), .Z(n6773) );
  XOR U10628 ( .A(n6776), .B(n6777), .Z(n6775) );
  XOR U10629 ( .A(DB[2160]), .B(DB[2129]), .Z(n6777) );
  AND U10630 ( .A(n240), .B(n6778), .Z(n6776) );
  XOR U10631 ( .A(n6779), .B(n6780), .Z(n6778) );
  XOR U10632 ( .A(DB[2129]), .B(DB[2098]), .Z(n6780) );
  AND U10633 ( .A(n244), .B(n6781), .Z(n6779) );
  XOR U10634 ( .A(n6782), .B(n6783), .Z(n6781) );
  XOR U10635 ( .A(DB[2098]), .B(DB[2067]), .Z(n6783) );
  AND U10636 ( .A(n248), .B(n6784), .Z(n6782) );
  XOR U10637 ( .A(n6785), .B(n6786), .Z(n6784) );
  XOR U10638 ( .A(DB[2067]), .B(DB[2036]), .Z(n6786) );
  AND U10639 ( .A(n252), .B(n6787), .Z(n6785) );
  XOR U10640 ( .A(n6788), .B(n6789), .Z(n6787) );
  XOR U10641 ( .A(DB[2036]), .B(DB[2005]), .Z(n6789) );
  AND U10642 ( .A(n256), .B(n6790), .Z(n6788) );
  XOR U10643 ( .A(n6791), .B(n6792), .Z(n6790) );
  XOR U10644 ( .A(DB[2005]), .B(DB[1974]), .Z(n6792) );
  AND U10645 ( .A(n260), .B(n6793), .Z(n6791) );
  XOR U10646 ( .A(n6794), .B(n6795), .Z(n6793) );
  XOR U10647 ( .A(DB[1974]), .B(DB[1943]), .Z(n6795) );
  AND U10648 ( .A(n264), .B(n6796), .Z(n6794) );
  XOR U10649 ( .A(n6797), .B(n6798), .Z(n6796) );
  XOR U10650 ( .A(DB[1943]), .B(DB[1912]), .Z(n6798) );
  AND U10651 ( .A(n268), .B(n6799), .Z(n6797) );
  XOR U10652 ( .A(n6800), .B(n6801), .Z(n6799) );
  XOR U10653 ( .A(DB[1912]), .B(DB[1881]), .Z(n6801) );
  AND U10654 ( .A(n272), .B(n6802), .Z(n6800) );
  XOR U10655 ( .A(n6803), .B(n6804), .Z(n6802) );
  XOR U10656 ( .A(DB[1881]), .B(DB[1850]), .Z(n6804) );
  AND U10657 ( .A(n276), .B(n6805), .Z(n6803) );
  XOR U10658 ( .A(n6806), .B(n6807), .Z(n6805) );
  XOR U10659 ( .A(DB[1850]), .B(DB[1819]), .Z(n6807) );
  AND U10660 ( .A(n280), .B(n6808), .Z(n6806) );
  XOR U10661 ( .A(n6809), .B(n6810), .Z(n6808) );
  XOR U10662 ( .A(DB[1819]), .B(DB[1788]), .Z(n6810) );
  AND U10663 ( .A(n284), .B(n6811), .Z(n6809) );
  XOR U10664 ( .A(n6812), .B(n6813), .Z(n6811) );
  XOR U10665 ( .A(DB[1788]), .B(DB[1757]), .Z(n6813) );
  AND U10666 ( .A(n288), .B(n6814), .Z(n6812) );
  XOR U10667 ( .A(n6815), .B(n6816), .Z(n6814) );
  XOR U10668 ( .A(DB[1757]), .B(DB[1726]), .Z(n6816) );
  AND U10669 ( .A(n292), .B(n6817), .Z(n6815) );
  XOR U10670 ( .A(n6818), .B(n6819), .Z(n6817) );
  XOR U10671 ( .A(DB[1726]), .B(DB[1695]), .Z(n6819) );
  AND U10672 ( .A(n296), .B(n6820), .Z(n6818) );
  XOR U10673 ( .A(n6821), .B(n6822), .Z(n6820) );
  XOR U10674 ( .A(DB[1695]), .B(DB[1664]), .Z(n6822) );
  AND U10675 ( .A(n300), .B(n6823), .Z(n6821) );
  XOR U10676 ( .A(n6824), .B(n6825), .Z(n6823) );
  XOR U10677 ( .A(DB[1664]), .B(DB[1633]), .Z(n6825) );
  AND U10678 ( .A(n304), .B(n6826), .Z(n6824) );
  XOR U10679 ( .A(n6827), .B(n6828), .Z(n6826) );
  XOR U10680 ( .A(DB[1633]), .B(DB[1602]), .Z(n6828) );
  AND U10681 ( .A(n308), .B(n6829), .Z(n6827) );
  XOR U10682 ( .A(n6830), .B(n6831), .Z(n6829) );
  XOR U10683 ( .A(DB[1602]), .B(DB[1571]), .Z(n6831) );
  AND U10684 ( .A(n312), .B(n6832), .Z(n6830) );
  XOR U10685 ( .A(n6833), .B(n6834), .Z(n6832) );
  XOR U10686 ( .A(DB[1571]), .B(DB[1540]), .Z(n6834) );
  AND U10687 ( .A(n316), .B(n6835), .Z(n6833) );
  XOR U10688 ( .A(n6836), .B(n6837), .Z(n6835) );
  XOR U10689 ( .A(DB[1540]), .B(DB[1509]), .Z(n6837) );
  AND U10690 ( .A(n320), .B(n6838), .Z(n6836) );
  XOR U10691 ( .A(n6839), .B(n6840), .Z(n6838) );
  XOR U10692 ( .A(DB[1509]), .B(DB[1478]), .Z(n6840) );
  AND U10693 ( .A(n324), .B(n6841), .Z(n6839) );
  XOR U10694 ( .A(n6842), .B(n6843), .Z(n6841) );
  XOR U10695 ( .A(DB[1478]), .B(DB[1447]), .Z(n6843) );
  AND U10696 ( .A(n328), .B(n6844), .Z(n6842) );
  XOR U10697 ( .A(n6845), .B(n6846), .Z(n6844) );
  XOR U10698 ( .A(DB[1447]), .B(DB[1416]), .Z(n6846) );
  AND U10699 ( .A(n332), .B(n6847), .Z(n6845) );
  XOR U10700 ( .A(n6848), .B(n6849), .Z(n6847) );
  XOR U10701 ( .A(DB[1416]), .B(DB[1385]), .Z(n6849) );
  AND U10702 ( .A(n336), .B(n6850), .Z(n6848) );
  XOR U10703 ( .A(n6851), .B(n6852), .Z(n6850) );
  XOR U10704 ( .A(DB[1385]), .B(DB[1354]), .Z(n6852) );
  AND U10705 ( .A(n340), .B(n6853), .Z(n6851) );
  XOR U10706 ( .A(n6854), .B(n6855), .Z(n6853) );
  XOR U10707 ( .A(DB[1354]), .B(DB[1323]), .Z(n6855) );
  AND U10708 ( .A(n344), .B(n6856), .Z(n6854) );
  XOR U10709 ( .A(n6857), .B(n6858), .Z(n6856) );
  XOR U10710 ( .A(DB[1323]), .B(DB[1292]), .Z(n6858) );
  AND U10711 ( .A(n348), .B(n6859), .Z(n6857) );
  XOR U10712 ( .A(n6860), .B(n6861), .Z(n6859) );
  XOR U10713 ( .A(DB[1292]), .B(DB[1261]), .Z(n6861) );
  AND U10714 ( .A(n352), .B(n6862), .Z(n6860) );
  XOR U10715 ( .A(n6863), .B(n6864), .Z(n6862) );
  XOR U10716 ( .A(DB[1261]), .B(DB[1230]), .Z(n6864) );
  AND U10717 ( .A(n356), .B(n6865), .Z(n6863) );
  XOR U10718 ( .A(n6866), .B(n6867), .Z(n6865) );
  XOR U10719 ( .A(DB[1230]), .B(DB[1199]), .Z(n6867) );
  AND U10720 ( .A(n360), .B(n6868), .Z(n6866) );
  XOR U10721 ( .A(n6869), .B(n6870), .Z(n6868) );
  XOR U10722 ( .A(DB[1199]), .B(DB[1168]), .Z(n6870) );
  AND U10723 ( .A(n364), .B(n6871), .Z(n6869) );
  XOR U10724 ( .A(n6872), .B(n6873), .Z(n6871) );
  XOR U10725 ( .A(DB[1168]), .B(DB[1137]), .Z(n6873) );
  AND U10726 ( .A(n368), .B(n6874), .Z(n6872) );
  XOR U10727 ( .A(n6875), .B(n6876), .Z(n6874) );
  XOR U10728 ( .A(DB[1137]), .B(DB[1106]), .Z(n6876) );
  AND U10729 ( .A(n372), .B(n6877), .Z(n6875) );
  XOR U10730 ( .A(n6878), .B(n6879), .Z(n6877) );
  XOR U10731 ( .A(DB[1106]), .B(DB[1075]), .Z(n6879) );
  AND U10732 ( .A(n376), .B(n6880), .Z(n6878) );
  XOR U10733 ( .A(n6881), .B(n6882), .Z(n6880) );
  XOR U10734 ( .A(DB[1075]), .B(DB[1044]), .Z(n6882) );
  AND U10735 ( .A(n380), .B(n6883), .Z(n6881) );
  XOR U10736 ( .A(n6884), .B(n6885), .Z(n6883) );
  XOR U10737 ( .A(DB[1044]), .B(DB[1013]), .Z(n6885) );
  AND U10738 ( .A(n384), .B(n6886), .Z(n6884) );
  XOR U10739 ( .A(n6887), .B(n6888), .Z(n6886) );
  XOR U10740 ( .A(DB[982]), .B(DB[1013]), .Z(n6888) );
  AND U10741 ( .A(n388), .B(n6889), .Z(n6887) );
  XOR U10742 ( .A(n6890), .B(n6891), .Z(n6889) );
  XOR U10743 ( .A(DB[982]), .B(DB[951]), .Z(n6891) );
  AND U10744 ( .A(n392), .B(n6892), .Z(n6890) );
  XOR U10745 ( .A(n6893), .B(n6894), .Z(n6892) );
  XOR U10746 ( .A(DB[951]), .B(DB[920]), .Z(n6894) );
  AND U10747 ( .A(n396), .B(n6895), .Z(n6893) );
  XOR U10748 ( .A(n6896), .B(n6897), .Z(n6895) );
  XOR U10749 ( .A(DB[920]), .B(DB[889]), .Z(n6897) );
  AND U10750 ( .A(n400), .B(n6898), .Z(n6896) );
  XOR U10751 ( .A(n6899), .B(n6900), .Z(n6898) );
  XOR U10752 ( .A(DB[889]), .B(DB[858]), .Z(n6900) );
  AND U10753 ( .A(n404), .B(n6901), .Z(n6899) );
  XOR U10754 ( .A(n6902), .B(n6903), .Z(n6901) );
  XOR U10755 ( .A(DB[858]), .B(DB[827]), .Z(n6903) );
  AND U10756 ( .A(n408), .B(n6904), .Z(n6902) );
  XOR U10757 ( .A(n6905), .B(n6906), .Z(n6904) );
  XOR U10758 ( .A(DB[827]), .B(DB[796]), .Z(n6906) );
  AND U10759 ( .A(n412), .B(n6907), .Z(n6905) );
  XOR U10760 ( .A(n6908), .B(n6909), .Z(n6907) );
  XOR U10761 ( .A(DB[796]), .B(DB[765]), .Z(n6909) );
  AND U10762 ( .A(n416), .B(n6910), .Z(n6908) );
  XOR U10763 ( .A(n6911), .B(n6912), .Z(n6910) );
  XOR U10764 ( .A(DB[765]), .B(DB[734]), .Z(n6912) );
  AND U10765 ( .A(n420), .B(n6913), .Z(n6911) );
  XOR U10766 ( .A(n6914), .B(n6915), .Z(n6913) );
  XOR U10767 ( .A(DB[734]), .B(DB[703]), .Z(n6915) );
  AND U10768 ( .A(n424), .B(n6916), .Z(n6914) );
  XOR U10769 ( .A(n6917), .B(n6918), .Z(n6916) );
  XOR U10770 ( .A(DB[703]), .B(DB[672]), .Z(n6918) );
  AND U10771 ( .A(n428), .B(n6919), .Z(n6917) );
  XOR U10772 ( .A(n6920), .B(n6921), .Z(n6919) );
  XOR U10773 ( .A(DB[672]), .B(DB[641]), .Z(n6921) );
  AND U10774 ( .A(n432), .B(n6922), .Z(n6920) );
  XOR U10775 ( .A(n6923), .B(n6924), .Z(n6922) );
  XOR U10776 ( .A(DB[641]), .B(DB[610]), .Z(n6924) );
  AND U10777 ( .A(n436), .B(n6925), .Z(n6923) );
  XOR U10778 ( .A(n6926), .B(n6927), .Z(n6925) );
  XOR U10779 ( .A(DB[610]), .B(DB[579]), .Z(n6927) );
  AND U10780 ( .A(n440), .B(n6928), .Z(n6926) );
  XOR U10781 ( .A(n6929), .B(n6930), .Z(n6928) );
  XOR U10782 ( .A(DB[579]), .B(DB[548]), .Z(n6930) );
  AND U10783 ( .A(n444), .B(n6931), .Z(n6929) );
  XOR U10784 ( .A(n6932), .B(n6933), .Z(n6931) );
  XOR U10785 ( .A(DB[548]), .B(DB[517]), .Z(n6933) );
  AND U10786 ( .A(n448), .B(n6934), .Z(n6932) );
  XOR U10787 ( .A(n6935), .B(n6936), .Z(n6934) );
  XOR U10788 ( .A(DB[517]), .B(DB[486]), .Z(n6936) );
  AND U10789 ( .A(n452), .B(n6937), .Z(n6935) );
  XOR U10790 ( .A(n6938), .B(n6939), .Z(n6937) );
  XOR U10791 ( .A(DB[486]), .B(DB[455]), .Z(n6939) );
  AND U10792 ( .A(n456), .B(n6940), .Z(n6938) );
  XOR U10793 ( .A(n6941), .B(n6942), .Z(n6940) );
  XOR U10794 ( .A(DB[455]), .B(DB[424]), .Z(n6942) );
  AND U10795 ( .A(n460), .B(n6943), .Z(n6941) );
  XOR U10796 ( .A(n6944), .B(n6945), .Z(n6943) );
  XOR U10797 ( .A(DB[424]), .B(DB[393]), .Z(n6945) );
  AND U10798 ( .A(n464), .B(n6946), .Z(n6944) );
  XOR U10799 ( .A(n6947), .B(n6948), .Z(n6946) );
  XOR U10800 ( .A(DB[393]), .B(DB[362]), .Z(n6948) );
  AND U10801 ( .A(n468), .B(n6949), .Z(n6947) );
  XOR U10802 ( .A(n6950), .B(n6951), .Z(n6949) );
  XOR U10803 ( .A(DB[362]), .B(DB[331]), .Z(n6951) );
  AND U10804 ( .A(n472), .B(n6952), .Z(n6950) );
  XOR U10805 ( .A(n6953), .B(n6954), .Z(n6952) );
  XOR U10806 ( .A(DB[331]), .B(DB[300]), .Z(n6954) );
  AND U10807 ( .A(n476), .B(n6955), .Z(n6953) );
  XOR U10808 ( .A(n6956), .B(n6957), .Z(n6955) );
  XOR U10809 ( .A(DB[300]), .B(DB[269]), .Z(n6957) );
  AND U10810 ( .A(n480), .B(n6958), .Z(n6956) );
  XOR U10811 ( .A(n6959), .B(n6960), .Z(n6958) );
  XOR U10812 ( .A(DB[269]), .B(DB[238]), .Z(n6960) );
  AND U10813 ( .A(n484), .B(n6961), .Z(n6959) );
  XOR U10814 ( .A(n6962), .B(n6963), .Z(n6961) );
  XOR U10815 ( .A(DB[238]), .B(DB[207]), .Z(n6963) );
  AND U10816 ( .A(n488), .B(n6964), .Z(n6962) );
  XOR U10817 ( .A(n6965), .B(n6966), .Z(n6964) );
  XOR U10818 ( .A(DB[207]), .B(DB[176]), .Z(n6966) );
  AND U10819 ( .A(n492), .B(n6967), .Z(n6965) );
  XOR U10820 ( .A(n6968), .B(n6969), .Z(n6967) );
  XOR U10821 ( .A(DB[176]), .B(DB[145]), .Z(n6969) );
  AND U10822 ( .A(n496), .B(n6970), .Z(n6968) );
  XOR U10823 ( .A(n6971), .B(n6972), .Z(n6970) );
  XOR U10824 ( .A(DB[145]), .B(DB[114]), .Z(n6972) );
  AND U10825 ( .A(n500), .B(n6973), .Z(n6971) );
  XOR U10826 ( .A(n6974), .B(n6975), .Z(n6973) );
  XOR U10827 ( .A(DB[83]), .B(DB[114]), .Z(n6975) );
  AND U10828 ( .A(n504), .B(n6976), .Z(n6974) );
  XOR U10829 ( .A(n6977), .B(n6978), .Z(n6976) );
  XOR U10830 ( .A(DB[83]), .B(DB[52]), .Z(n6978) );
  AND U10831 ( .A(n508), .B(n6979), .Z(n6977) );
  XOR U10832 ( .A(DB[52]), .B(DB[21]), .Z(n6979) );
  XOR U10833 ( .A(DB[3957]), .B(n6980), .Z(min_val_out[20]) );
  AND U10834 ( .A(n2), .B(n6981), .Z(n6980) );
  XOR U10835 ( .A(n6982), .B(n6983), .Z(n6981) );
  XOR U10836 ( .A(n6984), .B(n6985), .Z(n6983) );
  IV U10837 ( .A(DB[3957]), .Z(n6984) );
  AND U10838 ( .A(n8), .B(n6986), .Z(n6982) );
  XOR U10839 ( .A(n6987), .B(n6988), .Z(n6986) );
  XOR U10840 ( .A(DB[3926]), .B(DB[3895]), .Z(n6988) );
  AND U10841 ( .A(n12), .B(n6989), .Z(n6987) );
  XOR U10842 ( .A(n6990), .B(n6991), .Z(n6989) );
  XOR U10843 ( .A(DB[3895]), .B(DB[3864]), .Z(n6991) );
  AND U10844 ( .A(n16), .B(n6992), .Z(n6990) );
  XOR U10845 ( .A(n6993), .B(n6994), .Z(n6992) );
  XOR U10846 ( .A(DB[3864]), .B(DB[3833]), .Z(n6994) );
  AND U10847 ( .A(n20), .B(n6995), .Z(n6993) );
  XOR U10848 ( .A(n6996), .B(n6997), .Z(n6995) );
  XOR U10849 ( .A(DB[3833]), .B(DB[3802]), .Z(n6997) );
  AND U10850 ( .A(n24), .B(n6998), .Z(n6996) );
  XOR U10851 ( .A(n6999), .B(n7000), .Z(n6998) );
  XOR U10852 ( .A(DB[3802]), .B(DB[3771]), .Z(n7000) );
  AND U10853 ( .A(n28), .B(n7001), .Z(n6999) );
  XOR U10854 ( .A(n7002), .B(n7003), .Z(n7001) );
  XOR U10855 ( .A(DB[3771]), .B(DB[3740]), .Z(n7003) );
  AND U10856 ( .A(n32), .B(n7004), .Z(n7002) );
  XOR U10857 ( .A(n7005), .B(n7006), .Z(n7004) );
  XOR U10858 ( .A(DB[3740]), .B(DB[3709]), .Z(n7006) );
  AND U10859 ( .A(n36), .B(n7007), .Z(n7005) );
  XOR U10860 ( .A(n7008), .B(n7009), .Z(n7007) );
  XOR U10861 ( .A(DB[3709]), .B(DB[3678]), .Z(n7009) );
  AND U10862 ( .A(n40), .B(n7010), .Z(n7008) );
  XOR U10863 ( .A(n7011), .B(n7012), .Z(n7010) );
  XOR U10864 ( .A(DB[3678]), .B(DB[3647]), .Z(n7012) );
  AND U10865 ( .A(n44), .B(n7013), .Z(n7011) );
  XOR U10866 ( .A(n7014), .B(n7015), .Z(n7013) );
  XOR U10867 ( .A(DB[3647]), .B(DB[3616]), .Z(n7015) );
  AND U10868 ( .A(n48), .B(n7016), .Z(n7014) );
  XOR U10869 ( .A(n7017), .B(n7018), .Z(n7016) );
  XOR U10870 ( .A(DB[3616]), .B(DB[3585]), .Z(n7018) );
  AND U10871 ( .A(n52), .B(n7019), .Z(n7017) );
  XOR U10872 ( .A(n7020), .B(n7021), .Z(n7019) );
  XOR U10873 ( .A(DB[3585]), .B(DB[3554]), .Z(n7021) );
  AND U10874 ( .A(n56), .B(n7022), .Z(n7020) );
  XOR U10875 ( .A(n7023), .B(n7024), .Z(n7022) );
  XOR U10876 ( .A(DB[3554]), .B(DB[3523]), .Z(n7024) );
  AND U10877 ( .A(n60), .B(n7025), .Z(n7023) );
  XOR U10878 ( .A(n7026), .B(n7027), .Z(n7025) );
  XOR U10879 ( .A(DB[3523]), .B(DB[3492]), .Z(n7027) );
  AND U10880 ( .A(n64), .B(n7028), .Z(n7026) );
  XOR U10881 ( .A(n7029), .B(n7030), .Z(n7028) );
  XOR U10882 ( .A(DB[3492]), .B(DB[3461]), .Z(n7030) );
  AND U10883 ( .A(n68), .B(n7031), .Z(n7029) );
  XOR U10884 ( .A(n7032), .B(n7033), .Z(n7031) );
  XOR U10885 ( .A(DB[3461]), .B(DB[3430]), .Z(n7033) );
  AND U10886 ( .A(n72), .B(n7034), .Z(n7032) );
  XOR U10887 ( .A(n7035), .B(n7036), .Z(n7034) );
  XOR U10888 ( .A(DB[3430]), .B(DB[3399]), .Z(n7036) );
  AND U10889 ( .A(n76), .B(n7037), .Z(n7035) );
  XOR U10890 ( .A(n7038), .B(n7039), .Z(n7037) );
  XOR U10891 ( .A(DB[3399]), .B(DB[3368]), .Z(n7039) );
  AND U10892 ( .A(n80), .B(n7040), .Z(n7038) );
  XOR U10893 ( .A(n7041), .B(n7042), .Z(n7040) );
  XOR U10894 ( .A(DB[3368]), .B(DB[3337]), .Z(n7042) );
  AND U10895 ( .A(n84), .B(n7043), .Z(n7041) );
  XOR U10896 ( .A(n7044), .B(n7045), .Z(n7043) );
  XOR U10897 ( .A(DB[3337]), .B(DB[3306]), .Z(n7045) );
  AND U10898 ( .A(n88), .B(n7046), .Z(n7044) );
  XOR U10899 ( .A(n7047), .B(n7048), .Z(n7046) );
  XOR U10900 ( .A(DB[3306]), .B(DB[3275]), .Z(n7048) );
  AND U10901 ( .A(n92), .B(n7049), .Z(n7047) );
  XOR U10902 ( .A(n7050), .B(n7051), .Z(n7049) );
  XOR U10903 ( .A(DB[3275]), .B(DB[3244]), .Z(n7051) );
  AND U10904 ( .A(n96), .B(n7052), .Z(n7050) );
  XOR U10905 ( .A(n7053), .B(n7054), .Z(n7052) );
  XOR U10906 ( .A(DB[3244]), .B(DB[3213]), .Z(n7054) );
  AND U10907 ( .A(n100), .B(n7055), .Z(n7053) );
  XOR U10908 ( .A(n7056), .B(n7057), .Z(n7055) );
  XOR U10909 ( .A(DB[3213]), .B(DB[3182]), .Z(n7057) );
  AND U10910 ( .A(n104), .B(n7058), .Z(n7056) );
  XOR U10911 ( .A(n7059), .B(n7060), .Z(n7058) );
  XOR U10912 ( .A(DB[3182]), .B(DB[3151]), .Z(n7060) );
  AND U10913 ( .A(n108), .B(n7061), .Z(n7059) );
  XOR U10914 ( .A(n7062), .B(n7063), .Z(n7061) );
  XOR U10915 ( .A(DB[3151]), .B(DB[3120]), .Z(n7063) );
  AND U10916 ( .A(n112), .B(n7064), .Z(n7062) );
  XOR U10917 ( .A(n7065), .B(n7066), .Z(n7064) );
  XOR U10918 ( .A(DB[3120]), .B(DB[3089]), .Z(n7066) );
  AND U10919 ( .A(n116), .B(n7067), .Z(n7065) );
  XOR U10920 ( .A(n7068), .B(n7069), .Z(n7067) );
  XOR U10921 ( .A(DB[3089]), .B(DB[3058]), .Z(n7069) );
  AND U10922 ( .A(n120), .B(n7070), .Z(n7068) );
  XOR U10923 ( .A(n7071), .B(n7072), .Z(n7070) );
  XOR U10924 ( .A(DB[3058]), .B(DB[3027]), .Z(n7072) );
  AND U10925 ( .A(n124), .B(n7073), .Z(n7071) );
  XOR U10926 ( .A(n7074), .B(n7075), .Z(n7073) );
  XOR U10927 ( .A(DB[3027]), .B(DB[2996]), .Z(n7075) );
  AND U10928 ( .A(n128), .B(n7076), .Z(n7074) );
  XOR U10929 ( .A(n7077), .B(n7078), .Z(n7076) );
  XOR U10930 ( .A(DB[2996]), .B(DB[2965]), .Z(n7078) );
  AND U10931 ( .A(n132), .B(n7079), .Z(n7077) );
  XOR U10932 ( .A(n7080), .B(n7081), .Z(n7079) );
  XOR U10933 ( .A(DB[2965]), .B(DB[2934]), .Z(n7081) );
  AND U10934 ( .A(n136), .B(n7082), .Z(n7080) );
  XOR U10935 ( .A(n7083), .B(n7084), .Z(n7082) );
  XOR U10936 ( .A(DB[2934]), .B(DB[2903]), .Z(n7084) );
  AND U10937 ( .A(n140), .B(n7085), .Z(n7083) );
  XOR U10938 ( .A(n7086), .B(n7087), .Z(n7085) );
  XOR U10939 ( .A(DB[2903]), .B(DB[2872]), .Z(n7087) );
  AND U10940 ( .A(n144), .B(n7088), .Z(n7086) );
  XOR U10941 ( .A(n7089), .B(n7090), .Z(n7088) );
  XOR U10942 ( .A(DB[2872]), .B(DB[2841]), .Z(n7090) );
  AND U10943 ( .A(n148), .B(n7091), .Z(n7089) );
  XOR U10944 ( .A(n7092), .B(n7093), .Z(n7091) );
  XOR U10945 ( .A(DB[2841]), .B(DB[2810]), .Z(n7093) );
  AND U10946 ( .A(n152), .B(n7094), .Z(n7092) );
  XOR U10947 ( .A(n7095), .B(n7096), .Z(n7094) );
  XOR U10948 ( .A(DB[2810]), .B(DB[2779]), .Z(n7096) );
  AND U10949 ( .A(n156), .B(n7097), .Z(n7095) );
  XOR U10950 ( .A(n7098), .B(n7099), .Z(n7097) );
  XOR U10951 ( .A(DB[2779]), .B(DB[2748]), .Z(n7099) );
  AND U10952 ( .A(n160), .B(n7100), .Z(n7098) );
  XOR U10953 ( .A(n7101), .B(n7102), .Z(n7100) );
  XOR U10954 ( .A(DB[2748]), .B(DB[2717]), .Z(n7102) );
  AND U10955 ( .A(n164), .B(n7103), .Z(n7101) );
  XOR U10956 ( .A(n7104), .B(n7105), .Z(n7103) );
  XOR U10957 ( .A(DB[2717]), .B(DB[2686]), .Z(n7105) );
  AND U10958 ( .A(n168), .B(n7106), .Z(n7104) );
  XOR U10959 ( .A(n7107), .B(n7108), .Z(n7106) );
  XOR U10960 ( .A(DB[2686]), .B(DB[2655]), .Z(n7108) );
  AND U10961 ( .A(n172), .B(n7109), .Z(n7107) );
  XOR U10962 ( .A(n7110), .B(n7111), .Z(n7109) );
  XOR U10963 ( .A(DB[2655]), .B(DB[2624]), .Z(n7111) );
  AND U10964 ( .A(n176), .B(n7112), .Z(n7110) );
  XOR U10965 ( .A(n7113), .B(n7114), .Z(n7112) );
  XOR U10966 ( .A(DB[2624]), .B(DB[2593]), .Z(n7114) );
  AND U10967 ( .A(n180), .B(n7115), .Z(n7113) );
  XOR U10968 ( .A(n7116), .B(n7117), .Z(n7115) );
  XOR U10969 ( .A(DB[2593]), .B(DB[2562]), .Z(n7117) );
  AND U10970 ( .A(n184), .B(n7118), .Z(n7116) );
  XOR U10971 ( .A(n7119), .B(n7120), .Z(n7118) );
  XOR U10972 ( .A(DB[2562]), .B(DB[2531]), .Z(n7120) );
  AND U10973 ( .A(n188), .B(n7121), .Z(n7119) );
  XOR U10974 ( .A(n7122), .B(n7123), .Z(n7121) );
  XOR U10975 ( .A(DB[2531]), .B(DB[2500]), .Z(n7123) );
  AND U10976 ( .A(n192), .B(n7124), .Z(n7122) );
  XOR U10977 ( .A(n7125), .B(n7126), .Z(n7124) );
  XOR U10978 ( .A(DB[2500]), .B(DB[2469]), .Z(n7126) );
  AND U10979 ( .A(n196), .B(n7127), .Z(n7125) );
  XOR U10980 ( .A(n7128), .B(n7129), .Z(n7127) );
  XOR U10981 ( .A(DB[2469]), .B(DB[2438]), .Z(n7129) );
  AND U10982 ( .A(n200), .B(n7130), .Z(n7128) );
  XOR U10983 ( .A(n7131), .B(n7132), .Z(n7130) );
  XOR U10984 ( .A(DB[2438]), .B(DB[2407]), .Z(n7132) );
  AND U10985 ( .A(n204), .B(n7133), .Z(n7131) );
  XOR U10986 ( .A(n7134), .B(n7135), .Z(n7133) );
  XOR U10987 ( .A(DB[2407]), .B(DB[2376]), .Z(n7135) );
  AND U10988 ( .A(n208), .B(n7136), .Z(n7134) );
  XOR U10989 ( .A(n7137), .B(n7138), .Z(n7136) );
  XOR U10990 ( .A(DB[2376]), .B(DB[2345]), .Z(n7138) );
  AND U10991 ( .A(n212), .B(n7139), .Z(n7137) );
  XOR U10992 ( .A(n7140), .B(n7141), .Z(n7139) );
  XOR U10993 ( .A(DB[2345]), .B(DB[2314]), .Z(n7141) );
  AND U10994 ( .A(n216), .B(n7142), .Z(n7140) );
  XOR U10995 ( .A(n7143), .B(n7144), .Z(n7142) );
  XOR U10996 ( .A(DB[2314]), .B(DB[2283]), .Z(n7144) );
  AND U10997 ( .A(n220), .B(n7145), .Z(n7143) );
  XOR U10998 ( .A(n7146), .B(n7147), .Z(n7145) );
  XOR U10999 ( .A(DB[2283]), .B(DB[2252]), .Z(n7147) );
  AND U11000 ( .A(n224), .B(n7148), .Z(n7146) );
  XOR U11001 ( .A(n7149), .B(n7150), .Z(n7148) );
  XOR U11002 ( .A(DB[2252]), .B(DB[2221]), .Z(n7150) );
  AND U11003 ( .A(n228), .B(n7151), .Z(n7149) );
  XOR U11004 ( .A(n7152), .B(n7153), .Z(n7151) );
  XOR U11005 ( .A(DB[2221]), .B(DB[2190]), .Z(n7153) );
  AND U11006 ( .A(n232), .B(n7154), .Z(n7152) );
  XOR U11007 ( .A(n7155), .B(n7156), .Z(n7154) );
  XOR U11008 ( .A(DB[2190]), .B(DB[2159]), .Z(n7156) );
  AND U11009 ( .A(n236), .B(n7157), .Z(n7155) );
  XOR U11010 ( .A(n7158), .B(n7159), .Z(n7157) );
  XOR U11011 ( .A(DB[2159]), .B(DB[2128]), .Z(n7159) );
  AND U11012 ( .A(n240), .B(n7160), .Z(n7158) );
  XOR U11013 ( .A(n7161), .B(n7162), .Z(n7160) );
  XOR U11014 ( .A(DB[2128]), .B(DB[2097]), .Z(n7162) );
  AND U11015 ( .A(n244), .B(n7163), .Z(n7161) );
  XOR U11016 ( .A(n7164), .B(n7165), .Z(n7163) );
  XOR U11017 ( .A(DB[2097]), .B(DB[2066]), .Z(n7165) );
  AND U11018 ( .A(n248), .B(n7166), .Z(n7164) );
  XOR U11019 ( .A(n7167), .B(n7168), .Z(n7166) );
  XOR U11020 ( .A(DB[2066]), .B(DB[2035]), .Z(n7168) );
  AND U11021 ( .A(n252), .B(n7169), .Z(n7167) );
  XOR U11022 ( .A(n7170), .B(n7171), .Z(n7169) );
  XOR U11023 ( .A(DB[2035]), .B(DB[2004]), .Z(n7171) );
  AND U11024 ( .A(n256), .B(n7172), .Z(n7170) );
  XOR U11025 ( .A(n7173), .B(n7174), .Z(n7172) );
  XOR U11026 ( .A(DB[2004]), .B(DB[1973]), .Z(n7174) );
  AND U11027 ( .A(n260), .B(n7175), .Z(n7173) );
  XOR U11028 ( .A(n7176), .B(n7177), .Z(n7175) );
  XOR U11029 ( .A(DB[1973]), .B(DB[1942]), .Z(n7177) );
  AND U11030 ( .A(n264), .B(n7178), .Z(n7176) );
  XOR U11031 ( .A(n7179), .B(n7180), .Z(n7178) );
  XOR U11032 ( .A(DB[1942]), .B(DB[1911]), .Z(n7180) );
  AND U11033 ( .A(n268), .B(n7181), .Z(n7179) );
  XOR U11034 ( .A(n7182), .B(n7183), .Z(n7181) );
  XOR U11035 ( .A(DB[1911]), .B(DB[1880]), .Z(n7183) );
  AND U11036 ( .A(n272), .B(n7184), .Z(n7182) );
  XOR U11037 ( .A(n7185), .B(n7186), .Z(n7184) );
  XOR U11038 ( .A(DB[1880]), .B(DB[1849]), .Z(n7186) );
  AND U11039 ( .A(n276), .B(n7187), .Z(n7185) );
  XOR U11040 ( .A(n7188), .B(n7189), .Z(n7187) );
  XOR U11041 ( .A(DB[1849]), .B(DB[1818]), .Z(n7189) );
  AND U11042 ( .A(n280), .B(n7190), .Z(n7188) );
  XOR U11043 ( .A(n7191), .B(n7192), .Z(n7190) );
  XOR U11044 ( .A(DB[1818]), .B(DB[1787]), .Z(n7192) );
  AND U11045 ( .A(n284), .B(n7193), .Z(n7191) );
  XOR U11046 ( .A(n7194), .B(n7195), .Z(n7193) );
  XOR U11047 ( .A(DB[1787]), .B(DB[1756]), .Z(n7195) );
  AND U11048 ( .A(n288), .B(n7196), .Z(n7194) );
  XOR U11049 ( .A(n7197), .B(n7198), .Z(n7196) );
  XOR U11050 ( .A(DB[1756]), .B(DB[1725]), .Z(n7198) );
  AND U11051 ( .A(n292), .B(n7199), .Z(n7197) );
  XOR U11052 ( .A(n7200), .B(n7201), .Z(n7199) );
  XOR U11053 ( .A(DB[1725]), .B(DB[1694]), .Z(n7201) );
  AND U11054 ( .A(n296), .B(n7202), .Z(n7200) );
  XOR U11055 ( .A(n7203), .B(n7204), .Z(n7202) );
  XOR U11056 ( .A(DB[1694]), .B(DB[1663]), .Z(n7204) );
  AND U11057 ( .A(n300), .B(n7205), .Z(n7203) );
  XOR U11058 ( .A(n7206), .B(n7207), .Z(n7205) );
  XOR U11059 ( .A(DB[1663]), .B(DB[1632]), .Z(n7207) );
  AND U11060 ( .A(n304), .B(n7208), .Z(n7206) );
  XOR U11061 ( .A(n7209), .B(n7210), .Z(n7208) );
  XOR U11062 ( .A(DB[1632]), .B(DB[1601]), .Z(n7210) );
  AND U11063 ( .A(n308), .B(n7211), .Z(n7209) );
  XOR U11064 ( .A(n7212), .B(n7213), .Z(n7211) );
  XOR U11065 ( .A(DB[1601]), .B(DB[1570]), .Z(n7213) );
  AND U11066 ( .A(n312), .B(n7214), .Z(n7212) );
  XOR U11067 ( .A(n7215), .B(n7216), .Z(n7214) );
  XOR U11068 ( .A(DB[1570]), .B(DB[1539]), .Z(n7216) );
  AND U11069 ( .A(n316), .B(n7217), .Z(n7215) );
  XOR U11070 ( .A(n7218), .B(n7219), .Z(n7217) );
  XOR U11071 ( .A(DB[1539]), .B(DB[1508]), .Z(n7219) );
  AND U11072 ( .A(n320), .B(n7220), .Z(n7218) );
  XOR U11073 ( .A(n7221), .B(n7222), .Z(n7220) );
  XOR U11074 ( .A(DB[1508]), .B(DB[1477]), .Z(n7222) );
  AND U11075 ( .A(n324), .B(n7223), .Z(n7221) );
  XOR U11076 ( .A(n7224), .B(n7225), .Z(n7223) );
  XOR U11077 ( .A(DB[1477]), .B(DB[1446]), .Z(n7225) );
  AND U11078 ( .A(n328), .B(n7226), .Z(n7224) );
  XOR U11079 ( .A(n7227), .B(n7228), .Z(n7226) );
  XOR U11080 ( .A(DB[1446]), .B(DB[1415]), .Z(n7228) );
  AND U11081 ( .A(n332), .B(n7229), .Z(n7227) );
  XOR U11082 ( .A(n7230), .B(n7231), .Z(n7229) );
  XOR U11083 ( .A(DB[1415]), .B(DB[1384]), .Z(n7231) );
  AND U11084 ( .A(n336), .B(n7232), .Z(n7230) );
  XOR U11085 ( .A(n7233), .B(n7234), .Z(n7232) );
  XOR U11086 ( .A(DB[1384]), .B(DB[1353]), .Z(n7234) );
  AND U11087 ( .A(n340), .B(n7235), .Z(n7233) );
  XOR U11088 ( .A(n7236), .B(n7237), .Z(n7235) );
  XOR U11089 ( .A(DB[1353]), .B(DB[1322]), .Z(n7237) );
  AND U11090 ( .A(n344), .B(n7238), .Z(n7236) );
  XOR U11091 ( .A(n7239), .B(n7240), .Z(n7238) );
  XOR U11092 ( .A(DB[1322]), .B(DB[1291]), .Z(n7240) );
  AND U11093 ( .A(n348), .B(n7241), .Z(n7239) );
  XOR U11094 ( .A(n7242), .B(n7243), .Z(n7241) );
  XOR U11095 ( .A(DB[1291]), .B(DB[1260]), .Z(n7243) );
  AND U11096 ( .A(n352), .B(n7244), .Z(n7242) );
  XOR U11097 ( .A(n7245), .B(n7246), .Z(n7244) );
  XOR U11098 ( .A(DB[1260]), .B(DB[1229]), .Z(n7246) );
  AND U11099 ( .A(n356), .B(n7247), .Z(n7245) );
  XOR U11100 ( .A(n7248), .B(n7249), .Z(n7247) );
  XOR U11101 ( .A(DB[1229]), .B(DB[1198]), .Z(n7249) );
  AND U11102 ( .A(n360), .B(n7250), .Z(n7248) );
  XOR U11103 ( .A(n7251), .B(n7252), .Z(n7250) );
  XOR U11104 ( .A(DB[1198]), .B(DB[1167]), .Z(n7252) );
  AND U11105 ( .A(n364), .B(n7253), .Z(n7251) );
  XOR U11106 ( .A(n7254), .B(n7255), .Z(n7253) );
  XOR U11107 ( .A(DB[1167]), .B(DB[1136]), .Z(n7255) );
  AND U11108 ( .A(n368), .B(n7256), .Z(n7254) );
  XOR U11109 ( .A(n7257), .B(n7258), .Z(n7256) );
  XOR U11110 ( .A(DB[1136]), .B(DB[1105]), .Z(n7258) );
  AND U11111 ( .A(n372), .B(n7259), .Z(n7257) );
  XOR U11112 ( .A(n7260), .B(n7261), .Z(n7259) );
  XOR U11113 ( .A(DB[1105]), .B(DB[1074]), .Z(n7261) );
  AND U11114 ( .A(n376), .B(n7262), .Z(n7260) );
  XOR U11115 ( .A(n7263), .B(n7264), .Z(n7262) );
  XOR U11116 ( .A(DB[1074]), .B(DB[1043]), .Z(n7264) );
  AND U11117 ( .A(n380), .B(n7265), .Z(n7263) );
  XOR U11118 ( .A(n7266), .B(n7267), .Z(n7265) );
  XOR U11119 ( .A(DB[1043]), .B(DB[1012]), .Z(n7267) );
  AND U11120 ( .A(n384), .B(n7268), .Z(n7266) );
  XOR U11121 ( .A(n7269), .B(n7270), .Z(n7268) );
  XOR U11122 ( .A(DB[981]), .B(DB[1012]), .Z(n7270) );
  AND U11123 ( .A(n388), .B(n7271), .Z(n7269) );
  XOR U11124 ( .A(n7272), .B(n7273), .Z(n7271) );
  XOR U11125 ( .A(DB[981]), .B(DB[950]), .Z(n7273) );
  AND U11126 ( .A(n392), .B(n7274), .Z(n7272) );
  XOR U11127 ( .A(n7275), .B(n7276), .Z(n7274) );
  XOR U11128 ( .A(DB[950]), .B(DB[919]), .Z(n7276) );
  AND U11129 ( .A(n396), .B(n7277), .Z(n7275) );
  XOR U11130 ( .A(n7278), .B(n7279), .Z(n7277) );
  XOR U11131 ( .A(DB[919]), .B(DB[888]), .Z(n7279) );
  AND U11132 ( .A(n400), .B(n7280), .Z(n7278) );
  XOR U11133 ( .A(n7281), .B(n7282), .Z(n7280) );
  XOR U11134 ( .A(DB[888]), .B(DB[857]), .Z(n7282) );
  AND U11135 ( .A(n404), .B(n7283), .Z(n7281) );
  XOR U11136 ( .A(n7284), .B(n7285), .Z(n7283) );
  XOR U11137 ( .A(DB[857]), .B(DB[826]), .Z(n7285) );
  AND U11138 ( .A(n408), .B(n7286), .Z(n7284) );
  XOR U11139 ( .A(n7287), .B(n7288), .Z(n7286) );
  XOR U11140 ( .A(DB[826]), .B(DB[795]), .Z(n7288) );
  AND U11141 ( .A(n412), .B(n7289), .Z(n7287) );
  XOR U11142 ( .A(n7290), .B(n7291), .Z(n7289) );
  XOR U11143 ( .A(DB[795]), .B(DB[764]), .Z(n7291) );
  AND U11144 ( .A(n416), .B(n7292), .Z(n7290) );
  XOR U11145 ( .A(n7293), .B(n7294), .Z(n7292) );
  XOR U11146 ( .A(DB[764]), .B(DB[733]), .Z(n7294) );
  AND U11147 ( .A(n420), .B(n7295), .Z(n7293) );
  XOR U11148 ( .A(n7296), .B(n7297), .Z(n7295) );
  XOR U11149 ( .A(DB[733]), .B(DB[702]), .Z(n7297) );
  AND U11150 ( .A(n424), .B(n7298), .Z(n7296) );
  XOR U11151 ( .A(n7299), .B(n7300), .Z(n7298) );
  XOR U11152 ( .A(DB[702]), .B(DB[671]), .Z(n7300) );
  AND U11153 ( .A(n428), .B(n7301), .Z(n7299) );
  XOR U11154 ( .A(n7302), .B(n7303), .Z(n7301) );
  XOR U11155 ( .A(DB[671]), .B(DB[640]), .Z(n7303) );
  AND U11156 ( .A(n432), .B(n7304), .Z(n7302) );
  XOR U11157 ( .A(n7305), .B(n7306), .Z(n7304) );
  XOR U11158 ( .A(DB[640]), .B(DB[609]), .Z(n7306) );
  AND U11159 ( .A(n436), .B(n7307), .Z(n7305) );
  XOR U11160 ( .A(n7308), .B(n7309), .Z(n7307) );
  XOR U11161 ( .A(DB[609]), .B(DB[578]), .Z(n7309) );
  AND U11162 ( .A(n440), .B(n7310), .Z(n7308) );
  XOR U11163 ( .A(n7311), .B(n7312), .Z(n7310) );
  XOR U11164 ( .A(DB[578]), .B(DB[547]), .Z(n7312) );
  AND U11165 ( .A(n444), .B(n7313), .Z(n7311) );
  XOR U11166 ( .A(n7314), .B(n7315), .Z(n7313) );
  XOR U11167 ( .A(DB[547]), .B(DB[516]), .Z(n7315) );
  AND U11168 ( .A(n448), .B(n7316), .Z(n7314) );
  XOR U11169 ( .A(n7317), .B(n7318), .Z(n7316) );
  XOR U11170 ( .A(DB[516]), .B(DB[485]), .Z(n7318) );
  AND U11171 ( .A(n452), .B(n7319), .Z(n7317) );
  XOR U11172 ( .A(n7320), .B(n7321), .Z(n7319) );
  XOR U11173 ( .A(DB[485]), .B(DB[454]), .Z(n7321) );
  AND U11174 ( .A(n456), .B(n7322), .Z(n7320) );
  XOR U11175 ( .A(n7323), .B(n7324), .Z(n7322) );
  XOR U11176 ( .A(DB[454]), .B(DB[423]), .Z(n7324) );
  AND U11177 ( .A(n460), .B(n7325), .Z(n7323) );
  XOR U11178 ( .A(n7326), .B(n7327), .Z(n7325) );
  XOR U11179 ( .A(DB[423]), .B(DB[392]), .Z(n7327) );
  AND U11180 ( .A(n464), .B(n7328), .Z(n7326) );
  XOR U11181 ( .A(n7329), .B(n7330), .Z(n7328) );
  XOR U11182 ( .A(DB[392]), .B(DB[361]), .Z(n7330) );
  AND U11183 ( .A(n468), .B(n7331), .Z(n7329) );
  XOR U11184 ( .A(n7332), .B(n7333), .Z(n7331) );
  XOR U11185 ( .A(DB[361]), .B(DB[330]), .Z(n7333) );
  AND U11186 ( .A(n472), .B(n7334), .Z(n7332) );
  XOR U11187 ( .A(n7335), .B(n7336), .Z(n7334) );
  XOR U11188 ( .A(DB[330]), .B(DB[299]), .Z(n7336) );
  AND U11189 ( .A(n476), .B(n7337), .Z(n7335) );
  XOR U11190 ( .A(n7338), .B(n7339), .Z(n7337) );
  XOR U11191 ( .A(DB[299]), .B(DB[268]), .Z(n7339) );
  AND U11192 ( .A(n480), .B(n7340), .Z(n7338) );
  XOR U11193 ( .A(n7341), .B(n7342), .Z(n7340) );
  XOR U11194 ( .A(DB[268]), .B(DB[237]), .Z(n7342) );
  AND U11195 ( .A(n484), .B(n7343), .Z(n7341) );
  XOR U11196 ( .A(n7344), .B(n7345), .Z(n7343) );
  XOR U11197 ( .A(DB[237]), .B(DB[206]), .Z(n7345) );
  AND U11198 ( .A(n488), .B(n7346), .Z(n7344) );
  XOR U11199 ( .A(n7347), .B(n7348), .Z(n7346) );
  XOR U11200 ( .A(DB[206]), .B(DB[175]), .Z(n7348) );
  AND U11201 ( .A(n492), .B(n7349), .Z(n7347) );
  XOR U11202 ( .A(n7350), .B(n7351), .Z(n7349) );
  XOR U11203 ( .A(DB[175]), .B(DB[144]), .Z(n7351) );
  AND U11204 ( .A(n496), .B(n7352), .Z(n7350) );
  XOR U11205 ( .A(n7353), .B(n7354), .Z(n7352) );
  XOR U11206 ( .A(DB[144]), .B(DB[113]), .Z(n7354) );
  AND U11207 ( .A(n500), .B(n7355), .Z(n7353) );
  XOR U11208 ( .A(n7356), .B(n7357), .Z(n7355) );
  XOR U11209 ( .A(DB[82]), .B(DB[113]), .Z(n7357) );
  AND U11210 ( .A(n504), .B(n7358), .Z(n7356) );
  XOR U11211 ( .A(n7359), .B(n7360), .Z(n7358) );
  XOR U11212 ( .A(DB[82]), .B(DB[51]), .Z(n7360) );
  AND U11213 ( .A(n508), .B(n7361), .Z(n7359) );
  XOR U11214 ( .A(DB[51]), .B(DB[20]), .Z(n7361) );
  XOR U11215 ( .A(DB[3938]), .B(n7362), .Z(min_val_out[1]) );
  AND U11216 ( .A(n2), .B(n7363), .Z(n7362) );
  XOR U11217 ( .A(n7364), .B(n7365), .Z(n7363) );
  XOR U11218 ( .A(DB[3938]), .B(DB[3907]), .Z(n7365) );
  AND U11219 ( .A(n8), .B(n7366), .Z(n7364) );
  XOR U11220 ( .A(n7367), .B(n7368), .Z(n7366) );
  XOR U11221 ( .A(DB[3907]), .B(DB[3876]), .Z(n7368) );
  AND U11222 ( .A(n12), .B(n7369), .Z(n7367) );
  XOR U11223 ( .A(n7370), .B(n7371), .Z(n7369) );
  XOR U11224 ( .A(DB[3876]), .B(DB[3845]), .Z(n7371) );
  AND U11225 ( .A(n16), .B(n7372), .Z(n7370) );
  XOR U11226 ( .A(n7373), .B(n7374), .Z(n7372) );
  XOR U11227 ( .A(DB[3845]), .B(DB[3814]), .Z(n7374) );
  AND U11228 ( .A(n20), .B(n7375), .Z(n7373) );
  XOR U11229 ( .A(n7376), .B(n7377), .Z(n7375) );
  XOR U11230 ( .A(DB[3814]), .B(DB[3783]), .Z(n7377) );
  AND U11231 ( .A(n24), .B(n7378), .Z(n7376) );
  XOR U11232 ( .A(n7379), .B(n7380), .Z(n7378) );
  XOR U11233 ( .A(DB[3783]), .B(DB[3752]), .Z(n7380) );
  AND U11234 ( .A(n28), .B(n7381), .Z(n7379) );
  XOR U11235 ( .A(n7382), .B(n7383), .Z(n7381) );
  XOR U11236 ( .A(DB[3752]), .B(DB[3721]), .Z(n7383) );
  AND U11237 ( .A(n32), .B(n7384), .Z(n7382) );
  XOR U11238 ( .A(n7385), .B(n7386), .Z(n7384) );
  XOR U11239 ( .A(DB[3721]), .B(DB[3690]), .Z(n7386) );
  AND U11240 ( .A(n36), .B(n7387), .Z(n7385) );
  XOR U11241 ( .A(n7388), .B(n7389), .Z(n7387) );
  XOR U11242 ( .A(DB[3690]), .B(DB[3659]), .Z(n7389) );
  AND U11243 ( .A(n40), .B(n7390), .Z(n7388) );
  XOR U11244 ( .A(n7391), .B(n7392), .Z(n7390) );
  XOR U11245 ( .A(DB[3659]), .B(DB[3628]), .Z(n7392) );
  AND U11246 ( .A(n44), .B(n7393), .Z(n7391) );
  XOR U11247 ( .A(n7394), .B(n7395), .Z(n7393) );
  XOR U11248 ( .A(DB[3628]), .B(DB[3597]), .Z(n7395) );
  AND U11249 ( .A(n48), .B(n7396), .Z(n7394) );
  XOR U11250 ( .A(n7397), .B(n7398), .Z(n7396) );
  XOR U11251 ( .A(DB[3597]), .B(DB[3566]), .Z(n7398) );
  AND U11252 ( .A(n52), .B(n7399), .Z(n7397) );
  XOR U11253 ( .A(n7400), .B(n7401), .Z(n7399) );
  XOR U11254 ( .A(DB[3566]), .B(DB[3535]), .Z(n7401) );
  AND U11255 ( .A(n56), .B(n7402), .Z(n7400) );
  XOR U11256 ( .A(n7403), .B(n7404), .Z(n7402) );
  XOR U11257 ( .A(DB[3535]), .B(DB[3504]), .Z(n7404) );
  AND U11258 ( .A(n60), .B(n7405), .Z(n7403) );
  XOR U11259 ( .A(n7406), .B(n7407), .Z(n7405) );
  XOR U11260 ( .A(DB[3504]), .B(DB[3473]), .Z(n7407) );
  AND U11261 ( .A(n64), .B(n7408), .Z(n7406) );
  XOR U11262 ( .A(n7409), .B(n7410), .Z(n7408) );
  XOR U11263 ( .A(DB[3473]), .B(DB[3442]), .Z(n7410) );
  AND U11264 ( .A(n68), .B(n7411), .Z(n7409) );
  XOR U11265 ( .A(n7412), .B(n7413), .Z(n7411) );
  XOR U11266 ( .A(DB[3442]), .B(DB[3411]), .Z(n7413) );
  AND U11267 ( .A(n72), .B(n7414), .Z(n7412) );
  XOR U11268 ( .A(n7415), .B(n7416), .Z(n7414) );
  XOR U11269 ( .A(DB[3411]), .B(DB[3380]), .Z(n7416) );
  AND U11270 ( .A(n76), .B(n7417), .Z(n7415) );
  XOR U11271 ( .A(n7418), .B(n7419), .Z(n7417) );
  XOR U11272 ( .A(DB[3380]), .B(DB[3349]), .Z(n7419) );
  AND U11273 ( .A(n80), .B(n7420), .Z(n7418) );
  XOR U11274 ( .A(n7421), .B(n7422), .Z(n7420) );
  XOR U11275 ( .A(DB[3349]), .B(DB[3318]), .Z(n7422) );
  AND U11276 ( .A(n84), .B(n7423), .Z(n7421) );
  XOR U11277 ( .A(n7424), .B(n7425), .Z(n7423) );
  XOR U11278 ( .A(DB[3318]), .B(DB[3287]), .Z(n7425) );
  AND U11279 ( .A(n88), .B(n7426), .Z(n7424) );
  XOR U11280 ( .A(n7427), .B(n7428), .Z(n7426) );
  XOR U11281 ( .A(DB[3287]), .B(DB[3256]), .Z(n7428) );
  AND U11282 ( .A(n92), .B(n7429), .Z(n7427) );
  XOR U11283 ( .A(n7430), .B(n7431), .Z(n7429) );
  XOR U11284 ( .A(DB[3256]), .B(DB[3225]), .Z(n7431) );
  AND U11285 ( .A(n96), .B(n7432), .Z(n7430) );
  XOR U11286 ( .A(n7433), .B(n7434), .Z(n7432) );
  XOR U11287 ( .A(DB[3225]), .B(DB[3194]), .Z(n7434) );
  AND U11288 ( .A(n100), .B(n7435), .Z(n7433) );
  XOR U11289 ( .A(n7436), .B(n7437), .Z(n7435) );
  XOR U11290 ( .A(DB[3194]), .B(DB[3163]), .Z(n7437) );
  AND U11291 ( .A(n104), .B(n7438), .Z(n7436) );
  XOR U11292 ( .A(n7439), .B(n7440), .Z(n7438) );
  XOR U11293 ( .A(DB[3163]), .B(DB[3132]), .Z(n7440) );
  AND U11294 ( .A(n108), .B(n7441), .Z(n7439) );
  XOR U11295 ( .A(n7442), .B(n7443), .Z(n7441) );
  XOR U11296 ( .A(DB[3132]), .B(DB[3101]), .Z(n7443) );
  AND U11297 ( .A(n112), .B(n7444), .Z(n7442) );
  XOR U11298 ( .A(n7445), .B(n7446), .Z(n7444) );
  XOR U11299 ( .A(DB[3101]), .B(DB[3070]), .Z(n7446) );
  AND U11300 ( .A(n116), .B(n7447), .Z(n7445) );
  XOR U11301 ( .A(n7448), .B(n7449), .Z(n7447) );
  XOR U11302 ( .A(DB[3070]), .B(DB[3039]), .Z(n7449) );
  AND U11303 ( .A(n120), .B(n7450), .Z(n7448) );
  XOR U11304 ( .A(n7451), .B(n7452), .Z(n7450) );
  XOR U11305 ( .A(DB[3039]), .B(DB[3008]), .Z(n7452) );
  AND U11306 ( .A(n124), .B(n7453), .Z(n7451) );
  XOR U11307 ( .A(n7454), .B(n7455), .Z(n7453) );
  XOR U11308 ( .A(DB[3008]), .B(DB[2977]), .Z(n7455) );
  AND U11309 ( .A(n128), .B(n7456), .Z(n7454) );
  XOR U11310 ( .A(n7457), .B(n7458), .Z(n7456) );
  XOR U11311 ( .A(DB[2977]), .B(DB[2946]), .Z(n7458) );
  AND U11312 ( .A(n132), .B(n7459), .Z(n7457) );
  XOR U11313 ( .A(n7460), .B(n7461), .Z(n7459) );
  XOR U11314 ( .A(DB[2946]), .B(DB[2915]), .Z(n7461) );
  AND U11315 ( .A(n136), .B(n7462), .Z(n7460) );
  XOR U11316 ( .A(n7463), .B(n7464), .Z(n7462) );
  XOR U11317 ( .A(DB[2915]), .B(DB[2884]), .Z(n7464) );
  AND U11318 ( .A(n140), .B(n7465), .Z(n7463) );
  XOR U11319 ( .A(n7466), .B(n7467), .Z(n7465) );
  XOR U11320 ( .A(DB[2884]), .B(DB[2853]), .Z(n7467) );
  AND U11321 ( .A(n144), .B(n7468), .Z(n7466) );
  XOR U11322 ( .A(n7469), .B(n7470), .Z(n7468) );
  XOR U11323 ( .A(DB[2853]), .B(DB[2822]), .Z(n7470) );
  AND U11324 ( .A(n148), .B(n7471), .Z(n7469) );
  XOR U11325 ( .A(n7472), .B(n7473), .Z(n7471) );
  XOR U11326 ( .A(DB[2822]), .B(DB[2791]), .Z(n7473) );
  AND U11327 ( .A(n152), .B(n7474), .Z(n7472) );
  XOR U11328 ( .A(n7475), .B(n7476), .Z(n7474) );
  XOR U11329 ( .A(DB[2791]), .B(DB[2760]), .Z(n7476) );
  AND U11330 ( .A(n156), .B(n7477), .Z(n7475) );
  XOR U11331 ( .A(n7478), .B(n7479), .Z(n7477) );
  XOR U11332 ( .A(DB[2760]), .B(DB[2729]), .Z(n7479) );
  AND U11333 ( .A(n160), .B(n7480), .Z(n7478) );
  XOR U11334 ( .A(n7481), .B(n7482), .Z(n7480) );
  XOR U11335 ( .A(DB[2729]), .B(DB[2698]), .Z(n7482) );
  AND U11336 ( .A(n164), .B(n7483), .Z(n7481) );
  XOR U11337 ( .A(n7484), .B(n7485), .Z(n7483) );
  XOR U11338 ( .A(DB[2698]), .B(DB[2667]), .Z(n7485) );
  AND U11339 ( .A(n168), .B(n7486), .Z(n7484) );
  XOR U11340 ( .A(n7487), .B(n7488), .Z(n7486) );
  XOR U11341 ( .A(DB[2667]), .B(DB[2636]), .Z(n7488) );
  AND U11342 ( .A(n172), .B(n7489), .Z(n7487) );
  XOR U11343 ( .A(n7490), .B(n7491), .Z(n7489) );
  XOR U11344 ( .A(DB[2636]), .B(DB[2605]), .Z(n7491) );
  AND U11345 ( .A(n176), .B(n7492), .Z(n7490) );
  XOR U11346 ( .A(n7493), .B(n7494), .Z(n7492) );
  XOR U11347 ( .A(DB[2605]), .B(DB[2574]), .Z(n7494) );
  AND U11348 ( .A(n180), .B(n7495), .Z(n7493) );
  XOR U11349 ( .A(n7496), .B(n7497), .Z(n7495) );
  XOR U11350 ( .A(DB[2574]), .B(DB[2543]), .Z(n7497) );
  AND U11351 ( .A(n184), .B(n7498), .Z(n7496) );
  XOR U11352 ( .A(n7499), .B(n7500), .Z(n7498) );
  XOR U11353 ( .A(DB[2543]), .B(DB[2512]), .Z(n7500) );
  AND U11354 ( .A(n188), .B(n7501), .Z(n7499) );
  XOR U11355 ( .A(n7502), .B(n7503), .Z(n7501) );
  XOR U11356 ( .A(DB[2512]), .B(DB[2481]), .Z(n7503) );
  AND U11357 ( .A(n192), .B(n7504), .Z(n7502) );
  XOR U11358 ( .A(n7505), .B(n7506), .Z(n7504) );
  XOR U11359 ( .A(DB[2481]), .B(DB[2450]), .Z(n7506) );
  AND U11360 ( .A(n196), .B(n7507), .Z(n7505) );
  XOR U11361 ( .A(n7508), .B(n7509), .Z(n7507) );
  XOR U11362 ( .A(DB[2450]), .B(DB[2419]), .Z(n7509) );
  AND U11363 ( .A(n200), .B(n7510), .Z(n7508) );
  XOR U11364 ( .A(n7511), .B(n7512), .Z(n7510) );
  XOR U11365 ( .A(DB[2419]), .B(DB[2388]), .Z(n7512) );
  AND U11366 ( .A(n204), .B(n7513), .Z(n7511) );
  XOR U11367 ( .A(n7514), .B(n7515), .Z(n7513) );
  XOR U11368 ( .A(DB[2388]), .B(DB[2357]), .Z(n7515) );
  AND U11369 ( .A(n208), .B(n7516), .Z(n7514) );
  XOR U11370 ( .A(n7517), .B(n7518), .Z(n7516) );
  XOR U11371 ( .A(DB[2357]), .B(DB[2326]), .Z(n7518) );
  AND U11372 ( .A(n212), .B(n7519), .Z(n7517) );
  XOR U11373 ( .A(n7520), .B(n7521), .Z(n7519) );
  XOR U11374 ( .A(DB[2326]), .B(DB[2295]), .Z(n7521) );
  AND U11375 ( .A(n216), .B(n7522), .Z(n7520) );
  XOR U11376 ( .A(n7523), .B(n7524), .Z(n7522) );
  XOR U11377 ( .A(DB[2295]), .B(DB[2264]), .Z(n7524) );
  AND U11378 ( .A(n220), .B(n7525), .Z(n7523) );
  XOR U11379 ( .A(n7526), .B(n7527), .Z(n7525) );
  XOR U11380 ( .A(DB[2264]), .B(DB[2233]), .Z(n7527) );
  AND U11381 ( .A(n224), .B(n7528), .Z(n7526) );
  XOR U11382 ( .A(n7529), .B(n7530), .Z(n7528) );
  XOR U11383 ( .A(DB[2233]), .B(DB[2202]), .Z(n7530) );
  AND U11384 ( .A(n228), .B(n7531), .Z(n7529) );
  XOR U11385 ( .A(n7532), .B(n7533), .Z(n7531) );
  XOR U11386 ( .A(DB[2202]), .B(DB[2171]), .Z(n7533) );
  AND U11387 ( .A(n232), .B(n7534), .Z(n7532) );
  XOR U11388 ( .A(n7535), .B(n7536), .Z(n7534) );
  XOR U11389 ( .A(DB[2171]), .B(DB[2140]), .Z(n7536) );
  AND U11390 ( .A(n236), .B(n7537), .Z(n7535) );
  XOR U11391 ( .A(n7538), .B(n7539), .Z(n7537) );
  XOR U11392 ( .A(DB[2140]), .B(DB[2109]), .Z(n7539) );
  AND U11393 ( .A(n240), .B(n7540), .Z(n7538) );
  XOR U11394 ( .A(n7541), .B(n7542), .Z(n7540) );
  XOR U11395 ( .A(DB[2109]), .B(DB[2078]), .Z(n7542) );
  AND U11396 ( .A(n244), .B(n7543), .Z(n7541) );
  XOR U11397 ( .A(n7544), .B(n7545), .Z(n7543) );
  XOR U11398 ( .A(DB[2078]), .B(DB[2047]), .Z(n7545) );
  AND U11399 ( .A(n248), .B(n7546), .Z(n7544) );
  XOR U11400 ( .A(n7547), .B(n7548), .Z(n7546) );
  XOR U11401 ( .A(DB[2047]), .B(DB[2016]), .Z(n7548) );
  AND U11402 ( .A(n252), .B(n7549), .Z(n7547) );
  XOR U11403 ( .A(n7550), .B(n7551), .Z(n7549) );
  XOR U11404 ( .A(DB[2016]), .B(DB[1985]), .Z(n7551) );
  AND U11405 ( .A(n256), .B(n7552), .Z(n7550) );
  XOR U11406 ( .A(n7553), .B(n7554), .Z(n7552) );
  XOR U11407 ( .A(DB[1985]), .B(DB[1954]), .Z(n7554) );
  AND U11408 ( .A(n260), .B(n7555), .Z(n7553) );
  XOR U11409 ( .A(n7556), .B(n7557), .Z(n7555) );
  XOR U11410 ( .A(DB[1954]), .B(DB[1923]), .Z(n7557) );
  AND U11411 ( .A(n264), .B(n7558), .Z(n7556) );
  XOR U11412 ( .A(n7559), .B(n7560), .Z(n7558) );
  XOR U11413 ( .A(DB[1923]), .B(DB[1892]), .Z(n7560) );
  AND U11414 ( .A(n268), .B(n7561), .Z(n7559) );
  XOR U11415 ( .A(n7562), .B(n7563), .Z(n7561) );
  XOR U11416 ( .A(DB[1892]), .B(DB[1861]), .Z(n7563) );
  AND U11417 ( .A(n272), .B(n7564), .Z(n7562) );
  XOR U11418 ( .A(n7565), .B(n7566), .Z(n7564) );
  XOR U11419 ( .A(DB[1861]), .B(DB[1830]), .Z(n7566) );
  AND U11420 ( .A(n276), .B(n7567), .Z(n7565) );
  XOR U11421 ( .A(n7568), .B(n7569), .Z(n7567) );
  XOR U11422 ( .A(DB[1830]), .B(DB[1799]), .Z(n7569) );
  AND U11423 ( .A(n280), .B(n7570), .Z(n7568) );
  XOR U11424 ( .A(n7571), .B(n7572), .Z(n7570) );
  XOR U11425 ( .A(DB[1799]), .B(DB[1768]), .Z(n7572) );
  AND U11426 ( .A(n284), .B(n7573), .Z(n7571) );
  XOR U11427 ( .A(n7574), .B(n7575), .Z(n7573) );
  XOR U11428 ( .A(DB[1768]), .B(DB[1737]), .Z(n7575) );
  AND U11429 ( .A(n288), .B(n7576), .Z(n7574) );
  XOR U11430 ( .A(n7577), .B(n7578), .Z(n7576) );
  XOR U11431 ( .A(DB[1737]), .B(DB[1706]), .Z(n7578) );
  AND U11432 ( .A(n292), .B(n7579), .Z(n7577) );
  XOR U11433 ( .A(n7580), .B(n7581), .Z(n7579) );
  XOR U11434 ( .A(DB[1706]), .B(DB[1675]), .Z(n7581) );
  AND U11435 ( .A(n296), .B(n7582), .Z(n7580) );
  XOR U11436 ( .A(n7583), .B(n7584), .Z(n7582) );
  XOR U11437 ( .A(DB[1675]), .B(DB[1644]), .Z(n7584) );
  AND U11438 ( .A(n300), .B(n7585), .Z(n7583) );
  XOR U11439 ( .A(n7586), .B(n7587), .Z(n7585) );
  XOR U11440 ( .A(DB[1644]), .B(DB[1613]), .Z(n7587) );
  AND U11441 ( .A(n304), .B(n7588), .Z(n7586) );
  XOR U11442 ( .A(n7589), .B(n7590), .Z(n7588) );
  XOR U11443 ( .A(DB[1613]), .B(DB[1582]), .Z(n7590) );
  AND U11444 ( .A(n308), .B(n7591), .Z(n7589) );
  XOR U11445 ( .A(n7592), .B(n7593), .Z(n7591) );
  XOR U11446 ( .A(DB[1582]), .B(DB[1551]), .Z(n7593) );
  AND U11447 ( .A(n312), .B(n7594), .Z(n7592) );
  XOR U11448 ( .A(n7595), .B(n7596), .Z(n7594) );
  XOR U11449 ( .A(DB[1551]), .B(DB[1520]), .Z(n7596) );
  AND U11450 ( .A(n316), .B(n7597), .Z(n7595) );
  XOR U11451 ( .A(n7598), .B(n7599), .Z(n7597) );
  XOR U11452 ( .A(DB[1520]), .B(DB[1489]), .Z(n7599) );
  AND U11453 ( .A(n320), .B(n7600), .Z(n7598) );
  XOR U11454 ( .A(n7601), .B(n7602), .Z(n7600) );
  XOR U11455 ( .A(DB[1489]), .B(DB[1458]), .Z(n7602) );
  AND U11456 ( .A(n324), .B(n7603), .Z(n7601) );
  XOR U11457 ( .A(n7604), .B(n7605), .Z(n7603) );
  XOR U11458 ( .A(DB[1458]), .B(DB[1427]), .Z(n7605) );
  AND U11459 ( .A(n328), .B(n7606), .Z(n7604) );
  XOR U11460 ( .A(n7607), .B(n7608), .Z(n7606) );
  XOR U11461 ( .A(DB[1427]), .B(DB[1396]), .Z(n7608) );
  AND U11462 ( .A(n332), .B(n7609), .Z(n7607) );
  XOR U11463 ( .A(n7610), .B(n7611), .Z(n7609) );
  XOR U11464 ( .A(DB[1396]), .B(DB[1365]), .Z(n7611) );
  AND U11465 ( .A(n336), .B(n7612), .Z(n7610) );
  XOR U11466 ( .A(n7613), .B(n7614), .Z(n7612) );
  XOR U11467 ( .A(DB[1365]), .B(DB[1334]), .Z(n7614) );
  AND U11468 ( .A(n340), .B(n7615), .Z(n7613) );
  XOR U11469 ( .A(n7616), .B(n7617), .Z(n7615) );
  XOR U11470 ( .A(DB[1334]), .B(DB[1303]), .Z(n7617) );
  AND U11471 ( .A(n344), .B(n7618), .Z(n7616) );
  XOR U11472 ( .A(n7619), .B(n7620), .Z(n7618) );
  XOR U11473 ( .A(DB[1303]), .B(DB[1272]), .Z(n7620) );
  AND U11474 ( .A(n348), .B(n7621), .Z(n7619) );
  XOR U11475 ( .A(n7622), .B(n7623), .Z(n7621) );
  XOR U11476 ( .A(DB[1272]), .B(DB[1241]), .Z(n7623) );
  AND U11477 ( .A(n352), .B(n7624), .Z(n7622) );
  XOR U11478 ( .A(n7625), .B(n7626), .Z(n7624) );
  XOR U11479 ( .A(DB[1241]), .B(DB[1210]), .Z(n7626) );
  AND U11480 ( .A(n356), .B(n7627), .Z(n7625) );
  XOR U11481 ( .A(n7628), .B(n7629), .Z(n7627) );
  XOR U11482 ( .A(DB[1210]), .B(DB[1179]), .Z(n7629) );
  AND U11483 ( .A(n360), .B(n7630), .Z(n7628) );
  XOR U11484 ( .A(n7631), .B(n7632), .Z(n7630) );
  XOR U11485 ( .A(DB[1179]), .B(DB[1148]), .Z(n7632) );
  AND U11486 ( .A(n364), .B(n7633), .Z(n7631) );
  XOR U11487 ( .A(n7634), .B(n7635), .Z(n7633) );
  XOR U11488 ( .A(DB[1148]), .B(DB[1117]), .Z(n7635) );
  AND U11489 ( .A(n368), .B(n7636), .Z(n7634) );
  XOR U11490 ( .A(n7637), .B(n7638), .Z(n7636) );
  XOR U11491 ( .A(DB[1117]), .B(DB[1086]), .Z(n7638) );
  AND U11492 ( .A(n372), .B(n7639), .Z(n7637) );
  XOR U11493 ( .A(n7640), .B(n7641), .Z(n7639) );
  XOR U11494 ( .A(DB[1086]), .B(DB[1055]), .Z(n7641) );
  AND U11495 ( .A(n376), .B(n7642), .Z(n7640) );
  XOR U11496 ( .A(n7643), .B(n7644), .Z(n7642) );
  XOR U11497 ( .A(DB[1055]), .B(DB[1024]), .Z(n7644) );
  AND U11498 ( .A(n380), .B(n7645), .Z(n7643) );
  XOR U11499 ( .A(n7646), .B(n7647), .Z(n7645) );
  XOR U11500 ( .A(DB[993]), .B(DB[1024]), .Z(n7647) );
  AND U11501 ( .A(n384), .B(n7648), .Z(n7646) );
  XOR U11502 ( .A(n7649), .B(n7650), .Z(n7648) );
  XOR U11503 ( .A(DB[993]), .B(DB[962]), .Z(n7650) );
  AND U11504 ( .A(n388), .B(n7651), .Z(n7649) );
  XOR U11505 ( .A(n7652), .B(n7653), .Z(n7651) );
  XOR U11506 ( .A(DB[962]), .B(DB[931]), .Z(n7653) );
  AND U11507 ( .A(n392), .B(n7654), .Z(n7652) );
  XOR U11508 ( .A(n7655), .B(n7656), .Z(n7654) );
  XOR U11509 ( .A(DB[931]), .B(DB[900]), .Z(n7656) );
  AND U11510 ( .A(n396), .B(n7657), .Z(n7655) );
  XOR U11511 ( .A(n7658), .B(n7659), .Z(n7657) );
  XOR U11512 ( .A(DB[900]), .B(DB[869]), .Z(n7659) );
  AND U11513 ( .A(n400), .B(n7660), .Z(n7658) );
  XOR U11514 ( .A(n7661), .B(n7662), .Z(n7660) );
  XOR U11515 ( .A(DB[869]), .B(DB[838]), .Z(n7662) );
  AND U11516 ( .A(n404), .B(n7663), .Z(n7661) );
  XOR U11517 ( .A(n7664), .B(n7665), .Z(n7663) );
  XOR U11518 ( .A(DB[838]), .B(DB[807]), .Z(n7665) );
  AND U11519 ( .A(n408), .B(n7666), .Z(n7664) );
  XOR U11520 ( .A(n7667), .B(n7668), .Z(n7666) );
  XOR U11521 ( .A(DB[807]), .B(DB[776]), .Z(n7668) );
  AND U11522 ( .A(n412), .B(n7669), .Z(n7667) );
  XOR U11523 ( .A(n7670), .B(n7671), .Z(n7669) );
  XOR U11524 ( .A(DB[776]), .B(DB[745]), .Z(n7671) );
  AND U11525 ( .A(n416), .B(n7672), .Z(n7670) );
  XOR U11526 ( .A(n7673), .B(n7674), .Z(n7672) );
  XOR U11527 ( .A(DB[745]), .B(DB[714]), .Z(n7674) );
  AND U11528 ( .A(n420), .B(n7675), .Z(n7673) );
  XOR U11529 ( .A(n7676), .B(n7677), .Z(n7675) );
  XOR U11530 ( .A(DB[714]), .B(DB[683]), .Z(n7677) );
  AND U11531 ( .A(n424), .B(n7678), .Z(n7676) );
  XOR U11532 ( .A(n7679), .B(n7680), .Z(n7678) );
  XOR U11533 ( .A(DB[683]), .B(DB[652]), .Z(n7680) );
  AND U11534 ( .A(n428), .B(n7681), .Z(n7679) );
  XOR U11535 ( .A(n7682), .B(n7683), .Z(n7681) );
  XOR U11536 ( .A(DB[652]), .B(DB[621]), .Z(n7683) );
  AND U11537 ( .A(n432), .B(n7684), .Z(n7682) );
  XOR U11538 ( .A(n7685), .B(n7686), .Z(n7684) );
  XOR U11539 ( .A(DB[621]), .B(DB[590]), .Z(n7686) );
  AND U11540 ( .A(n436), .B(n7687), .Z(n7685) );
  XOR U11541 ( .A(n7688), .B(n7689), .Z(n7687) );
  XOR U11542 ( .A(DB[590]), .B(DB[559]), .Z(n7689) );
  AND U11543 ( .A(n440), .B(n7690), .Z(n7688) );
  XOR U11544 ( .A(n7691), .B(n7692), .Z(n7690) );
  XOR U11545 ( .A(DB[559]), .B(DB[528]), .Z(n7692) );
  AND U11546 ( .A(n444), .B(n7693), .Z(n7691) );
  XOR U11547 ( .A(n7694), .B(n7695), .Z(n7693) );
  XOR U11548 ( .A(DB[528]), .B(DB[497]), .Z(n7695) );
  AND U11549 ( .A(n448), .B(n7696), .Z(n7694) );
  XOR U11550 ( .A(n7697), .B(n7698), .Z(n7696) );
  XOR U11551 ( .A(DB[497]), .B(DB[466]), .Z(n7698) );
  AND U11552 ( .A(n452), .B(n7699), .Z(n7697) );
  XOR U11553 ( .A(n7700), .B(n7701), .Z(n7699) );
  XOR U11554 ( .A(DB[466]), .B(DB[435]), .Z(n7701) );
  AND U11555 ( .A(n456), .B(n7702), .Z(n7700) );
  XOR U11556 ( .A(n7703), .B(n7704), .Z(n7702) );
  XOR U11557 ( .A(DB[435]), .B(DB[404]), .Z(n7704) );
  AND U11558 ( .A(n460), .B(n7705), .Z(n7703) );
  XOR U11559 ( .A(n7706), .B(n7707), .Z(n7705) );
  XOR U11560 ( .A(DB[404]), .B(DB[373]), .Z(n7707) );
  AND U11561 ( .A(n464), .B(n7708), .Z(n7706) );
  XOR U11562 ( .A(n7709), .B(n7710), .Z(n7708) );
  XOR U11563 ( .A(DB[373]), .B(DB[342]), .Z(n7710) );
  AND U11564 ( .A(n468), .B(n7711), .Z(n7709) );
  XOR U11565 ( .A(n7712), .B(n7713), .Z(n7711) );
  XOR U11566 ( .A(DB[342]), .B(DB[311]), .Z(n7713) );
  AND U11567 ( .A(n472), .B(n7714), .Z(n7712) );
  XOR U11568 ( .A(n7715), .B(n7716), .Z(n7714) );
  XOR U11569 ( .A(DB[311]), .B(DB[280]), .Z(n7716) );
  AND U11570 ( .A(n476), .B(n7717), .Z(n7715) );
  XOR U11571 ( .A(n7718), .B(n7719), .Z(n7717) );
  XOR U11572 ( .A(DB[280]), .B(DB[249]), .Z(n7719) );
  AND U11573 ( .A(n480), .B(n7720), .Z(n7718) );
  XOR U11574 ( .A(n7721), .B(n7722), .Z(n7720) );
  XOR U11575 ( .A(DB[249]), .B(DB[218]), .Z(n7722) );
  AND U11576 ( .A(n484), .B(n7723), .Z(n7721) );
  XOR U11577 ( .A(n7724), .B(n7725), .Z(n7723) );
  XOR U11578 ( .A(DB[218]), .B(DB[187]), .Z(n7725) );
  AND U11579 ( .A(n488), .B(n7726), .Z(n7724) );
  XOR U11580 ( .A(n7727), .B(n7728), .Z(n7726) );
  XOR U11581 ( .A(DB[187]), .B(DB[156]), .Z(n7728) );
  AND U11582 ( .A(n492), .B(n7729), .Z(n7727) );
  XOR U11583 ( .A(n7730), .B(n7731), .Z(n7729) );
  XOR U11584 ( .A(DB[156]), .B(DB[125]), .Z(n7731) );
  AND U11585 ( .A(n496), .B(n7732), .Z(n7730) );
  XOR U11586 ( .A(n7733), .B(n7734), .Z(n7732) );
  XOR U11587 ( .A(DB[94]), .B(DB[125]), .Z(n7734) );
  AND U11588 ( .A(n500), .B(n7735), .Z(n7733) );
  XOR U11589 ( .A(n7736), .B(n7737), .Z(n7735) );
  XOR U11590 ( .A(DB[94]), .B(DB[63]), .Z(n7737) );
  AND U11591 ( .A(n504), .B(n7738), .Z(n7736) );
  XOR U11592 ( .A(n7739), .B(n7740), .Z(n7738) );
  XOR U11593 ( .A(DB[63]), .B(DB[32]), .Z(n7740) );
  AND U11594 ( .A(n508), .B(n7741), .Z(n7739) );
  XOR U11595 ( .A(DB[32]), .B(DB[1]), .Z(n7741) );
  XOR U11596 ( .A(DB[3956]), .B(n7742), .Z(min_val_out[19]) );
  AND U11597 ( .A(n2), .B(n7743), .Z(n7742) );
  XOR U11598 ( .A(n7744), .B(n7745), .Z(n7743) );
  XOR U11599 ( .A(DB[3956]), .B(DB[3925]), .Z(n7745) );
  AND U11600 ( .A(n8), .B(n7746), .Z(n7744) );
  XOR U11601 ( .A(n7747), .B(n7748), .Z(n7746) );
  XOR U11602 ( .A(DB[3925]), .B(DB[3894]), .Z(n7748) );
  AND U11603 ( .A(n12), .B(n7749), .Z(n7747) );
  XOR U11604 ( .A(n7750), .B(n7751), .Z(n7749) );
  XOR U11605 ( .A(DB[3894]), .B(DB[3863]), .Z(n7751) );
  AND U11606 ( .A(n16), .B(n7752), .Z(n7750) );
  XOR U11607 ( .A(n7753), .B(n7754), .Z(n7752) );
  XOR U11608 ( .A(DB[3863]), .B(DB[3832]), .Z(n7754) );
  AND U11609 ( .A(n20), .B(n7755), .Z(n7753) );
  XOR U11610 ( .A(n7756), .B(n7757), .Z(n7755) );
  XOR U11611 ( .A(DB[3832]), .B(DB[3801]), .Z(n7757) );
  AND U11612 ( .A(n24), .B(n7758), .Z(n7756) );
  XOR U11613 ( .A(n7759), .B(n7760), .Z(n7758) );
  XOR U11614 ( .A(DB[3801]), .B(DB[3770]), .Z(n7760) );
  AND U11615 ( .A(n28), .B(n7761), .Z(n7759) );
  XOR U11616 ( .A(n7762), .B(n7763), .Z(n7761) );
  XOR U11617 ( .A(DB[3770]), .B(DB[3739]), .Z(n7763) );
  AND U11618 ( .A(n32), .B(n7764), .Z(n7762) );
  XOR U11619 ( .A(n7765), .B(n7766), .Z(n7764) );
  XOR U11620 ( .A(DB[3739]), .B(DB[3708]), .Z(n7766) );
  AND U11621 ( .A(n36), .B(n7767), .Z(n7765) );
  XOR U11622 ( .A(n7768), .B(n7769), .Z(n7767) );
  XOR U11623 ( .A(DB[3708]), .B(DB[3677]), .Z(n7769) );
  AND U11624 ( .A(n40), .B(n7770), .Z(n7768) );
  XOR U11625 ( .A(n7771), .B(n7772), .Z(n7770) );
  XOR U11626 ( .A(DB[3677]), .B(DB[3646]), .Z(n7772) );
  AND U11627 ( .A(n44), .B(n7773), .Z(n7771) );
  XOR U11628 ( .A(n7774), .B(n7775), .Z(n7773) );
  XOR U11629 ( .A(DB[3646]), .B(DB[3615]), .Z(n7775) );
  AND U11630 ( .A(n48), .B(n7776), .Z(n7774) );
  XOR U11631 ( .A(n7777), .B(n7778), .Z(n7776) );
  XOR U11632 ( .A(DB[3615]), .B(DB[3584]), .Z(n7778) );
  AND U11633 ( .A(n52), .B(n7779), .Z(n7777) );
  XOR U11634 ( .A(n7780), .B(n7781), .Z(n7779) );
  XOR U11635 ( .A(DB[3584]), .B(DB[3553]), .Z(n7781) );
  AND U11636 ( .A(n56), .B(n7782), .Z(n7780) );
  XOR U11637 ( .A(n7783), .B(n7784), .Z(n7782) );
  XOR U11638 ( .A(DB[3553]), .B(DB[3522]), .Z(n7784) );
  AND U11639 ( .A(n60), .B(n7785), .Z(n7783) );
  XOR U11640 ( .A(n7786), .B(n7787), .Z(n7785) );
  XOR U11641 ( .A(DB[3522]), .B(DB[3491]), .Z(n7787) );
  AND U11642 ( .A(n64), .B(n7788), .Z(n7786) );
  XOR U11643 ( .A(n7789), .B(n7790), .Z(n7788) );
  XOR U11644 ( .A(DB[3491]), .B(DB[3460]), .Z(n7790) );
  AND U11645 ( .A(n68), .B(n7791), .Z(n7789) );
  XOR U11646 ( .A(n7792), .B(n7793), .Z(n7791) );
  XOR U11647 ( .A(DB[3460]), .B(DB[3429]), .Z(n7793) );
  AND U11648 ( .A(n72), .B(n7794), .Z(n7792) );
  XOR U11649 ( .A(n7795), .B(n7796), .Z(n7794) );
  XOR U11650 ( .A(DB[3429]), .B(DB[3398]), .Z(n7796) );
  AND U11651 ( .A(n76), .B(n7797), .Z(n7795) );
  XOR U11652 ( .A(n7798), .B(n7799), .Z(n7797) );
  XOR U11653 ( .A(DB[3398]), .B(DB[3367]), .Z(n7799) );
  AND U11654 ( .A(n80), .B(n7800), .Z(n7798) );
  XOR U11655 ( .A(n7801), .B(n7802), .Z(n7800) );
  XOR U11656 ( .A(DB[3367]), .B(DB[3336]), .Z(n7802) );
  AND U11657 ( .A(n84), .B(n7803), .Z(n7801) );
  XOR U11658 ( .A(n7804), .B(n7805), .Z(n7803) );
  XOR U11659 ( .A(DB[3336]), .B(DB[3305]), .Z(n7805) );
  AND U11660 ( .A(n88), .B(n7806), .Z(n7804) );
  XOR U11661 ( .A(n7807), .B(n7808), .Z(n7806) );
  XOR U11662 ( .A(DB[3305]), .B(DB[3274]), .Z(n7808) );
  AND U11663 ( .A(n92), .B(n7809), .Z(n7807) );
  XOR U11664 ( .A(n7810), .B(n7811), .Z(n7809) );
  XOR U11665 ( .A(DB[3274]), .B(DB[3243]), .Z(n7811) );
  AND U11666 ( .A(n96), .B(n7812), .Z(n7810) );
  XOR U11667 ( .A(n7813), .B(n7814), .Z(n7812) );
  XOR U11668 ( .A(DB[3243]), .B(DB[3212]), .Z(n7814) );
  AND U11669 ( .A(n100), .B(n7815), .Z(n7813) );
  XOR U11670 ( .A(n7816), .B(n7817), .Z(n7815) );
  XOR U11671 ( .A(DB[3212]), .B(DB[3181]), .Z(n7817) );
  AND U11672 ( .A(n104), .B(n7818), .Z(n7816) );
  XOR U11673 ( .A(n7819), .B(n7820), .Z(n7818) );
  XOR U11674 ( .A(DB[3181]), .B(DB[3150]), .Z(n7820) );
  AND U11675 ( .A(n108), .B(n7821), .Z(n7819) );
  XOR U11676 ( .A(n7822), .B(n7823), .Z(n7821) );
  XOR U11677 ( .A(DB[3150]), .B(DB[3119]), .Z(n7823) );
  AND U11678 ( .A(n112), .B(n7824), .Z(n7822) );
  XOR U11679 ( .A(n7825), .B(n7826), .Z(n7824) );
  XOR U11680 ( .A(DB[3119]), .B(DB[3088]), .Z(n7826) );
  AND U11681 ( .A(n116), .B(n7827), .Z(n7825) );
  XOR U11682 ( .A(n7828), .B(n7829), .Z(n7827) );
  XOR U11683 ( .A(DB[3088]), .B(DB[3057]), .Z(n7829) );
  AND U11684 ( .A(n120), .B(n7830), .Z(n7828) );
  XOR U11685 ( .A(n7831), .B(n7832), .Z(n7830) );
  XOR U11686 ( .A(DB[3057]), .B(DB[3026]), .Z(n7832) );
  AND U11687 ( .A(n124), .B(n7833), .Z(n7831) );
  XOR U11688 ( .A(n7834), .B(n7835), .Z(n7833) );
  XOR U11689 ( .A(DB[3026]), .B(DB[2995]), .Z(n7835) );
  AND U11690 ( .A(n128), .B(n7836), .Z(n7834) );
  XOR U11691 ( .A(n7837), .B(n7838), .Z(n7836) );
  XOR U11692 ( .A(DB[2995]), .B(DB[2964]), .Z(n7838) );
  AND U11693 ( .A(n132), .B(n7839), .Z(n7837) );
  XOR U11694 ( .A(n7840), .B(n7841), .Z(n7839) );
  XOR U11695 ( .A(DB[2964]), .B(DB[2933]), .Z(n7841) );
  AND U11696 ( .A(n136), .B(n7842), .Z(n7840) );
  XOR U11697 ( .A(n7843), .B(n7844), .Z(n7842) );
  XOR U11698 ( .A(DB[2933]), .B(DB[2902]), .Z(n7844) );
  AND U11699 ( .A(n140), .B(n7845), .Z(n7843) );
  XOR U11700 ( .A(n7846), .B(n7847), .Z(n7845) );
  XOR U11701 ( .A(DB[2902]), .B(DB[2871]), .Z(n7847) );
  AND U11702 ( .A(n144), .B(n7848), .Z(n7846) );
  XOR U11703 ( .A(n7849), .B(n7850), .Z(n7848) );
  XOR U11704 ( .A(DB[2871]), .B(DB[2840]), .Z(n7850) );
  AND U11705 ( .A(n148), .B(n7851), .Z(n7849) );
  XOR U11706 ( .A(n7852), .B(n7853), .Z(n7851) );
  XOR U11707 ( .A(DB[2840]), .B(DB[2809]), .Z(n7853) );
  AND U11708 ( .A(n152), .B(n7854), .Z(n7852) );
  XOR U11709 ( .A(n7855), .B(n7856), .Z(n7854) );
  XOR U11710 ( .A(DB[2809]), .B(DB[2778]), .Z(n7856) );
  AND U11711 ( .A(n156), .B(n7857), .Z(n7855) );
  XOR U11712 ( .A(n7858), .B(n7859), .Z(n7857) );
  XOR U11713 ( .A(DB[2778]), .B(DB[2747]), .Z(n7859) );
  AND U11714 ( .A(n160), .B(n7860), .Z(n7858) );
  XOR U11715 ( .A(n7861), .B(n7862), .Z(n7860) );
  XOR U11716 ( .A(DB[2747]), .B(DB[2716]), .Z(n7862) );
  AND U11717 ( .A(n164), .B(n7863), .Z(n7861) );
  XOR U11718 ( .A(n7864), .B(n7865), .Z(n7863) );
  XOR U11719 ( .A(DB[2716]), .B(DB[2685]), .Z(n7865) );
  AND U11720 ( .A(n168), .B(n7866), .Z(n7864) );
  XOR U11721 ( .A(n7867), .B(n7868), .Z(n7866) );
  XOR U11722 ( .A(DB[2685]), .B(DB[2654]), .Z(n7868) );
  AND U11723 ( .A(n172), .B(n7869), .Z(n7867) );
  XOR U11724 ( .A(n7870), .B(n7871), .Z(n7869) );
  XOR U11725 ( .A(DB[2654]), .B(DB[2623]), .Z(n7871) );
  AND U11726 ( .A(n176), .B(n7872), .Z(n7870) );
  XOR U11727 ( .A(n7873), .B(n7874), .Z(n7872) );
  XOR U11728 ( .A(DB[2623]), .B(DB[2592]), .Z(n7874) );
  AND U11729 ( .A(n180), .B(n7875), .Z(n7873) );
  XOR U11730 ( .A(n7876), .B(n7877), .Z(n7875) );
  XOR U11731 ( .A(DB[2592]), .B(DB[2561]), .Z(n7877) );
  AND U11732 ( .A(n184), .B(n7878), .Z(n7876) );
  XOR U11733 ( .A(n7879), .B(n7880), .Z(n7878) );
  XOR U11734 ( .A(DB[2561]), .B(DB[2530]), .Z(n7880) );
  AND U11735 ( .A(n188), .B(n7881), .Z(n7879) );
  XOR U11736 ( .A(n7882), .B(n7883), .Z(n7881) );
  XOR U11737 ( .A(DB[2530]), .B(DB[2499]), .Z(n7883) );
  AND U11738 ( .A(n192), .B(n7884), .Z(n7882) );
  XOR U11739 ( .A(n7885), .B(n7886), .Z(n7884) );
  XOR U11740 ( .A(DB[2499]), .B(DB[2468]), .Z(n7886) );
  AND U11741 ( .A(n196), .B(n7887), .Z(n7885) );
  XOR U11742 ( .A(n7888), .B(n7889), .Z(n7887) );
  XOR U11743 ( .A(DB[2468]), .B(DB[2437]), .Z(n7889) );
  AND U11744 ( .A(n200), .B(n7890), .Z(n7888) );
  XOR U11745 ( .A(n7891), .B(n7892), .Z(n7890) );
  XOR U11746 ( .A(DB[2437]), .B(DB[2406]), .Z(n7892) );
  AND U11747 ( .A(n204), .B(n7893), .Z(n7891) );
  XOR U11748 ( .A(n7894), .B(n7895), .Z(n7893) );
  XOR U11749 ( .A(DB[2406]), .B(DB[2375]), .Z(n7895) );
  AND U11750 ( .A(n208), .B(n7896), .Z(n7894) );
  XOR U11751 ( .A(n7897), .B(n7898), .Z(n7896) );
  XOR U11752 ( .A(DB[2375]), .B(DB[2344]), .Z(n7898) );
  AND U11753 ( .A(n212), .B(n7899), .Z(n7897) );
  XOR U11754 ( .A(n7900), .B(n7901), .Z(n7899) );
  XOR U11755 ( .A(DB[2344]), .B(DB[2313]), .Z(n7901) );
  AND U11756 ( .A(n216), .B(n7902), .Z(n7900) );
  XOR U11757 ( .A(n7903), .B(n7904), .Z(n7902) );
  XOR U11758 ( .A(DB[2313]), .B(DB[2282]), .Z(n7904) );
  AND U11759 ( .A(n220), .B(n7905), .Z(n7903) );
  XOR U11760 ( .A(n7906), .B(n7907), .Z(n7905) );
  XOR U11761 ( .A(DB[2282]), .B(DB[2251]), .Z(n7907) );
  AND U11762 ( .A(n224), .B(n7908), .Z(n7906) );
  XOR U11763 ( .A(n7909), .B(n7910), .Z(n7908) );
  XOR U11764 ( .A(DB[2251]), .B(DB[2220]), .Z(n7910) );
  AND U11765 ( .A(n228), .B(n7911), .Z(n7909) );
  XOR U11766 ( .A(n7912), .B(n7913), .Z(n7911) );
  XOR U11767 ( .A(DB[2220]), .B(DB[2189]), .Z(n7913) );
  AND U11768 ( .A(n232), .B(n7914), .Z(n7912) );
  XOR U11769 ( .A(n7915), .B(n7916), .Z(n7914) );
  XOR U11770 ( .A(DB[2189]), .B(DB[2158]), .Z(n7916) );
  AND U11771 ( .A(n236), .B(n7917), .Z(n7915) );
  XOR U11772 ( .A(n7918), .B(n7919), .Z(n7917) );
  XOR U11773 ( .A(DB[2158]), .B(DB[2127]), .Z(n7919) );
  AND U11774 ( .A(n240), .B(n7920), .Z(n7918) );
  XOR U11775 ( .A(n7921), .B(n7922), .Z(n7920) );
  XOR U11776 ( .A(DB[2127]), .B(DB[2096]), .Z(n7922) );
  AND U11777 ( .A(n244), .B(n7923), .Z(n7921) );
  XOR U11778 ( .A(n7924), .B(n7925), .Z(n7923) );
  XOR U11779 ( .A(DB[2096]), .B(DB[2065]), .Z(n7925) );
  AND U11780 ( .A(n248), .B(n7926), .Z(n7924) );
  XOR U11781 ( .A(n7927), .B(n7928), .Z(n7926) );
  XOR U11782 ( .A(DB[2065]), .B(DB[2034]), .Z(n7928) );
  AND U11783 ( .A(n252), .B(n7929), .Z(n7927) );
  XOR U11784 ( .A(n7930), .B(n7931), .Z(n7929) );
  XOR U11785 ( .A(DB[2034]), .B(DB[2003]), .Z(n7931) );
  AND U11786 ( .A(n256), .B(n7932), .Z(n7930) );
  XOR U11787 ( .A(n7933), .B(n7934), .Z(n7932) );
  XOR U11788 ( .A(DB[2003]), .B(DB[1972]), .Z(n7934) );
  AND U11789 ( .A(n260), .B(n7935), .Z(n7933) );
  XOR U11790 ( .A(n7936), .B(n7937), .Z(n7935) );
  XOR U11791 ( .A(DB[1972]), .B(DB[1941]), .Z(n7937) );
  AND U11792 ( .A(n264), .B(n7938), .Z(n7936) );
  XOR U11793 ( .A(n7939), .B(n7940), .Z(n7938) );
  XOR U11794 ( .A(DB[1941]), .B(DB[1910]), .Z(n7940) );
  AND U11795 ( .A(n268), .B(n7941), .Z(n7939) );
  XOR U11796 ( .A(n7942), .B(n7943), .Z(n7941) );
  XOR U11797 ( .A(DB[1910]), .B(DB[1879]), .Z(n7943) );
  AND U11798 ( .A(n272), .B(n7944), .Z(n7942) );
  XOR U11799 ( .A(n7945), .B(n7946), .Z(n7944) );
  XOR U11800 ( .A(DB[1879]), .B(DB[1848]), .Z(n7946) );
  AND U11801 ( .A(n276), .B(n7947), .Z(n7945) );
  XOR U11802 ( .A(n7948), .B(n7949), .Z(n7947) );
  XOR U11803 ( .A(DB[1848]), .B(DB[1817]), .Z(n7949) );
  AND U11804 ( .A(n280), .B(n7950), .Z(n7948) );
  XOR U11805 ( .A(n7951), .B(n7952), .Z(n7950) );
  XOR U11806 ( .A(DB[1817]), .B(DB[1786]), .Z(n7952) );
  AND U11807 ( .A(n284), .B(n7953), .Z(n7951) );
  XOR U11808 ( .A(n7954), .B(n7955), .Z(n7953) );
  XOR U11809 ( .A(DB[1786]), .B(DB[1755]), .Z(n7955) );
  AND U11810 ( .A(n288), .B(n7956), .Z(n7954) );
  XOR U11811 ( .A(n7957), .B(n7958), .Z(n7956) );
  XOR U11812 ( .A(DB[1755]), .B(DB[1724]), .Z(n7958) );
  AND U11813 ( .A(n292), .B(n7959), .Z(n7957) );
  XOR U11814 ( .A(n7960), .B(n7961), .Z(n7959) );
  XOR U11815 ( .A(DB[1724]), .B(DB[1693]), .Z(n7961) );
  AND U11816 ( .A(n296), .B(n7962), .Z(n7960) );
  XOR U11817 ( .A(n7963), .B(n7964), .Z(n7962) );
  XOR U11818 ( .A(DB[1693]), .B(DB[1662]), .Z(n7964) );
  AND U11819 ( .A(n300), .B(n7965), .Z(n7963) );
  XOR U11820 ( .A(n7966), .B(n7967), .Z(n7965) );
  XOR U11821 ( .A(DB[1662]), .B(DB[1631]), .Z(n7967) );
  AND U11822 ( .A(n304), .B(n7968), .Z(n7966) );
  XOR U11823 ( .A(n7969), .B(n7970), .Z(n7968) );
  XOR U11824 ( .A(DB[1631]), .B(DB[1600]), .Z(n7970) );
  AND U11825 ( .A(n308), .B(n7971), .Z(n7969) );
  XOR U11826 ( .A(n7972), .B(n7973), .Z(n7971) );
  XOR U11827 ( .A(DB[1600]), .B(DB[1569]), .Z(n7973) );
  AND U11828 ( .A(n312), .B(n7974), .Z(n7972) );
  XOR U11829 ( .A(n7975), .B(n7976), .Z(n7974) );
  XOR U11830 ( .A(DB[1569]), .B(DB[1538]), .Z(n7976) );
  AND U11831 ( .A(n316), .B(n7977), .Z(n7975) );
  XOR U11832 ( .A(n7978), .B(n7979), .Z(n7977) );
  XOR U11833 ( .A(DB[1538]), .B(DB[1507]), .Z(n7979) );
  AND U11834 ( .A(n320), .B(n7980), .Z(n7978) );
  XOR U11835 ( .A(n7981), .B(n7982), .Z(n7980) );
  XOR U11836 ( .A(DB[1507]), .B(DB[1476]), .Z(n7982) );
  AND U11837 ( .A(n324), .B(n7983), .Z(n7981) );
  XOR U11838 ( .A(n7984), .B(n7985), .Z(n7983) );
  XOR U11839 ( .A(DB[1476]), .B(DB[1445]), .Z(n7985) );
  AND U11840 ( .A(n328), .B(n7986), .Z(n7984) );
  XOR U11841 ( .A(n7987), .B(n7988), .Z(n7986) );
  XOR U11842 ( .A(DB[1445]), .B(DB[1414]), .Z(n7988) );
  AND U11843 ( .A(n332), .B(n7989), .Z(n7987) );
  XOR U11844 ( .A(n7990), .B(n7991), .Z(n7989) );
  XOR U11845 ( .A(DB[1414]), .B(DB[1383]), .Z(n7991) );
  AND U11846 ( .A(n336), .B(n7992), .Z(n7990) );
  XOR U11847 ( .A(n7993), .B(n7994), .Z(n7992) );
  XOR U11848 ( .A(DB[1383]), .B(DB[1352]), .Z(n7994) );
  AND U11849 ( .A(n340), .B(n7995), .Z(n7993) );
  XOR U11850 ( .A(n7996), .B(n7997), .Z(n7995) );
  XOR U11851 ( .A(DB[1352]), .B(DB[1321]), .Z(n7997) );
  AND U11852 ( .A(n344), .B(n7998), .Z(n7996) );
  XOR U11853 ( .A(n7999), .B(n8000), .Z(n7998) );
  XOR U11854 ( .A(DB[1321]), .B(DB[1290]), .Z(n8000) );
  AND U11855 ( .A(n348), .B(n8001), .Z(n7999) );
  XOR U11856 ( .A(n8002), .B(n8003), .Z(n8001) );
  XOR U11857 ( .A(DB[1290]), .B(DB[1259]), .Z(n8003) );
  AND U11858 ( .A(n352), .B(n8004), .Z(n8002) );
  XOR U11859 ( .A(n8005), .B(n8006), .Z(n8004) );
  XOR U11860 ( .A(DB[1259]), .B(DB[1228]), .Z(n8006) );
  AND U11861 ( .A(n356), .B(n8007), .Z(n8005) );
  XOR U11862 ( .A(n8008), .B(n8009), .Z(n8007) );
  XOR U11863 ( .A(DB[1228]), .B(DB[1197]), .Z(n8009) );
  AND U11864 ( .A(n360), .B(n8010), .Z(n8008) );
  XOR U11865 ( .A(n8011), .B(n8012), .Z(n8010) );
  XOR U11866 ( .A(DB[1197]), .B(DB[1166]), .Z(n8012) );
  AND U11867 ( .A(n364), .B(n8013), .Z(n8011) );
  XOR U11868 ( .A(n8014), .B(n8015), .Z(n8013) );
  XOR U11869 ( .A(DB[1166]), .B(DB[1135]), .Z(n8015) );
  AND U11870 ( .A(n368), .B(n8016), .Z(n8014) );
  XOR U11871 ( .A(n8017), .B(n8018), .Z(n8016) );
  XOR U11872 ( .A(DB[1135]), .B(DB[1104]), .Z(n8018) );
  AND U11873 ( .A(n372), .B(n8019), .Z(n8017) );
  XOR U11874 ( .A(n8020), .B(n8021), .Z(n8019) );
  XOR U11875 ( .A(DB[1104]), .B(DB[1073]), .Z(n8021) );
  AND U11876 ( .A(n376), .B(n8022), .Z(n8020) );
  XOR U11877 ( .A(n8023), .B(n8024), .Z(n8022) );
  XOR U11878 ( .A(DB[1073]), .B(DB[1042]), .Z(n8024) );
  AND U11879 ( .A(n380), .B(n8025), .Z(n8023) );
  XOR U11880 ( .A(n8026), .B(n8027), .Z(n8025) );
  XOR U11881 ( .A(DB[1042]), .B(DB[1011]), .Z(n8027) );
  AND U11882 ( .A(n384), .B(n8028), .Z(n8026) );
  XOR U11883 ( .A(n8029), .B(n8030), .Z(n8028) );
  XOR U11884 ( .A(DB[980]), .B(DB[1011]), .Z(n8030) );
  AND U11885 ( .A(n388), .B(n8031), .Z(n8029) );
  XOR U11886 ( .A(n8032), .B(n8033), .Z(n8031) );
  XOR U11887 ( .A(DB[980]), .B(DB[949]), .Z(n8033) );
  AND U11888 ( .A(n392), .B(n8034), .Z(n8032) );
  XOR U11889 ( .A(n8035), .B(n8036), .Z(n8034) );
  XOR U11890 ( .A(DB[949]), .B(DB[918]), .Z(n8036) );
  AND U11891 ( .A(n396), .B(n8037), .Z(n8035) );
  XOR U11892 ( .A(n8038), .B(n8039), .Z(n8037) );
  XOR U11893 ( .A(DB[918]), .B(DB[887]), .Z(n8039) );
  AND U11894 ( .A(n400), .B(n8040), .Z(n8038) );
  XOR U11895 ( .A(n8041), .B(n8042), .Z(n8040) );
  XOR U11896 ( .A(DB[887]), .B(DB[856]), .Z(n8042) );
  AND U11897 ( .A(n404), .B(n8043), .Z(n8041) );
  XOR U11898 ( .A(n8044), .B(n8045), .Z(n8043) );
  XOR U11899 ( .A(DB[856]), .B(DB[825]), .Z(n8045) );
  AND U11900 ( .A(n408), .B(n8046), .Z(n8044) );
  XOR U11901 ( .A(n8047), .B(n8048), .Z(n8046) );
  XOR U11902 ( .A(DB[825]), .B(DB[794]), .Z(n8048) );
  AND U11903 ( .A(n412), .B(n8049), .Z(n8047) );
  XOR U11904 ( .A(n8050), .B(n8051), .Z(n8049) );
  XOR U11905 ( .A(DB[794]), .B(DB[763]), .Z(n8051) );
  AND U11906 ( .A(n416), .B(n8052), .Z(n8050) );
  XOR U11907 ( .A(n8053), .B(n8054), .Z(n8052) );
  XOR U11908 ( .A(DB[763]), .B(DB[732]), .Z(n8054) );
  AND U11909 ( .A(n420), .B(n8055), .Z(n8053) );
  XOR U11910 ( .A(n8056), .B(n8057), .Z(n8055) );
  XOR U11911 ( .A(DB[732]), .B(DB[701]), .Z(n8057) );
  AND U11912 ( .A(n424), .B(n8058), .Z(n8056) );
  XOR U11913 ( .A(n8059), .B(n8060), .Z(n8058) );
  XOR U11914 ( .A(DB[701]), .B(DB[670]), .Z(n8060) );
  AND U11915 ( .A(n428), .B(n8061), .Z(n8059) );
  XOR U11916 ( .A(n8062), .B(n8063), .Z(n8061) );
  XOR U11917 ( .A(DB[670]), .B(DB[639]), .Z(n8063) );
  AND U11918 ( .A(n432), .B(n8064), .Z(n8062) );
  XOR U11919 ( .A(n8065), .B(n8066), .Z(n8064) );
  XOR U11920 ( .A(DB[639]), .B(DB[608]), .Z(n8066) );
  AND U11921 ( .A(n436), .B(n8067), .Z(n8065) );
  XOR U11922 ( .A(n8068), .B(n8069), .Z(n8067) );
  XOR U11923 ( .A(DB[608]), .B(DB[577]), .Z(n8069) );
  AND U11924 ( .A(n440), .B(n8070), .Z(n8068) );
  XOR U11925 ( .A(n8071), .B(n8072), .Z(n8070) );
  XOR U11926 ( .A(DB[577]), .B(DB[546]), .Z(n8072) );
  AND U11927 ( .A(n444), .B(n8073), .Z(n8071) );
  XOR U11928 ( .A(n8074), .B(n8075), .Z(n8073) );
  XOR U11929 ( .A(DB[546]), .B(DB[515]), .Z(n8075) );
  AND U11930 ( .A(n448), .B(n8076), .Z(n8074) );
  XOR U11931 ( .A(n8077), .B(n8078), .Z(n8076) );
  XOR U11932 ( .A(DB[515]), .B(DB[484]), .Z(n8078) );
  AND U11933 ( .A(n452), .B(n8079), .Z(n8077) );
  XOR U11934 ( .A(n8080), .B(n8081), .Z(n8079) );
  XOR U11935 ( .A(DB[484]), .B(DB[453]), .Z(n8081) );
  AND U11936 ( .A(n456), .B(n8082), .Z(n8080) );
  XOR U11937 ( .A(n8083), .B(n8084), .Z(n8082) );
  XOR U11938 ( .A(DB[453]), .B(DB[422]), .Z(n8084) );
  AND U11939 ( .A(n460), .B(n8085), .Z(n8083) );
  XOR U11940 ( .A(n8086), .B(n8087), .Z(n8085) );
  XOR U11941 ( .A(DB[422]), .B(DB[391]), .Z(n8087) );
  AND U11942 ( .A(n464), .B(n8088), .Z(n8086) );
  XOR U11943 ( .A(n8089), .B(n8090), .Z(n8088) );
  XOR U11944 ( .A(DB[391]), .B(DB[360]), .Z(n8090) );
  AND U11945 ( .A(n468), .B(n8091), .Z(n8089) );
  XOR U11946 ( .A(n8092), .B(n8093), .Z(n8091) );
  XOR U11947 ( .A(DB[360]), .B(DB[329]), .Z(n8093) );
  AND U11948 ( .A(n472), .B(n8094), .Z(n8092) );
  XOR U11949 ( .A(n8095), .B(n8096), .Z(n8094) );
  XOR U11950 ( .A(DB[329]), .B(DB[298]), .Z(n8096) );
  AND U11951 ( .A(n476), .B(n8097), .Z(n8095) );
  XOR U11952 ( .A(n8098), .B(n8099), .Z(n8097) );
  XOR U11953 ( .A(DB[298]), .B(DB[267]), .Z(n8099) );
  AND U11954 ( .A(n480), .B(n8100), .Z(n8098) );
  XOR U11955 ( .A(n8101), .B(n8102), .Z(n8100) );
  XOR U11956 ( .A(DB[267]), .B(DB[236]), .Z(n8102) );
  AND U11957 ( .A(n484), .B(n8103), .Z(n8101) );
  XOR U11958 ( .A(n8104), .B(n8105), .Z(n8103) );
  XOR U11959 ( .A(DB[236]), .B(DB[205]), .Z(n8105) );
  AND U11960 ( .A(n488), .B(n8106), .Z(n8104) );
  XOR U11961 ( .A(n8107), .B(n8108), .Z(n8106) );
  XOR U11962 ( .A(DB[205]), .B(DB[174]), .Z(n8108) );
  AND U11963 ( .A(n492), .B(n8109), .Z(n8107) );
  XOR U11964 ( .A(n8110), .B(n8111), .Z(n8109) );
  XOR U11965 ( .A(DB[174]), .B(DB[143]), .Z(n8111) );
  AND U11966 ( .A(n496), .B(n8112), .Z(n8110) );
  XOR U11967 ( .A(n8113), .B(n8114), .Z(n8112) );
  XOR U11968 ( .A(DB[143]), .B(DB[112]), .Z(n8114) );
  AND U11969 ( .A(n500), .B(n8115), .Z(n8113) );
  XOR U11970 ( .A(n8116), .B(n8117), .Z(n8115) );
  XOR U11971 ( .A(DB[81]), .B(DB[112]), .Z(n8117) );
  AND U11972 ( .A(n504), .B(n8118), .Z(n8116) );
  XOR U11973 ( .A(n8119), .B(n8120), .Z(n8118) );
  XOR U11974 ( .A(DB[81]), .B(DB[50]), .Z(n8120) );
  AND U11975 ( .A(n508), .B(n8121), .Z(n8119) );
  XOR U11976 ( .A(DB[50]), .B(DB[19]), .Z(n8121) );
  XOR U11977 ( .A(DB[3955]), .B(n8122), .Z(min_val_out[18]) );
  AND U11978 ( .A(n2), .B(n8123), .Z(n8122) );
  XOR U11979 ( .A(n8124), .B(n8125), .Z(n8123) );
  XOR U11980 ( .A(n8126), .B(n8127), .Z(n8125) );
  IV U11981 ( .A(DB[3955]), .Z(n8126) );
  AND U11982 ( .A(n8), .B(n8128), .Z(n8124) );
  XOR U11983 ( .A(n8129), .B(n8130), .Z(n8128) );
  XOR U11984 ( .A(DB[3924]), .B(DB[3893]), .Z(n8130) );
  AND U11985 ( .A(n12), .B(n8131), .Z(n8129) );
  XOR U11986 ( .A(n8132), .B(n8133), .Z(n8131) );
  XOR U11987 ( .A(DB[3893]), .B(DB[3862]), .Z(n8133) );
  AND U11988 ( .A(n16), .B(n8134), .Z(n8132) );
  XOR U11989 ( .A(n8135), .B(n8136), .Z(n8134) );
  XOR U11990 ( .A(DB[3862]), .B(DB[3831]), .Z(n8136) );
  AND U11991 ( .A(n20), .B(n8137), .Z(n8135) );
  XOR U11992 ( .A(n8138), .B(n8139), .Z(n8137) );
  XOR U11993 ( .A(DB[3831]), .B(DB[3800]), .Z(n8139) );
  AND U11994 ( .A(n24), .B(n8140), .Z(n8138) );
  XOR U11995 ( .A(n8141), .B(n8142), .Z(n8140) );
  XOR U11996 ( .A(DB[3800]), .B(DB[3769]), .Z(n8142) );
  AND U11997 ( .A(n28), .B(n8143), .Z(n8141) );
  XOR U11998 ( .A(n8144), .B(n8145), .Z(n8143) );
  XOR U11999 ( .A(DB[3769]), .B(DB[3738]), .Z(n8145) );
  AND U12000 ( .A(n32), .B(n8146), .Z(n8144) );
  XOR U12001 ( .A(n8147), .B(n8148), .Z(n8146) );
  XOR U12002 ( .A(DB[3738]), .B(DB[3707]), .Z(n8148) );
  AND U12003 ( .A(n36), .B(n8149), .Z(n8147) );
  XOR U12004 ( .A(n8150), .B(n8151), .Z(n8149) );
  XOR U12005 ( .A(DB[3707]), .B(DB[3676]), .Z(n8151) );
  AND U12006 ( .A(n40), .B(n8152), .Z(n8150) );
  XOR U12007 ( .A(n8153), .B(n8154), .Z(n8152) );
  XOR U12008 ( .A(DB[3676]), .B(DB[3645]), .Z(n8154) );
  AND U12009 ( .A(n44), .B(n8155), .Z(n8153) );
  XOR U12010 ( .A(n8156), .B(n8157), .Z(n8155) );
  XOR U12011 ( .A(DB[3645]), .B(DB[3614]), .Z(n8157) );
  AND U12012 ( .A(n48), .B(n8158), .Z(n8156) );
  XOR U12013 ( .A(n8159), .B(n8160), .Z(n8158) );
  XOR U12014 ( .A(DB[3614]), .B(DB[3583]), .Z(n8160) );
  AND U12015 ( .A(n52), .B(n8161), .Z(n8159) );
  XOR U12016 ( .A(n8162), .B(n8163), .Z(n8161) );
  XOR U12017 ( .A(DB[3583]), .B(DB[3552]), .Z(n8163) );
  AND U12018 ( .A(n56), .B(n8164), .Z(n8162) );
  XOR U12019 ( .A(n8165), .B(n8166), .Z(n8164) );
  XOR U12020 ( .A(DB[3552]), .B(DB[3521]), .Z(n8166) );
  AND U12021 ( .A(n60), .B(n8167), .Z(n8165) );
  XOR U12022 ( .A(n8168), .B(n8169), .Z(n8167) );
  XOR U12023 ( .A(DB[3521]), .B(DB[3490]), .Z(n8169) );
  AND U12024 ( .A(n64), .B(n8170), .Z(n8168) );
  XOR U12025 ( .A(n8171), .B(n8172), .Z(n8170) );
  XOR U12026 ( .A(DB[3490]), .B(DB[3459]), .Z(n8172) );
  AND U12027 ( .A(n68), .B(n8173), .Z(n8171) );
  XOR U12028 ( .A(n8174), .B(n8175), .Z(n8173) );
  XOR U12029 ( .A(DB[3459]), .B(DB[3428]), .Z(n8175) );
  AND U12030 ( .A(n72), .B(n8176), .Z(n8174) );
  XOR U12031 ( .A(n8177), .B(n8178), .Z(n8176) );
  XOR U12032 ( .A(DB[3428]), .B(DB[3397]), .Z(n8178) );
  AND U12033 ( .A(n76), .B(n8179), .Z(n8177) );
  XOR U12034 ( .A(n8180), .B(n8181), .Z(n8179) );
  XOR U12035 ( .A(DB[3397]), .B(DB[3366]), .Z(n8181) );
  AND U12036 ( .A(n80), .B(n8182), .Z(n8180) );
  XOR U12037 ( .A(n8183), .B(n8184), .Z(n8182) );
  XOR U12038 ( .A(DB[3366]), .B(DB[3335]), .Z(n8184) );
  AND U12039 ( .A(n84), .B(n8185), .Z(n8183) );
  XOR U12040 ( .A(n8186), .B(n8187), .Z(n8185) );
  XOR U12041 ( .A(DB[3335]), .B(DB[3304]), .Z(n8187) );
  AND U12042 ( .A(n88), .B(n8188), .Z(n8186) );
  XOR U12043 ( .A(n8189), .B(n8190), .Z(n8188) );
  XOR U12044 ( .A(DB[3304]), .B(DB[3273]), .Z(n8190) );
  AND U12045 ( .A(n92), .B(n8191), .Z(n8189) );
  XOR U12046 ( .A(n8192), .B(n8193), .Z(n8191) );
  XOR U12047 ( .A(DB[3273]), .B(DB[3242]), .Z(n8193) );
  AND U12048 ( .A(n96), .B(n8194), .Z(n8192) );
  XOR U12049 ( .A(n8195), .B(n8196), .Z(n8194) );
  XOR U12050 ( .A(DB[3242]), .B(DB[3211]), .Z(n8196) );
  AND U12051 ( .A(n100), .B(n8197), .Z(n8195) );
  XOR U12052 ( .A(n8198), .B(n8199), .Z(n8197) );
  XOR U12053 ( .A(DB[3211]), .B(DB[3180]), .Z(n8199) );
  AND U12054 ( .A(n104), .B(n8200), .Z(n8198) );
  XOR U12055 ( .A(n8201), .B(n8202), .Z(n8200) );
  XOR U12056 ( .A(DB[3180]), .B(DB[3149]), .Z(n8202) );
  AND U12057 ( .A(n108), .B(n8203), .Z(n8201) );
  XOR U12058 ( .A(n8204), .B(n8205), .Z(n8203) );
  XOR U12059 ( .A(DB[3149]), .B(DB[3118]), .Z(n8205) );
  AND U12060 ( .A(n112), .B(n8206), .Z(n8204) );
  XOR U12061 ( .A(n8207), .B(n8208), .Z(n8206) );
  XOR U12062 ( .A(DB[3118]), .B(DB[3087]), .Z(n8208) );
  AND U12063 ( .A(n116), .B(n8209), .Z(n8207) );
  XOR U12064 ( .A(n8210), .B(n8211), .Z(n8209) );
  XOR U12065 ( .A(DB[3087]), .B(DB[3056]), .Z(n8211) );
  AND U12066 ( .A(n120), .B(n8212), .Z(n8210) );
  XOR U12067 ( .A(n8213), .B(n8214), .Z(n8212) );
  XOR U12068 ( .A(DB[3056]), .B(DB[3025]), .Z(n8214) );
  AND U12069 ( .A(n124), .B(n8215), .Z(n8213) );
  XOR U12070 ( .A(n8216), .B(n8217), .Z(n8215) );
  XOR U12071 ( .A(DB[3025]), .B(DB[2994]), .Z(n8217) );
  AND U12072 ( .A(n128), .B(n8218), .Z(n8216) );
  XOR U12073 ( .A(n8219), .B(n8220), .Z(n8218) );
  XOR U12074 ( .A(DB[2994]), .B(DB[2963]), .Z(n8220) );
  AND U12075 ( .A(n132), .B(n8221), .Z(n8219) );
  XOR U12076 ( .A(n8222), .B(n8223), .Z(n8221) );
  XOR U12077 ( .A(DB[2963]), .B(DB[2932]), .Z(n8223) );
  AND U12078 ( .A(n136), .B(n8224), .Z(n8222) );
  XOR U12079 ( .A(n8225), .B(n8226), .Z(n8224) );
  XOR U12080 ( .A(DB[2932]), .B(DB[2901]), .Z(n8226) );
  AND U12081 ( .A(n140), .B(n8227), .Z(n8225) );
  XOR U12082 ( .A(n8228), .B(n8229), .Z(n8227) );
  XOR U12083 ( .A(DB[2901]), .B(DB[2870]), .Z(n8229) );
  AND U12084 ( .A(n144), .B(n8230), .Z(n8228) );
  XOR U12085 ( .A(n8231), .B(n8232), .Z(n8230) );
  XOR U12086 ( .A(DB[2870]), .B(DB[2839]), .Z(n8232) );
  AND U12087 ( .A(n148), .B(n8233), .Z(n8231) );
  XOR U12088 ( .A(n8234), .B(n8235), .Z(n8233) );
  XOR U12089 ( .A(DB[2839]), .B(DB[2808]), .Z(n8235) );
  AND U12090 ( .A(n152), .B(n8236), .Z(n8234) );
  XOR U12091 ( .A(n8237), .B(n8238), .Z(n8236) );
  XOR U12092 ( .A(DB[2808]), .B(DB[2777]), .Z(n8238) );
  AND U12093 ( .A(n156), .B(n8239), .Z(n8237) );
  XOR U12094 ( .A(n8240), .B(n8241), .Z(n8239) );
  XOR U12095 ( .A(DB[2777]), .B(DB[2746]), .Z(n8241) );
  AND U12096 ( .A(n160), .B(n8242), .Z(n8240) );
  XOR U12097 ( .A(n8243), .B(n8244), .Z(n8242) );
  XOR U12098 ( .A(DB[2746]), .B(DB[2715]), .Z(n8244) );
  AND U12099 ( .A(n164), .B(n8245), .Z(n8243) );
  XOR U12100 ( .A(n8246), .B(n8247), .Z(n8245) );
  XOR U12101 ( .A(DB[2715]), .B(DB[2684]), .Z(n8247) );
  AND U12102 ( .A(n168), .B(n8248), .Z(n8246) );
  XOR U12103 ( .A(n8249), .B(n8250), .Z(n8248) );
  XOR U12104 ( .A(DB[2684]), .B(DB[2653]), .Z(n8250) );
  AND U12105 ( .A(n172), .B(n8251), .Z(n8249) );
  XOR U12106 ( .A(n8252), .B(n8253), .Z(n8251) );
  XOR U12107 ( .A(DB[2653]), .B(DB[2622]), .Z(n8253) );
  AND U12108 ( .A(n176), .B(n8254), .Z(n8252) );
  XOR U12109 ( .A(n8255), .B(n8256), .Z(n8254) );
  XOR U12110 ( .A(DB[2622]), .B(DB[2591]), .Z(n8256) );
  AND U12111 ( .A(n180), .B(n8257), .Z(n8255) );
  XOR U12112 ( .A(n8258), .B(n8259), .Z(n8257) );
  XOR U12113 ( .A(DB[2591]), .B(DB[2560]), .Z(n8259) );
  AND U12114 ( .A(n184), .B(n8260), .Z(n8258) );
  XOR U12115 ( .A(n8261), .B(n8262), .Z(n8260) );
  XOR U12116 ( .A(DB[2560]), .B(DB[2529]), .Z(n8262) );
  AND U12117 ( .A(n188), .B(n8263), .Z(n8261) );
  XOR U12118 ( .A(n8264), .B(n8265), .Z(n8263) );
  XOR U12119 ( .A(DB[2529]), .B(DB[2498]), .Z(n8265) );
  AND U12120 ( .A(n192), .B(n8266), .Z(n8264) );
  XOR U12121 ( .A(n8267), .B(n8268), .Z(n8266) );
  XOR U12122 ( .A(DB[2498]), .B(DB[2467]), .Z(n8268) );
  AND U12123 ( .A(n196), .B(n8269), .Z(n8267) );
  XOR U12124 ( .A(n8270), .B(n8271), .Z(n8269) );
  XOR U12125 ( .A(DB[2467]), .B(DB[2436]), .Z(n8271) );
  AND U12126 ( .A(n200), .B(n8272), .Z(n8270) );
  XOR U12127 ( .A(n8273), .B(n8274), .Z(n8272) );
  XOR U12128 ( .A(DB[2436]), .B(DB[2405]), .Z(n8274) );
  AND U12129 ( .A(n204), .B(n8275), .Z(n8273) );
  XOR U12130 ( .A(n8276), .B(n8277), .Z(n8275) );
  XOR U12131 ( .A(DB[2405]), .B(DB[2374]), .Z(n8277) );
  AND U12132 ( .A(n208), .B(n8278), .Z(n8276) );
  XOR U12133 ( .A(n8279), .B(n8280), .Z(n8278) );
  XOR U12134 ( .A(DB[2374]), .B(DB[2343]), .Z(n8280) );
  AND U12135 ( .A(n212), .B(n8281), .Z(n8279) );
  XOR U12136 ( .A(n8282), .B(n8283), .Z(n8281) );
  XOR U12137 ( .A(DB[2343]), .B(DB[2312]), .Z(n8283) );
  AND U12138 ( .A(n216), .B(n8284), .Z(n8282) );
  XOR U12139 ( .A(n8285), .B(n8286), .Z(n8284) );
  XOR U12140 ( .A(DB[2312]), .B(DB[2281]), .Z(n8286) );
  AND U12141 ( .A(n220), .B(n8287), .Z(n8285) );
  XOR U12142 ( .A(n8288), .B(n8289), .Z(n8287) );
  XOR U12143 ( .A(DB[2281]), .B(DB[2250]), .Z(n8289) );
  AND U12144 ( .A(n224), .B(n8290), .Z(n8288) );
  XOR U12145 ( .A(n8291), .B(n8292), .Z(n8290) );
  XOR U12146 ( .A(DB[2250]), .B(DB[2219]), .Z(n8292) );
  AND U12147 ( .A(n228), .B(n8293), .Z(n8291) );
  XOR U12148 ( .A(n8294), .B(n8295), .Z(n8293) );
  XOR U12149 ( .A(DB[2219]), .B(DB[2188]), .Z(n8295) );
  AND U12150 ( .A(n232), .B(n8296), .Z(n8294) );
  XOR U12151 ( .A(n8297), .B(n8298), .Z(n8296) );
  XOR U12152 ( .A(DB[2188]), .B(DB[2157]), .Z(n8298) );
  AND U12153 ( .A(n236), .B(n8299), .Z(n8297) );
  XOR U12154 ( .A(n8300), .B(n8301), .Z(n8299) );
  XOR U12155 ( .A(DB[2157]), .B(DB[2126]), .Z(n8301) );
  AND U12156 ( .A(n240), .B(n8302), .Z(n8300) );
  XOR U12157 ( .A(n8303), .B(n8304), .Z(n8302) );
  XOR U12158 ( .A(DB[2126]), .B(DB[2095]), .Z(n8304) );
  AND U12159 ( .A(n244), .B(n8305), .Z(n8303) );
  XOR U12160 ( .A(n8306), .B(n8307), .Z(n8305) );
  XOR U12161 ( .A(DB[2095]), .B(DB[2064]), .Z(n8307) );
  AND U12162 ( .A(n248), .B(n8308), .Z(n8306) );
  XOR U12163 ( .A(n8309), .B(n8310), .Z(n8308) );
  XOR U12164 ( .A(DB[2064]), .B(DB[2033]), .Z(n8310) );
  AND U12165 ( .A(n252), .B(n8311), .Z(n8309) );
  XOR U12166 ( .A(n8312), .B(n8313), .Z(n8311) );
  XOR U12167 ( .A(DB[2033]), .B(DB[2002]), .Z(n8313) );
  AND U12168 ( .A(n256), .B(n8314), .Z(n8312) );
  XOR U12169 ( .A(n8315), .B(n8316), .Z(n8314) );
  XOR U12170 ( .A(DB[2002]), .B(DB[1971]), .Z(n8316) );
  AND U12171 ( .A(n260), .B(n8317), .Z(n8315) );
  XOR U12172 ( .A(n8318), .B(n8319), .Z(n8317) );
  XOR U12173 ( .A(DB[1971]), .B(DB[1940]), .Z(n8319) );
  AND U12174 ( .A(n264), .B(n8320), .Z(n8318) );
  XOR U12175 ( .A(n8321), .B(n8322), .Z(n8320) );
  XOR U12176 ( .A(DB[1940]), .B(DB[1909]), .Z(n8322) );
  AND U12177 ( .A(n268), .B(n8323), .Z(n8321) );
  XOR U12178 ( .A(n8324), .B(n8325), .Z(n8323) );
  XOR U12179 ( .A(DB[1909]), .B(DB[1878]), .Z(n8325) );
  AND U12180 ( .A(n272), .B(n8326), .Z(n8324) );
  XOR U12181 ( .A(n8327), .B(n8328), .Z(n8326) );
  XOR U12182 ( .A(DB[1878]), .B(DB[1847]), .Z(n8328) );
  AND U12183 ( .A(n276), .B(n8329), .Z(n8327) );
  XOR U12184 ( .A(n8330), .B(n8331), .Z(n8329) );
  XOR U12185 ( .A(DB[1847]), .B(DB[1816]), .Z(n8331) );
  AND U12186 ( .A(n280), .B(n8332), .Z(n8330) );
  XOR U12187 ( .A(n8333), .B(n8334), .Z(n8332) );
  XOR U12188 ( .A(DB[1816]), .B(DB[1785]), .Z(n8334) );
  AND U12189 ( .A(n284), .B(n8335), .Z(n8333) );
  XOR U12190 ( .A(n8336), .B(n8337), .Z(n8335) );
  XOR U12191 ( .A(DB[1785]), .B(DB[1754]), .Z(n8337) );
  AND U12192 ( .A(n288), .B(n8338), .Z(n8336) );
  XOR U12193 ( .A(n8339), .B(n8340), .Z(n8338) );
  XOR U12194 ( .A(DB[1754]), .B(DB[1723]), .Z(n8340) );
  AND U12195 ( .A(n292), .B(n8341), .Z(n8339) );
  XOR U12196 ( .A(n8342), .B(n8343), .Z(n8341) );
  XOR U12197 ( .A(DB[1723]), .B(DB[1692]), .Z(n8343) );
  AND U12198 ( .A(n296), .B(n8344), .Z(n8342) );
  XOR U12199 ( .A(n8345), .B(n8346), .Z(n8344) );
  XOR U12200 ( .A(DB[1692]), .B(DB[1661]), .Z(n8346) );
  AND U12201 ( .A(n300), .B(n8347), .Z(n8345) );
  XOR U12202 ( .A(n8348), .B(n8349), .Z(n8347) );
  XOR U12203 ( .A(DB[1661]), .B(DB[1630]), .Z(n8349) );
  AND U12204 ( .A(n304), .B(n8350), .Z(n8348) );
  XOR U12205 ( .A(n8351), .B(n8352), .Z(n8350) );
  XOR U12206 ( .A(DB[1630]), .B(DB[1599]), .Z(n8352) );
  AND U12207 ( .A(n308), .B(n8353), .Z(n8351) );
  XOR U12208 ( .A(n8354), .B(n8355), .Z(n8353) );
  XOR U12209 ( .A(DB[1599]), .B(DB[1568]), .Z(n8355) );
  AND U12210 ( .A(n312), .B(n8356), .Z(n8354) );
  XOR U12211 ( .A(n8357), .B(n8358), .Z(n8356) );
  XOR U12212 ( .A(DB[1568]), .B(DB[1537]), .Z(n8358) );
  AND U12213 ( .A(n316), .B(n8359), .Z(n8357) );
  XOR U12214 ( .A(n8360), .B(n8361), .Z(n8359) );
  XOR U12215 ( .A(DB[1537]), .B(DB[1506]), .Z(n8361) );
  AND U12216 ( .A(n320), .B(n8362), .Z(n8360) );
  XOR U12217 ( .A(n8363), .B(n8364), .Z(n8362) );
  XOR U12218 ( .A(DB[1506]), .B(DB[1475]), .Z(n8364) );
  AND U12219 ( .A(n324), .B(n8365), .Z(n8363) );
  XOR U12220 ( .A(n8366), .B(n8367), .Z(n8365) );
  XOR U12221 ( .A(DB[1475]), .B(DB[1444]), .Z(n8367) );
  AND U12222 ( .A(n328), .B(n8368), .Z(n8366) );
  XOR U12223 ( .A(n8369), .B(n8370), .Z(n8368) );
  XOR U12224 ( .A(DB[1444]), .B(DB[1413]), .Z(n8370) );
  AND U12225 ( .A(n332), .B(n8371), .Z(n8369) );
  XOR U12226 ( .A(n8372), .B(n8373), .Z(n8371) );
  XOR U12227 ( .A(DB[1413]), .B(DB[1382]), .Z(n8373) );
  AND U12228 ( .A(n336), .B(n8374), .Z(n8372) );
  XOR U12229 ( .A(n8375), .B(n8376), .Z(n8374) );
  XOR U12230 ( .A(DB[1382]), .B(DB[1351]), .Z(n8376) );
  AND U12231 ( .A(n340), .B(n8377), .Z(n8375) );
  XOR U12232 ( .A(n8378), .B(n8379), .Z(n8377) );
  XOR U12233 ( .A(DB[1351]), .B(DB[1320]), .Z(n8379) );
  AND U12234 ( .A(n344), .B(n8380), .Z(n8378) );
  XOR U12235 ( .A(n8381), .B(n8382), .Z(n8380) );
  XOR U12236 ( .A(DB[1320]), .B(DB[1289]), .Z(n8382) );
  AND U12237 ( .A(n348), .B(n8383), .Z(n8381) );
  XOR U12238 ( .A(n8384), .B(n8385), .Z(n8383) );
  XOR U12239 ( .A(DB[1289]), .B(DB[1258]), .Z(n8385) );
  AND U12240 ( .A(n352), .B(n8386), .Z(n8384) );
  XOR U12241 ( .A(n8387), .B(n8388), .Z(n8386) );
  XOR U12242 ( .A(DB[1258]), .B(DB[1227]), .Z(n8388) );
  AND U12243 ( .A(n356), .B(n8389), .Z(n8387) );
  XOR U12244 ( .A(n8390), .B(n8391), .Z(n8389) );
  XOR U12245 ( .A(DB[1227]), .B(DB[1196]), .Z(n8391) );
  AND U12246 ( .A(n360), .B(n8392), .Z(n8390) );
  XOR U12247 ( .A(n8393), .B(n8394), .Z(n8392) );
  XOR U12248 ( .A(DB[1196]), .B(DB[1165]), .Z(n8394) );
  AND U12249 ( .A(n364), .B(n8395), .Z(n8393) );
  XOR U12250 ( .A(n8396), .B(n8397), .Z(n8395) );
  XOR U12251 ( .A(DB[1165]), .B(DB[1134]), .Z(n8397) );
  AND U12252 ( .A(n368), .B(n8398), .Z(n8396) );
  XOR U12253 ( .A(n8399), .B(n8400), .Z(n8398) );
  XOR U12254 ( .A(DB[1134]), .B(DB[1103]), .Z(n8400) );
  AND U12255 ( .A(n372), .B(n8401), .Z(n8399) );
  XOR U12256 ( .A(n8402), .B(n8403), .Z(n8401) );
  XOR U12257 ( .A(DB[1103]), .B(DB[1072]), .Z(n8403) );
  AND U12258 ( .A(n376), .B(n8404), .Z(n8402) );
  XOR U12259 ( .A(n8405), .B(n8406), .Z(n8404) );
  XOR U12260 ( .A(DB[1072]), .B(DB[1041]), .Z(n8406) );
  AND U12261 ( .A(n380), .B(n8407), .Z(n8405) );
  XOR U12262 ( .A(n8408), .B(n8409), .Z(n8407) );
  XOR U12263 ( .A(DB[1041]), .B(DB[1010]), .Z(n8409) );
  AND U12264 ( .A(n384), .B(n8410), .Z(n8408) );
  XOR U12265 ( .A(n8411), .B(n8412), .Z(n8410) );
  XOR U12266 ( .A(DB[979]), .B(DB[1010]), .Z(n8412) );
  AND U12267 ( .A(n388), .B(n8413), .Z(n8411) );
  XOR U12268 ( .A(n8414), .B(n8415), .Z(n8413) );
  XOR U12269 ( .A(DB[979]), .B(DB[948]), .Z(n8415) );
  AND U12270 ( .A(n392), .B(n8416), .Z(n8414) );
  XOR U12271 ( .A(n8417), .B(n8418), .Z(n8416) );
  XOR U12272 ( .A(DB[948]), .B(DB[917]), .Z(n8418) );
  AND U12273 ( .A(n396), .B(n8419), .Z(n8417) );
  XOR U12274 ( .A(n8420), .B(n8421), .Z(n8419) );
  XOR U12275 ( .A(DB[917]), .B(DB[886]), .Z(n8421) );
  AND U12276 ( .A(n400), .B(n8422), .Z(n8420) );
  XOR U12277 ( .A(n8423), .B(n8424), .Z(n8422) );
  XOR U12278 ( .A(DB[886]), .B(DB[855]), .Z(n8424) );
  AND U12279 ( .A(n404), .B(n8425), .Z(n8423) );
  XOR U12280 ( .A(n8426), .B(n8427), .Z(n8425) );
  XOR U12281 ( .A(DB[855]), .B(DB[824]), .Z(n8427) );
  AND U12282 ( .A(n408), .B(n8428), .Z(n8426) );
  XOR U12283 ( .A(n8429), .B(n8430), .Z(n8428) );
  XOR U12284 ( .A(DB[824]), .B(DB[793]), .Z(n8430) );
  AND U12285 ( .A(n412), .B(n8431), .Z(n8429) );
  XOR U12286 ( .A(n8432), .B(n8433), .Z(n8431) );
  XOR U12287 ( .A(DB[793]), .B(DB[762]), .Z(n8433) );
  AND U12288 ( .A(n416), .B(n8434), .Z(n8432) );
  XOR U12289 ( .A(n8435), .B(n8436), .Z(n8434) );
  XOR U12290 ( .A(DB[762]), .B(DB[731]), .Z(n8436) );
  AND U12291 ( .A(n420), .B(n8437), .Z(n8435) );
  XOR U12292 ( .A(n8438), .B(n8439), .Z(n8437) );
  XOR U12293 ( .A(DB[731]), .B(DB[700]), .Z(n8439) );
  AND U12294 ( .A(n424), .B(n8440), .Z(n8438) );
  XOR U12295 ( .A(n8441), .B(n8442), .Z(n8440) );
  XOR U12296 ( .A(DB[700]), .B(DB[669]), .Z(n8442) );
  AND U12297 ( .A(n428), .B(n8443), .Z(n8441) );
  XOR U12298 ( .A(n8444), .B(n8445), .Z(n8443) );
  XOR U12299 ( .A(DB[669]), .B(DB[638]), .Z(n8445) );
  AND U12300 ( .A(n432), .B(n8446), .Z(n8444) );
  XOR U12301 ( .A(n8447), .B(n8448), .Z(n8446) );
  XOR U12302 ( .A(DB[638]), .B(DB[607]), .Z(n8448) );
  AND U12303 ( .A(n436), .B(n8449), .Z(n8447) );
  XOR U12304 ( .A(n8450), .B(n8451), .Z(n8449) );
  XOR U12305 ( .A(DB[607]), .B(DB[576]), .Z(n8451) );
  AND U12306 ( .A(n440), .B(n8452), .Z(n8450) );
  XOR U12307 ( .A(n8453), .B(n8454), .Z(n8452) );
  XOR U12308 ( .A(DB[576]), .B(DB[545]), .Z(n8454) );
  AND U12309 ( .A(n444), .B(n8455), .Z(n8453) );
  XOR U12310 ( .A(n8456), .B(n8457), .Z(n8455) );
  XOR U12311 ( .A(DB[545]), .B(DB[514]), .Z(n8457) );
  AND U12312 ( .A(n448), .B(n8458), .Z(n8456) );
  XOR U12313 ( .A(n8459), .B(n8460), .Z(n8458) );
  XOR U12314 ( .A(DB[514]), .B(DB[483]), .Z(n8460) );
  AND U12315 ( .A(n452), .B(n8461), .Z(n8459) );
  XOR U12316 ( .A(n8462), .B(n8463), .Z(n8461) );
  XOR U12317 ( .A(DB[483]), .B(DB[452]), .Z(n8463) );
  AND U12318 ( .A(n456), .B(n8464), .Z(n8462) );
  XOR U12319 ( .A(n8465), .B(n8466), .Z(n8464) );
  XOR U12320 ( .A(DB[452]), .B(DB[421]), .Z(n8466) );
  AND U12321 ( .A(n460), .B(n8467), .Z(n8465) );
  XOR U12322 ( .A(n8468), .B(n8469), .Z(n8467) );
  XOR U12323 ( .A(DB[421]), .B(DB[390]), .Z(n8469) );
  AND U12324 ( .A(n464), .B(n8470), .Z(n8468) );
  XOR U12325 ( .A(n8471), .B(n8472), .Z(n8470) );
  XOR U12326 ( .A(DB[390]), .B(DB[359]), .Z(n8472) );
  AND U12327 ( .A(n468), .B(n8473), .Z(n8471) );
  XOR U12328 ( .A(n8474), .B(n8475), .Z(n8473) );
  XOR U12329 ( .A(DB[359]), .B(DB[328]), .Z(n8475) );
  AND U12330 ( .A(n472), .B(n8476), .Z(n8474) );
  XOR U12331 ( .A(n8477), .B(n8478), .Z(n8476) );
  XOR U12332 ( .A(DB[328]), .B(DB[297]), .Z(n8478) );
  AND U12333 ( .A(n476), .B(n8479), .Z(n8477) );
  XOR U12334 ( .A(n8480), .B(n8481), .Z(n8479) );
  XOR U12335 ( .A(DB[297]), .B(DB[266]), .Z(n8481) );
  AND U12336 ( .A(n480), .B(n8482), .Z(n8480) );
  XOR U12337 ( .A(n8483), .B(n8484), .Z(n8482) );
  XOR U12338 ( .A(DB[266]), .B(DB[235]), .Z(n8484) );
  AND U12339 ( .A(n484), .B(n8485), .Z(n8483) );
  XOR U12340 ( .A(n8486), .B(n8487), .Z(n8485) );
  XOR U12341 ( .A(DB[235]), .B(DB[204]), .Z(n8487) );
  AND U12342 ( .A(n488), .B(n8488), .Z(n8486) );
  XOR U12343 ( .A(n8489), .B(n8490), .Z(n8488) );
  XOR U12344 ( .A(DB[204]), .B(DB[173]), .Z(n8490) );
  AND U12345 ( .A(n492), .B(n8491), .Z(n8489) );
  XOR U12346 ( .A(n8492), .B(n8493), .Z(n8491) );
  XOR U12347 ( .A(DB[173]), .B(DB[142]), .Z(n8493) );
  AND U12348 ( .A(n496), .B(n8494), .Z(n8492) );
  XOR U12349 ( .A(n8495), .B(n8496), .Z(n8494) );
  XOR U12350 ( .A(DB[142]), .B(DB[111]), .Z(n8496) );
  AND U12351 ( .A(n500), .B(n8497), .Z(n8495) );
  XOR U12352 ( .A(n8498), .B(n8499), .Z(n8497) );
  XOR U12353 ( .A(DB[80]), .B(DB[111]), .Z(n8499) );
  AND U12354 ( .A(n504), .B(n8500), .Z(n8498) );
  XOR U12355 ( .A(n8501), .B(n8502), .Z(n8500) );
  XOR U12356 ( .A(DB[80]), .B(DB[49]), .Z(n8502) );
  AND U12357 ( .A(n508), .B(n8503), .Z(n8501) );
  XOR U12358 ( .A(DB[49]), .B(DB[18]), .Z(n8503) );
  XOR U12359 ( .A(DB[3954]), .B(n8504), .Z(min_val_out[17]) );
  AND U12360 ( .A(n2), .B(n8505), .Z(n8504) );
  XOR U12361 ( .A(n8506), .B(n8507), .Z(n8505) );
  XOR U12362 ( .A(n8508), .B(n8509), .Z(n8507) );
  IV U12363 ( .A(DB[3954]), .Z(n8508) );
  AND U12364 ( .A(n8), .B(n8510), .Z(n8506) );
  XOR U12365 ( .A(n8511), .B(n8512), .Z(n8510) );
  XOR U12366 ( .A(DB[3923]), .B(DB[3892]), .Z(n8512) );
  AND U12367 ( .A(n12), .B(n8513), .Z(n8511) );
  XOR U12368 ( .A(n8514), .B(n8515), .Z(n8513) );
  XOR U12369 ( .A(DB[3892]), .B(DB[3861]), .Z(n8515) );
  AND U12370 ( .A(n16), .B(n8516), .Z(n8514) );
  XOR U12371 ( .A(n8517), .B(n8518), .Z(n8516) );
  XOR U12372 ( .A(DB[3861]), .B(DB[3830]), .Z(n8518) );
  AND U12373 ( .A(n20), .B(n8519), .Z(n8517) );
  XOR U12374 ( .A(n8520), .B(n8521), .Z(n8519) );
  XOR U12375 ( .A(DB[3830]), .B(DB[3799]), .Z(n8521) );
  AND U12376 ( .A(n24), .B(n8522), .Z(n8520) );
  XOR U12377 ( .A(n8523), .B(n8524), .Z(n8522) );
  XOR U12378 ( .A(DB[3799]), .B(DB[3768]), .Z(n8524) );
  AND U12379 ( .A(n28), .B(n8525), .Z(n8523) );
  XOR U12380 ( .A(n8526), .B(n8527), .Z(n8525) );
  XOR U12381 ( .A(DB[3768]), .B(DB[3737]), .Z(n8527) );
  AND U12382 ( .A(n32), .B(n8528), .Z(n8526) );
  XOR U12383 ( .A(n8529), .B(n8530), .Z(n8528) );
  XOR U12384 ( .A(DB[3737]), .B(DB[3706]), .Z(n8530) );
  AND U12385 ( .A(n36), .B(n8531), .Z(n8529) );
  XOR U12386 ( .A(n8532), .B(n8533), .Z(n8531) );
  XOR U12387 ( .A(DB[3706]), .B(DB[3675]), .Z(n8533) );
  AND U12388 ( .A(n40), .B(n8534), .Z(n8532) );
  XOR U12389 ( .A(n8535), .B(n8536), .Z(n8534) );
  XOR U12390 ( .A(DB[3675]), .B(DB[3644]), .Z(n8536) );
  AND U12391 ( .A(n44), .B(n8537), .Z(n8535) );
  XOR U12392 ( .A(n8538), .B(n8539), .Z(n8537) );
  XOR U12393 ( .A(DB[3644]), .B(DB[3613]), .Z(n8539) );
  AND U12394 ( .A(n48), .B(n8540), .Z(n8538) );
  XOR U12395 ( .A(n8541), .B(n8542), .Z(n8540) );
  XOR U12396 ( .A(DB[3613]), .B(DB[3582]), .Z(n8542) );
  AND U12397 ( .A(n52), .B(n8543), .Z(n8541) );
  XOR U12398 ( .A(n8544), .B(n8545), .Z(n8543) );
  XOR U12399 ( .A(DB[3582]), .B(DB[3551]), .Z(n8545) );
  AND U12400 ( .A(n56), .B(n8546), .Z(n8544) );
  XOR U12401 ( .A(n8547), .B(n8548), .Z(n8546) );
  XOR U12402 ( .A(DB[3551]), .B(DB[3520]), .Z(n8548) );
  AND U12403 ( .A(n60), .B(n8549), .Z(n8547) );
  XOR U12404 ( .A(n8550), .B(n8551), .Z(n8549) );
  XOR U12405 ( .A(DB[3520]), .B(DB[3489]), .Z(n8551) );
  AND U12406 ( .A(n64), .B(n8552), .Z(n8550) );
  XOR U12407 ( .A(n8553), .B(n8554), .Z(n8552) );
  XOR U12408 ( .A(DB[3489]), .B(DB[3458]), .Z(n8554) );
  AND U12409 ( .A(n68), .B(n8555), .Z(n8553) );
  XOR U12410 ( .A(n8556), .B(n8557), .Z(n8555) );
  XOR U12411 ( .A(DB[3458]), .B(DB[3427]), .Z(n8557) );
  AND U12412 ( .A(n72), .B(n8558), .Z(n8556) );
  XOR U12413 ( .A(n8559), .B(n8560), .Z(n8558) );
  XOR U12414 ( .A(DB[3427]), .B(DB[3396]), .Z(n8560) );
  AND U12415 ( .A(n76), .B(n8561), .Z(n8559) );
  XOR U12416 ( .A(n8562), .B(n8563), .Z(n8561) );
  XOR U12417 ( .A(DB[3396]), .B(DB[3365]), .Z(n8563) );
  AND U12418 ( .A(n80), .B(n8564), .Z(n8562) );
  XOR U12419 ( .A(n8565), .B(n8566), .Z(n8564) );
  XOR U12420 ( .A(DB[3365]), .B(DB[3334]), .Z(n8566) );
  AND U12421 ( .A(n84), .B(n8567), .Z(n8565) );
  XOR U12422 ( .A(n8568), .B(n8569), .Z(n8567) );
  XOR U12423 ( .A(DB[3334]), .B(DB[3303]), .Z(n8569) );
  AND U12424 ( .A(n88), .B(n8570), .Z(n8568) );
  XOR U12425 ( .A(n8571), .B(n8572), .Z(n8570) );
  XOR U12426 ( .A(DB[3303]), .B(DB[3272]), .Z(n8572) );
  AND U12427 ( .A(n92), .B(n8573), .Z(n8571) );
  XOR U12428 ( .A(n8574), .B(n8575), .Z(n8573) );
  XOR U12429 ( .A(DB[3272]), .B(DB[3241]), .Z(n8575) );
  AND U12430 ( .A(n96), .B(n8576), .Z(n8574) );
  XOR U12431 ( .A(n8577), .B(n8578), .Z(n8576) );
  XOR U12432 ( .A(DB[3241]), .B(DB[3210]), .Z(n8578) );
  AND U12433 ( .A(n100), .B(n8579), .Z(n8577) );
  XOR U12434 ( .A(n8580), .B(n8581), .Z(n8579) );
  XOR U12435 ( .A(DB[3210]), .B(DB[3179]), .Z(n8581) );
  AND U12436 ( .A(n104), .B(n8582), .Z(n8580) );
  XOR U12437 ( .A(n8583), .B(n8584), .Z(n8582) );
  XOR U12438 ( .A(DB[3179]), .B(DB[3148]), .Z(n8584) );
  AND U12439 ( .A(n108), .B(n8585), .Z(n8583) );
  XOR U12440 ( .A(n8586), .B(n8587), .Z(n8585) );
  XOR U12441 ( .A(DB[3148]), .B(DB[3117]), .Z(n8587) );
  AND U12442 ( .A(n112), .B(n8588), .Z(n8586) );
  XOR U12443 ( .A(n8589), .B(n8590), .Z(n8588) );
  XOR U12444 ( .A(DB[3117]), .B(DB[3086]), .Z(n8590) );
  AND U12445 ( .A(n116), .B(n8591), .Z(n8589) );
  XOR U12446 ( .A(n8592), .B(n8593), .Z(n8591) );
  XOR U12447 ( .A(DB[3086]), .B(DB[3055]), .Z(n8593) );
  AND U12448 ( .A(n120), .B(n8594), .Z(n8592) );
  XOR U12449 ( .A(n8595), .B(n8596), .Z(n8594) );
  XOR U12450 ( .A(DB[3055]), .B(DB[3024]), .Z(n8596) );
  AND U12451 ( .A(n124), .B(n8597), .Z(n8595) );
  XOR U12452 ( .A(n8598), .B(n8599), .Z(n8597) );
  XOR U12453 ( .A(DB[3024]), .B(DB[2993]), .Z(n8599) );
  AND U12454 ( .A(n128), .B(n8600), .Z(n8598) );
  XOR U12455 ( .A(n8601), .B(n8602), .Z(n8600) );
  XOR U12456 ( .A(DB[2993]), .B(DB[2962]), .Z(n8602) );
  AND U12457 ( .A(n132), .B(n8603), .Z(n8601) );
  XOR U12458 ( .A(n8604), .B(n8605), .Z(n8603) );
  XOR U12459 ( .A(DB[2962]), .B(DB[2931]), .Z(n8605) );
  AND U12460 ( .A(n136), .B(n8606), .Z(n8604) );
  XOR U12461 ( .A(n8607), .B(n8608), .Z(n8606) );
  XOR U12462 ( .A(DB[2931]), .B(DB[2900]), .Z(n8608) );
  AND U12463 ( .A(n140), .B(n8609), .Z(n8607) );
  XOR U12464 ( .A(n8610), .B(n8611), .Z(n8609) );
  XOR U12465 ( .A(DB[2900]), .B(DB[2869]), .Z(n8611) );
  AND U12466 ( .A(n144), .B(n8612), .Z(n8610) );
  XOR U12467 ( .A(n8613), .B(n8614), .Z(n8612) );
  XOR U12468 ( .A(DB[2869]), .B(DB[2838]), .Z(n8614) );
  AND U12469 ( .A(n148), .B(n8615), .Z(n8613) );
  XOR U12470 ( .A(n8616), .B(n8617), .Z(n8615) );
  XOR U12471 ( .A(DB[2838]), .B(DB[2807]), .Z(n8617) );
  AND U12472 ( .A(n152), .B(n8618), .Z(n8616) );
  XOR U12473 ( .A(n8619), .B(n8620), .Z(n8618) );
  XOR U12474 ( .A(DB[2807]), .B(DB[2776]), .Z(n8620) );
  AND U12475 ( .A(n156), .B(n8621), .Z(n8619) );
  XOR U12476 ( .A(n8622), .B(n8623), .Z(n8621) );
  XOR U12477 ( .A(DB[2776]), .B(DB[2745]), .Z(n8623) );
  AND U12478 ( .A(n160), .B(n8624), .Z(n8622) );
  XOR U12479 ( .A(n8625), .B(n8626), .Z(n8624) );
  XOR U12480 ( .A(DB[2745]), .B(DB[2714]), .Z(n8626) );
  AND U12481 ( .A(n164), .B(n8627), .Z(n8625) );
  XOR U12482 ( .A(n8628), .B(n8629), .Z(n8627) );
  XOR U12483 ( .A(DB[2714]), .B(DB[2683]), .Z(n8629) );
  AND U12484 ( .A(n168), .B(n8630), .Z(n8628) );
  XOR U12485 ( .A(n8631), .B(n8632), .Z(n8630) );
  XOR U12486 ( .A(DB[2683]), .B(DB[2652]), .Z(n8632) );
  AND U12487 ( .A(n172), .B(n8633), .Z(n8631) );
  XOR U12488 ( .A(n8634), .B(n8635), .Z(n8633) );
  XOR U12489 ( .A(DB[2652]), .B(DB[2621]), .Z(n8635) );
  AND U12490 ( .A(n176), .B(n8636), .Z(n8634) );
  XOR U12491 ( .A(n8637), .B(n8638), .Z(n8636) );
  XOR U12492 ( .A(DB[2621]), .B(DB[2590]), .Z(n8638) );
  AND U12493 ( .A(n180), .B(n8639), .Z(n8637) );
  XOR U12494 ( .A(n8640), .B(n8641), .Z(n8639) );
  XOR U12495 ( .A(DB[2590]), .B(DB[2559]), .Z(n8641) );
  AND U12496 ( .A(n184), .B(n8642), .Z(n8640) );
  XOR U12497 ( .A(n8643), .B(n8644), .Z(n8642) );
  XOR U12498 ( .A(DB[2559]), .B(DB[2528]), .Z(n8644) );
  AND U12499 ( .A(n188), .B(n8645), .Z(n8643) );
  XOR U12500 ( .A(n8646), .B(n8647), .Z(n8645) );
  XOR U12501 ( .A(DB[2528]), .B(DB[2497]), .Z(n8647) );
  AND U12502 ( .A(n192), .B(n8648), .Z(n8646) );
  XOR U12503 ( .A(n8649), .B(n8650), .Z(n8648) );
  XOR U12504 ( .A(DB[2497]), .B(DB[2466]), .Z(n8650) );
  AND U12505 ( .A(n196), .B(n8651), .Z(n8649) );
  XOR U12506 ( .A(n8652), .B(n8653), .Z(n8651) );
  XOR U12507 ( .A(DB[2466]), .B(DB[2435]), .Z(n8653) );
  AND U12508 ( .A(n200), .B(n8654), .Z(n8652) );
  XOR U12509 ( .A(n8655), .B(n8656), .Z(n8654) );
  XOR U12510 ( .A(DB[2435]), .B(DB[2404]), .Z(n8656) );
  AND U12511 ( .A(n204), .B(n8657), .Z(n8655) );
  XOR U12512 ( .A(n8658), .B(n8659), .Z(n8657) );
  XOR U12513 ( .A(DB[2404]), .B(DB[2373]), .Z(n8659) );
  AND U12514 ( .A(n208), .B(n8660), .Z(n8658) );
  XOR U12515 ( .A(n8661), .B(n8662), .Z(n8660) );
  XOR U12516 ( .A(DB[2373]), .B(DB[2342]), .Z(n8662) );
  AND U12517 ( .A(n212), .B(n8663), .Z(n8661) );
  XOR U12518 ( .A(n8664), .B(n8665), .Z(n8663) );
  XOR U12519 ( .A(DB[2342]), .B(DB[2311]), .Z(n8665) );
  AND U12520 ( .A(n216), .B(n8666), .Z(n8664) );
  XOR U12521 ( .A(n8667), .B(n8668), .Z(n8666) );
  XOR U12522 ( .A(DB[2311]), .B(DB[2280]), .Z(n8668) );
  AND U12523 ( .A(n220), .B(n8669), .Z(n8667) );
  XOR U12524 ( .A(n8670), .B(n8671), .Z(n8669) );
  XOR U12525 ( .A(DB[2280]), .B(DB[2249]), .Z(n8671) );
  AND U12526 ( .A(n224), .B(n8672), .Z(n8670) );
  XOR U12527 ( .A(n8673), .B(n8674), .Z(n8672) );
  XOR U12528 ( .A(DB[2249]), .B(DB[2218]), .Z(n8674) );
  AND U12529 ( .A(n228), .B(n8675), .Z(n8673) );
  XOR U12530 ( .A(n8676), .B(n8677), .Z(n8675) );
  XOR U12531 ( .A(DB[2218]), .B(DB[2187]), .Z(n8677) );
  AND U12532 ( .A(n232), .B(n8678), .Z(n8676) );
  XOR U12533 ( .A(n8679), .B(n8680), .Z(n8678) );
  XOR U12534 ( .A(DB[2187]), .B(DB[2156]), .Z(n8680) );
  AND U12535 ( .A(n236), .B(n8681), .Z(n8679) );
  XOR U12536 ( .A(n8682), .B(n8683), .Z(n8681) );
  XOR U12537 ( .A(DB[2156]), .B(DB[2125]), .Z(n8683) );
  AND U12538 ( .A(n240), .B(n8684), .Z(n8682) );
  XOR U12539 ( .A(n8685), .B(n8686), .Z(n8684) );
  XOR U12540 ( .A(DB[2125]), .B(DB[2094]), .Z(n8686) );
  AND U12541 ( .A(n244), .B(n8687), .Z(n8685) );
  XOR U12542 ( .A(n8688), .B(n8689), .Z(n8687) );
  XOR U12543 ( .A(DB[2094]), .B(DB[2063]), .Z(n8689) );
  AND U12544 ( .A(n248), .B(n8690), .Z(n8688) );
  XOR U12545 ( .A(n8691), .B(n8692), .Z(n8690) );
  XOR U12546 ( .A(DB[2063]), .B(DB[2032]), .Z(n8692) );
  AND U12547 ( .A(n252), .B(n8693), .Z(n8691) );
  XOR U12548 ( .A(n8694), .B(n8695), .Z(n8693) );
  XOR U12549 ( .A(DB[2032]), .B(DB[2001]), .Z(n8695) );
  AND U12550 ( .A(n256), .B(n8696), .Z(n8694) );
  XOR U12551 ( .A(n8697), .B(n8698), .Z(n8696) );
  XOR U12552 ( .A(DB[2001]), .B(DB[1970]), .Z(n8698) );
  AND U12553 ( .A(n260), .B(n8699), .Z(n8697) );
  XOR U12554 ( .A(n8700), .B(n8701), .Z(n8699) );
  XOR U12555 ( .A(DB[1970]), .B(DB[1939]), .Z(n8701) );
  AND U12556 ( .A(n264), .B(n8702), .Z(n8700) );
  XOR U12557 ( .A(n8703), .B(n8704), .Z(n8702) );
  XOR U12558 ( .A(DB[1939]), .B(DB[1908]), .Z(n8704) );
  AND U12559 ( .A(n268), .B(n8705), .Z(n8703) );
  XOR U12560 ( .A(n8706), .B(n8707), .Z(n8705) );
  XOR U12561 ( .A(DB[1908]), .B(DB[1877]), .Z(n8707) );
  AND U12562 ( .A(n272), .B(n8708), .Z(n8706) );
  XOR U12563 ( .A(n8709), .B(n8710), .Z(n8708) );
  XOR U12564 ( .A(DB[1877]), .B(DB[1846]), .Z(n8710) );
  AND U12565 ( .A(n276), .B(n8711), .Z(n8709) );
  XOR U12566 ( .A(n8712), .B(n8713), .Z(n8711) );
  XOR U12567 ( .A(DB[1846]), .B(DB[1815]), .Z(n8713) );
  AND U12568 ( .A(n280), .B(n8714), .Z(n8712) );
  XOR U12569 ( .A(n8715), .B(n8716), .Z(n8714) );
  XOR U12570 ( .A(DB[1815]), .B(DB[1784]), .Z(n8716) );
  AND U12571 ( .A(n284), .B(n8717), .Z(n8715) );
  XOR U12572 ( .A(n8718), .B(n8719), .Z(n8717) );
  XOR U12573 ( .A(DB[1784]), .B(DB[1753]), .Z(n8719) );
  AND U12574 ( .A(n288), .B(n8720), .Z(n8718) );
  XOR U12575 ( .A(n8721), .B(n8722), .Z(n8720) );
  XOR U12576 ( .A(DB[1753]), .B(DB[1722]), .Z(n8722) );
  AND U12577 ( .A(n292), .B(n8723), .Z(n8721) );
  XOR U12578 ( .A(n8724), .B(n8725), .Z(n8723) );
  XOR U12579 ( .A(DB[1722]), .B(DB[1691]), .Z(n8725) );
  AND U12580 ( .A(n296), .B(n8726), .Z(n8724) );
  XOR U12581 ( .A(n8727), .B(n8728), .Z(n8726) );
  XOR U12582 ( .A(DB[1691]), .B(DB[1660]), .Z(n8728) );
  AND U12583 ( .A(n300), .B(n8729), .Z(n8727) );
  XOR U12584 ( .A(n8730), .B(n8731), .Z(n8729) );
  XOR U12585 ( .A(DB[1660]), .B(DB[1629]), .Z(n8731) );
  AND U12586 ( .A(n304), .B(n8732), .Z(n8730) );
  XOR U12587 ( .A(n8733), .B(n8734), .Z(n8732) );
  XOR U12588 ( .A(DB[1629]), .B(DB[1598]), .Z(n8734) );
  AND U12589 ( .A(n308), .B(n8735), .Z(n8733) );
  XOR U12590 ( .A(n8736), .B(n8737), .Z(n8735) );
  XOR U12591 ( .A(DB[1598]), .B(DB[1567]), .Z(n8737) );
  AND U12592 ( .A(n312), .B(n8738), .Z(n8736) );
  XOR U12593 ( .A(n8739), .B(n8740), .Z(n8738) );
  XOR U12594 ( .A(DB[1567]), .B(DB[1536]), .Z(n8740) );
  AND U12595 ( .A(n316), .B(n8741), .Z(n8739) );
  XOR U12596 ( .A(n8742), .B(n8743), .Z(n8741) );
  XOR U12597 ( .A(DB[1536]), .B(DB[1505]), .Z(n8743) );
  AND U12598 ( .A(n320), .B(n8744), .Z(n8742) );
  XOR U12599 ( .A(n8745), .B(n8746), .Z(n8744) );
  XOR U12600 ( .A(DB[1505]), .B(DB[1474]), .Z(n8746) );
  AND U12601 ( .A(n324), .B(n8747), .Z(n8745) );
  XOR U12602 ( .A(n8748), .B(n8749), .Z(n8747) );
  XOR U12603 ( .A(DB[1474]), .B(DB[1443]), .Z(n8749) );
  AND U12604 ( .A(n328), .B(n8750), .Z(n8748) );
  XOR U12605 ( .A(n8751), .B(n8752), .Z(n8750) );
  XOR U12606 ( .A(DB[1443]), .B(DB[1412]), .Z(n8752) );
  AND U12607 ( .A(n332), .B(n8753), .Z(n8751) );
  XOR U12608 ( .A(n8754), .B(n8755), .Z(n8753) );
  XOR U12609 ( .A(DB[1412]), .B(DB[1381]), .Z(n8755) );
  AND U12610 ( .A(n336), .B(n8756), .Z(n8754) );
  XOR U12611 ( .A(n8757), .B(n8758), .Z(n8756) );
  XOR U12612 ( .A(DB[1381]), .B(DB[1350]), .Z(n8758) );
  AND U12613 ( .A(n340), .B(n8759), .Z(n8757) );
  XOR U12614 ( .A(n8760), .B(n8761), .Z(n8759) );
  XOR U12615 ( .A(DB[1350]), .B(DB[1319]), .Z(n8761) );
  AND U12616 ( .A(n344), .B(n8762), .Z(n8760) );
  XOR U12617 ( .A(n8763), .B(n8764), .Z(n8762) );
  XOR U12618 ( .A(DB[1319]), .B(DB[1288]), .Z(n8764) );
  AND U12619 ( .A(n348), .B(n8765), .Z(n8763) );
  XOR U12620 ( .A(n8766), .B(n8767), .Z(n8765) );
  XOR U12621 ( .A(DB[1288]), .B(DB[1257]), .Z(n8767) );
  AND U12622 ( .A(n352), .B(n8768), .Z(n8766) );
  XOR U12623 ( .A(n8769), .B(n8770), .Z(n8768) );
  XOR U12624 ( .A(DB[1257]), .B(DB[1226]), .Z(n8770) );
  AND U12625 ( .A(n356), .B(n8771), .Z(n8769) );
  XOR U12626 ( .A(n8772), .B(n8773), .Z(n8771) );
  XOR U12627 ( .A(DB[1226]), .B(DB[1195]), .Z(n8773) );
  AND U12628 ( .A(n360), .B(n8774), .Z(n8772) );
  XOR U12629 ( .A(n8775), .B(n8776), .Z(n8774) );
  XOR U12630 ( .A(DB[1195]), .B(DB[1164]), .Z(n8776) );
  AND U12631 ( .A(n364), .B(n8777), .Z(n8775) );
  XOR U12632 ( .A(n8778), .B(n8779), .Z(n8777) );
  XOR U12633 ( .A(DB[1164]), .B(DB[1133]), .Z(n8779) );
  AND U12634 ( .A(n368), .B(n8780), .Z(n8778) );
  XOR U12635 ( .A(n8781), .B(n8782), .Z(n8780) );
  XOR U12636 ( .A(DB[1133]), .B(DB[1102]), .Z(n8782) );
  AND U12637 ( .A(n372), .B(n8783), .Z(n8781) );
  XOR U12638 ( .A(n8784), .B(n8785), .Z(n8783) );
  XOR U12639 ( .A(DB[1102]), .B(DB[1071]), .Z(n8785) );
  AND U12640 ( .A(n376), .B(n8786), .Z(n8784) );
  XOR U12641 ( .A(n8787), .B(n8788), .Z(n8786) );
  XOR U12642 ( .A(DB[1071]), .B(DB[1040]), .Z(n8788) );
  AND U12643 ( .A(n380), .B(n8789), .Z(n8787) );
  XOR U12644 ( .A(n8790), .B(n8791), .Z(n8789) );
  XOR U12645 ( .A(DB[1040]), .B(DB[1009]), .Z(n8791) );
  AND U12646 ( .A(n384), .B(n8792), .Z(n8790) );
  XOR U12647 ( .A(n8793), .B(n8794), .Z(n8792) );
  XOR U12648 ( .A(DB[978]), .B(DB[1009]), .Z(n8794) );
  AND U12649 ( .A(n388), .B(n8795), .Z(n8793) );
  XOR U12650 ( .A(n8796), .B(n8797), .Z(n8795) );
  XOR U12651 ( .A(DB[978]), .B(DB[947]), .Z(n8797) );
  AND U12652 ( .A(n392), .B(n8798), .Z(n8796) );
  XOR U12653 ( .A(n8799), .B(n8800), .Z(n8798) );
  XOR U12654 ( .A(DB[947]), .B(DB[916]), .Z(n8800) );
  AND U12655 ( .A(n396), .B(n8801), .Z(n8799) );
  XOR U12656 ( .A(n8802), .B(n8803), .Z(n8801) );
  XOR U12657 ( .A(DB[916]), .B(DB[885]), .Z(n8803) );
  AND U12658 ( .A(n400), .B(n8804), .Z(n8802) );
  XOR U12659 ( .A(n8805), .B(n8806), .Z(n8804) );
  XOR U12660 ( .A(DB[885]), .B(DB[854]), .Z(n8806) );
  AND U12661 ( .A(n404), .B(n8807), .Z(n8805) );
  XOR U12662 ( .A(n8808), .B(n8809), .Z(n8807) );
  XOR U12663 ( .A(DB[854]), .B(DB[823]), .Z(n8809) );
  AND U12664 ( .A(n408), .B(n8810), .Z(n8808) );
  XOR U12665 ( .A(n8811), .B(n8812), .Z(n8810) );
  XOR U12666 ( .A(DB[823]), .B(DB[792]), .Z(n8812) );
  AND U12667 ( .A(n412), .B(n8813), .Z(n8811) );
  XOR U12668 ( .A(n8814), .B(n8815), .Z(n8813) );
  XOR U12669 ( .A(DB[792]), .B(DB[761]), .Z(n8815) );
  AND U12670 ( .A(n416), .B(n8816), .Z(n8814) );
  XOR U12671 ( .A(n8817), .B(n8818), .Z(n8816) );
  XOR U12672 ( .A(DB[761]), .B(DB[730]), .Z(n8818) );
  AND U12673 ( .A(n420), .B(n8819), .Z(n8817) );
  XOR U12674 ( .A(n8820), .B(n8821), .Z(n8819) );
  XOR U12675 ( .A(DB[730]), .B(DB[699]), .Z(n8821) );
  AND U12676 ( .A(n424), .B(n8822), .Z(n8820) );
  XOR U12677 ( .A(n8823), .B(n8824), .Z(n8822) );
  XOR U12678 ( .A(DB[699]), .B(DB[668]), .Z(n8824) );
  AND U12679 ( .A(n428), .B(n8825), .Z(n8823) );
  XOR U12680 ( .A(n8826), .B(n8827), .Z(n8825) );
  XOR U12681 ( .A(DB[668]), .B(DB[637]), .Z(n8827) );
  AND U12682 ( .A(n432), .B(n8828), .Z(n8826) );
  XOR U12683 ( .A(n8829), .B(n8830), .Z(n8828) );
  XOR U12684 ( .A(DB[637]), .B(DB[606]), .Z(n8830) );
  AND U12685 ( .A(n436), .B(n8831), .Z(n8829) );
  XOR U12686 ( .A(n8832), .B(n8833), .Z(n8831) );
  XOR U12687 ( .A(DB[606]), .B(DB[575]), .Z(n8833) );
  AND U12688 ( .A(n440), .B(n8834), .Z(n8832) );
  XOR U12689 ( .A(n8835), .B(n8836), .Z(n8834) );
  XOR U12690 ( .A(DB[575]), .B(DB[544]), .Z(n8836) );
  AND U12691 ( .A(n444), .B(n8837), .Z(n8835) );
  XOR U12692 ( .A(n8838), .B(n8839), .Z(n8837) );
  XOR U12693 ( .A(DB[544]), .B(DB[513]), .Z(n8839) );
  AND U12694 ( .A(n448), .B(n8840), .Z(n8838) );
  XOR U12695 ( .A(n8841), .B(n8842), .Z(n8840) );
  XOR U12696 ( .A(DB[513]), .B(DB[482]), .Z(n8842) );
  AND U12697 ( .A(n452), .B(n8843), .Z(n8841) );
  XOR U12698 ( .A(n8844), .B(n8845), .Z(n8843) );
  XOR U12699 ( .A(DB[482]), .B(DB[451]), .Z(n8845) );
  AND U12700 ( .A(n456), .B(n8846), .Z(n8844) );
  XOR U12701 ( .A(n8847), .B(n8848), .Z(n8846) );
  XOR U12702 ( .A(DB[451]), .B(DB[420]), .Z(n8848) );
  AND U12703 ( .A(n460), .B(n8849), .Z(n8847) );
  XOR U12704 ( .A(n8850), .B(n8851), .Z(n8849) );
  XOR U12705 ( .A(DB[420]), .B(DB[389]), .Z(n8851) );
  AND U12706 ( .A(n464), .B(n8852), .Z(n8850) );
  XOR U12707 ( .A(n8853), .B(n8854), .Z(n8852) );
  XOR U12708 ( .A(DB[389]), .B(DB[358]), .Z(n8854) );
  AND U12709 ( .A(n468), .B(n8855), .Z(n8853) );
  XOR U12710 ( .A(n8856), .B(n8857), .Z(n8855) );
  XOR U12711 ( .A(DB[358]), .B(DB[327]), .Z(n8857) );
  AND U12712 ( .A(n472), .B(n8858), .Z(n8856) );
  XOR U12713 ( .A(n8859), .B(n8860), .Z(n8858) );
  XOR U12714 ( .A(DB[327]), .B(DB[296]), .Z(n8860) );
  AND U12715 ( .A(n476), .B(n8861), .Z(n8859) );
  XOR U12716 ( .A(n8862), .B(n8863), .Z(n8861) );
  XOR U12717 ( .A(DB[296]), .B(DB[265]), .Z(n8863) );
  AND U12718 ( .A(n480), .B(n8864), .Z(n8862) );
  XOR U12719 ( .A(n8865), .B(n8866), .Z(n8864) );
  XOR U12720 ( .A(DB[265]), .B(DB[234]), .Z(n8866) );
  AND U12721 ( .A(n484), .B(n8867), .Z(n8865) );
  XOR U12722 ( .A(n8868), .B(n8869), .Z(n8867) );
  XOR U12723 ( .A(DB[234]), .B(DB[203]), .Z(n8869) );
  AND U12724 ( .A(n488), .B(n8870), .Z(n8868) );
  XOR U12725 ( .A(n8871), .B(n8872), .Z(n8870) );
  XOR U12726 ( .A(DB[203]), .B(DB[172]), .Z(n8872) );
  AND U12727 ( .A(n492), .B(n8873), .Z(n8871) );
  XOR U12728 ( .A(n8874), .B(n8875), .Z(n8873) );
  XOR U12729 ( .A(DB[172]), .B(DB[141]), .Z(n8875) );
  AND U12730 ( .A(n496), .B(n8876), .Z(n8874) );
  XOR U12731 ( .A(n8877), .B(n8878), .Z(n8876) );
  XOR U12732 ( .A(DB[141]), .B(DB[110]), .Z(n8878) );
  AND U12733 ( .A(n500), .B(n8879), .Z(n8877) );
  XOR U12734 ( .A(n8880), .B(n8881), .Z(n8879) );
  XOR U12735 ( .A(DB[79]), .B(DB[110]), .Z(n8881) );
  AND U12736 ( .A(n504), .B(n8882), .Z(n8880) );
  XOR U12737 ( .A(n8883), .B(n8884), .Z(n8882) );
  XOR U12738 ( .A(DB[79]), .B(DB[48]), .Z(n8884) );
  AND U12739 ( .A(n508), .B(n8885), .Z(n8883) );
  XOR U12740 ( .A(DB[48]), .B(DB[17]), .Z(n8885) );
  XOR U12741 ( .A(DB[3953]), .B(n8886), .Z(min_val_out[16]) );
  AND U12742 ( .A(n2), .B(n8887), .Z(n8886) );
  XOR U12743 ( .A(n8888), .B(n8889), .Z(n8887) );
  XOR U12744 ( .A(n8890), .B(n8891), .Z(n8889) );
  IV U12745 ( .A(DB[3953]), .Z(n8890) );
  AND U12746 ( .A(n8), .B(n8892), .Z(n8888) );
  XOR U12747 ( .A(n8893), .B(n8894), .Z(n8892) );
  XOR U12748 ( .A(DB[3922]), .B(DB[3891]), .Z(n8894) );
  AND U12749 ( .A(n12), .B(n8895), .Z(n8893) );
  XOR U12750 ( .A(n8896), .B(n8897), .Z(n8895) );
  XOR U12751 ( .A(DB[3891]), .B(DB[3860]), .Z(n8897) );
  AND U12752 ( .A(n16), .B(n8898), .Z(n8896) );
  XOR U12753 ( .A(n8899), .B(n8900), .Z(n8898) );
  XOR U12754 ( .A(DB[3860]), .B(DB[3829]), .Z(n8900) );
  AND U12755 ( .A(n20), .B(n8901), .Z(n8899) );
  XOR U12756 ( .A(n8902), .B(n8903), .Z(n8901) );
  XOR U12757 ( .A(DB[3829]), .B(DB[3798]), .Z(n8903) );
  AND U12758 ( .A(n24), .B(n8904), .Z(n8902) );
  XOR U12759 ( .A(n8905), .B(n8906), .Z(n8904) );
  XOR U12760 ( .A(DB[3798]), .B(DB[3767]), .Z(n8906) );
  AND U12761 ( .A(n28), .B(n8907), .Z(n8905) );
  XOR U12762 ( .A(n8908), .B(n8909), .Z(n8907) );
  XOR U12763 ( .A(DB[3767]), .B(DB[3736]), .Z(n8909) );
  AND U12764 ( .A(n32), .B(n8910), .Z(n8908) );
  XOR U12765 ( .A(n8911), .B(n8912), .Z(n8910) );
  XOR U12766 ( .A(DB[3736]), .B(DB[3705]), .Z(n8912) );
  AND U12767 ( .A(n36), .B(n8913), .Z(n8911) );
  XOR U12768 ( .A(n8914), .B(n8915), .Z(n8913) );
  XOR U12769 ( .A(DB[3705]), .B(DB[3674]), .Z(n8915) );
  AND U12770 ( .A(n40), .B(n8916), .Z(n8914) );
  XOR U12771 ( .A(n8917), .B(n8918), .Z(n8916) );
  XOR U12772 ( .A(DB[3674]), .B(DB[3643]), .Z(n8918) );
  AND U12773 ( .A(n44), .B(n8919), .Z(n8917) );
  XOR U12774 ( .A(n8920), .B(n8921), .Z(n8919) );
  XOR U12775 ( .A(DB[3643]), .B(DB[3612]), .Z(n8921) );
  AND U12776 ( .A(n48), .B(n8922), .Z(n8920) );
  XOR U12777 ( .A(n8923), .B(n8924), .Z(n8922) );
  XOR U12778 ( .A(DB[3612]), .B(DB[3581]), .Z(n8924) );
  AND U12779 ( .A(n52), .B(n8925), .Z(n8923) );
  XOR U12780 ( .A(n8926), .B(n8927), .Z(n8925) );
  XOR U12781 ( .A(DB[3581]), .B(DB[3550]), .Z(n8927) );
  AND U12782 ( .A(n56), .B(n8928), .Z(n8926) );
  XOR U12783 ( .A(n8929), .B(n8930), .Z(n8928) );
  XOR U12784 ( .A(DB[3550]), .B(DB[3519]), .Z(n8930) );
  AND U12785 ( .A(n60), .B(n8931), .Z(n8929) );
  XOR U12786 ( .A(n8932), .B(n8933), .Z(n8931) );
  XOR U12787 ( .A(DB[3519]), .B(DB[3488]), .Z(n8933) );
  AND U12788 ( .A(n64), .B(n8934), .Z(n8932) );
  XOR U12789 ( .A(n8935), .B(n8936), .Z(n8934) );
  XOR U12790 ( .A(DB[3488]), .B(DB[3457]), .Z(n8936) );
  AND U12791 ( .A(n68), .B(n8937), .Z(n8935) );
  XOR U12792 ( .A(n8938), .B(n8939), .Z(n8937) );
  XOR U12793 ( .A(DB[3457]), .B(DB[3426]), .Z(n8939) );
  AND U12794 ( .A(n72), .B(n8940), .Z(n8938) );
  XOR U12795 ( .A(n8941), .B(n8942), .Z(n8940) );
  XOR U12796 ( .A(DB[3426]), .B(DB[3395]), .Z(n8942) );
  AND U12797 ( .A(n76), .B(n8943), .Z(n8941) );
  XOR U12798 ( .A(n8944), .B(n8945), .Z(n8943) );
  XOR U12799 ( .A(DB[3395]), .B(DB[3364]), .Z(n8945) );
  AND U12800 ( .A(n80), .B(n8946), .Z(n8944) );
  XOR U12801 ( .A(n8947), .B(n8948), .Z(n8946) );
  XOR U12802 ( .A(DB[3364]), .B(DB[3333]), .Z(n8948) );
  AND U12803 ( .A(n84), .B(n8949), .Z(n8947) );
  XOR U12804 ( .A(n8950), .B(n8951), .Z(n8949) );
  XOR U12805 ( .A(DB[3333]), .B(DB[3302]), .Z(n8951) );
  AND U12806 ( .A(n88), .B(n8952), .Z(n8950) );
  XOR U12807 ( .A(n8953), .B(n8954), .Z(n8952) );
  XOR U12808 ( .A(DB[3302]), .B(DB[3271]), .Z(n8954) );
  AND U12809 ( .A(n92), .B(n8955), .Z(n8953) );
  XOR U12810 ( .A(n8956), .B(n8957), .Z(n8955) );
  XOR U12811 ( .A(DB[3271]), .B(DB[3240]), .Z(n8957) );
  AND U12812 ( .A(n96), .B(n8958), .Z(n8956) );
  XOR U12813 ( .A(n8959), .B(n8960), .Z(n8958) );
  XOR U12814 ( .A(DB[3240]), .B(DB[3209]), .Z(n8960) );
  AND U12815 ( .A(n100), .B(n8961), .Z(n8959) );
  XOR U12816 ( .A(n8962), .B(n8963), .Z(n8961) );
  XOR U12817 ( .A(DB[3209]), .B(DB[3178]), .Z(n8963) );
  AND U12818 ( .A(n104), .B(n8964), .Z(n8962) );
  XOR U12819 ( .A(n8965), .B(n8966), .Z(n8964) );
  XOR U12820 ( .A(DB[3178]), .B(DB[3147]), .Z(n8966) );
  AND U12821 ( .A(n108), .B(n8967), .Z(n8965) );
  XOR U12822 ( .A(n8968), .B(n8969), .Z(n8967) );
  XOR U12823 ( .A(DB[3147]), .B(DB[3116]), .Z(n8969) );
  AND U12824 ( .A(n112), .B(n8970), .Z(n8968) );
  XOR U12825 ( .A(n8971), .B(n8972), .Z(n8970) );
  XOR U12826 ( .A(DB[3116]), .B(DB[3085]), .Z(n8972) );
  AND U12827 ( .A(n116), .B(n8973), .Z(n8971) );
  XOR U12828 ( .A(n8974), .B(n8975), .Z(n8973) );
  XOR U12829 ( .A(DB[3085]), .B(DB[3054]), .Z(n8975) );
  AND U12830 ( .A(n120), .B(n8976), .Z(n8974) );
  XOR U12831 ( .A(n8977), .B(n8978), .Z(n8976) );
  XOR U12832 ( .A(DB[3054]), .B(DB[3023]), .Z(n8978) );
  AND U12833 ( .A(n124), .B(n8979), .Z(n8977) );
  XOR U12834 ( .A(n8980), .B(n8981), .Z(n8979) );
  XOR U12835 ( .A(DB[3023]), .B(DB[2992]), .Z(n8981) );
  AND U12836 ( .A(n128), .B(n8982), .Z(n8980) );
  XOR U12837 ( .A(n8983), .B(n8984), .Z(n8982) );
  XOR U12838 ( .A(DB[2992]), .B(DB[2961]), .Z(n8984) );
  AND U12839 ( .A(n132), .B(n8985), .Z(n8983) );
  XOR U12840 ( .A(n8986), .B(n8987), .Z(n8985) );
  XOR U12841 ( .A(DB[2961]), .B(DB[2930]), .Z(n8987) );
  AND U12842 ( .A(n136), .B(n8988), .Z(n8986) );
  XOR U12843 ( .A(n8989), .B(n8990), .Z(n8988) );
  XOR U12844 ( .A(DB[2930]), .B(DB[2899]), .Z(n8990) );
  AND U12845 ( .A(n140), .B(n8991), .Z(n8989) );
  XOR U12846 ( .A(n8992), .B(n8993), .Z(n8991) );
  XOR U12847 ( .A(DB[2899]), .B(DB[2868]), .Z(n8993) );
  AND U12848 ( .A(n144), .B(n8994), .Z(n8992) );
  XOR U12849 ( .A(n8995), .B(n8996), .Z(n8994) );
  XOR U12850 ( .A(DB[2868]), .B(DB[2837]), .Z(n8996) );
  AND U12851 ( .A(n148), .B(n8997), .Z(n8995) );
  XOR U12852 ( .A(n8998), .B(n8999), .Z(n8997) );
  XOR U12853 ( .A(DB[2837]), .B(DB[2806]), .Z(n8999) );
  AND U12854 ( .A(n152), .B(n9000), .Z(n8998) );
  XOR U12855 ( .A(n9001), .B(n9002), .Z(n9000) );
  XOR U12856 ( .A(DB[2806]), .B(DB[2775]), .Z(n9002) );
  AND U12857 ( .A(n156), .B(n9003), .Z(n9001) );
  XOR U12858 ( .A(n9004), .B(n9005), .Z(n9003) );
  XOR U12859 ( .A(DB[2775]), .B(DB[2744]), .Z(n9005) );
  AND U12860 ( .A(n160), .B(n9006), .Z(n9004) );
  XOR U12861 ( .A(n9007), .B(n9008), .Z(n9006) );
  XOR U12862 ( .A(DB[2744]), .B(DB[2713]), .Z(n9008) );
  AND U12863 ( .A(n164), .B(n9009), .Z(n9007) );
  XOR U12864 ( .A(n9010), .B(n9011), .Z(n9009) );
  XOR U12865 ( .A(DB[2713]), .B(DB[2682]), .Z(n9011) );
  AND U12866 ( .A(n168), .B(n9012), .Z(n9010) );
  XOR U12867 ( .A(n9013), .B(n9014), .Z(n9012) );
  XOR U12868 ( .A(DB[2682]), .B(DB[2651]), .Z(n9014) );
  AND U12869 ( .A(n172), .B(n9015), .Z(n9013) );
  XOR U12870 ( .A(n9016), .B(n9017), .Z(n9015) );
  XOR U12871 ( .A(DB[2651]), .B(DB[2620]), .Z(n9017) );
  AND U12872 ( .A(n176), .B(n9018), .Z(n9016) );
  XOR U12873 ( .A(n9019), .B(n9020), .Z(n9018) );
  XOR U12874 ( .A(DB[2620]), .B(DB[2589]), .Z(n9020) );
  AND U12875 ( .A(n180), .B(n9021), .Z(n9019) );
  XOR U12876 ( .A(n9022), .B(n9023), .Z(n9021) );
  XOR U12877 ( .A(DB[2589]), .B(DB[2558]), .Z(n9023) );
  AND U12878 ( .A(n184), .B(n9024), .Z(n9022) );
  XOR U12879 ( .A(n9025), .B(n9026), .Z(n9024) );
  XOR U12880 ( .A(DB[2558]), .B(DB[2527]), .Z(n9026) );
  AND U12881 ( .A(n188), .B(n9027), .Z(n9025) );
  XOR U12882 ( .A(n9028), .B(n9029), .Z(n9027) );
  XOR U12883 ( .A(DB[2527]), .B(DB[2496]), .Z(n9029) );
  AND U12884 ( .A(n192), .B(n9030), .Z(n9028) );
  XOR U12885 ( .A(n9031), .B(n9032), .Z(n9030) );
  XOR U12886 ( .A(DB[2496]), .B(DB[2465]), .Z(n9032) );
  AND U12887 ( .A(n196), .B(n9033), .Z(n9031) );
  XOR U12888 ( .A(n9034), .B(n9035), .Z(n9033) );
  XOR U12889 ( .A(DB[2465]), .B(DB[2434]), .Z(n9035) );
  AND U12890 ( .A(n200), .B(n9036), .Z(n9034) );
  XOR U12891 ( .A(n9037), .B(n9038), .Z(n9036) );
  XOR U12892 ( .A(DB[2434]), .B(DB[2403]), .Z(n9038) );
  AND U12893 ( .A(n204), .B(n9039), .Z(n9037) );
  XOR U12894 ( .A(n9040), .B(n9041), .Z(n9039) );
  XOR U12895 ( .A(DB[2403]), .B(DB[2372]), .Z(n9041) );
  AND U12896 ( .A(n208), .B(n9042), .Z(n9040) );
  XOR U12897 ( .A(n9043), .B(n9044), .Z(n9042) );
  XOR U12898 ( .A(DB[2372]), .B(DB[2341]), .Z(n9044) );
  AND U12899 ( .A(n212), .B(n9045), .Z(n9043) );
  XOR U12900 ( .A(n9046), .B(n9047), .Z(n9045) );
  XOR U12901 ( .A(DB[2341]), .B(DB[2310]), .Z(n9047) );
  AND U12902 ( .A(n216), .B(n9048), .Z(n9046) );
  XOR U12903 ( .A(n9049), .B(n9050), .Z(n9048) );
  XOR U12904 ( .A(DB[2310]), .B(DB[2279]), .Z(n9050) );
  AND U12905 ( .A(n220), .B(n9051), .Z(n9049) );
  XOR U12906 ( .A(n9052), .B(n9053), .Z(n9051) );
  XOR U12907 ( .A(DB[2279]), .B(DB[2248]), .Z(n9053) );
  AND U12908 ( .A(n224), .B(n9054), .Z(n9052) );
  XOR U12909 ( .A(n9055), .B(n9056), .Z(n9054) );
  XOR U12910 ( .A(DB[2248]), .B(DB[2217]), .Z(n9056) );
  AND U12911 ( .A(n228), .B(n9057), .Z(n9055) );
  XOR U12912 ( .A(n9058), .B(n9059), .Z(n9057) );
  XOR U12913 ( .A(DB[2217]), .B(DB[2186]), .Z(n9059) );
  AND U12914 ( .A(n232), .B(n9060), .Z(n9058) );
  XOR U12915 ( .A(n9061), .B(n9062), .Z(n9060) );
  XOR U12916 ( .A(DB[2186]), .B(DB[2155]), .Z(n9062) );
  AND U12917 ( .A(n236), .B(n9063), .Z(n9061) );
  XOR U12918 ( .A(n9064), .B(n9065), .Z(n9063) );
  XOR U12919 ( .A(DB[2155]), .B(DB[2124]), .Z(n9065) );
  AND U12920 ( .A(n240), .B(n9066), .Z(n9064) );
  XOR U12921 ( .A(n9067), .B(n9068), .Z(n9066) );
  XOR U12922 ( .A(DB[2124]), .B(DB[2093]), .Z(n9068) );
  AND U12923 ( .A(n244), .B(n9069), .Z(n9067) );
  XOR U12924 ( .A(n9070), .B(n9071), .Z(n9069) );
  XOR U12925 ( .A(DB[2093]), .B(DB[2062]), .Z(n9071) );
  AND U12926 ( .A(n248), .B(n9072), .Z(n9070) );
  XOR U12927 ( .A(n9073), .B(n9074), .Z(n9072) );
  XOR U12928 ( .A(DB[2062]), .B(DB[2031]), .Z(n9074) );
  AND U12929 ( .A(n252), .B(n9075), .Z(n9073) );
  XOR U12930 ( .A(n9076), .B(n9077), .Z(n9075) );
  XOR U12931 ( .A(DB[2031]), .B(DB[2000]), .Z(n9077) );
  AND U12932 ( .A(n256), .B(n9078), .Z(n9076) );
  XOR U12933 ( .A(n9079), .B(n9080), .Z(n9078) );
  XOR U12934 ( .A(DB[2000]), .B(DB[1969]), .Z(n9080) );
  AND U12935 ( .A(n260), .B(n9081), .Z(n9079) );
  XOR U12936 ( .A(n9082), .B(n9083), .Z(n9081) );
  XOR U12937 ( .A(DB[1969]), .B(DB[1938]), .Z(n9083) );
  AND U12938 ( .A(n264), .B(n9084), .Z(n9082) );
  XOR U12939 ( .A(n9085), .B(n9086), .Z(n9084) );
  XOR U12940 ( .A(DB[1938]), .B(DB[1907]), .Z(n9086) );
  AND U12941 ( .A(n268), .B(n9087), .Z(n9085) );
  XOR U12942 ( .A(n9088), .B(n9089), .Z(n9087) );
  XOR U12943 ( .A(DB[1907]), .B(DB[1876]), .Z(n9089) );
  AND U12944 ( .A(n272), .B(n9090), .Z(n9088) );
  XOR U12945 ( .A(n9091), .B(n9092), .Z(n9090) );
  XOR U12946 ( .A(DB[1876]), .B(DB[1845]), .Z(n9092) );
  AND U12947 ( .A(n276), .B(n9093), .Z(n9091) );
  XOR U12948 ( .A(n9094), .B(n9095), .Z(n9093) );
  XOR U12949 ( .A(DB[1845]), .B(DB[1814]), .Z(n9095) );
  AND U12950 ( .A(n280), .B(n9096), .Z(n9094) );
  XOR U12951 ( .A(n9097), .B(n9098), .Z(n9096) );
  XOR U12952 ( .A(DB[1814]), .B(DB[1783]), .Z(n9098) );
  AND U12953 ( .A(n284), .B(n9099), .Z(n9097) );
  XOR U12954 ( .A(n9100), .B(n9101), .Z(n9099) );
  XOR U12955 ( .A(DB[1783]), .B(DB[1752]), .Z(n9101) );
  AND U12956 ( .A(n288), .B(n9102), .Z(n9100) );
  XOR U12957 ( .A(n9103), .B(n9104), .Z(n9102) );
  XOR U12958 ( .A(DB[1752]), .B(DB[1721]), .Z(n9104) );
  AND U12959 ( .A(n292), .B(n9105), .Z(n9103) );
  XOR U12960 ( .A(n9106), .B(n9107), .Z(n9105) );
  XOR U12961 ( .A(DB[1721]), .B(DB[1690]), .Z(n9107) );
  AND U12962 ( .A(n296), .B(n9108), .Z(n9106) );
  XOR U12963 ( .A(n9109), .B(n9110), .Z(n9108) );
  XOR U12964 ( .A(DB[1690]), .B(DB[1659]), .Z(n9110) );
  AND U12965 ( .A(n300), .B(n9111), .Z(n9109) );
  XOR U12966 ( .A(n9112), .B(n9113), .Z(n9111) );
  XOR U12967 ( .A(DB[1659]), .B(DB[1628]), .Z(n9113) );
  AND U12968 ( .A(n304), .B(n9114), .Z(n9112) );
  XOR U12969 ( .A(n9115), .B(n9116), .Z(n9114) );
  XOR U12970 ( .A(DB[1628]), .B(DB[1597]), .Z(n9116) );
  AND U12971 ( .A(n308), .B(n9117), .Z(n9115) );
  XOR U12972 ( .A(n9118), .B(n9119), .Z(n9117) );
  XOR U12973 ( .A(DB[1597]), .B(DB[1566]), .Z(n9119) );
  AND U12974 ( .A(n312), .B(n9120), .Z(n9118) );
  XOR U12975 ( .A(n9121), .B(n9122), .Z(n9120) );
  XOR U12976 ( .A(DB[1566]), .B(DB[1535]), .Z(n9122) );
  AND U12977 ( .A(n316), .B(n9123), .Z(n9121) );
  XOR U12978 ( .A(n9124), .B(n9125), .Z(n9123) );
  XOR U12979 ( .A(DB[1535]), .B(DB[1504]), .Z(n9125) );
  AND U12980 ( .A(n320), .B(n9126), .Z(n9124) );
  XOR U12981 ( .A(n9127), .B(n9128), .Z(n9126) );
  XOR U12982 ( .A(DB[1504]), .B(DB[1473]), .Z(n9128) );
  AND U12983 ( .A(n324), .B(n9129), .Z(n9127) );
  XOR U12984 ( .A(n9130), .B(n9131), .Z(n9129) );
  XOR U12985 ( .A(DB[1473]), .B(DB[1442]), .Z(n9131) );
  AND U12986 ( .A(n328), .B(n9132), .Z(n9130) );
  XOR U12987 ( .A(n9133), .B(n9134), .Z(n9132) );
  XOR U12988 ( .A(DB[1442]), .B(DB[1411]), .Z(n9134) );
  AND U12989 ( .A(n332), .B(n9135), .Z(n9133) );
  XOR U12990 ( .A(n9136), .B(n9137), .Z(n9135) );
  XOR U12991 ( .A(DB[1411]), .B(DB[1380]), .Z(n9137) );
  AND U12992 ( .A(n336), .B(n9138), .Z(n9136) );
  XOR U12993 ( .A(n9139), .B(n9140), .Z(n9138) );
  XOR U12994 ( .A(DB[1380]), .B(DB[1349]), .Z(n9140) );
  AND U12995 ( .A(n340), .B(n9141), .Z(n9139) );
  XOR U12996 ( .A(n9142), .B(n9143), .Z(n9141) );
  XOR U12997 ( .A(DB[1349]), .B(DB[1318]), .Z(n9143) );
  AND U12998 ( .A(n344), .B(n9144), .Z(n9142) );
  XOR U12999 ( .A(n9145), .B(n9146), .Z(n9144) );
  XOR U13000 ( .A(DB[1318]), .B(DB[1287]), .Z(n9146) );
  AND U13001 ( .A(n348), .B(n9147), .Z(n9145) );
  XOR U13002 ( .A(n9148), .B(n9149), .Z(n9147) );
  XOR U13003 ( .A(DB[1287]), .B(DB[1256]), .Z(n9149) );
  AND U13004 ( .A(n352), .B(n9150), .Z(n9148) );
  XOR U13005 ( .A(n9151), .B(n9152), .Z(n9150) );
  XOR U13006 ( .A(DB[1256]), .B(DB[1225]), .Z(n9152) );
  AND U13007 ( .A(n356), .B(n9153), .Z(n9151) );
  XOR U13008 ( .A(n9154), .B(n9155), .Z(n9153) );
  XOR U13009 ( .A(DB[1225]), .B(DB[1194]), .Z(n9155) );
  AND U13010 ( .A(n360), .B(n9156), .Z(n9154) );
  XOR U13011 ( .A(n9157), .B(n9158), .Z(n9156) );
  XOR U13012 ( .A(DB[1194]), .B(DB[1163]), .Z(n9158) );
  AND U13013 ( .A(n364), .B(n9159), .Z(n9157) );
  XOR U13014 ( .A(n9160), .B(n9161), .Z(n9159) );
  XOR U13015 ( .A(DB[1163]), .B(DB[1132]), .Z(n9161) );
  AND U13016 ( .A(n368), .B(n9162), .Z(n9160) );
  XOR U13017 ( .A(n9163), .B(n9164), .Z(n9162) );
  XOR U13018 ( .A(DB[1132]), .B(DB[1101]), .Z(n9164) );
  AND U13019 ( .A(n372), .B(n9165), .Z(n9163) );
  XOR U13020 ( .A(n9166), .B(n9167), .Z(n9165) );
  XOR U13021 ( .A(DB[1101]), .B(DB[1070]), .Z(n9167) );
  AND U13022 ( .A(n376), .B(n9168), .Z(n9166) );
  XOR U13023 ( .A(n9169), .B(n9170), .Z(n9168) );
  XOR U13024 ( .A(DB[1070]), .B(DB[1039]), .Z(n9170) );
  AND U13025 ( .A(n380), .B(n9171), .Z(n9169) );
  XOR U13026 ( .A(n9172), .B(n9173), .Z(n9171) );
  XOR U13027 ( .A(DB[1039]), .B(DB[1008]), .Z(n9173) );
  AND U13028 ( .A(n384), .B(n9174), .Z(n9172) );
  XOR U13029 ( .A(n9175), .B(n9176), .Z(n9174) );
  XOR U13030 ( .A(DB[977]), .B(DB[1008]), .Z(n9176) );
  AND U13031 ( .A(n388), .B(n9177), .Z(n9175) );
  XOR U13032 ( .A(n9178), .B(n9179), .Z(n9177) );
  XOR U13033 ( .A(DB[977]), .B(DB[946]), .Z(n9179) );
  AND U13034 ( .A(n392), .B(n9180), .Z(n9178) );
  XOR U13035 ( .A(n9181), .B(n9182), .Z(n9180) );
  XOR U13036 ( .A(DB[946]), .B(DB[915]), .Z(n9182) );
  AND U13037 ( .A(n396), .B(n9183), .Z(n9181) );
  XOR U13038 ( .A(n9184), .B(n9185), .Z(n9183) );
  XOR U13039 ( .A(DB[915]), .B(DB[884]), .Z(n9185) );
  AND U13040 ( .A(n400), .B(n9186), .Z(n9184) );
  XOR U13041 ( .A(n9187), .B(n9188), .Z(n9186) );
  XOR U13042 ( .A(DB[884]), .B(DB[853]), .Z(n9188) );
  AND U13043 ( .A(n404), .B(n9189), .Z(n9187) );
  XOR U13044 ( .A(n9190), .B(n9191), .Z(n9189) );
  XOR U13045 ( .A(DB[853]), .B(DB[822]), .Z(n9191) );
  AND U13046 ( .A(n408), .B(n9192), .Z(n9190) );
  XOR U13047 ( .A(n9193), .B(n9194), .Z(n9192) );
  XOR U13048 ( .A(DB[822]), .B(DB[791]), .Z(n9194) );
  AND U13049 ( .A(n412), .B(n9195), .Z(n9193) );
  XOR U13050 ( .A(n9196), .B(n9197), .Z(n9195) );
  XOR U13051 ( .A(DB[791]), .B(DB[760]), .Z(n9197) );
  AND U13052 ( .A(n416), .B(n9198), .Z(n9196) );
  XOR U13053 ( .A(n9199), .B(n9200), .Z(n9198) );
  XOR U13054 ( .A(DB[760]), .B(DB[729]), .Z(n9200) );
  AND U13055 ( .A(n420), .B(n9201), .Z(n9199) );
  XOR U13056 ( .A(n9202), .B(n9203), .Z(n9201) );
  XOR U13057 ( .A(DB[729]), .B(DB[698]), .Z(n9203) );
  AND U13058 ( .A(n424), .B(n9204), .Z(n9202) );
  XOR U13059 ( .A(n9205), .B(n9206), .Z(n9204) );
  XOR U13060 ( .A(DB[698]), .B(DB[667]), .Z(n9206) );
  AND U13061 ( .A(n428), .B(n9207), .Z(n9205) );
  XOR U13062 ( .A(n9208), .B(n9209), .Z(n9207) );
  XOR U13063 ( .A(DB[667]), .B(DB[636]), .Z(n9209) );
  AND U13064 ( .A(n432), .B(n9210), .Z(n9208) );
  XOR U13065 ( .A(n9211), .B(n9212), .Z(n9210) );
  XOR U13066 ( .A(DB[636]), .B(DB[605]), .Z(n9212) );
  AND U13067 ( .A(n436), .B(n9213), .Z(n9211) );
  XOR U13068 ( .A(n9214), .B(n9215), .Z(n9213) );
  XOR U13069 ( .A(DB[605]), .B(DB[574]), .Z(n9215) );
  AND U13070 ( .A(n440), .B(n9216), .Z(n9214) );
  XOR U13071 ( .A(n9217), .B(n9218), .Z(n9216) );
  XOR U13072 ( .A(DB[574]), .B(DB[543]), .Z(n9218) );
  AND U13073 ( .A(n444), .B(n9219), .Z(n9217) );
  XOR U13074 ( .A(n9220), .B(n9221), .Z(n9219) );
  XOR U13075 ( .A(DB[543]), .B(DB[512]), .Z(n9221) );
  AND U13076 ( .A(n448), .B(n9222), .Z(n9220) );
  XOR U13077 ( .A(n9223), .B(n9224), .Z(n9222) );
  XOR U13078 ( .A(DB[512]), .B(DB[481]), .Z(n9224) );
  AND U13079 ( .A(n452), .B(n9225), .Z(n9223) );
  XOR U13080 ( .A(n9226), .B(n9227), .Z(n9225) );
  XOR U13081 ( .A(DB[481]), .B(DB[450]), .Z(n9227) );
  AND U13082 ( .A(n456), .B(n9228), .Z(n9226) );
  XOR U13083 ( .A(n9229), .B(n9230), .Z(n9228) );
  XOR U13084 ( .A(DB[450]), .B(DB[419]), .Z(n9230) );
  AND U13085 ( .A(n460), .B(n9231), .Z(n9229) );
  XOR U13086 ( .A(n9232), .B(n9233), .Z(n9231) );
  XOR U13087 ( .A(DB[419]), .B(DB[388]), .Z(n9233) );
  AND U13088 ( .A(n464), .B(n9234), .Z(n9232) );
  XOR U13089 ( .A(n9235), .B(n9236), .Z(n9234) );
  XOR U13090 ( .A(DB[388]), .B(DB[357]), .Z(n9236) );
  AND U13091 ( .A(n468), .B(n9237), .Z(n9235) );
  XOR U13092 ( .A(n9238), .B(n9239), .Z(n9237) );
  XOR U13093 ( .A(DB[357]), .B(DB[326]), .Z(n9239) );
  AND U13094 ( .A(n472), .B(n9240), .Z(n9238) );
  XOR U13095 ( .A(n9241), .B(n9242), .Z(n9240) );
  XOR U13096 ( .A(DB[326]), .B(DB[295]), .Z(n9242) );
  AND U13097 ( .A(n476), .B(n9243), .Z(n9241) );
  XOR U13098 ( .A(n9244), .B(n9245), .Z(n9243) );
  XOR U13099 ( .A(DB[295]), .B(DB[264]), .Z(n9245) );
  AND U13100 ( .A(n480), .B(n9246), .Z(n9244) );
  XOR U13101 ( .A(n9247), .B(n9248), .Z(n9246) );
  XOR U13102 ( .A(DB[264]), .B(DB[233]), .Z(n9248) );
  AND U13103 ( .A(n484), .B(n9249), .Z(n9247) );
  XOR U13104 ( .A(n9250), .B(n9251), .Z(n9249) );
  XOR U13105 ( .A(DB[233]), .B(DB[202]), .Z(n9251) );
  AND U13106 ( .A(n488), .B(n9252), .Z(n9250) );
  XOR U13107 ( .A(n9253), .B(n9254), .Z(n9252) );
  XOR U13108 ( .A(DB[202]), .B(DB[171]), .Z(n9254) );
  AND U13109 ( .A(n492), .B(n9255), .Z(n9253) );
  XOR U13110 ( .A(n9256), .B(n9257), .Z(n9255) );
  XOR U13111 ( .A(DB[171]), .B(DB[140]), .Z(n9257) );
  AND U13112 ( .A(n496), .B(n9258), .Z(n9256) );
  XOR U13113 ( .A(n9259), .B(n9260), .Z(n9258) );
  XOR U13114 ( .A(DB[140]), .B(DB[109]), .Z(n9260) );
  AND U13115 ( .A(n500), .B(n9261), .Z(n9259) );
  XOR U13116 ( .A(n9262), .B(n9263), .Z(n9261) );
  XOR U13117 ( .A(DB[78]), .B(DB[109]), .Z(n9263) );
  AND U13118 ( .A(n504), .B(n9264), .Z(n9262) );
  XOR U13119 ( .A(n9265), .B(n9266), .Z(n9264) );
  XOR U13120 ( .A(DB[78]), .B(DB[47]), .Z(n9266) );
  AND U13121 ( .A(n508), .B(n9267), .Z(n9265) );
  XOR U13122 ( .A(DB[47]), .B(DB[16]), .Z(n9267) );
  XOR U13123 ( .A(DB[3952]), .B(n9268), .Z(min_val_out[15]) );
  AND U13124 ( .A(n2), .B(n9269), .Z(n9268) );
  XOR U13125 ( .A(n9270), .B(n9271), .Z(n9269) );
  XOR U13126 ( .A(DB[3952]), .B(DB[3921]), .Z(n9271) );
  AND U13127 ( .A(n8), .B(n9272), .Z(n9270) );
  XOR U13128 ( .A(n9273), .B(n9274), .Z(n9272) );
  XOR U13129 ( .A(DB[3921]), .B(DB[3890]), .Z(n9274) );
  AND U13130 ( .A(n12), .B(n9275), .Z(n9273) );
  XOR U13131 ( .A(n9276), .B(n9277), .Z(n9275) );
  XOR U13132 ( .A(DB[3890]), .B(DB[3859]), .Z(n9277) );
  AND U13133 ( .A(n16), .B(n9278), .Z(n9276) );
  XOR U13134 ( .A(n9279), .B(n9280), .Z(n9278) );
  XOR U13135 ( .A(DB[3859]), .B(DB[3828]), .Z(n9280) );
  AND U13136 ( .A(n20), .B(n9281), .Z(n9279) );
  XOR U13137 ( .A(n9282), .B(n9283), .Z(n9281) );
  XOR U13138 ( .A(DB[3828]), .B(DB[3797]), .Z(n9283) );
  AND U13139 ( .A(n24), .B(n9284), .Z(n9282) );
  XOR U13140 ( .A(n9285), .B(n9286), .Z(n9284) );
  XOR U13141 ( .A(DB[3797]), .B(DB[3766]), .Z(n9286) );
  AND U13142 ( .A(n28), .B(n9287), .Z(n9285) );
  XOR U13143 ( .A(n9288), .B(n9289), .Z(n9287) );
  XOR U13144 ( .A(DB[3766]), .B(DB[3735]), .Z(n9289) );
  AND U13145 ( .A(n32), .B(n9290), .Z(n9288) );
  XOR U13146 ( .A(n9291), .B(n9292), .Z(n9290) );
  XOR U13147 ( .A(DB[3735]), .B(DB[3704]), .Z(n9292) );
  AND U13148 ( .A(n36), .B(n9293), .Z(n9291) );
  XOR U13149 ( .A(n9294), .B(n9295), .Z(n9293) );
  XOR U13150 ( .A(DB[3704]), .B(DB[3673]), .Z(n9295) );
  AND U13151 ( .A(n40), .B(n9296), .Z(n9294) );
  XOR U13152 ( .A(n9297), .B(n9298), .Z(n9296) );
  XOR U13153 ( .A(DB[3673]), .B(DB[3642]), .Z(n9298) );
  AND U13154 ( .A(n44), .B(n9299), .Z(n9297) );
  XOR U13155 ( .A(n9300), .B(n9301), .Z(n9299) );
  XOR U13156 ( .A(DB[3642]), .B(DB[3611]), .Z(n9301) );
  AND U13157 ( .A(n48), .B(n9302), .Z(n9300) );
  XOR U13158 ( .A(n9303), .B(n9304), .Z(n9302) );
  XOR U13159 ( .A(DB[3611]), .B(DB[3580]), .Z(n9304) );
  AND U13160 ( .A(n52), .B(n9305), .Z(n9303) );
  XOR U13161 ( .A(n9306), .B(n9307), .Z(n9305) );
  XOR U13162 ( .A(DB[3580]), .B(DB[3549]), .Z(n9307) );
  AND U13163 ( .A(n56), .B(n9308), .Z(n9306) );
  XOR U13164 ( .A(n9309), .B(n9310), .Z(n9308) );
  XOR U13165 ( .A(DB[3549]), .B(DB[3518]), .Z(n9310) );
  AND U13166 ( .A(n60), .B(n9311), .Z(n9309) );
  XOR U13167 ( .A(n9312), .B(n9313), .Z(n9311) );
  XOR U13168 ( .A(DB[3518]), .B(DB[3487]), .Z(n9313) );
  AND U13169 ( .A(n64), .B(n9314), .Z(n9312) );
  XOR U13170 ( .A(n9315), .B(n9316), .Z(n9314) );
  XOR U13171 ( .A(DB[3487]), .B(DB[3456]), .Z(n9316) );
  AND U13172 ( .A(n68), .B(n9317), .Z(n9315) );
  XOR U13173 ( .A(n9318), .B(n9319), .Z(n9317) );
  XOR U13174 ( .A(DB[3456]), .B(DB[3425]), .Z(n9319) );
  AND U13175 ( .A(n72), .B(n9320), .Z(n9318) );
  XOR U13176 ( .A(n9321), .B(n9322), .Z(n9320) );
  XOR U13177 ( .A(DB[3425]), .B(DB[3394]), .Z(n9322) );
  AND U13178 ( .A(n76), .B(n9323), .Z(n9321) );
  XOR U13179 ( .A(n9324), .B(n9325), .Z(n9323) );
  XOR U13180 ( .A(DB[3394]), .B(DB[3363]), .Z(n9325) );
  AND U13181 ( .A(n80), .B(n9326), .Z(n9324) );
  XOR U13182 ( .A(n9327), .B(n9328), .Z(n9326) );
  XOR U13183 ( .A(DB[3363]), .B(DB[3332]), .Z(n9328) );
  AND U13184 ( .A(n84), .B(n9329), .Z(n9327) );
  XOR U13185 ( .A(n9330), .B(n9331), .Z(n9329) );
  XOR U13186 ( .A(DB[3332]), .B(DB[3301]), .Z(n9331) );
  AND U13187 ( .A(n88), .B(n9332), .Z(n9330) );
  XOR U13188 ( .A(n9333), .B(n9334), .Z(n9332) );
  XOR U13189 ( .A(DB[3301]), .B(DB[3270]), .Z(n9334) );
  AND U13190 ( .A(n92), .B(n9335), .Z(n9333) );
  XOR U13191 ( .A(n9336), .B(n9337), .Z(n9335) );
  XOR U13192 ( .A(DB[3270]), .B(DB[3239]), .Z(n9337) );
  AND U13193 ( .A(n96), .B(n9338), .Z(n9336) );
  XOR U13194 ( .A(n9339), .B(n9340), .Z(n9338) );
  XOR U13195 ( .A(DB[3239]), .B(DB[3208]), .Z(n9340) );
  AND U13196 ( .A(n100), .B(n9341), .Z(n9339) );
  XOR U13197 ( .A(n9342), .B(n9343), .Z(n9341) );
  XOR U13198 ( .A(DB[3208]), .B(DB[3177]), .Z(n9343) );
  AND U13199 ( .A(n104), .B(n9344), .Z(n9342) );
  XOR U13200 ( .A(n9345), .B(n9346), .Z(n9344) );
  XOR U13201 ( .A(DB[3177]), .B(DB[3146]), .Z(n9346) );
  AND U13202 ( .A(n108), .B(n9347), .Z(n9345) );
  XOR U13203 ( .A(n9348), .B(n9349), .Z(n9347) );
  XOR U13204 ( .A(DB[3146]), .B(DB[3115]), .Z(n9349) );
  AND U13205 ( .A(n112), .B(n9350), .Z(n9348) );
  XOR U13206 ( .A(n9351), .B(n9352), .Z(n9350) );
  XOR U13207 ( .A(DB[3115]), .B(DB[3084]), .Z(n9352) );
  AND U13208 ( .A(n116), .B(n9353), .Z(n9351) );
  XOR U13209 ( .A(n9354), .B(n9355), .Z(n9353) );
  XOR U13210 ( .A(DB[3084]), .B(DB[3053]), .Z(n9355) );
  AND U13211 ( .A(n120), .B(n9356), .Z(n9354) );
  XOR U13212 ( .A(n9357), .B(n9358), .Z(n9356) );
  XOR U13213 ( .A(DB[3053]), .B(DB[3022]), .Z(n9358) );
  AND U13214 ( .A(n124), .B(n9359), .Z(n9357) );
  XOR U13215 ( .A(n9360), .B(n9361), .Z(n9359) );
  XOR U13216 ( .A(DB[3022]), .B(DB[2991]), .Z(n9361) );
  AND U13217 ( .A(n128), .B(n9362), .Z(n9360) );
  XOR U13218 ( .A(n9363), .B(n9364), .Z(n9362) );
  XOR U13219 ( .A(DB[2991]), .B(DB[2960]), .Z(n9364) );
  AND U13220 ( .A(n132), .B(n9365), .Z(n9363) );
  XOR U13221 ( .A(n9366), .B(n9367), .Z(n9365) );
  XOR U13222 ( .A(DB[2960]), .B(DB[2929]), .Z(n9367) );
  AND U13223 ( .A(n136), .B(n9368), .Z(n9366) );
  XOR U13224 ( .A(n9369), .B(n9370), .Z(n9368) );
  XOR U13225 ( .A(DB[2929]), .B(DB[2898]), .Z(n9370) );
  AND U13226 ( .A(n140), .B(n9371), .Z(n9369) );
  XOR U13227 ( .A(n9372), .B(n9373), .Z(n9371) );
  XOR U13228 ( .A(DB[2898]), .B(DB[2867]), .Z(n9373) );
  AND U13229 ( .A(n144), .B(n9374), .Z(n9372) );
  XOR U13230 ( .A(n9375), .B(n9376), .Z(n9374) );
  XOR U13231 ( .A(DB[2867]), .B(DB[2836]), .Z(n9376) );
  AND U13232 ( .A(n148), .B(n9377), .Z(n9375) );
  XOR U13233 ( .A(n9378), .B(n9379), .Z(n9377) );
  XOR U13234 ( .A(DB[2836]), .B(DB[2805]), .Z(n9379) );
  AND U13235 ( .A(n152), .B(n9380), .Z(n9378) );
  XOR U13236 ( .A(n9381), .B(n9382), .Z(n9380) );
  XOR U13237 ( .A(DB[2805]), .B(DB[2774]), .Z(n9382) );
  AND U13238 ( .A(n156), .B(n9383), .Z(n9381) );
  XOR U13239 ( .A(n9384), .B(n9385), .Z(n9383) );
  XOR U13240 ( .A(DB[2774]), .B(DB[2743]), .Z(n9385) );
  AND U13241 ( .A(n160), .B(n9386), .Z(n9384) );
  XOR U13242 ( .A(n9387), .B(n9388), .Z(n9386) );
  XOR U13243 ( .A(DB[2743]), .B(DB[2712]), .Z(n9388) );
  AND U13244 ( .A(n164), .B(n9389), .Z(n9387) );
  XOR U13245 ( .A(n9390), .B(n9391), .Z(n9389) );
  XOR U13246 ( .A(DB[2712]), .B(DB[2681]), .Z(n9391) );
  AND U13247 ( .A(n168), .B(n9392), .Z(n9390) );
  XOR U13248 ( .A(n9393), .B(n9394), .Z(n9392) );
  XOR U13249 ( .A(DB[2681]), .B(DB[2650]), .Z(n9394) );
  AND U13250 ( .A(n172), .B(n9395), .Z(n9393) );
  XOR U13251 ( .A(n9396), .B(n9397), .Z(n9395) );
  XOR U13252 ( .A(DB[2650]), .B(DB[2619]), .Z(n9397) );
  AND U13253 ( .A(n176), .B(n9398), .Z(n9396) );
  XOR U13254 ( .A(n9399), .B(n9400), .Z(n9398) );
  XOR U13255 ( .A(DB[2619]), .B(DB[2588]), .Z(n9400) );
  AND U13256 ( .A(n180), .B(n9401), .Z(n9399) );
  XOR U13257 ( .A(n9402), .B(n9403), .Z(n9401) );
  XOR U13258 ( .A(DB[2588]), .B(DB[2557]), .Z(n9403) );
  AND U13259 ( .A(n184), .B(n9404), .Z(n9402) );
  XOR U13260 ( .A(n9405), .B(n9406), .Z(n9404) );
  XOR U13261 ( .A(DB[2557]), .B(DB[2526]), .Z(n9406) );
  AND U13262 ( .A(n188), .B(n9407), .Z(n9405) );
  XOR U13263 ( .A(n9408), .B(n9409), .Z(n9407) );
  XOR U13264 ( .A(DB[2526]), .B(DB[2495]), .Z(n9409) );
  AND U13265 ( .A(n192), .B(n9410), .Z(n9408) );
  XOR U13266 ( .A(n9411), .B(n9412), .Z(n9410) );
  XOR U13267 ( .A(DB[2495]), .B(DB[2464]), .Z(n9412) );
  AND U13268 ( .A(n196), .B(n9413), .Z(n9411) );
  XOR U13269 ( .A(n9414), .B(n9415), .Z(n9413) );
  XOR U13270 ( .A(DB[2464]), .B(DB[2433]), .Z(n9415) );
  AND U13271 ( .A(n200), .B(n9416), .Z(n9414) );
  XOR U13272 ( .A(n9417), .B(n9418), .Z(n9416) );
  XOR U13273 ( .A(DB[2433]), .B(DB[2402]), .Z(n9418) );
  AND U13274 ( .A(n204), .B(n9419), .Z(n9417) );
  XOR U13275 ( .A(n9420), .B(n9421), .Z(n9419) );
  XOR U13276 ( .A(DB[2402]), .B(DB[2371]), .Z(n9421) );
  AND U13277 ( .A(n208), .B(n9422), .Z(n9420) );
  XOR U13278 ( .A(n9423), .B(n9424), .Z(n9422) );
  XOR U13279 ( .A(DB[2371]), .B(DB[2340]), .Z(n9424) );
  AND U13280 ( .A(n212), .B(n9425), .Z(n9423) );
  XOR U13281 ( .A(n9426), .B(n9427), .Z(n9425) );
  XOR U13282 ( .A(DB[2340]), .B(DB[2309]), .Z(n9427) );
  AND U13283 ( .A(n216), .B(n9428), .Z(n9426) );
  XOR U13284 ( .A(n9429), .B(n9430), .Z(n9428) );
  XOR U13285 ( .A(DB[2309]), .B(DB[2278]), .Z(n9430) );
  AND U13286 ( .A(n220), .B(n9431), .Z(n9429) );
  XOR U13287 ( .A(n9432), .B(n9433), .Z(n9431) );
  XOR U13288 ( .A(DB[2278]), .B(DB[2247]), .Z(n9433) );
  AND U13289 ( .A(n224), .B(n9434), .Z(n9432) );
  XOR U13290 ( .A(n9435), .B(n9436), .Z(n9434) );
  XOR U13291 ( .A(DB[2247]), .B(DB[2216]), .Z(n9436) );
  AND U13292 ( .A(n228), .B(n9437), .Z(n9435) );
  XOR U13293 ( .A(n9438), .B(n9439), .Z(n9437) );
  XOR U13294 ( .A(DB[2216]), .B(DB[2185]), .Z(n9439) );
  AND U13295 ( .A(n232), .B(n9440), .Z(n9438) );
  XOR U13296 ( .A(n9441), .B(n9442), .Z(n9440) );
  XOR U13297 ( .A(DB[2185]), .B(DB[2154]), .Z(n9442) );
  AND U13298 ( .A(n236), .B(n9443), .Z(n9441) );
  XOR U13299 ( .A(n9444), .B(n9445), .Z(n9443) );
  XOR U13300 ( .A(DB[2154]), .B(DB[2123]), .Z(n9445) );
  AND U13301 ( .A(n240), .B(n9446), .Z(n9444) );
  XOR U13302 ( .A(n9447), .B(n9448), .Z(n9446) );
  XOR U13303 ( .A(DB[2123]), .B(DB[2092]), .Z(n9448) );
  AND U13304 ( .A(n244), .B(n9449), .Z(n9447) );
  XOR U13305 ( .A(n9450), .B(n9451), .Z(n9449) );
  XOR U13306 ( .A(DB[2092]), .B(DB[2061]), .Z(n9451) );
  AND U13307 ( .A(n248), .B(n9452), .Z(n9450) );
  XOR U13308 ( .A(n9453), .B(n9454), .Z(n9452) );
  XOR U13309 ( .A(DB[2061]), .B(DB[2030]), .Z(n9454) );
  AND U13310 ( .A(n252), .B(n9455), .Z(n9453) );
  XOR U13311 ( .A(n9456), .B(n9457), .Z(n9455) );
  XOR U13312 ( .A(DB[2030]), .B(DB[1999]), .Z(n9457) );
  AND U13313 ( .A(n256), .B(n9458), .Z(n9456) );
  XOR U13314 ( .A(n9459), .B(n9460), .Z(n9458) );
  XOR U13315 ( .A(DB[1999]), .B(DB[1968]), .Z(n9460) );
  AND U13316 ( .A(n260), .B(n9461), .Z(n9459) );
  XOR U13317 ( .A(n9462), .B(n9463), .Z(n9461) );
  XOR U13318 ( .A(DB[1968]), .B(DB[1937]), .Z(n9463) );
  AND U13319 ( .A(n264), .B(n9464), .Z(n9462) );
  XOR U13320 ( .A(n9465), .B(n9466), .Z(n9464) );
  XOR U13321 ( .A(DB[1937]), .B(DB[1906]), .Z(n9466) );
  AND U13322 ( .A(n268), .B(n9467), .Z(n9465) );
  XOR U13323 ( .A(n9468), .B(n9469), .Z(n9467) );
  XOR U13324 ( .A(DB[1906]), .B(DB[1875]), .Z(n9469) );
  AND U13325 ( .A(n272), .B(n9470), .Z(n9468) );
  XOR U13326 ( .A(n9471), .B(n9472), .Z(n9470) );
  XOR U13327 ( .A(DB[1875]), .B(DB[1844]), .Z(n9472) );
  AND U13328 ( .A(n276), .B(n9473), .Z(n9471) );
  XOR U13329 ( .A(n9474), .B(n9475), .Z(n9473) );
  XOR U13330 ( .A(DB[1844]), .B(DB[1813]), .Z(n9475) );
  AND U13331 ( .A(n280), .B(n9476), .Z(n9474) );
  XOR U13332 ( .A(n9477), .B(n9478), .Z(n9476) );
  XOR U13333 ( .A(DB[1813]), .B(DB[1782]), .Z(n9478) );
  AND U13334 ( .A(n284), .B(n9479), .Z(n9477) );
  XOR U13335 ( .A(n9480), .B(n9481), .Z(n9479) );
  XOR U13336 ( .A(DB[1782]), .B(DB[1751]), .Z(n9481) );
  AND U13337 ( .A(n288), .B(n9482), .Z(n9480) );
  XOR U13338 ( .A(n9483), .B(n9484), .Z(n9482) );
  XOR U13339 ( .A(DB[1751]), .B(DB[1720]), .Z(n9484) );
  AND U13340 ( .A(n292), .B(n9485), .Z(n9483) );
  XOR U13341 ( .A(n9486), .B(n9487), .Z(n9485) );
  XOR U13342 ( .A(DB[1720]), .B(DB[1689]), .Z(n9487) );
  AND U13343 ( .A(n296), .B(n9488), .Z(n9486) );
  XOR U13344 ( .A(n9489), .B(n9490), .Z(n9488) );
  XOR U13345 ( .A(DB[1689]), .B(DB[1658]), .Z(n9490) );
  AND U13346 ( .A(n300), .B(n9491), .Z(n9489) );
  XOR U13347 ( .A(n9492), .B(n9493), .Z(n9491) );
  XOR U13348 ( .A(DB[1658]), .B(DB[1627]), .Z(n9493) );
  AND U13349 ( .A(n304), .B(n9494), .Z(n9492) );
  XOR U13350 ( .A(n9495), .B(n9496), .Z(n9494) );
  XOR U13351 ( .A(DB[1627]), .B(DB[1596]), .Z(n9496) );
  AND U13352 ( .A(n308), .B(n9497), .Z(n9495) );
  XOR U13353 ( .A(n9498), .B(n9499), .Z(n9497) );
  XOR U13354 ( .A(DB[1596]), .B(DB[1565]), .Z(n9499) );
  AND U13355 ( .A(n312), .B(n9500), .Z(n9498) );
  XOR U13356 ( .A(n9501), .B(n9502), .Z(n9500) );
  XOR U13357 ( .A(DB[1565]), .B(DB[1534]), .Z(n9502) );
  AND U13358 ( .A(n316), .B(n9503), .Z(n9501) );
  XOR U13359 ( .A(n9504), .B(n9505), .Z(n9503) );
  XOR U13360 ( .A(DB[1534]), .B(DB[1503]), .Z(n9505) );
  AND U13361 ( .A(n320), .B(n9506), .Z(n9504) );
  XOR U13362 ( .A(n9507), .B(n9508), .Z(n9506) );
  XOR U13363 ( .A(DB[1503]), .B(DB[1472]), .Z(n9508) );
  AND U13364 ( .A(n324), .B(n9509), .Z(n9507) );
  XOR U13365 ( .A(n9510), .B(n9511), .Z(n9509) );
  XOR U13366 ( .A(DB[1472]), .B(DB[1441]), .Z(n9511) );
  AND U13367 ( .A(n328), .B(n9512), .Z(n9510) );
  XOR U13368 ( .A(n9513), .B(n9514), .Z(n9512) );
  XOR U13369 ( .A(DB[1441]), .B(DB[1410]), .Z(n9514) );
  AND U13370 ( .A(n332), .B(n9515), .Z(n9513) );
  XOR U13371 ( .A(n9516), .B(n9517), .Z(n9515) );
  XOR U13372 ( .A(DB[1410]), .B(DB[1379]), .Z(n9517) );
  AND U13373 ( .A(n336), .B(n9518), .Z(n9516) );
  XOR U13374 ( .A(n9519), .B(n9520), .Z(n9518) );
  XOR U13375 ( .A(DB[1379]), .B(DB[1348]), .Z(n9520) );
  AND U13376 ( .A(n340), .B(n9521), .Z(n9519) );
  XOR U13377 ( .A(n9522), .B(n9523), .Z(n9521) );
  XOR U13378 ( .A(DB[1348]), .B(DB[1317]), .Z(n9523) );
  AND U13379 ( .A(n344), .B(n9524), .Z(n9522) );
  XOR U13380 ( .A(n9525), .B(n9526), .Z(n9524) );
  XOR U13381 ( .A(DB[1317]), .B(DB[1286]), .Z(n9526) );
  AND U13382 ( .A(n348), .B(n9527), .Z(n9525) );
  XOR U13383 ( .A(n9528), .B(n9529), .Z(n9527) );
  XOR U13384 ( .A(DB[1286]), .B(DB[1255]), .Z(n9529) );
  AND U13385 ( .A(n352), .B(n9530), .Z(n9528) );
  XOR U13386 ( .A(n9531), .B(n9532), .Z(n9530) );
  XOR U13387 ( .A(DB[1255]), .B(DB[1224]), .Z(n9532) );
  AND U13388 ( .A(n356), .B(n9533), .Z(n9531) );
  XOR U13389 ( .A(n9534), .B(n9535), .Z(n9533) );
  XOR U13390 ( .A(DB[1224]), .B(DB[1193]), .Z(n9535) );
  AND U13391 ( .A(n360), .B(n9536), .Z(n9534) );
  XOR U13392 ( .A(n9537), .B(n9538), .Z(n9536) );
  XOR U13393 ( .A(DB[1193]), .B(DB[1162]), .Z(n9538) );
  AND U13394 ( .A(n364), .B(n9539), .Z(n9537) );
  XOR U13395 ( .A(n9540), .B(n9541), .Z(n9539) );
  XOR U13396 ( .A(DB[1162]), .B(DB[1131]), .Z(n9541) );
  AND U13397 ( .A(n368), .B(n9542), .Z(n9540) );
  XOR U13398 ( .A(n9543), .B(n9544), .Z(n9542) );
  XOR U13399 ( .A(DB[1131]), .B(DB[1100]), .Z(n9544) );
  AND U13400 ( .A(n372), .B(n9545), .Z(n9543) );
  XOR U13401 ( .A(n9546), .B(n9547), .Z(n9545) );
  XOR U13402 ( .A(DB[1100]), .B(DB[1069]), .Z(n9547) );
  AND U13403 ( .A(n376), .B(n9548), .Z(n9546) );
  XOR U13404 ( .A(n9549), .B(n9550), .Z(n9548) );
  XOR U13405 ( .A(DB[1069]), .B(DB[1038]), .Z(n9550) );
  AND U13406 ( .A(n380), .B(n9551), .Z(n9549) );
  XOR U13407 ( .A(n9552), .B(n9553), .Z(n9551) );
  XOR U13408 ( .A(DB[1038]), .B(DB[1007]), .Z(n9553) );
  AND U13409 ( .A(n384), .B(n9554), .Z(n9552) );
  XOR U13410 ( .A(n9555), .B(n9556), .Z(n9554) );
  XOR U13411 ( .A(DB[976]), .B(DB[1007]), .Z(n9556) );
  AND U13412 ( .A(n388), .B(n9557), .Z(n9555) );
  XOR U13413 ( .A(n9558), .B(n9559), .Z(n9557) );
  XOR U13414 ( .A(DB[976]), .B(DB[945]), .Z(n9559) );
  AND U13415 ( .A(n392), .B(n9560), .Z(n9558) );
  XOR U13416 ( .A(n9561), .B(n9562), .Z(n9560) );
  XOR U13417 ( .A(DB[945]), .B(DB[914]), .Z(n9562) );
  AND U13418 ( .A(n396), .B(n9563), .Z(n9561) );
  XOR U13419 ( .A(n9564), .B(n9565), .Z(n9563) );
  XOR U13420 ( .A(DB[914]), .B(DB[883]), .Z(n9565) );
  AND U13421 ( .A(n400), .B(n9566), .Z(n9564) );
  XOR U13422 ( .A(n9567), .B(n9568), .Z(n9566) );
  XOR U13423 ( .A(DB[883]), .B(DB[852]), .Z(n9568) );
  AND U13424 ( .A(n404), .B(n9569), .Z(n9567) );
  XOR U13425 ( .A(n9570), .B(n9571), .Z(n9569) );
  XOR U13426 ( .A(DB[852]), .B(DB[821]), .Z(n9571) );
  AND U13427 ( .A(n408), .B(n9572), .Z(n9570) );
  XOR U13428 ( .A(n9573), .B(n9574), .Z(n9572) );
  XOR U13429 ( .A(DB[821]), .B(DB[790]), .Z(n9574) );
  AND U13430 ( .A(n412), .B(n9575), .Z(n9573) );
  XOR U13431 ( .A(n9576), .B(n9577), .Z(n9575) );
  XOR U13432 ( .A(DB[790]), .B(DB[759]), .Z(n9577) );
  AND U13433 ( .A(n416), .B(n9578), .Z(n9576) );
  XOR U13434 ( .A(n9579), .B(n9580), .Z(n9578) );
  XOR U13435 ( .A(DB[759]), .B(DB[728]), .Z(n9580) );
  AND U13436 ( .A(n420), .B(n9581), .Z(n9579) );
  XOR U13437 ( .A(n9582), .B(n9583), .Z(n9581) );
  XOR U13438 ( .A(DB[728]), .B(DB[697]), .Z(n9583) );
  AND U13439 ( .A(n424), .B(n9584), .Z(n9582) );
  XOR U13440 ( .A(n9585), .B(n9586), .Z(n9584) );
  XOR U13441 ( .A(DB[697]), .B(DB[666]), .Z(n9586) );
  AND U13442 ( .A(n428), .B(n9587), .Z(n9585) );
  XOR U13443 ( .A(n9588), .B(n9589), .Z(n9587) );
  XOR U13444 ( .A(DB[666]), .B(DB[635]), .Z(n9589) );
  AND U13445 ( .A(n432), .B(n9590), .Z(n9588) );
  XOR U13446 ( .A(n9591), .B(n9592), .Z(n9590) );
  XOR U13447 ( .A(DB[635]), .B(DB[604]), .Z(n9592) );
  AND U13448 ( .A(n436), .B(n9593), .Z(n9591) );
  XOR U13449 ( .A(n9594), .B(n9595), .Z(n9593) );
  XOR U13450 ( .A(DB[604]), .B(DB[573]), .Z(n9595) );
  AND U13451 ( .A(n440), .B(n9596), .Z(n9594) );
  XOR U13452 ( .A(n9597), .B(n9598), .Z(n9596) );
  XOR U13453 ( .A(DB[573]), .B(DB[542]), .Z(n9598) );
  AND U13454 ( .A(n444), .B(n9599), .Z(n9597) );
  XOR U13455 ( .A(n9600), .B(n9601), .Z(n9599) );
  XOR U13456 ( .A(DB[542]), .B(DB[511]), .Z(n9601) );
  AND U13457 ( .A(n448), .B(n9602), .Z(n9600) );
  XOR U13458 ( .A(n9603), .B(n9604), .Z(n9602) );
  XOR U13459 ( .A(DB[511]), .B(DB[480]), .Z(n9604) );
  AND U13460 ( .A(n452), .B(n9605), .Z(n9603) );
  XOR U13461 ( .A(n9606), .B(n9607), .Z(n9605) );
  XOR U13462 ( .A(DB[480]), .B(DB[449]), .Z(n9607) );
  AND U13463 ( .A(n456), .B(n9608), .Z(n9606) );
  XOR U13464 ( .A(n9609), .B(n9610), .Z(n9608) );
  XOR U13465 ( .A(DB[449]), .B(DB[418]), .Z(n9610) );
  AND U13466 ( .A(n460), .B(n9611), .Z(n9609) );
  XOR U13467 ( .A(n9612), .B(n9613), .Z(n9611) );
  XOR U13468 ( .A(DB[418]), .B(DB[387]), .Z(n9613) );
  AND U13469 ( .A(n464), .B(n9614), .Z(n9612) );
  XOR U13470 ( .A(n9615), .B(n9616), .Z(n9614) );
  XOR U13471 ( .A(DB[387]), .B(DB[356]), .Z(n9616) );
  AND U13472 ( .A(n468), .B(n9617), .Z(n9615) );
  XOR U13473 ( .A(n9618), .B(n9619), .Z(n9617) );
  XOR U13474 ( .A(DB[356]), .B(DB[325]), .Z(n9619) );
  AND U13475 ( .A(n472), .B(n9620), .Z(n9618) );
  XOR U13476 ( .A(n9621), .B(n9622), .Z(n9620) );
  XOR U13477 ( .A(DB[325]), .B(DB[294]), .Z(n9622) );
  AND U13478 ( .A(n476), .B(n9623), .Z(n9621) );
  XOR U13479 ( .A(n9624), .B(n9625), .Z(n9623) );
  XOR U13480 ( .A(DB[294]), .B(DB[263]), .Z(n9625) );
  AND U13481 ( .A(n480), .B(n9626), .Z(n9624) );
  XOR U13482 ( .A(n9627), .B(n9628), .Z(n9626) );
  XOR U13483 ( .A(DB[263]), .B(DB[232]), .Z(n9628) );
  AND U13484 ( .A(n484), .B(n9629), .Z(n9627) );
  XOR U13485 ( .A(n9630), .B(n9631), .Z(n9629) );
  XOR U13486 ( .A(DB[232]), .B(DB[201]), .Z(n9631) );
  AND U13487 ( .A(n488), .B(n9632), .Z(n9630) );
  XOR U13488 ( .A(n9633), .B(n9634), .Z(n9632) );
  XOR U13489 ( .A(DB[201]), .B(DB[170]), .Z(n9634) );
  AND U13490 ( .A(n492), .B(n9635), .Z(n9633) );
  XOR U13491 ( .A(n9636), .B(n9637), .Z(n9635) );
  XOR U13492 ( .A(DB[170]), .B(DB[139]), .Z(n9637) );
  AND U13493 ( .A(n496), .B(n9638), .Z(n9636) );
  XOR U13494 ( .A(n9639), .B(n9640), .Z(n9638) );
  XOR U13495 ( .A(DB[139]), .B(DB[108]), .Z(n9640) );
  AND U13496 ( .A(n500), .B(n9641), .Z(n9639) );
  XOR U13497 ( .A(n9642), .B(n9643), .Z(n9641) );
  XOR U13498 ( .A(DB[77]), .B(DB[108]), .Z(n9643) );
  AND U13499 ( .A(n504), .B(n9644), .Z(n9642) );
  XOR U13500 ( .A(n9645), .B(n9646), .Z(n9644) );
  XOR U13501 ( .A(DB[77]), .B(DB[46]), .Z(n9646) );
  AND U13502 ( .A(n508), .B(n9647), .Z(n9645) );
  XOR U13503 ( .A(DB[46]), .B(DB[15]), .Z(n9647) );
  XOR U13504 ( .A(DB[3951]), .B(n9648), .Z(min_val_out[14]) );
  AND U13505 ( .A(n2), .B(n9649), .Z(n9648) );
  XOR U13506 ( .A(n9650), .B(n9651), .Z(n9649) );
  XOR U13507 ( .A(DB[3951]), .B(DB[3920]), .Z(n9651) );
  AND U13508 ( .A(n8), .B(n9652), .Z(n9650) );
  XOR U13509 ( .A(n9653), .B(n9654), .Z(n9652) );
  XOR U13510 ( .A(DB[3920]), .B(DB[3889]), .Z(n9654) );
  AND U13511 ( .A(n12), .B(n9655), .Z(n9653) );
  XOR U13512 ( .A(n9656), .B(n9657), .Z(n9655) );
  XOR U13513 ( .A(DB[3889]), .B(DB[3858]), .Z(n9657) );
  AND U13514 ( .A(n16), .B(n9658), .Z(n9656) );
  XOR U13515 ( .A(n9659), .B(n9660), .Z(n9658) );
  XOR U13516 ( .A(DB[3858]), .B(DB[3827]), .Z(n9660) );
  AND U13517 ( .A(n20), .B(n9661), .Z(n9659) );
  XOR U13518 ( .A(n9662), .B(n9663), .Z(n9661) );
  XOR U13519 ( .A(DB[3827]), .B(DB[3796]), .Z(n9663) );
  AND U13520 ( .A(n24), .B(n9664), .Z(n9662) );
  XOR U13521 ( .A(n9665), .B(n9666), .Z(n9664) );
  XOR U13522 ( .A(DB[3796]), .B(DB[3765]), .Z(n9666) );
  AND U13523 ( .A(n28), .B(n9667), .Z(n9665) );
  XOR U13524 ( .A(n9668), .B(n9669), .Z(n9667) );
  XOR U13525 ( .A(DB[3765]), .B(DB[3734]), .Z(n9669) );
  AND U13526 ( .A(n32), .B(n9670), .Z(n9668) );
  XOR U13527 ( .A(n9671), .B(n9672), .Z(n9670) );
  XOR U13528 ( .A(DB[3734]), .B(DB[3703]), .Z(n9672) );
  AND U13529 ( .A(n36), .B(n9673), .Z(n9671) );
  XOR U13530 ( .A(n9674), .B(n9675), .Z(n9673) );
  XOR U13531 ( .A(DB[3703]), .B(DB[3672]), .Z(n9675) );
  AND U13532 ( .A(n40), .B(n9676), .Z(n9674) );
  XOR U13533 ( .A(n9677), .B(n9678), .Z(n9676) );
  XOR U13534 ( .A(DB[3672]), .B(DB[3641]), .Z(n9678) );
  AND U13535 ( .A(n44), .B(n9679), .Z(n9677) );
  XOR U13536 ( .A(n9680), .B(n9681), .Z(n9679) );
  XOR U13537 ( .A(DB[3641]), .B(DB[3610]), .Z(n9681) );
  AND U13538 ( .A(n48), .B(n9682), .Z(n9680) );
  XOR U13539 ( .A(n9683), .B(n9684), .Z(n9682) );
  XOR U13540 ( .A(DB[3610]), .B(DB[3579]), .Z(n9684) );
  AND U13541 ( .A(n52), .B(n9685), .Z(n9683) );
  XOR U13542 ( .A(n9686), .B(n9687), .Z(n9685) );
  XOR U13543 ( .A(DB[3579]), .B(DB[3548]), .Z(n9687) );
  AND U13544 ( .A(n56), .B(n9688), .Z(n9686) );
  XOR U13545 ( .A(n9689), .B(n9690), .Z(n9688) );
  XOR U13546 ( .A(DB[3548]), .B(DB[3517]), .Z(n9690) );
  AND U13547 ( .A(n60), .B(n9691), .Z(n9689) );
  XOR U13548 ( .A(n9692), .B(n9693), .Z(n9691) );
  XOR U13549 ( .A(DB[3517]), .B(DB[3486]), .Z(n9693) );
  AND U13550 ( .A(n64), .B(n9694), .Z(n9692) );
  XOR U13551 ( .A(n9695), .B(n9696), .Z(n9694) );
  XOR U13552 ( .A(DB[3486]), .B(DB[3455]), .Z(n9696) );
  AND U13553 ( .A(n68), .B(n9697), .Z(n9695) );
  XOR U13554 ( .A(n9698), .B(n9699), .Z(n9697) );
  XOR U13555 ( .A(DB[3455]), .B(DB[3424]), .Z(n9699) );
  AND U13556 ( .A(n72), .B(n9700), .Z(n9698) );
  XOR U13557 ( .A(n9701), .B(n9702), .Z(n9700) );
  XOR U13558 ( .A(DB[3424]), .B(DB[3393]), .Z(n9702) );
  AND U13559 ( .A(n76), .B(n9703), .Z(n9701) );
  XOR U13560 ( .A(n9704), .B(n9705), .Z(n9703) );
  XOR U13561 ( .A(DB[3393]), .B(DB[3362]), .Z(n9705) );
  AND U13562 ( .A(n80), .B(n9706), .Z(n9704) );
  XOR U13563 ( .A(n9707), .B(n9708), .Z(n9706) );
  XOR U13564 ( .A(DB[3362]), .B(DB[3331]), .Z(n9708) );
  AND U13565 ( .A(n84), .B(n9709), .Z(n9707) );
  XOR U13566 ( .A(n9710), .B(n9711), .Z(n9709) );
  XOR U13567 ( .A(DB[3331]), .B(DB[3300]), .Z(n9711) );
  AND U13568 ( .A(n88), .B(n9712), .Z(n9710) );
  XOR U13569 ( .A(n9713), .B(n9714), .Z(n9712) );
  XOR U13570 ( .A(DB[3300]), .B(DB[3269]), .Z(n9714) );
  AND U13571 ( .A(n92), .B(n9715), .Z(n9713) );
  XOR U13572 ( .A(n9716), .B(n9717), .Z(n9715) );
  XOR U13573 ( .A(DB[3269]), .B(DB[3238]), .Z(n9717) );
  AND U13574 ( .A(n96), .B(n9718), .Z(n9716) );
  XOR U13575 ( .A(n9719), .B(n9720), .Z(n9718) );
  XOR U13576 ( .A(DB[3238]), .B(DB[3207]), .Z(n9720) );
  AND U13577 ( .A(n100), .B(n9721), .Z(n9719) );
  XOR U13578 ( .A(n9722), .B(n9723), .Z(n9721) );
  XOR U13579 ( .A(DB[3207]), .B(DB[3176]), .Z(n9723) );
  AND U13580 ( .A(n104), .B(n9724), .Z(n9722) );
  XOR U13581 ( .A(n9725), .B(n9726), .Z(n9724) );
  XOR U13582 ( .A(DB[3176]), .B(DB[3145]), .Z(n9726) );
  AND U13583 ( .A(n108), .B(n9727), .Z(n9725) );
  XOR U13584 ( .A(n9728), .B(n9729), .Z(n9727) );
  XOR U13585 ( .A(DB[3145]), .B(DB[3114]), .Z(n9729) );
  AND U13586 ( .A(n112), .B(n9730), .Z(n9728) );
  XOR U13587 ( .A(n9731), .B(n9732), .Z(n9730) );
  XOR U13588 ( .A(DB[3114]), .B(DB[3083]), .Z(n9732) );
  AND U13589 ( .A(n116), .B(n9733), .Z(n9731) );
  XOR U13590 ( .A(n9734), .B(n9735), .Z(n9733) );
  XOR U13591 ( .A(DB[3083]), .B(DB[3052]), .Z(n9735) );
  AND U13592 ( .A(n120), .B(n9736), .Z(n9734) );
  XOR U13593 ( .A(n9737), .B(n9738), .Z(n9736) );
  XOR U13594 ( .A(DB[3052]), .B(DB[3021]), .Z(n9738) );
  AND U13595 ( .A(n124), .B(n9739), .Z(n9737) );
  XOR U13596 ( .A(n9740), .B(n9741), .Z(n9739) );
  XOR U13597 ( .A(DB[3021]), .B(DB[2990]), .Z(n9741) );
  AND U13598 ( .A(n128), .B(n9742), .Z(n9740) );
  XOR U13599 ( .A(n9743), .B(n9744), .Z(n9742) );
  XOR U13600 ( .A(DB[2990]), .B(DB[2959]), .Z(n9744) );
  AND U13601 ( .A(n132), .B(n9745), .Z(n9743) );
  XOR U13602 ( .A(n9746), .B(n9747), .Z(n9745) );
  XOR U13603 ( .A(DB[2959]), .B(DB[2928]), .Z(n9747) );
  AND U13604 ( .A(n136), .B(n9748), .Z(n9746) );
  XOR U13605 ( .A(n9749), .B(n9750), .Z(n9748) );
  XOR U13606 ( .A(DB[2928]), .B(DB[2897]), .Z(n9750) );
  AND U13607 ( .A(n140), .B(n9751), .Z(n9749) );
  XOR U13608 ( .A(n9752), .B(n9753), .Z(n9751) );
  XOR U13609 ( .A(DB[2897]), .B(DB[2866]), .Z(n9753) );
  AND U13610 ( .A(n144), .B(n9754), .Z(n9752) );
  XOR U13611 ( .A(n9755), .B(n9756), .Z(n9754) );
  XOR U13612 ( .A(DB[2866]), .B(DB[2835]), .Z(n9756) );
  AND U13613 ( .A(n148), .B(n9757), .Z(n9755) );
  XOR U13614 ( .A(n9758), .B(n9759), .Z(n9757) );
  XOR U13615 ( .A(DB[2835]), .B(DB[2804]), .Z(n9759) );
  AND U13616 ( .A(n152), .B(n9760), .Z(n9758) );
  XOR U13617 ( .A(n9761), .B(n9762), .Z(n9760) );
  XOR U13618 ( .A(DB[2804]), .B(DB[2773]), .Z(n9762) );
  AND U13619 ( .A(n156), .B(n9763), .Z(n9761) );
  XOR U13620 ( .A(n9764), .B(n9765), .Z(n9763) );
  XOR U13621 ( .A(DB[2773]), .B(DB[2742]), .Z(n9765) );
  AND U13622 ( .A(n160), .B(n9766), .Z(n9764) );
  XOR U13623 ( .A(n9767), .B(n9768), .Z(n9766) );
  XOR U13624 ( .A(DB[2742]), .B(DB[2711]), .Z(n9768) );
  AND U13625 ( .A(n164), .B(n9769), .Z(n9767) );
  XOR U13626 ( .A(n9770), .B(n9771), .Z(n9769) );
  XOR U13627 ( .A(DB[2711]), .B(DB[2680]), .Z(n9771) );
  AND U13628 ( .A(n168), .B(n9772), .Z(n9770) );
  XOR U13629 ( .A(n9773), .B(n9774), .Z(n9772) );
  XOR U13630 ( .A(DB[2680]), .B(DB[2649]), .Z(n9774) );
  AND U13631 ( .A(n172), .B(n9775), .Z(n9773) );
  XOR U13632 ( .A(n9776), .B(n9777), .Z(n9775) );
  XOR U13633 ( .A(DB[2649]), .B(DB[2618]), .Z(n9777) );
  AND U13634 ( .A(n176), .B(n9778), .Z(n9776) );
  XOR U13635 ( .A(n9779), .B(n9780), .Z(n9778) );
  XOR U13636 ( .A(DB[2618]), .B(DB[2587]), .Z(n9780) );
  AND U13637 ( .A(n180), .B(n9781), .Z(n9779) );
  XOR U13638 ( .A(n9782), .B(n9783), .Z(n9781) );
  XOR U13639 ( .A(DB[2587]), .B(DB[2556]), .Z(n9783) );
  AND U13640 ( .A(n184), .B(n9784), .Z(n9782) );
  XOR U13641 ( .A(n9785), .B(n9786), .Z(n9784) );
  XOR U13642 ( .A(DB[2556]), .B(DB[2525]), .Z(n9786) );
  AND U13643 ( .A(n188), .B(n9787), .Z(n9785) );
  XOR U13644 ( .A(n9788), .B(n9789), .Z(n9787) );
  XOR U13645 ( .A(DB[2525]), .B(DB[2494]), .Z(n9789) );
  AND U13646 ( .A(n192), .B(n9790), .Z(n9788) );
  XOR U13647 ( .A(n9791), .B(n9792), .Z(n9790) );
  XOR U13648 ( .A(DB[2494]), .B(DB[2463]), .Z(n9792) );
  AND U13649 ( .A(n196), .B(n9793), .Z(n9791) );
  XOR U13650 ( .A(n9794), .B(n9795), .Z(n9793) );
  XOR U13651 ( .A(DB[2463]), .B(DB[2432]), .Z(n9795) );
  AND U13652 ( .A(n200), .B(n9796), .Z(n9794) );
  XOR U13653 ( .A(n9797), .B(n9798), .Z(n9796) );
  XOR U13654 ( .A(DB[2432]), .B(DB[2401]), .Z(n9798) );
  AND U13655 ( .A(n204), .B(n9799), .Z(n9797) );
  XOR U13656 ( .A(n9800), .B(n9801), .Z(n9799) );
  XOR U13657 ( .A(DB[2401]), .B(DB[2370]), .Z(n9801) );
  AND U13658 ( .A(n208), .B(n9802), .Z(n9800) );
  XOR U13659 ( .A(n9803), .B(n9804), .Z(n9802) );
  XOR U13660 ( .A(DB[2370]), .B(DB[2339]), .Z(n9804) );
  AND U13661 ( .A(n212), .B(n9805), .Z(n9803) );
  XOR U13662 ( .A(n9806), .B(n9807), .Z(n9805) );
  XOR U13663 ( .A(DB[2339]), .B(DB[2308]), .Z(n9807) );
  AND U13664 ( .A(n216), .B(n9808), .Z(n9806) );
  XOR U13665 ( .A(n9809), .B(n9810), .Z(n9808) );
  XOR U13666 ( .A(DB[2308]), .B(DB[2277]), .Z(n9810) );
  AND U13667 ( .A(n220), .B(n9811), .Z(n9809) );
  XOR U13668 ( .A(n9812), .B(n9813), .Z(n9811) );
  XOR U13669 ( .A(DB[2277]), .B(DB[2246]), .Z(n9813) );
  AND U13670 ( .A(n224), .B(n9814), .Z(n9812) );
  XOR U13671 ( .A(n9815), .B(n9816), .Z(n9814) );
  XOR U13672 ( .A(DB[2246]), .B(DB[2215]), .Z(n9816) );
  AND U13673 ( .A(n228), .B(n9817), .Z(n9815) );
  XOR U13674 ( .A(n9818), .B(n9819), .Z(n9817) );
  XOR U13675 ( .A(DB[2215]), .B(DB[2184]), .Z(n9819) );
  AND U13676 ( .A(n232), .B(n9820), .Z(n9818) );
  XOR U13677 ( .A(n9821), .B(n9822), .Z(n9820) );
  XOR U13678 ( .A(DB[2184]), .B(DB[2153]), .Z(n9822) );
  AND U13679 ( .A(n236), .B(n9823), .Z(n9821) );
  XOR U13680 ( .A(n9824), .B(n9825), .Z(n9823) );
  XOR U13681 ( .A(DB[2153]), .B(DB[2122]), .Z(n9825) );
  AND U13682 ( .A(n240), .B(n9826), .Z(n9824) );
  XOR U13683 ( .A(n9827), .B(n9828), .Z(n9826) );
  XOR U13684 ( .A(DB[2122]), .B(DB[2091]), .Z(n9828) );
  AND U13685 ( .A(n244), .B(n9829), .Z(n9827) );
  XOR U13686 ( .A(n9830), .B(n9831), .Z(n9829) );
  XOR U13687 ( .A(DB[2091]), .B(DB[2060]), .Z(n9831) );
  AND U13688 ( .A(n248), .B(n9832), .Z(n9830) );
  XOR U13689 ( .A(n9833), .B(n9834), .Z(n9832) );
  XOR U13690 ( .A(DB[2060]), .B(DB[2029]), .Z(n9834) );
  AND U13691 ( .A(n252), .B(n9835), .Z(n9833) );
  XOR U13692 ( .A(n9836), .B(n9837), .Z(n9835) );
  XOR U13693 ( .A(DB[2029]), .B(DB[1998]), .Z(n9837) );
  AND U13694 ( .A(n256), .B(n9838), .Z(n9836) );
  XOR U13695 ( .A(n9839), .B(n9840), .Z(n9838) );
  XOR U13696 ( .A(DB[1998]), .B(DB[1967]), .Z(n9840) );
  AND U13697 ( .A(n260), .B(n9841), .Z(n9839) );
  XOR U13698 ( .A(n9842), .B(n9843), .Z(n9841) );
  XOR U13699 ( .A(DB[1967]), .B(DB[1936]), .Z(n9843) );
  AND U13700 ( .A(n264), .B(n9844), .Z(n9842) );
  XOR U13701 ( .A(n9845), .B(n9846), .Z(n9844) );
  XOR U13702 ( .A(DB[1936]), .B(DB[1905]), .Z(n9846) );
  AND U13703 ( .A(n268), .B(n9847), .Z(n9845) );
  XOR U13704 ( .A(n9848), .B(n9849), .Z(n9847) );
  XOR U13705 ( .A(DB[1905]), .B(DB[1874]), .Z(n9849) );
  AND U13706 ( .A(n272), .B(n9850), .Z(n9848) );
  XOR U13707 ( .A(n9851), .B(n9852), .Z(n9850) );
  XOR U13708 ( .A(DB[1874]), .B(DB[1843]), .Z(n9852) );
  AND U13709 ( .A(n276), .B(n9853), .Z(n9851) );
  XOR U13710 ( .A(n9854), .B(n9855), .Z(n9853) );
  XOR U13711 ( .A(DB[1843]), .B(DB[1812]), .Z(n9855) );
  AND U13712 ( .A(n280), .B(n9856), .Z(n9854) );
  XOR U13713 ( .A(n9857), .B(n9858), .Z(n9856) );
  XOR U13714 ( .A(DB[1812]), .B(DB[1781]), .Z(n9858) );
  AND U13715 ( .A(n284), .B(n9859), .Z(n9857) );
  XOR U13716 ( .A(n9860), .B(n9861), .Z(n9859) );
  XOR U13717 ( .A(DB[1781]), .B(DB[1750]), .Z(n9861) );
  AND U13718 ( .A(n288), .B(n9862), .Z(n9860) );
  XOR U13719 ( .A(n9863), .B(n9864), .Z(n9862) );
  XOR U13720 ( .A(DB[1750]), .B(DB[1719]), .Z(n9864) );
  AND U13721 ( .A(n292), .B(n9865), .Z(n9863) );
  XOR U13722 ( .A(n9866), .B(n9867), .Z(n9865) );
  XOR U13723 ( .A(DB[1719]), .B(DB[1688]), .Z(n9867) );
  AND U13724 ( .A(n296), .B(n9868), .Z(n9866) );
  XOR U13725 ( .A(n9869), .B(n9870), .Z(n9868) );
  XOR U13726 ( .A(DB[1688]), .B(DB[1657]), .Z(n9870) );
  AND U13727 ( .A(n300), .B(n9871), .Z(n9869) );
  XOR U13728 ( .A(n9872), .B(n9873), .Z(n9871) );
  XOR U13729 ( .A(DB[1657]), .B(DB[1626]), .Z(n9873) );
  AND U13730 ( .A(n304), .B(n9874), .Z(n9872) );
  XOR U13731 ( .A(n9875), .B(n9876), .Z(n9874) );
  XOR U13732 ( .A(DB[1626]), .B(DB[1595]), .Z(n9876) );
  AND U13733 ( .A(n308), .B(n9877), .Z(n9875) );
  XOR U13734 ( .A(n9878), .B(n9879), .Z(n9877) );
  XOR U13735 ( .A(DB[1595]), .B(DB[1564]), .Z(n9879) );
  AND U13736 ( .A(n312), .B(n9880), .Z(n9878) );
  XOR U13737 ( .A(n9881), .B(n9882), .Z(n9880) );
  XOR U13738 ( .A(DB[1564]), .B(DB[1533]), .Z(n9882) );
  AND U13739 ( .A(n316), .B(n9883), .Z(n9881) );
  XOR U13740 ( .A(n9884), .B(n9885), .Z(n9883) );
  XOR U13741 ( .A(DB[1533]), .B(DB[1502]), .Z(n9885) );
  AND U13742 ( .A(n320), .B(n9886), .Z(n9884) );
  XOR U13743 ( .A(n9887), .B(n9888), .Z(n9886) );
  XOR U13744 ( .A(DB[1502]), .B(DB[1471]), .Z(n9888) );
  AND U13745 ( .A(n324), .B(n9889), .Z(n9887) );
  XOR U13746 ( .A(n9890), .B(n9891), .Z(n9889) );
  XOR U13747 ( .A(DB[1471]), .B(DB[1440]), .Z(n9891) );
  AND U13748 ( .A(n328), .B(n9892), .Z(n9890) );
  XOR U13749 ( .A(n9893), .B(n9894), .Z(n9892) );
  XOR U13750 ( .A(DB[1440]), .B(DB[1409]), .Z(n9894) );
  AND U13751 ( .A(n332), .B(n9895), .Z(n9893) );
  XOR U13752 ( .A(n9896), .B(n9897), .Z(n9895) );
  XOR U13753 ( .A(DB[1409]), .B(DB[1378]), .Z(n9897) );
  AND U13754 ( .A(n336), .B(n9898), .Z(n9896) );
  XOR U13755 ( .A(n9899), .B(n9900), .Z(n9898) );
  XOR U13756 ( .A(DB[1378]), .B(DB[1347]), .Z(n9900) );
  AND U13757 ( .A(n340), .B(n9901), .Z(n9899) );
  XOR U13758 ( .A(n9902), .B(n9903), .Z(n9901) );
  XOR U13759 ( .A(DB[1347]), .B(DB[1316]), .Z(n9903) );
  AND U13760 ( .A(n344), .B(n9904), .Z(n9902) );
  XOR U13761 ( .A(n9905), .B(n9906), .Z(n9904) );
  XOR U13762 ( .A(DB[1316]), .B(DB[1285]), .Z(n9906) );
  AND U13763 ( .A(n348), .B(n9907), .Z(n9905) );
  XOR U13764 ( .A(n9908), .B(n9909), .Z(n9907) );
  XOR U13765 ( .A(DB[1285]), .B(DB[1254]), .Z(n9909) );
  AND U13766 ( .A(n352), .B(n9910), .Z(n9908) );
  XOR U13767 ( .A(n9911), .B(n9912), .Z(n9910) );
  XOR U13768 ( .A(DB[1254]), .B(DB[1223]), .Z(n9912) );
  AND U13769 ( .A(n356), .B(n9913), .Z(n9911) );
  XOR U13770 ( .A(n9914), .B(n9915), .Z(n9913) );
  XOR U13771 ( .A(DB[1223]), .B(DB[1192]), .Z(n9915) );
  AND U13772 ( .A(n360), .B(n9916), .Z(n9914) );
  XOR U13773 ( .A(n9917), .B(n9918), .Z(n9916) );
  XOR U13774 ( .A(DB[1192]), .B(DB[1161]), .Z(n9918) );
  AND U13775 ( .A(n364), .B(n9919), .Z(n9917) );
  XOR U13776 ( .A(n9920), .B(n9921), .Z(n9919) );
  XOR U13777 ( .A(DB[1161]), .B(DB[1130]), .Z(n9921) );
  AND U13778 ( .A(n368), .B(n9922), .Z(n9920) );
  XOR U13779 ( .A(n9923), .B(n9924), .Z(n9922) );
  XOR U13780 ( .A(DB[1130]), .B(DB[1099]), .Z(n9924) );
  AND U13781 ( .A(n372), .B(n9925), .Z(n9923) );
  XOR U13782 ( .A(n9926), .B(n9927), .Z(n9925) );
  XOR U13783 ( .A(DB[1099]), .B(DB[1068]), .Z(n9927) );
  AND U13784 ( .A(n376), .B(n9928), .Z(n9926) );
  XOR U13785 ( .A(n9929), .B(n9930), .Z(n9928) );
  XOR U13786 ( .A(DB[1068]), .B(DB[1037]), .Z(n9930) );
  AND U13787 ( .A(n380), .B(n9931), .Z(n9929) );
  XOR U13788 ( .A(n9932), .B(n9933), .Z(n9931) );
  XOR U13789 ( .A(DB[1037]), .B(DB[1006]), .Z(n9933) );
  AND U13790 ( .A(n384), .B(n9934), .Z(n9932) );
  XOR U13791 ( .A(n9935), .B(n9936), .Z(n9934) );
  XOR U13792 ( .A(DB[975]), .B(DB[1006]), .Z(n9936) );
  AND U13793 ( .A(n388), .B(n9937), .Z(n9935) );
  XOR U13794 ( .A(n9938), .B(n9939), .Z(n9937) );
  XOR U13795 ( .A(DB[975]), .B(DB[944]), .Z(n9939) );
  AND U13796 ( .A(n392), .B(n9940), .Z(n9938) );
  XOR U13797 ( .A(n9941), .B(n9942), .Z(n9940) );
  XOR U13798 ( .A(DB[944]), .B(DB[913]), .Z(n9942) );
  AND U13799 ( .A(n396), .B(n9943), .Z(n9941) );
  XOR U13800 ( .A(n9944), .B(n9945), .Z(n9943) );
  XOR U13801 ( .A(DB[913]), .B(DB[882]), .Z(n9945) );
  AND U13802 ( .A(n400), .B(n9946), .Z(n9944) );
  XOR U13803 ( .A(n9947), .B(n9948), .Z(n9946) );
  XOR U13804 ( .A(DB[882]), .B(DB[851]), .Z(n9948) );
  AND U13805 ( .A(n404), .B(n9949), .Z(n9947) );
  XOR U13806 ( .A(n9950), .B(n9951), .Z(n9949) );
  XOR U13807 ( .A(DB[851]), .B(DB[820]), .Z(n9951) );
  AND U13808 ( .A(n408), .B(n9952), .Z(n9950) );
  XOR U13809 ( .A(n9953), .B(n9954), .Z(n9952) );
  XOR U13810 ( .A(DB[820]), .B(DB[789]), .Z(n9954) );
  AND U13811 ( .A(n412), .B(n9955), .Z(n9953) );
  XOR U13812 ( .A(n9956), .B(n9957), .Z(n9955) );
  XOR U13813 ( .A(DB[789]), .B(DB[758]), .Z(n9957) );
  AND U13814 ( .A(n416), .B(n9958), .Z(n9956) );
  XOR U13815 ( .A(n9959), .B(n9960), .Z(n9958) );
  XOR U13816 ( .A(DB[758]), .B(DB[727]), .Z(n9960) );
  AND U13817 ( .A(n420), .B(n9961), .Z(n9959) );
  XOR U13818 ( .A(n9962), .B(n9963), .Z(n9961) );
  XOR U13819 ( .A(DB[727]), .B(DB[696]), .Z(n9963) );
  AND U13820 ( .A(n424), .B(n9964), .Z(n9962) );
  XOR U13821 ( .A(n9965), .B(n9966), .Z(n9964) );
  XOR U13822 ( .A(DB[696]), .B(DB[665]), .Z(n9966) );
  AND U13823 ( .A(n428), .B(n9967), .Z(n9965) );
  XOR U13824 ( .A(n9968), .B(n9969), .Z(n9967) );
  XOR U13825 ( .A(DB[665]), .B(DB[634]), .Z(n9969) );
  AND U13826 ( .A(n432), .B(n9970), .Z(n9968) );
  XOR U13827 ( .A(n9971), .B(n9972), .Z(n9970) );
  XOR U13828 ( .A(DB[634]), .B(DB[603]), .Z(n9972) );
  AND U13829 ( .A(n436), .B(n9973), .Z(n9971) );
  XOR U13830 ( .A(n9974), .B(n9975), .Z(n9973) );
  XOR U13831 ( .A(DB[603]), .B(DB[572]), .Z(n9975) );
  AND U13832 ( .A(n440), .B(n9976), .Z(n9974) );
  XOR U13833 ( .A(n9977), .B(n9978), .Z(n9976) );
  XOR U13834 ( .A(DB[572]), .B(DB[541]), .Z(n9978) );
  AND U13835 ( .A(n444), .B(n9979), .Z(n9977) );
  XOR U13836 ( .A(n9980), .B(n9981), .Z(n9979) );
  XOR U13837 ( .A(DB[541]), .B(DB[510]), .Z(n9981) );
  AND U13838 ( .A(n448), .B(n9982), .Z(n9980) );
  XOR U13839 ( .A(n9983), .B(n9984), .Z(n9982) );
  XOR U13840 ( .A(DB[510]), .B(DB[479]), .Z(n9984) );
  AND U13841 ( .A(n452), .B(n9985), .Z(n9983) );
  XOR U13842 ( .A(n9986), .B(n9987), .Z(n9985) );
  XOR U13843 ( .A(DB[479]), .B(DB[448]), .Z(n9987) );
  AND U13844 ( .A(n456), .B(n9988), .Z(n9986) );
  XOR U13845 ( .A(n9989), .B(n9990), .Z(n9988) );
  XOR U13846 ( .A(DB[448]), .B(DB[417]), .Z(n9990) );
  AND U13847 ( .A(n460), .B(n9991), .Z(n9989) );
  XOR U13848 ( .A(n9992), .B(n9993), .Z(n9991) );
  XOR U13849 ( .A(DB[417]), .B(DB[386]), .Z(n9993) );
  AND U13850 ( .A(n464), .B(n9994), .Z(n9992) );
  XOR U13851 ( .A(n9995), .B(n9996), .Z(n9994) );
  XOR U13852 ( .A(DB[386]), .B(DB[355]), .Z(n9996) );
  AND U13853 ( .A(n468), .B(n9997), .Z(n9995) );
  XOR U13854 ( .A(n9998), .B(n9999), .Z(n9997) );
  XOR U13855 ( .A(DB[355]), .B(DB[324]), .Z(n9999) );
  AND U13856 ( .A(n472), .B(n10000), .Z(n9998) );
  XOR U13857 ( .A(n10001), .B(n10002), .Z(n10000) );
  XOR U13858 ( .A(DB[324]), .B(DB[293]), .Z(n10002) );
  AND U13859 ( .A(n476), .B(n10003), .Z(n10001) );
  XOR U13860 ( .A(n10004), .B(n10005), .Z(n10003) );
  XOR U13861 ( .A(DB[293]), .B(DB[262]), .Z(n10005) );
  AND U13862 ( .A(n480), .B(n10006), .Z(n10004) );
  XOR U13863 ( .A(n10007), .B(n10008), .Z(n10006) );
  XOR U13864 ( .A(DB[262]), .B(DB[231]), .Z(n10008) );
  AND U13865 ( .A(n484), .B(n10009), .Z(n10007) );
  XOR U13866 ( .A(n10010), .B(n10011), .Z(n10009) );
  XOR U13867 ( .A(DB[231]), .B(DB[200]), .Z(n10011) );
  AND U13868 ( .A(n488), .B(n10012), .Z(n10010) );
  XOR U13869 ( .A(n10013), .B(n10014), .Z(n10012) );
  XOR U13870 ( .A(DB[200]), .B(DB[169]), .Z(n10014) );
  AND U13871 ( .A(n492), .B(n10015), .Z(n10013) );
  XOR U13872 ( .A(n10016), .B(n10017), .Z(n10015) );
  XOR U13873 ( .A(DB[169]), .B(DB[138]), .Z(n10017) );
  AND U13874 ( .A(n496), .B(n10018), .Z(n10016) );
  XOR U13875 ( .A(n10019), .B(n10020), .Z(n10018) );
  XOR U13876 ( .A(DB[138]), .B(DB[107]), .Z(n10020) );
  AND U13877 ( .A(n500), .B(n10021), .Z(n10019) );
  XOR U13878 ( .A(n10022), .B(n10023), .Z(n10021) );
  XOR U13879 ( .A(DB[76]), .B(DB[107]), .Z(n10023) );
  AND U13880 ( .A(n504), .B(n10024), .Z(n10022) );
  XOR U13881 ( .A(n10025), .B(n10026), .Z(n10024) );
  XOR U13882 ( .A(DB[76]), .B(DB[45]), .Z(n10026) );
  AND U13883 ( .A(n508), .B(n10027), .Z(n10025) );
  XOR U13884 ( .A(DB[45]), .B(DB[14]), .Z(n10027) );
  XOR U13885 ( .A(DB[3950]), .B(n10028), .Z(min_val_out[13]) );
  AND U13886 ( .A(n2), .B(n10029), .Z(n10028) );
  XOR U13887 ( .A(n10030), .B(n10031), .Z(n10029) );
  XOR U13888 ( .A(n10032), .B(n10033), .Z(n10031) );
  IV U13889 ( .A(DB[3950]), .Z(n10032) );
  AND U13890 ( .A(n8), .B(n10034), .Z(n10030) );
  XOR U13891 ( .A(n10035), .B(n10036), .Z(n10034) );
  XOR U13892 ( .A(DB[3919]), .B(DB[3888]), .Z(n10036) );
  AND U13893 ( .A(n12), .B(n10037), .Z(n10035) );
  XOR U13894 ( .A(n10038), .B(n10039), .Z(n10037) );
  XOR U13895 ( .A(DB[3888]), .B(DB[3857]), .Z(n10039) );
  AND U13896 ( .A(n16), .B(n10040), .Z(n10038) );
  XOR U13897 ( .A(n10041), .B(n10042), .Z(n10040) );
  XOR U13898 ( .A(DB[3857]), .B(DB[3826]), .Z(n10042) );
  AND U13899 ( .A(n20), .B(n10043), .Z(n10041) );
  XOR U13900 ( .A(n10044), .B(n10045), .Z(n10043) );
  XOR U13901 ( .A(DB[3826]), .B(DB[3795]), .Z(n10045) );
  AND U13902 ( .A(n24), .B(n10046), .Z(n10044) );
  XOR U13903 ( .A(n10047), .B(n10048), .Z(n10046) );
  XOR U13904 ( .A(DB[3795]), .B(DB[3764]), .Z(n10048) );
  AND U13905 ( .A(n28), .B(n10049), .Z(n10047) );
  XOR U13906 ( .A(n10050), .B(n10051), .Z(n10049) );
  XOR U13907 ( .A(DB[3764]), .B(DB[3733]), .Z(n10051) );
  AND U13908 ( .A(n32), .B(n10052), .Z(n10050) );
  XOR U13909 ( .A(n10053), .B(n10054), .Z(n10052) );
  XOR U13910 ( .A(DB[3733]), .B(DB[3702]), .Z(n10054) );
  AND U13911 ( .A(n36), .B(n10055), .Z(n10053) );
  XOR U13912 ( .A(n10056), .B(n10057), .Z(n10055) );
  XOR U13913 ( .A(DB[3702]), .B(DB[3671]), .Z(n10057) );
  AND U13914 ( .A(n40), .B(n10058), .Z(n10056) );
  XOR U13915 ( .A(n10059), .B(n10060), .Z(n10058) );
  XOR U13916 ( .A(DB[3671]), .B(DB[3640]), .Z(n10060) );
  AND U13917 ( .A(n44), .B(n10061), .Z(n10059) );
  XOR U13918 ( .A(n10062), .B(n10063), .Z(n10061) );
  XOR U13919 ( .A(DB[3640]), .B(DB[3609]), .Z(n10063) );
  AND U13920 ( .A(n48), .B(n10064), .Z(n10062) );
  XOR U13921 ( .A(n10065), .B(n10066), .Z(n10064) );
  XOR U13922 ( .A(DB[3609]), .B(DB[3578]), .Z(n10066) );
  AND U13923 ( .A(n52), .B(n10067), .Z(n10065) );
  XOR U13924 ( .A(n10068), .B(n10069), .Z(n10067) );
  XOR U13925 ( .A(DB[3578]), .B(DB[3547]), .Z(n10069) );
  AND U13926 ( .A(n56), .B(n10070), .Z(n10068) );
  XOR U13927 ( .A(n10071), .B(n10072), .Z(n10070) );
  XOR U13928 ( .A(DB[3547]), .B(DB[3516]), .Z(n10072) );
  AND U13929 ( .A(n60), .B(n10073), .Z(n10071) );
  XOR U13930 ( .A(n10074), .B(n10075), .Z(n10073) );
  XOR U13931 ( .A(DB[3516]), .B(DB[3485]), .Z(n10075) );
  AND U13932 ( .A(n64), .B(n10076), .Z(n10074) );
  XOR U13933 ( .A(n10077), .B(n10078), .Z(n10076) );
  XOR U13934 ( .A(DB[3485]), .B(DB[3454]), .Z(n10078) );
  AND U13935 ( .A(n68), .B(n10079), .Z(n10077) );
  XOR U13936 ( .A(n10080), .B(n10081), .Z(n10079) );
  XOR U13937 ( .A(DB[3454]), .B(DB[3423]), .Z(n10081) );
  AND U13938 ( .A(n72), .B(n10082), .Z(n10080) );
  XOR U13939 ( .A(n10083), .B(n10084), .Z(n10082) );
  XOR U13940 ( .A(DB[3423]), .B(DB[3392]), .Z(n10084) );
  AND U13941 ( .A(n76), .B(n10085), .Z(n10083) );
  XOR U13942 ( .A(n10086), .B(n10087), .Z(n10085) );
  XOR U13943 ( .A(DB[3392]), .B(DB[3361]), .Z(n10087) );
  AND U13944 ( .A(n80), .B(n10088), .Z(n10086) );
  XOR U13945 ( .A(n10089), .B(n10090), .Z(n10088) );
  XOR U13946 ( .A(DB[3361]), .B(DB[3330]), .Z(n10090) );
  AND U13947 ( .A(n84), .B(n10091), .Z(n10089) );
  XOR U13948 ( .A(n10092), .B(n10093), .Z(n10091) );
  XOR U13949 ( .A(DB[3330]), .B(DB[3299]), .Z(n10093) );
  AND U13950 ( .A(n88), .B(n10094), .Z(n10092) );
  XOR U13951 ( .A(n10095), .B(n10096), .Z(n10094) );
  XOR U13952 ( .A(DB[3299]), .B(DB[3268]), .Z(n10096) );
  AND U13953 ( .A(n92), .B(n10097), .Z(n10095) );
  XOR U13954 ( .A(n10098), .B(n10099), .Z(n10097) );
  XOR U13955 ( .A(DB[3268]), .B(DB[3237]), .Z(n10099) );
  AND U13956 ( .A(n96), .B(n10100), .Z(n10098) );
  XOR U13957 ( .A(n10101), .B(n10102), .Z(n10100) );
  XOR U13958 ( .A(DB[3237]), .B(DB[3206]), .Z(n10102) );
  AND U13959 ( .A(n100), .B(n10103), .Z(n10101) );
  XOR U13960 ( .A(n10104), .B(n10105), .Z(n10103) );
  XOR U13961 ( .A(DB[3206]), .B(DB[3175]), .Z(n10105) );
  AND U13962 ( .A(n104), .B(n10106), .Z(n10104) );
  XOR U13963 ( .A(n10107), .B(n10108), .Z(n10106) );
  XOR U13964 ( .A(DB[3175]), .B(DB[3144]), .Z(n10108) );
  AND U13965 ( .A(n108), .B(n10109), .Z(n10107) );
  XOR U13966 ( .A(n10110), .B(n10111), .Z(n10109) );
  XOR U13967 ( .A(DB[3144]), .B(DB[3113]), .Z(n10111) );
  AND U13968 ( .A(n112), .B(n10112), .Z(n10110) );
  XOR U13969 ( .A(n10113), .B(n10114), .Z(n10112) );
  XOR U13970 ( .A(DB[3113]), .B(DB[3082]), .Z(n10114) );
  AND U13971 ( .A(n116), .B(n10115), .Z(n10113) );
  XOR U13972 ( .A(n10116), .B(n10117), .Z(n10115) );
  XOR U13973 ( .A(DB[3082]), .B(DB[3051]), .Z(n10117) );
  AND U13974 ( .A(n120), .B(n10118), .Z(n10116) );
  XOR U13975 ( .A(n10119), .B(n10120), .Z(n10118) );
  XOR U13976 ( .A(DB[3051]), .B(DB[3020]), .Z(n10120) );
  AND U13977 ( .A(n124), .B(n10121), .Z(n10119) );
  XOR U13978 ( .A(n10122), .B(n10123), .Z(n10121) );
  XOR U13979 ( .A(DB[3020]), .B(DB[2989]), .Z(n10123) );
  AND U13980 ( .A(n128), .B(n10124), .Z(n10122) );
  XOR U13981 ( .A(n10125), .B(n10126), .Z(n10124) );
  XOR U13982 ( .A(DB[2989]), .B(DB[2958]), .Z(n10126) );
  AND U13983 ( .A(n132), .B(n10127), .Z(n10125) );
  XOR U13984 ( .A(n10128), .B(n10129), .Z(n10127) );
  XOR U13985 ( .A(DB[2958]), .B(DB[2927]), .Z(n10129) );
  AND U13986 ( .A(n136), .B(n10130), .Z(n10128) );
  XOR U13987 ( .A(n10131), .B(n10132), .Z(n10130) );
  XOR U13988 ( .A(DB[2927]), .B(DB[2896]), .Z(n10132) );
  AND U13989 ( .A(n140), .B(n10133), .Z(n10131) );
  XOR U13990 ( .A(n10134), .B(n10135), .Z(n10133) );
  XOR U13991 ( .A(DB[2896]), .B(DB[2865]), .Z(n10135) );
  AND U13992 ( .A(n144), .B(n10136), .Z(n10134) );
  XOR U13993 ( .A(n10137), .B(n10138), .Z(n10136) );
  XOR U13994 ( .A(DB[2865]), .B(DB[2834]), .Z(n10138) );
  AND U13995 ( .A(n148), .B(n10139), .Z(n10137) );
  XOR U13996 ( .A(n10140), .B(n10141), .Z(n10139) );
  XOR U13997 ( .A(DB[2834]), .B(DB[2803]), .Z(n10141) );
  AND U13998 ( .A(n152), .B(n10142), .Z(n10140) );
  XOR U13999 ( .A(n10143), .B(n10144), .Z(n10142) );
  XOR U14000 ( .A(DB[2803]), .B(DB[2772]), .Z(n10144) );
  AND U14001 ( .A(n156), .B(n10145), .Z(n10143) );
  XOR U14002 ( .A(n10146), .B(n10147), .Z(n10145) );
  XOR U14003 ( .A(DB[2772]), .B(DB[2741]), .Z(n10147) );
  AND U14004 ( .A(n160), .B(n10148), .Z(n10146) );
  XOR U14005 ( .A(n10149), .B(n10150), .Z(n10148) );
  XOR U14006 ( .A(DB[2741]), .B(DB[2710]), .Z(n10150) );
  AND U14007 ( .A(n164), .B(n10151), .Z(n10149) );
  XOR U14008 ( .A(n10152), .B(n10153), .Z(n10151) );
  XOR U14009 ( .A(DB[2710]), .B(DB[2679]), .Z(n10153) );
  AND U14010 ( .A(n168), .B(n10154), .Z(n10152) );
  XOR U14011 ( .A(n10155), .B(n10156), .Z(n10154) );
  XOR U14012 ( .A(DB[2679]), .B(DB[2648]), .Z(n10156) );
  AND U14013 ( .A(n172), .B(n10157), .Z(n10155) );
  XOR U14014 ( .A(n10158), .B(n10159), .Z(n10157) );
  XOR U14015 ( .A(DB[2648]), .B(DB[2617]), .Z(n10159) );
  AND U14016 ( .A(n176), .B(n10160), .Z(n10158) );
  XOR U14017 ( .A(n10161), .B(n10162), .Z(n10160) );
  XOR U14018 ( .A(DB[2617]), .B(DB[2586]), .Z(n10162) );
  AND U14019 ( .A(n180), .B(n10163), .Z(n10161) );
  XOR U14020 ( .A(n10164), .B(n10165), .Z(n10163) );
  XOR U14021 ( .A(DB[2586]), .B(DB[2555]), .Z(n10165) );
  AND U14022 ( .A(n184), .B(n10166), .Z(n10164) );
  XOR U14023 ( .A(n10167), .B(n10168), .Z(n10166) );
  XOR U14024 ( .A(DB[2555]), .B(DB[2524]), .Z(n10168) );
  AND U14025 ( .A(n188), .B(n10169), .Z(n10167) );
  XOR U14026 ( .A(n10170), .B(n10171), .Z(n10169) );
  XOR U14027 ( .A(DB[2524]), .B(DB[2493]), .Z(n10171) );
  AND U14028 ( .A(n192), .B(n10172), .Z(n10170) );
  XOR U14029 ( .A(n10173), .B(n10174), .Z(n10172) );
  XOR U14030 ( .A(DB[2493]), .B(DB[2462]), .Z(n10174) );
  AND U14031 ( .A(n196), .B(n10175), .Z(n10173) );
  XOR U14032 ( .A(n10176), .B(n10177), .Z(n10175) );
  XOR U14033 ( .A(DB[2462]), .B(DB[2431]), .Z(n10177) );
  AND U14034 ( .A(n200), .B(n10178), .Z(n10176) );
  XOR U14035 ( .A(n10179), .B(n10180), .Z(n10178) );
  XOR U14036 ( .A(DB[2431]), .B(DB[2400]), .Z(n10180) );
  AND U14037 ( .A(n204), .B(n10181), .Z(n10179) );
  XOR U14038 ( .A(n10182), .B(n10183), .Z(n10181) );
  XOR U14039 ( .A(DB[2400]), .B(DB[2369]), .Z(n10183) );
  AND U14040 ( .A(n208), .B(n10184), .Z(n10182) );
  XOR U14041 ( .A(n10185), .B(n10186), .Z(n10184) );
  XOR U14042 ( .A(DB[2369]), .B(DB[2338]), .Z(n10186) );
  AND U14043 ( .A(n212), .B(n10187), .Z(n10185) );
  XOR U14044 ( .A(n10188), .B(n10189), .Z(n10187) );
  XOR U14045 ( .A(DB[2338]), .B(DB[2307]), .Z(n10189) );
  AND U14046 ( .A(n216), .B(n10190), .Z(n10188) );
  XOR U14047 ( .A(n10191), .B(n10192), .Z(n10190) );
  XOR U14048 ( .A(DB[2307]), .B(DB[2276]), .Z(n10192) );
  AND U14049 ( .A(n220), .B(n10193), .Z(n10191) );
  XOR U14050 ( .A(n10194), .B(n10195), .Z(n10193) );
  XOR U14051 ( .A(DB[2276]), .B(DB[2245]), .Z(n10195) );
  AND U14052 ( .A(n224), .B(n10196), .Z(n10194) );
  XOR U14053 ( .A(n10197), .B(n10198), .Z(n10196) );
  XOR U14054 ( .A(DB[2245]), .B(DB[2214]), .Z(n10198) );
  AND U14055 ( .A(n228), .B(n10199), .Z(n10197) );
  XOR U14056 ( .A(n10200), .B(n10201), .Z(n10199) );
  XOR U14057 ( .A(DB[2214]), .B(DB[2183]), .Z(n10201) );
  AND U14058 ( .A(n232), .B(n10202), .Z(n10200) );
  XOR U14059 ( .A(n10203), .B(n10204), .Z(n10202) );
  XOR U14060 ( .A(DB[2183]), .B(DB[2152]), .Z(n10204) );
  AND U14061 ( .A(n236), .B(n10205), .Z(n10203) );
  XOR U14062 ( .A(n10206), .B(n10207), .Z(n10205) );
  XOR U14063 ( .A(DB[2152]), .B(DB[2121]), .Z(n10207) );
  AND U14064 ( .A(n240), .B(n10208), .Z(n10206) );
  XOR U14065 ( .A(n10209), .B(n10210), .Z(n10208) );
  XOR U14066 ( .A(DB[2121]), .B(DB[2090]), .Z(n10210) );
  AND U14067 ( .A(n244), .B(n10211), .Z(n10209) );
  XOR U14068 ( .A(n10212), .B(n10213), .Z(n10211) );
  XOR U14069 ( .A(DB[2090]), .B(DB[2059]), .Z(n10213) );
  AND U14070 ( .A(n248), .B(n10214), .Z(n10212) );
  XOR U14071 ( .A(n10215), .B(n10216), .Z(n10214) );
  XOR U14072 ( .A(DB[2059]), .B(DB[2028]), .Z(n10216) );
  AND U14073 ( .A(n252), .B(n10217), .Z(n10215) );
  XOR U14074 ( .A(n10218), .B(n10219), .Z(n10217) );
  XOR U14075 ( .A(DB[2028]), .B(DB[1997]), .Z(n10219) );
  AND U14076 ( .A(n256), .B(n10220), .Z(n10218) );
  XOR U14077 ( .A(n10221), .B(n10222), .Z(n10220) );
  XOR U14078 ( .A(DB[1997]), .B(DB[1966]), .Z(n10222) );
  AND U14079 ( .A(n260), .B(n10223), .Z(n10221) );
  XOR U14080 ( .A(n10224), .B(n10225), .Z(n10223) );
  XOR U14081 ( .A(DB[1966]), .B(DB[1935]), .Z(n10225) );
  AND U14082 ( .A(n264), .B(n10226), .Z(n10224) );
  XOR U14083 ( .A(n10227), .B(n10228), .Z(n10226) );
  XOR U14084 ( .A(DB[1935]), .B(DB[1904]), .Z(n10228) );
  AND U14085 ( .A(n268), .B(n10229), .Z(n10227) );
  XOR U14086 ( .A(n10230), .B(n10231), .Z(n10229) );
  XOR U14087 ( .A(DB[1904]), .B(DB[1873]), .Z(n10231) );
  AND U14088 ( .A(n272), .B(n10232), .Z(n10230) );
  XOR U14089 ( .A(n10233), .B(n10234), .Z(n10232) );
  XOR U14090 ( .A(DB[1873]), .B(DB[1842]), .Z(n10234) );
  AND U14091 ( .A(n276), .B(n10235), .Z(n10233) );
  XOR U14092 ( .A(n10236), .B(n10237), .Z(n10235) );
  XOR U14093 ( .A(DB[1842]), .B(DB[1811]), .Z(n10237) );
  AND U14094 ( .A(n280), .B(n10238), .Z(n10236) );
  XOR U14095 ( .A(n10239), .B(n10240), .Z(n10238) );
  XOR U14096 ( .A(DB[1811]), .B(DB[1780]), .Z(n10240) );
  AND U14097 ( .A(n284), .B(n10241), .Z(n10239) );
  XOR U14098 ( .A(n10242), .B(n10243), .Z(n10241) );
  XOR U14099 ( .A(DB[1780]), .B(DB[1749]), .Z(n10243) );
  AND U14100 ( .A(n288), .B(n10244), .Z(n10242) );
  XOR U14101 ( .A(n10245), .B(n10246), .Z(n10244) );
  XOR U14102 ( .A(DB[1749]), .B(DB[1718]), .Z(n10246) );
  AND U14103 ( .A(n292), .B(n10247), .Z(n10245) );
  XOR U14104 ( .A(n10248), .B(n10249), .Z(n10247) );
  XOR U14105 ( .A(DB[1718]), .B(DB[1687]), .Z(n10249) );
  AND U14106 ( .A(n296), .B(n10250), .Z(n10248) );
  XOR U14107 ( .A(n10251), .B(n10252), .Z(n10250) );
  XOR U14108 ( .A(DB[1687]), .B(DB[1656]), .Z(n10252) );
  AND U14109 ( .A(n300), .B(n10253), .Z(n10251) );
  XOR U14110 ( .A(n10254), .B(n10255), .Z(n10253) );
  XOR U14111 ( .A(DB[1656]), .B(DB[1625]), .Z(n10255) );
  AND U14112 ( .A(n304), .B(n10256), .Z(n10254) );
  XOR U14113 ( .A(n10257), .B(n10258), .Z(n10256) );
  XOR U14114 ( .A(DB[1625]), .B(DB[1594]), .Z(n10258) );
  AND U14115 ( .A(n308), .B(n10259), .Z(n10257) );
  XOR U14116 ( .A(n10260), .B(n10261), .Z(n10259) );
  XOR U14117 ( .A(DB[1594]), .B(DB[1563]), .Z(n10261) );
  AND U14118 ( .A(n312), .B(n10262), .Z(n10260) );
  XOR U14119 ( .A(n10263), .B(n10264), .Z(n10262) );
  XOR U14120 ( .A(DB[1563]), .B(DB[1532]), .Z(n10264) );
  AND U14121 ( .A(n316), .B(n10265), .Z(n10263) );
  XOR U14122 ( .A(n10266), .B(n10267), .Z(n10265) );
  XOR U14123 ( .A(DB[1532]), .B(DB[1501]), .Z(n10267) );
  AND U14124 ( .A(n320), .B(n10268), .Z(n10266) );
  XOR U14125 ( .A(n10269), .B(n10270), .Z(n10268) );
  XOR U14126 ( .A(DB[1501]), .B(DB[1470]), .Z(n10270) );
  AND U14127 ( .A(n324), .B(n10271), .Z(n10269) );
  XOR U14128 ( .A(n10272), .B(n10273), .Z(n10271) );
  XOR U14129 ( .A(DB[1470]), .B(DB[1439]), .Z(n10273) );
  AND U14130 ( .A(n328), .B(n10274), .Z(n10272) );
  XOR U14131 ( .A(n10275), .B(n10276), .Z(n10274) );
  XOR U14132 ( .A(DB[1439]), .B(DB[1408]), .Z(n10276) );
  AND U14133 ( .A(n332), .B(n10277), .Z(n10275) );
  XOR U14134 ( .A(n10278), .B(n10279), .Z(n10277) );
  XOR U14135 ( .A(DB[1408]), .B(DB[1377]), .Z(n10279) );
  AND U14136 ( .A(n336), .B(n10280), .Z(n10278) );
  XOR U14137 ( .A(n10281), .B(n10282), .Z(n10280) );
  XOR U14138 ( .A(DB[1377]), .B(DB[1346]), .Z(n10282) );
  AND U14139 ( .A(n340), .B(n10283), .Z(n10281) );
  XOR U14140 ( .A(n10284), .B(n10285), .Z(n10283) );
  XOR U14141 ( .A(DB[1346]), .B(DB[1315]), .Z(n10285) );
  AND U14142 ( .A(n344), .B(n10286), .Z(n10284) );
  XOR U14143 ( .A(n10287), .B(n10288), .Z(n10286) );
  XOR U14144 ( .A(DB[1315]), .B(DB[1284]), .Z(n10288) );
  AND U14145 ( .A(n348), .B(n10289), .Z(n10287) );
  XOR U14146 ( .A(n10290), .B(n10291), .Z(n10289) );
  XOR U14147 ( .A(DB[1284]), .B(DB[1253]), .Z(n10291) );
  AND U14148 ( .A(n352), .B(n10292), .Z(n10290) );
  XOR U14149 ( .A(n10293), .B(n10294), .Z(n10292) );
  XOR U14150 ( .A(DB[1253]), .B(DB[1222]), .Z(n10294) );
  AND U14151 ( .A(n356), .B(n10295), .Z(n10293) );
  XOR U14152 ( .A(n10296), .B(n10297), .Z(n10295) );
  XOR U14153 ( .A(DB[1222]), .B(DB[1191]), .Z(n10297) );
  AND U14154 ( .A(n360), .B(n10298), .Z(n10296) );
  XOR U14155 ( .A(n10299), .B(n10300), .Z(n10298) );
  XOR U14156 ( .A(DB[1191]), .B(DB[1160]), .Z(n10300) );
  AND U14157 ( .A(n364), .B(n10301), .Z(n10299) );
  XOR U14158 ( .A(n10302), .B(n10303), .Z(n10301) );
  XOR U14159 ( .A(DB[1160]), .B(DB[1129]), .Z(n10303) );
  AND U14160 ( .A(n368), .B(n10304), .Z(n10302) );
  XOR U14161 ( .A(n10305), .B(n10306), .Z(n10304) );
  XOR U14162 ( .A(DB[1129]), .B(DB[1098]), .Z(n10306) );
  AND U14163 ( .A(n372), .B(n10307), .Z(n10305) );
  XOR U14164 ( .A(n10308), .B(n10309), .Z(n10307) );
  XOR U14165 ( .A(DB[1098]), .B(DB[1067]), .Z(n10309) );
  AND U14166 ( .A(n376), .B(n10310), .Z(n10308) );
  XOR U14167 ( .A(n10311), .B(n10312), .Z(n10310) );
  XOR U14168 ( .A(DB[1067]), .B(DB[1036]), .Z(n10312) );
  AND U14169 ( .A(n380), .B(n10313), .Z(n10311) );
  XOR U14170 ( .A(n10314), .B(n10315), .Z(n10313) );
  XOR U14171 ( .A(DB[1036]), .B(DB[1005]), .Z(n10315) );
  AND U14172 ( .A(n384), .B(n10316), .Z(n10314) );
  XOR U14173 ( .A(n10317), .B(n10318), .Z(n10316) );
  XOR U14174 ( .A(DB[974]), .B(DB[1005]), .Z(n10318) );
  AND U14175 ( .A(n388), .B(n10319), .Z(n10317) );
  XOR U14176 ( .A(n10320), .B(n10321), .Z(n10319) );
  XOR U14177 ( .A(DB[974]), .B(DB[943]), .Z(n10321) );
  AND U14178 ( .A(n392), .B(n10322), .Z(n10320) );
  XOR U14179 ( .A(n10323), .B(n10324), .Z(n10322) );
  XOR U14180 ( .A(DB[943]), .B(DB[912]), .Z(n10324) );
  AND U14181 ( .A(n396), .B(n10325), .Z(n10323) );
  XOR U14182 ( .A(n10326), .B(n10327), .Z(n10325) );
  XOR U14183 ( .A(DB[912]), .B(DB[881]), .Z(n10327) );
  AND U14184 ( .A(n400), .B(n10328), .Z(n10326) );
  XOR U14185 ( .A(n10329), .B(n10330), .Z(n10328) );
  XOR U14186 ( .A(DB[881]), .B(DB[850]), .Z(n10330) );
  AND U14187 ( .A(n404), .B(n10331), .Z(n10329) );
  XOR U14188 ( .A(n10332), .B(n10333), .Z(n10331) );
  XOR U14189 ( .A(DB[850]), .B(DB[819]), .Z(n10333) );
  AND U14190 ( .A(n408), .B(n10334), .Z(n10332) );
  XOR U14191 ( .A(n10335), .B(n10336), .Z(n10334) );
  XOR U14192 ( .A(DB[819]), .B(DB[788]), .Z(n10336) );
  AND U14193 ( .A(n412), .B(n10337), .Z(n10335) );
  XOR U14194 ( .A(n10338), .B(n10339), .Z(n10337) );
  XOR U14195 ( .A(DB[788]), .B(DB[757]), .Z(n10339) );
  AND U14196 ( .A(n416), .B(n10340), .Z(n10338) );
  XOR U14197 ( .A(n10341), .B(n10342), .Z(n10340) );
  XOR U14198 ( .A(DB[757]), .B(DB[726]), .Z(n10342) );
  AND U14199 ( .A(n420), .B(n10343), .Z(n10341) );
  XOR U14200 ( .A(n10344), .B(n10345), .Z(n10343) );
  XOR U14201 ( .A(DB[726]), .B(DB[695]), .Z(n10345) );
  AND U14202 ( .A(n424), .B(n10346), .Z(n10344) );
  XOR U14203 ( .A(n10347), .B(n10348), .Z(n10346) );
  XOR U14204 ( .A(DB[695]), .B(DB[664]), .Z(n10348) );
  AND U14205 ( .A(n428), .B(n10349), .Z(n10347) );
  XOR U14206 ( .A(n10350), .B(n10351), .Z(n10349) );
  XOR U14207 ( .A(DB[664]), .B(DB[633]), .Z(n10351) );
  AND U14208 ( .A(n432), .B(n10352), .Z(n10350) );
  XOR U14209 ( .A(n10353), .B(n10354), .Z(n10352) );
  XOR U14210 ( .A(DB[633]), .B(DB[602]), .Z(n10354) );
  AND U14211 ( .A(n436), .B(n10355), .Z(n10353) );
  XOR U14212 ( .A(n10356), .B(n10357), .Z(n10355) );
  XOR U14213 ( .A(DB[602]), .B(DB[571]), .Z(n10357) );
  AND U14214 ( .A(n440), .B(n10358), .Z(n10356) );
  XOR U14215 ( .A(n10359), .B(n10360), .Z(n10358) );
  XOR U14216 ( .A(DB[571]), .B(DB[540]), .Z(n10360) );
  AND U14217 ( .A(n444), .B(n10361), .Z(n10359) );
  XOR U14218 ( .A(n10362), .B(n10363), .Z(n10361) );
  XOR U14219 ( .A(DB[540]), .B(DB[509]), .Z(n10363) );
  AND U14220 ( .A(n448), .B(n10364), .Z(n10362) );
  XOR U14221 ( .A(n10365), .B(n10366), .Z(n10364) );
  XOR U14222 ( .A(DB[509]), .B(DB[478]), .Z(n10366) );
  AND U14223 ( .A(n452), .B(n10367), .Z(n10365) );
  XOR U14224 ( .A(n10368), .B(n10369), .Z(n10367) );
  XOR U14225 ( .A(DB[478]), .B(DB[447]), .Z(n10369) );
  AND U14226 ( .A(n456), .B(n10370), .Z(n10368) );
  XOR U14227 ( .A(n10371), .B(n10372), .Z(n10370) );
  XOR U14228 ( .A(DB[447]), .B(DB[416]), .Z(n10372) );
  AND U14229 ( .A(n460), .B(n10373), .Z(n10371) );
  XOR U14230 ( .A(n10374), .B(n10375), .Z(n10373) );
  XOR U14231 ( .A(DB[416]), .B(DB[385]), .Z(n10375) );
  AND U14232 ( .A(n464), .B(n10376), .Z(n10374) );
  XOR U14233 ( .A(n10377), .B(n10378), .Z(n10376) );
  XOR U14234 ( .A(DB[385]), .B(DB[354]), .Z(n10378) );
  AND U14235 ( .A(n468), .B(n10379), .Z(n10377) );
  XOR U14236 ( .A(n10380), .B(n10381), .Z(n10379) );
  XOR U14237 ( .A(DB[354]), .B(DB[323]), .Z(n10381) );
  AND U14238 ( .A(n472), .B(n10382), .Z(n10380) );
  XOR U14239 ( .A(n10383), .B(n10384), .Z(n10382) );
  XOR U14240 ( .A(DB[323]), .B(DB[292]), .Z(n10384) );
  AND U14241 ( .A(n476), .B(n10385), .Z(n10383) );
  XOR U14242 ( .A(n10386), .B(n10387), .Z(n10385) );
  XOR U14243 ( .A(DB[292]), .B(DB[261]), .Z(n10387) );
  AND U14244 ( .A(n480), .B(n10388), .Z(n10386) );
  XOR U14245 ( .A(n10389), .B(n10390), .Z(n10388) );
  XOR U14246 ( .A(DB[261]), .B(DB[230]), .Z(n10390) );
  AND U14247 ( .A(n484), .B(n10391), .Z(n10389) );
  XOR U14248 ( .A(n10392), .B(n10393), .Z(n10391) );
  XOR U14249 ( .A(DB[230]), .B(DB[199]), .Z(n10393) );
  AND U14250 ( .A(n488), .B(n10394), .Z(n10392) );
  XOR U14251 ( .A(n10395), .B(n10396), .Z(n10394) );
  XOR U14252 ( .A(DB[199]), .B(DB[168]), .Z(n10396) );
  AND U14253 ( .A(n492), .B(n10397), .Z(n10395) );
  XOR U14254 ( .A(n10398), .B(n10399), .Z(n10397) );
  XOR U14255 ( .A(DB[168]), .B(DB[137]), .Z(n10399) );
  AND U14256 ( .A(n496), .B(n10400), .Z(n10398) );
  XOR U14257 ( .A(n10401), .B(n10402), .Z(n10400) );
  XOR U14258 ( .A(DB[137]), .B(DB[106]), .Z(n10402) );
  AND U14259 ( .A(n500), .B(n10403), .Z(n10401) );
  XOR U14260 ( .A(n10404), .B(n10405), .Z(n10403) );
  XOR U14261 ( .A(DB[75]), .B(DB[106]), .Z(n10405) );
  AND U14262 ( .A(n504), .B(n10406), .Z(n10404) );
  XOR U14263 ( .A(n10407), .B(n10408), .Z(n10406) );
  XOR U14264 ( .A(DB[75]), .B(DB[44]), .Z(n10408) );
  AND U14265 ( .A(n508), .B(n10409), .Z(n10407) );
  XOR U14266 ( .A(DB[44]), .B(DB[13]), .Z(n10409) );
  XOR U14267 ( .A(DB[3949]), .B(n10410), .Z(min_val_out[12]) );
  AND U14268 ( .A(n2), .B(n10411), .Z(n10410) );
  XOR U14269 ( .A(n10412), .B(n10413), .Z(n10411) );
  XOR U14270 ( .A(n10414), .B(n10415), .Z(n10413) );
  IV U14271 ( .A(DB[3949]), .Z(n10414) );
  AND U14272 ( .A(n8), .B(n10416), .Z(n10412) );
  XOR U14273 ( .A(n10417), .B(n10418), .Z(n10416) );
  XOR U14274 ( .A(DB[3918]), .B(DB[3887]), .Z(n10418) );
  AND U14275 ( .A(n12), .B(n10419), .Z(n10417) );
  XOR U14276 ( .A(n10420), .B(n10421), .Z(n10419) );
  XOR U14277 ( .A(DB[3887]), .B(DB[3856]), .Z(n10421) );
  AND U14278 ( .A(n16), .B(n10422), .Z(n10420) );
  XOR U14279 ( .A(n10423), .B(n10424), .Z(n10422) );
  XOR U14280 ( .A(DB[3856]), .B(DB[3825]), .Z(n10424) );
  AND U14281 ( .A(n20), .B(n10425), .Z(n10423) );
  XOR U14282 ( .A(n10426), .B(n10427), .Z(n10425) );
  XOR U14283 ( .A(DB[3825]), .B(DB[3794]), .Z(n10427) );
  AND U14284 ( .A(n24), .B(n10428), .Z(n10426) );
  XOR U14285 ( .A(n10429), .B(n10430), .Z(n10428) );
  XOR U14286 ( .A(DB[3794]), .B(DB[3763]), .Z(n10430) );
  AND U14287 ( .A(n28), .B(n10431), .Z(n10429) );
  XOR U14288 ( .A(n10432), .B(n10433), .Z(n10431) );
  XOR U14289 ( .A(DB[3763]), .B(DB[3732]), .Z(n10433) );
  AND U14290 ( .A(n32), .B(n10434), .Z(n10432) );
  XOR U14291 ( .A(n10435), .B(n10436), .Z(n10434) );
  XOR U14292 ( .A(DB[3732]), .B(DB[3701]), .Z(n10436) );
  AND U14293 ( .A(n36), .B(n10437), .Z(n10435) );
  XOR U14294 ( .A(n10438), .B(n10439), .Z(n10437) );
  XOR U14295 ( .A(DB[3701]), .B(DB[3670]), .Z(n10439) );
  AND U14296 ( .A(n40), .B(n10440), .Z(n10438) );
  XOR U14297 ( .A(n10441), .B(n10442), .Z(n10440) );
  XOR U14298 ( .A(DB[3670]), .B(DB[3639]), .Z(n10442) );
  AND U14299 ( .A(n44), .B(n10443), .Z(n10441) );
  XOR U14300 ( .A(n10444), .B(n10445), .Z(n10443) );
  XOR U14301 ( .A(DB[3639]), .B(DB[3608]), .Z(n10445) );
  AND U14302 ( .A(n48), .B(n10446), .Z(n10444) );
  XOR U14303 ( .A(n10447), .B(n10448), .Z(n10446) );
  XOR U14304 ( .A(DB[3608]), .B(DB[3577]), .Z(n10448) );
  AND U14305 ( .A(n52), .B(n10449), .Z(n10447) );
  XOR U14306 ( .A(n10450), .B(n10451), .Z(n10449) );
  XOR U14307 ( .A(DB[3577]), .B(DB[3546]), .Z(n10451) );
  AND U14308 ( .A(n56), .B(n10452), .Z(n10450) );
  XOR U14309 ( .A(n10453), .B(n10454), .Z(n10452) );
  XOR U14310 ( .A(DB[3546]), .B(DB[3515]), .Z(n10454) );
  AND U14311 ( .A(n60), .B(n10455), .Z(n10453) );
  XOR U14312 ( .A(n10456), .B(n10457), .Z(n10455) );
  XOR U14313 ( .A(DB[3515]), .B(DB[3484]), .Z(n10457) );
  AND U14314 ( .A(n64), .B(n10458), .Z(n10456) );
  XOR U14315 ( .A(n10459), .B(n10460), .Z(n10458) );
  XOR U14316 ( .A(DB[3484]), .B(DB[3453]), .Z(n10460) );
  AND U14317 ( .A(n68), .B(n10461), .Z(n10459) );
  XOR U14318 ( .A(n10462), .B(n10463), .Z(n10461) );
  XOR U14319 ( .A(DB[3453]), .B(DB[3422]), .Z(n10463) );
  AND U14320 ( .A(n72), .B(n10464), .Z(n10462) );
  XOR U14321 ( .A(n10465), .B(n10466), .Z(n10464) );
  XOR U14322 ( .A(DB[3422]), .B(DB[3391]), .Z(n10466) );
  AND U14323 ( .A(n76), .B(n10467), .Z(n10465) );
  XOR U14324 ( .A(n10468), .B(n10469), .Z(n10467) );
  XOR U14325 ( .A(DB[3391]), .B(DB[3360]), .Z(n10469) );
  AND U14326 ( .A(n80), .B(n10470), .Z(n10468) );
  XOR U14327 ( .A(n10471), .B(n10472), .Z(n10470) );
  XOR U14328 ( .A(DB[3360]), .B(DB[3329]), .Z(n10472) );
  AND U14329 ( .A(n84), .B(n10473), .Z(n10471) );
  XOR U14330 ( .A(n10474), .B(n10475), .Z(n10473) );
  XOR U14331 ( .A(DB[3329]), .B(DB[3298]), .Z(n10475) );
  AND U14332 ( .A(n88), .B(n10476), .Z(n10474) );
  XOR U14333 ( .A(n10477), .B(n10478), .Z(n10476) );
  XOR U14334 ( .A(DB[3298]), .B(DB[3267]), .Z(n10478) );
  AND U14335 ( .A(n92), .B(n10479), .Z(n10477) );
  XOR U14336 ( .A(n10480), .B(n10481), .Z(n10479) );
  XOR U14337 ( .A(DB[3267]), .B(DB[3236]), .Z(n10481) );
  AND U14338 ( .A(n96), .B(n10482), .Z(n10480) );
  XOR U14339 ( .A(n10483), .B(n10484), .Z(n10482) );
  XOR U14340 ( .A(DB[3236]), .B(DB[3205]), .Z(n10484) );
  AND U14341 ( .A(n100), .B(n10485), .Z(n10483) );
  XOR U14342 ( .A(n10486), .B(n10487), .Z(n10485) );
  XOR U14343 ( .A(DB[3205]), .B(DB[3174]), .Z(n10487) );
  AND U14344 ( .A(n104), .B(n10488), .Z(n10486) );
  XOR U14345 ( .A(n10489), .B(n10490), .Z(n10488) );
  XOR U14346 ( .A(DB[3174]), .B(DB[3143]), .Z(n10490) );
  AND U14347 ( .A(n108), .B(n10491), .Z(n10489) );
  XOR U14348 ( .A(n10492), .B(n10493), .Z(n10491) );
  XOR U14349 ( .A(DB[3143]), .B(DB[3112]), .Z(n10493) );
  AND U14350 ( .A(n112), .B(n10494), .Z(n10492) );
  XOR U14351 ( .A(n10495), .B(n10496), .Z(n10494) );
  XOR U14352 ( .A(DB[3112]), .B(DB[3081]), .Z(n10496) );
  AND U14353 ( .A(n116), .B(n10497), .Z(n10495) );
  XOR U14354 ( .A(n10498), .B(n10499), .Z(n10497) );
  XOR U14355 ( .A(DB[3081]), .B(DB[3050]), .Z(n10499) );
  AND U14356 ( .A(n120), .B(n10500), .Z(n10498) );
  XOR U14357 ( .A(n10501), .B(n10502), .Z(n10500) );
  XOR U14358 ( .A(DB[3050]), .B(DB[3019]), .Z(n10502) );
  AND U14359 ( .A(n124), .B(n10503), .Z(n10501) );
  XOR U14360 ( .A(n10504), .B(n10505), .Z(n10503) );
  XOR U14361 ( .A(DB[3019]), .B(DB[2988]), .Z(n10505) );
  AND U14362 ( .A(n128), .B(n10506), .Z(n10504) );
  XOR U14363 ( .A(n10507), .B(n10508), .Z(n10506) );
  XOR U14364 ( .A(DB[2988]), .B(DB[2957]), .Z(n10508) );
  AND U14365 ( .A(n132), .B(n10509), .Z(n10507) );
  XOR U14366 ( .A(n10510), .B(n10511), .Z(n10509) );
  XOR U14367 ( .A(DB[2957]), .B(DB[2926]), .Z(n10511) );
  AND U14368 ( .A(n136), .B(n10512), .Z(n10510) );
  XOR U14369 ( .A(n10513), .B(n10514), .Z(n10512) );
  XOR U14370 ( .A(DB[2926]), .B(DB[2895]), .Z(n10514) );
  AND U14371 ( .A(n140), .B(n10515), .Z(n10513) );
  XOR U14372 ( .A(n10516), .B(n10517), .Z(n10515) );
  XOR U14373 ( .A(DB[2895]), .B(DB[2864]), .Z(n10517) );
  AND U14374 ( .A(n144), .B(n10518), .Z(n10516) );
  XOR U14375 ( .A(n10519), .B(n10520), .Z(n10518) );
  XOR U14376 ( .A(DB[2864]), .B(DB[2833]), .Z(n10520) );
  AND U14377 ( .A(n148), .B(n10521), .Z(n10519) );
  XOR U14378 ( .A(n10522), .B(n10523), .Z(n10521) );
  XOR U14379 ( .A(DB[2833]), .B(DB[2802]), .Z(n10523) );
  AND U14380 ( .A(n152), .B(n10524), .Z(n10522) );
  XOR U14381 ( .A(n10525), .B(n10526), .Z(n10524) );
  XOR U14382 ( .A(DB[2802]), .B(DB[2771]), .Z(n10526) );
  AND U14383 ( .A(n156), .B(n10527), .Z(n10525) );
  XOR U14384 ( .A(n10528), .B(n10529), .Z(n10527) );
  XOR U14385 ( .A(DB[2771]), .B(DB[2740]), .Z(n10529) );
  AND U14386 ( .A(n160), .B(n10530), .Z(n10528) );
  XOR U14387 ( .A(n10531), .B(n10532), .Z(n10530) );
  XOR U14388 ( .A(DB[2740]), .B(DB[2709]), .Z(n10532) );
  AND U14389 ( .A(n164), .B(n10533), .Z(n10531) );
  XOR U14390 ( .A(n10534), .B(n10535), .Z(n10533) );
  XOR U14391 ( .A(DB[2709]), .B(DB[2678]), .Z(n10535) );
  AND U14392 ( .A(n168), .B(n10536), .Z(n10534) );
  XOR U14393 ( .A(n10537), .B(n10538), .Z(n10536) );
  XOR U14394 ( .A(DB[2678]), .B(DB[2647]), .Z(n10538) );
  AND U14395 ( .A(n172), .B(n10539), .Z(n10537) );
  XOR U14396 ( .A(n10540), .B(n10541), .Z(n10539) );
  XOR U14397 ( .A(DB[2647]), .B(DB[2616]), .Z(n10541) );
  AND U14398 ( .A(n176), .B(n10542), .Z(n10540) );
  XOR U14399 ( .A(n10543), .B(n10544), .Z(n10542) );
  XOR U14400 ( .A(DB[2616]), .B(DB[2585]), .Z(n10544) );
  AND U14401 ( .A(n180), .B(n10545), .Z(n10543) );
  XOR U14402 ( .A(n10546), .B(n10547), .Z(n10545) );
  XOR U14403 ( .A(DB[2585]), .B(DB[2554]), .Z(n10547) );
  AND U14404 ( .A(n184), .B(n10548), .Z(n10546) );
  XOR U14405 ( .A(n10549), .B(n10550), .Z(n10548) );
  XOR U14406 ( .A(DB[2554]), .B(DB[2523]), .Z(n10550) );
  AND U14407 ( .A(n188), .B(n10551), .Z(n10549) );
  XOR U14408 ( .A(n10552), .B(n10553), .Z(n10551) );
  XOR U14409 ( .A(DB[2523]), .B(DB[2492]), .Z(n10553) );
  AND U14410 ( .A(n192), .B(n10554), .Z(n10552) );
  XOR U14411 ( .A(n10555), .B(n10556), .Z(n10554) );
  XOR U14412 ( .A(DB[2492]), .B(DB[2461]), .Z(n10556) );
  AND U14413 ( .A(n196), .B(n10557), .Z(n10555) );
  XOR U14414 ( .A(n10558), .B(n10559), .Z(n10557) );
  XOR U14415 ( .A(DB[2461]), .B(DB[2430]), .Z(n10559) );
  AND U14416 ( .A(n200), .B(n10560), .Z(n10558) );
  XOR U14417 ( .A(n10561), .B(n10562), .Z(n10560) );
  XOR U14418 ( .A(DB[2430]), .B(DB[2399]), .Z(n10562) );
  AND U14419 ( .A(n204), .B(n10563), .Z(n10561) );
  XOR U14420 ( .A(n10564), .B(n10565), .Z(n10563) );
  XOR U14421 ( .A(DB[2399]), .B(DB[2368]), .Z(n10565) );
  AND U14422 ( .A(n208), .B(n10566), .Z(n10564) );
  XOR U14423 ( .A(n10567), .B(n10568), .Z(n10566) );
  XOR U14424 ( .A(DB[2368]), .B(DB[2337]), .Z(n10568) );
  AND U14425 ( .A(n212), .B(n10569), .Z(n10567) );
  XOR U14426 ( .A(n10570), .B(n10571), .Z(n10569) );
  XOR U14427 ( .A(DB[2337]), .B(DB[2306]), .Z(n10571) );
  AND U14428 ( .A(n216), .B(n10572), .Z(n10570) );
  XOR U14429 ( .A(n10573), .B(n10574), .Z(n10572) );
  XOR U14430 ( .A(DB[2306]), .B(DB[2275]), .Z(n10574) );
  AND U14431 ( .A(n220), .B(n10575), .Z(n10573) );
  XOR U14432 ( .A(n10576), .B(n10577), .Z(n10575) );
  XOR U14433 ( .A(DB[2275]), .B(DB[2244]), .Z(n10577) );
  AND U14434 ( .A(n224), .B(n10578), .Z(n10576) );
  XOR U14435 ( .A(n10579), .B(n10580), .Z(n10578) );
  XOR U14436 ( .A(DB[2244]), .B(DB[2213]), .Z(n10580) );
  AND U14437 ( .A(n228), .B(n10581), .Z(n10579) );
  XOR U14438 ( .A(n10582), .B(n10583), .Z(n10581) );
  XOR U14439 ( .A(DB[2213]), .B(DB[2182]), .Z(n10583) );
  AND U14440 ( .A(n232), .B(n10584), .Z(n10582) );
  XOR U14441 ( .A(n10585), .B(n10586), .Z(n10584) );
  XOR U14442 ( .A(DB[2182]), .B(DB[2151]), .Z(n10586) );
  AND U14443 ( .A(n236), .B(n10587), .Z(n10585) );
  XOR U14444 ( .A(n10588), .B(n10589), .Z(n10587) );
  XOR U14445 ( .A(DB[2151]), .B(DB[2120]), .Z(n10589) );
  AND U14446 ( .A(n240), .B(n10590), .Z(n10588) );
  XOR U14447 ( .A(n10591), .B(n10592), .Z(n10590) );
  XOR U14448 ( .A(DB[2120]), .B(DB[2089]), .Z(n10592) );
  AND U14449 ( .A(n244), .B(n10593), .Z(n10591) );
  XOR U14450 ( .A(n10594), .B(n10595), .Z(n10593) );
  XOR U14451 ( .A(DB[2089]), .B(DB[2058]), .Z(n10595) );
  AND U14452 ( .A(n248), .B(n10596), .Z(n10594) );
  XOR U14453 ( .A(n10597), .B(n10598), .Z(n10596) );
  XOR U14454 ( .A(DB[2058]), .B(DB[2027]), .Z(n10598) );
  AND U14455 ( .A(n252), .B(n10599), .Z(n10597) );
  XOR U14456 ( .A(n10600), .B(n10601), .Z(n10599) );
  XOR U14457 ( .A(DB[2027]), .B(DB[1996]), .Z(n10601) );
  AND U14458 ( .A(n256), .B(n10602), .Z(n10600) );
  XOR U14459 ( .A(n10603), .B(n10604), .Z(n10602) );
  XOR U14460 ( .A(DB[1996]), .B(DB[1965]), .Z(n10604) );
  AND U14461 ( .A(n260), .B(n10605), .Z(n10603) );
  XOR U14462 ( .A(n10606), .B(n10607), .Z(n10605) );
  XOR U14463 ( .A(DB[1965]), .B(DB[1934]), .Z(n10607) );
  AND U14464 ( .A(n264), .B(n10608), .Z(n10606) );
  XOR U14465 ( .A(n10609), .B(n10610), .Z(n10608) );
  XOR U14466 ( .A(DB[1934]), .B(DB[1903]), .Z(n10610) );
  AND U14467 ( .A(n268), .B(n10611), .Z(n10609) );
  XOR U14468 ( .A(n10612), .B(n10613), .Z(n10611) );
  XOR U14469 ( .A(DB[1903]), .B(DB[1872]), .Z(n10613) );
  AND U14470 ( .A(n272), .B(n10614), .Z(n10612) );
  XOR U14471 ( .A(n10615), .B(n10616), .Z(n10614) );
  XOR U14472 ( .A(DB[1872]), .B(DB[1841]), .Z(n10616) );
  AND U14473 ( .A(n276), .B(n10617), .Z(n10615) );
  XOR U14474 ( .A(n10618), .B(n10619), .Z(n10617) );
  XOR U14475 ( .A(DB[1841]), .B(DB[1810]), .Z(n10619) );
  AND U14476 ( .A(n280), .B(n10620), .Z(n10618) );
  XOR U14477 ( .A(n10621), .B(n10622), .Z(n10620) );
  XOR U14478 ( .A(DB[1810]), .B(DB[1779]), .Z(n10622) );
  AND U14479 ( .A(n284), .B(n10623), .Z(n10621) );
  XOR U14480 ( .A(n10624), .B(n10625), .Z(n10623) );
  XOR U14481 ( .A(DB[1779]), .B(DB[1748]), .Z(n10625) );
  AND U14482 ( .A(n288), .B(n10626), .Z(n10624) );
  XOR U14483 ( .A(n10627), .B(n10628), .Z(n10626) );
  XOR U14484 ( .A(DB[1748]), .B(DB[1717]), .Z(n10628) );
  AND U14485 ( .A(n292), .B(n10629), .Z(n10627) );
  XOR U14486 ( .A(n10630), .B(n10631), .Z(n10629) );
  XOR U14487 ( .A(DB[1717]), .B(DB[1686]), .Z(n10631) );
  AND U14488 ( .A(n296), .B(n10632), .Z(n10630) );
  XOR U14489 ( .A(n10633), .B(n10634), .Z(n10632) );
  XOR U14490 ( .A(DB[1686]), .B(DB[1655]), .Z(n10634) );
  AND U14491 ( .A(n300), .B(n10635), .Z(n10633) );
  XOR U14492 ( .A(n10636), .B(n10637), .Z(n10635) );
  XOR U14493 ( .A(DB[1655]), .B(DB[1624]), .Z(n10637) );
  AND U14494 ( .A(n304), .B(n10638), .Z(n10636) );
  XOR U14495 ( .A(n10639), .B(n10640), .Z(n10638) );
  XOR U14496 ( .A(DB[1624]), .B(DB[1593]), .Z(n10640) );
  AND U14497 ( .A(n308), .B(n10641), .Z(n10639) );
  XOR U14498 ( .A(n10642), .B(n10643), .Z(n10641) );
  XOR U14499 ( .A(DB[1593]), .B(DB[1562]), .Z(n10643) );
  AND U14500 ( .A(n312), .B(n10644), .Z(n10642) );
  XOR U14501 ( .A(n10645), .B(n10646), .Z(n10644) );
  XOR U14502 ( .A(DB[1562]), .B(DB[1531]), .Z(n10646) );
  AND U14503 ( .A(n316), .B(n10647), .Z(n10645) );
  XOR U14504 ( .A(n10648), .B(n10649), .Z(n10647) );
  XOR U14505 ( .A(DB[1531]), .B(DB[1500]), .Z(n10649) );
  AND U14506 ( .A(n320), .B(n10650), .Z(n10648) );
  XOR U14507 ( .A(n10651), .B(n10652), .Z(n10650) );
  XOR U14508 ( .A(DB[1500]), .B(DB[1469]), .Z(n10652) );
  AND U14509 ( .A(n324), .B(n10653), .Z(n10651) );
  XOR U14510 ( .A(n10654), .B(n10655), .Z(n10653) );
  XOR U14511 ( .A(DB[1469]), .B(DB[1438]), .Z(n10655) );
  AND U14512 ( .A(n328), .B(n10656), .Z(n10654) );
  XOR U14513 ( .A(n10657), .B(n10658), .Z(n10656) );
  XOR U14514 ( .A(DB[1438]), .B(DB[1407]), .Z(n10658) );
  AND U14515 ( .A(n332), .B(n10659), .Z(n10657) );
  XOR U14516 ( .A(n10660), .B(n10661), .Z(n10659) );
  XOR U14517 ( .A(DB[1407]), .B(DB[1376]), .Z(n10661) );
  AND U14518 ( .A(n336), .B(n10662), .Z(n10660) );
  XOR U14519 ( .A(n10663), .B(n10664), .Z(n10662) );
  XOR U14520 ( .A(DB[1376]), .B(DB[1345]), .Z(n10664) );
  AND U14521 ( .A(n340), .B(n10665), .Z(n10663) );
  XOR U14522 ( .A(n10666), .B(n10667), .Z(n10665) );
  XOR U14523 ( .A(DB[1345]), .B(DB[1314]), .Z(n10667) );
  AND U14524 ( .A(n344), .B(n10668), .Z(n10666) );
  XOR U14525 ( .A(n10669), .B(n10670), .Z(n10668) );
  XOR U14526 ( .A(DB[1314]), .B(DB[1283]), .Z(n10670) );
  AND U14527 ( .A(n348), .B(n10671), .Z(n10669) );
  XOR U14528 ( .A(n10672), .B(n10673), .Z(n10671) );
  XOR U14529 ( .A(DB[1283]), .B(DB[1252]), .Z(n10673) );
  AND U14530 ( .A(n352), .B(n10674), .Z(n10672) );
  XOR U14531 ( .A(n10675), .B(n10676), .Z(n10674) );
  XOR U14532 ( .A(DB[1252]), .B(DB[1221]), .Z(n10676) );
  AND U14533 ( .A(n356), .B(n10677), .Z(n10675) );
  XOR U14534 ( .A(n10678), .B(n10679), .Z(n10677) );
  XOR U14535 ( .A(DB[1221]), .B(DB[1190]), .Z(n10679) );
  AND U14536 ( .A(n360), .B(n10680), .Z(n10678) );
  XOR U14537 ( .A(n10681), .B(n10682), .Z(n10680) );
  XOR U14538 ( .A(DB[1190]), .B(DB[1159]), .Z(n10682) );
  AND U14539 ( .A(n364), .B(n10683), .Z(n10681) );
  XOR U14540 ( .A(n10684), .B(n10685), .Z(n10683) );
  XOR U14541 ( .A(DB[1159]), .B(DB[1128]), .Z(n10685) );
  AND U14542 ( .A(n368), .B(n10686), .Z(n10684) );
  XOR U14543 ( .A(n10687), .B(n10688), .Z(n10686) );
  XOR U14544 ( .A(DB[1128]), .B(DB[1097]), .Z(n10688) );
  AND U14545 ( .A(n372), .B(n10689), .Z(n10687) );
  XOR U14546 ( .A(n10690), .B(n10691), .Z(n10689) );
  XOR U14547 ( .A(DB[1097]), .B(DB[1066]), .Z(n10691) );
  AND U14548 ( .A(n376), .B(n10692), .Z(n10690) );
  XOR U14549 ( .A(n10693), .B(n10694), .Z(n10692) );
  XOR U14550 ( .A(DB[1066]), .B(DB[1035]), .Z(n10694) );
  AND U14551 ( .A(n380), .B(n10695), .Z(n10693) );
  XOR U14552 ( .A(n10696), .B(n10697), .Z(n10695) );
  XOR U14553 ( .A(DB[1035]), .B(DB[1004]), .Z(n10697) );
  AND U14554 ( .A(n384), .B(n10698), .Z(n10696) );
  XOR U14555 ( .A(n10699), .B(n10700), .Z(n10698) );
  XOR U14556 ( .A(DB[973]), .B(DB[1004]), .Z(n10700) );
  AND U14557 ( .A(n388), .B(n10701), .Z(n10699) );
  XOR U14558 ( .A(n10702), .B(n10703), .Z(n10701) );
  XOR U14559 ( .A(DB[973]), .B(DB[942]), .Z(n10703) );
  AND U14560 ( .A(n392), .B(n10704), .Z(n10702) );
  XOR U14561 ( .A(n10705), .B(n10706), .Z(n10704) );
  XOR U14562 ( .A(DB[942]), .B(DB[911]), .Z(n10706) );
  AND U14563 ( .A(n396), .B(n10707), .Z(n10705) );
  XOR U14564 ( .A(n10708), .B(n10709), .Z(n10707) );
  XOR U14565 ( .A(DB[911]), .B(DB[880]), .Z(n10709) );
  AND U14566 ( .A(n400), .B(n10710), .Z(n10708) );
  XOR U14567 ( .A(n10711), .B(n10712), .Z(n10710) );
  XOR U14568 ( .A(DB[880]), .B(DB[849]), .Z(n10712) );
  AND U14569 ( .A(n404), .B(n10713), .Z(n10711) );
  XOR U14570 ( .A(n10714), .B(n10715), .Z(n10713) );
  XOR U14571 ( .A(DB[849]), .B(DB[818]), .Z(n10715) );
  AND U14572 ( .A(n408), .B(n10716), .Z(n10714) );
  XOR U14573 ( .A(n10717), .B(n10718), .Z(n10716) );
  XOR U14574 ( .A(DB[818]), .B(DB[787]), .Z(n10718) );
  AND U14575 ( .A(n412), .B(n10719), .Z(n10717) );
  XOR U14576 ( .A(n10720), .B(n10721), .Z(n10719) );
  XOR U14577 ( .A(DB[787]), .B(DB[756]), .Z(n10721) );
  AND U14578 ( .A(n416), .B(n10722), .Z(n10720) );
  XOR U14579 ( .A(n10723), .B(n10724), .Z(n10722) );
  XOR U14580 ( .A(DB[756]), .B(DB[725]), .Z(n10724) );
  AND U14581 ( .A(n420), .B(n10725), .Z(n10723) );
  XOR U14582 ( .A(n10726), .B(n10727), .Z(n10725) );
  XOR U14583 ( .A(DB[725]), .B(DB[694]), .Z(n10727) );
  AND U14584 ( .A(n424), .B(n10728), .Z(n10726) );
  XOR U14585 ( .A(n10729), .B(n10730), .Z(n10728) );
  XOR U14586 ( .A(DB[694]), .B(DB[663]), .Z(n10730) );
  AND U14587 ( .A(n428), .B(n10731), .Z(n10729) );
  XOR U14588 ( .A(n10732), .B(n10733), .Z(n10731) );
  XOR U14589 ( .A(DB[663]), .B(DB[632]), .Z(n10733) );
  AND U14590 ( .A(n432), .B(n10734), .Z(n10732) );
  XOR U14591 ( .A(n10735), .B(n10736), .Z(n10734) );
  XOR U14592 ( .A(DB[632]), .B(DB[601]), .Z(n10736) );
  AND U14593 ( .A(n436), .B(n10737), .Z(n10735) );
  XOR U14594 ( .A(n10738), .B(n10739), .Z(n10737) );
  XOR U14595 ( .A(DB[601]), .B(DB[570]), .Z(n10739) );
  AND U14596 ( .A(n440), .B(n10740), .Z(n10738) );
  XOR U14597 ( .A(n10741), .B(n10742), .Z(n10740) );
  XOR U14598 ( .A(DB[570]), .B(DB[539]), .Z(n10742) );
  AND U14599 ( .A(n444), .B(n10743), .Z(n10741) );
  XOR U14600 ( .A(n10744), .B(n10745), .Z(n10743) );
  XOR U14601 ( .A(DB[539]), .B(DB[508]), .Z(n10745) );
  AND U14602 ( .A(n448), .B(n10746), .Z(n10744) );
  XOR U14603 ( .A(n10747), .B(n10748), .Z(n10746) );
  XOR U14604 ( .A(DB[508]), .B(DB[477]), .Z(n10748) );
  AND U14605 ( .A(n452), .B(n10749), .Z(n10747) );
  XOR U14606 ( .A(n10750), .B(n10751), .Z(n10749) );
  XOR U14607 ( .A(DB[477]), .B(DB[446]), .Z(n10751) );
  AND U14608 ( .A(n456), .B(n10752), .Z(n10750) );
  XOR U14609 ( .A(n10753), .B(n10754), .Z(n10752) );
  XOR U14610 ( .A(DB[446]), .B(DB[415]), .Z(n10754) );
  AND U14611 ( .A(n460), .B(n10755), .Z(n10753) );
  XOR U14612 ( .A(n10756), .B(n10757), .Z(n10755) );
  XOR U14613 ( .A(DB[415]), .B(DB[384]), .Z(n10757) );
  AND U14614 ( .A(n464), .B(n10758), .Z(n10756) );
  XOR U14615 ( .A(n10759), .B(n10760), .Z(n10758) );
  XOR U14616 ( .A(DB[384]), .B(DB[353]), .Z(n10760) );
  AND U14617 ( .A(n468), .B(n10761), .Z(n10759) );
  XOR U14618 ( .A(n10762), .B(n10763), .Z(n10761) );
  XOR U14619 ( .A(DB[353]), .B(DB[322]), .Z(n10763) );
  AND U14620 ( .A(n472), .B(n10764), .Z(n10762) );
  XOR U14621 ( .A(n10765), .B(n10766), .Z(n10764) );
  XOR U14622 ( .A(DB[322]), .B(DB[291]), .Z(n10766) );
  AND U14623 ( .A(n476), .B(n10767), .Z(n10765) );
  XOR U14624 ( .A(n10768), .B(n10769), .Z(n10767) );
  XOR U14625 ( .A(DB[291]), .B(DB[260]), .Z(n10769) );
  AND U14626 ( .A(n480), .B(n10770), .Z(n10768) );
  XOR U14627 ( .A(n10771), .B(n10772), .Z(n10770) );
  XOR U14628 ( .A(DB[260]), .B(DB[229]), .Z(n10772) );
  AND U14629 ( .A(n484), .B(n10773), .Z(n10771) );
  XOR U14630 ( .A(n10774), .B(n10775), .Z(n10773) );
  XOR U14631 ( .A(DB[229]), .B(DB[198]), .Z(n10775) );
  AND U14632 ( .A(n488), .B(n10776), .Z(n10774) );
  XOR U14633 ( .A(n10777), .B(n10778), .Z(n10776) );
  XOR U14634 ( .A(DB[198]), .B(DB[167]), .Z(n10778) );
  AND U14635 ( .A(n492), .B(n10779), .Z(n10777) );
  XOR U14636 ( .A(n10780), .B(n10781), .Z(n10779) );
  XOR U14637 ( .A(DB[167]), .B(DB[136]), .Z(n10781) );
  AND U14638 ( .A(n496), .B(n10782), .Z(n10780) );
  XOR U14639 ( .A(n10783), .B(n10784), .Z(n10782) );
  XOR U14640 ( .A(DB[136]), .B(DB[105]), .Z(n10784) );
  AND U14641 ( .A(n500), .B(n10785), .Z(n10783) );
  XOR U14642 ( .A(n10786), .B(n10787), .Z(n10785) );
  XOR U14643 ( .A(DB[74]), .B(DB[105]), .Z(n10787) );
  AND U14644 ( .A(n504), .B(n10788), .Z(n10786) );
  XOR U14645 ( .A(n10789), .B(n10790), .Z(n10788) );
  XOR U14646 ( .A(DB[74]), .B(DB[43]), .Z(n10790) );
  AND U14647 ( .A(n508), .B(n10791), .Z(n10789) );
  XOR U14648 ( .A(DB[43]), .B(DB[12]), .Z(n10791) );
  XOR U14649 ( .A(DB[3948]), .B(n10792), .Z(min_val_out[11]) );
  AND U14650 ( .A(n2), .B(n10793), .Z(n10792) );
  XOR U14651 ( .A(n10794), .B(n10795), .Z(n10793) );
  XOR U14652 ( .A(DB[3948]), .B(DB[3917]), .Z(n10795) );
  AND U14653 ( .A(n8), .B(n10796), .Z(n10794) );
  XOR U14654 ( .A(n10797), .B(n10798), .Z(n10796) );
  XOR U14655 ( .A(DB[3917]), .B(DB[3886]), .Z(n10798) );
  AND U14656 ( .A(n12), .B(n10799), .Z(n10797) );
  XOR U14657 ( .A(n10800), .B(n10801), .Z(n10799) );
  XOR U14658 ( .A(DB[3886]), .B(DB[3855]), .Z(n10801) );
  AND U14659 ( .A(n16), .B(n10802), .Z(n10800) );
  XOR U14660 ( .A(n10803), .B(n10804), .Z(n10802) );
  XOR U14661 ( .A(DB[3855]), .B(DB[3824]), .Z(n10804) );
  AND U14662 ( .A(n20), .B(n10805), .Z(n10803) );
  XOR U14663 ( .A(n10806), .B(n10807), .Z(n10805) );
  XOR U14664 ( .A(DB[3824]), .B(DB[3793]), .Z(n10807) );
  AND U14665 ( .A(n24), .B(n10808), .Z(n10806) );
  XOR U14666 ( .A(n10809), .B(n10810), .Z(n10808) );
  XOR U14667 ( .A(DB[3793]), .B(DB[3762]), .Z(n10810) );
  AND U14668 ( .A(n28), .B(n10811), .Z(n10809) );
  XOR U14669 ( .A(n10812), .B(n10813), .Z(n10811) );
  XOR U14670 ( .A(DB[3762]), .B(DB[3731]), .Z(n10813) );
  AND U14671 ( .A(n32), .B(n10814), .Z(n10812) );
  XOR U14672 ( .A(n10815), .B(n10816), .Z(n10814) );
  XOR U14673 ( .A(DB[3731]), .B(DB[3700]), .Z(n10816) );
  AND U14674 ( .A(n36), .B(n10817), .Z(n10815) );
  XOR U14675 ( .A(n10818), .B(n10819), .Z(n10817) );
  XOR U14676 ( .A(DB[3700]), .B(DB[3669]), .Z(n10819) );
  AND U14677 ( .A(n40), .B(n10820), .Z(n10818) );
  XOR U14678 ( .A(n10821), .B(n10822), .Z(n10820) );
  XOR U14679 ( .A(DB[3669]), .B(DB[3638]), .Z(n10822) );
  AND U14680 ( .A(n44), .B(n10823), .Z(n10821) );
  XOR U14681 ( .A(n10824), .B(n10825), .Z(n10823) );
  XOR U14682 ( .A(DB[3638]), .B(DB[3607]), .Z(n10825) );
  AND U14683 ( .A(n48), .B(n10826), .Z(n10824) );
  XOR U14684 ( .A(n10827), .B(n10828), .Z(n10826) );
  XOR U14685 ( .A(DB[3607]), .B(DB[3576]), .Z(n10828) );
  AND U14686 ( .A(n52), .B(n10829), .Z(n10827) );
  XOR U14687 ( .A(n10830), .B(n10831), .Z(n10829) );
  XOR U14688 ( .A(DB[3576]), .B(DB[3545]), .Z(n10831) );
  AND U14689 ( .A(n56), .B(n10832), .Z(n10830) );
  XOR U14690 ( .A(n10833), .B(n10834), .Z(n10832) );
  XOR U14691 ( .A(DB[3545]), .B(DB[3514]), .Z(n10834) );
  AND U14692 ( .A(n60), .B(n10835), .Z(n10833) );
  XOR U14693 ( .A(n10836), .B(n10837), .Z(n10835) );
  XOR U14694 ( .A(DB[3514]), .B(DB[3483]), .Z(n10837) );
  AND U14695 ( .A(n64), .B(n10838), .Z(n10836) );
  XOR U14696 ( .A(n10839), .B(n10840), .Z(n10838) );
  XOR U14697 ( .A(DB[3483]), .B(DB[3452]), .Z(n10840) );
  AND U14698 ( .A(n68), .B(n10841), .Z(n10839) );
  XOR U14699 ( .A(n10842), .B(n10843), .Z(n10841) );
  XOR U14700 ( .A(DB[3452]), .B(DB[3421]), .Z(n10843) );
  AND U14701 ( .A(n72), .B(n10844), .Z(n10842) );
  XOR U14702 ( .A(n10845), .B(n10846), .Z(n10844) );
  XOR U14703 ( .A(DB[3421]), .B(DB[3390]), .Z(n10846) );
  AND U14704 ( .A(n76), .B(n10847), .Z(n10845) );
  XOR U14705 ( .A(n10848), .B(n10849), .Z(n10847) );
  XOR U14706 ( .A(DB[3390]), .B(DB[3359]), .Z(n10849) );
  AND U14707 ( .A(n80), .B(n10850), .Z(n10848) );
  XOR U14708 ( .A(n10851), .B(n10852), .Z(n10850) );
  XOR U14709 ( .A(DB[3359]), .B(DB[3328]), .Z(n10852) );
  AND U14710 ( .A(n84), .B(n10853), .Z(n10851) );
  XOR U14711 ( .A(n10854), .B(n10855), .Z(n10853) );
  XOR U14712 ( .A(DB[3328]), .B(DB[3297]), .Z(n10855) );
  AND U14713 ( .A(n88), .B(n10856), .Z(n10854) );
  XOR U14714 ( .A(n10857), .B(n10858), .Z(n10856) );
  XOR U14715 ( .A(DB[3297]), .B(DB[3266]), .Z(n10858) );
  AND U14716 ( .A(n92), .B(n10859), .Z(n10857) );
  XOR U14717 ( .A(n10860), .B(n10861), .Z(n10859) );
  XOR U14718 ( .A(DB[3266]), .B(DB[3235]), .Z(n10861) );
  AND U14719 ( .A(n96), .B(n10862), .Z(n10860) );
  XOR U14720 ( .A(n10863), .B(n10864), .Z(n10862) );
  XOR U14721 ( .A(DB[3235]), .B(DB[3204]), .Z(n10864) );
  AND U14722 ( .A(n100), .B(n10865), .Z(n10863) );
  XOR U14723 ( .A(n10866), .B(n10867), .Z(n10865) );
  XOR U14724 ( .A(DB[3204]), .B(DB[3173]), .Z(n10867) );
  AND U14725 ( .A(n104), .B(n10868), .Z(n10866) );
  XOR U14726 ( .A(n10869), .B(n10870), .Z(n10868) );
  XOR U14727 ( .A(DB[3173]), .B(DB[3142]), .Z(n10870) );
  AND U14728 ( .A(n108), .B(n10871), .Z(n10869) );
  XOR U14729 ( .A(n10872), .B(n10873), .Z(n10871) );
  XOR U14730 ( .A(DB[3142]), .B(DB[3111]), .Z(n10873) );
  AND U14731 ( .A(n112), .B(n10874), .Z(n10872) );
  XOR U14732 ( .A(n10875), .B(n10876), .Z(n10874) );
  XOR U14733 ( .A(DB[3111]), .B(DB[3080]), .Z(n10876) );
  AND U14734 ( .A(n116), .B(n10877), .Z(n10875) );
  XOR U14735 ( .A(n10878), .B(n10879), .Z(n10877) );
  XOR U14736 ( .A(DB[3080]), .B(DB[3049]), .Z(n10879) );
  AND U14737 ( .A(n120), .B(n10880), .Z(n10878) );
  XOR U14738 ( .A(n10881), .B(n10882), .Z(n10880) );
  XOR U14739 ( .A(DB[3049]), .B(DB[3018]), .Z(n10882) );
  AND U14740 ( .A(n124), .B(n10883), .Z(n10881) );
  XOR U14741 ( .A(n10884), .B(n10885), .Z(n10883) );
  XOR U14742 ( .A(DB[3018]), .B(DB[2987]), .Z(n10885) );
  AND U14743 ( .A(n128), .B(n10886), .Z(n10884) );
  XOR U14744 ( .A(n10887), .B(n10888), .Z(n10886) );
  XOR U14745 ( .A(DB[2987]), .B(DB[2956]), .Z(n10888) );
  AND U14746 ( .A(n132), .B(n10889), .Z(n10887) );
  XOR U14747 ( .A(n10890), .B(n10891), .Z(n10889) );
  XOR U14748 ( .A(DB[2956]), .B(DB[2925]), .Z(n10891) );
  AND U14749 ( .A(n136), .B(n10892), .Z(n10890) );
  XOR U14750 ( .A(n10893), .B(n10894), .Z(n10892) );
  XOR U14751 ( .A(DB[2925]), .B(DB[2894]), .Z(n10894) );
  AND U14752 ( .A(n140), .B(n10895), .Z(n10893) );
  XOR U14753 ( .A(n10896), .B(n10897), .Z(n10895) );
  XOR U14754 ( .A(DB[2894]), .B(DB[2863]), .Z(n10897) );
  AND U14755 ( .A(n144), .B(n10898), .Z(n10896) );
  XOR U14756 ( .A(n10899), .B(n10900), .Z(n10898) );
  XOR U14757 ( .A(DB[2863]), .B(DB[2832]), .Z(n10900) );
  AND U14758 ( .A(n148), .B(n10901), .Z(n10899) );
  XOR U14759 ( .A(n10902), .B(n10903), .Z(n10901) );
  XOR U14760 ( .A(DB[2832]), .B(DB[2801]), .Z(n10903) );
  AND U14761 ( .A(n152), .B(n10904), .Z(n10902) );
  XOR U14762 ( .A(n10905), .B(n10906), .Z(n10904) );
  XOR U14763 ( .A(DB[2801]), .B(DB[2770]), .Z(n10906) );
  AND U14764 ( .A(n156), .B(n10907), .Z(n10905) );
  XOR U14765 ( .A(n10908), .B(n10909), .Z(n10907) );
  XOR U14766 ( .A(DB[2770]), .B(DB[2739]), .Z(n10909) );
  AND U14767 ( .A(n160), .B(n10910), .Z(n10908) );
  XOR U14768 ( .A(n10911), .B(n10912), .Z(n10910) );
  XOR U14769 ( .A(DB[2739]), .B(DB[2708]), .Z(n10912) );
  AND U14770 ( .A(n164), .B(n10913), .Z(n10911) );
  XOR U14771 ( .A(n10914), .B(n10915), .Z(n10913) );
  XOR U14772 ( .A(DB[2708]), .B(DB[2677]), .Z(n10915) );
  AND U14773 ( .A(n168), .B(n10916), .Z(n10914) );
  XOR U14774 ( .A(n10917), .B(n10918), .Z(n10916) );
  XOR U14775 ( .A(DB[2677]), .B(DB[2646]), .Z(n10918) );
  AND U14776 ( .A(n172), .B(n10919), .Z(n10917) );
  XOR U14777 ( .A(n10920), .B(n10921), .Z(n10919) );
  XOR U14778 ( .A(DB[2646]), .B(DB[2615]), .Z(n10921) );
  AND U14779 ( .A(n176), .B(n10922), .Z(n10920) );
  XOR U14780 ( .A(n10923), .B(n10924), .Z(n10922) );
  XOR U14781 ( .A(DB[2615]), .B(DB[2584]), .Z(n10924) );
  AND U14782 ( .A(n180), .B(n10925), .Z(n10923) );
  XOR U14783 ( .A(n10926), .B(n10927), .Z(n10925) );
  XOR U14784 ( .A(DB[2584]), .B(DB[2553]), .Z(n10927) );
  AND U14785 ( .A(n184), .B(n10928), .Z(n10926) );
  XOR U14786 ( .A(n10929), .B(n10930), .Z(n10928) );
  XOR U14787 ( .A(DB[2553]), .B(DB[2522]), .Z(n10930) );
  AND U14788 ( .A(n188), .B(n10931), .Z(n10929) );
  XOR U14789 ( .A(n10932), .B(n10933), .Z(n10931) );
  XOR U14790 ( .A(DB[2522]), .B(DB[2491]), .Z(n10933) );
  AND U14791 ( .A(n192), .B(n10934), .Z(n10932) );
  XOR U14792 ( .A(n10935), .B(n10936), .Z(n10934) );
  XOR U14793 ( .A(DB[2491]), .B(DB[2460]), .Z(n10936) );
  AND U14794 ( .A(n196), .B(n10937), .Z(n10935) );
  XOR U14795 ( .A(n10938), .B(n10939), .Z(n10937) );
  XOR U14796 ( .A(DB[2460]), .B(DB[2429]), .Z(n10939) );
  AND U14797 ( .A(n200), .B(n10940), .Z(n10938) );
  XOR U14798 ( .A(n10941), .B(n10942), .Z(n10940) );
  XOR U14799 ( .A(DB[2429]), .B(DB[2398]), .Z(n10942) );
  AND U14800 ( .A(n204), .B(n10943), .Z(n10941) );
  XOR U14801 ( .A(n10944), .B(n10945), .Z(n10943) );
  XOR U14802 ( .A(DB[2398]), .B(DB[2367]), .Z(n10945) );
  AND U14803 ( .A(n208), .B(n10946), .Z(n10944) );
  XOR U14804 ( .A(n10947), .B(n10948), .Z(n10946) );
  XOR U14805 ( .A(DB[2367]), .B(DB[2336]), .Z(n10948) );
  AND U14806 ( .A(n212), .B(n10949), .Z(n10947) );
  XOR U14807 ( .A(n10950), .B(n10951), .Z(n10949) );
  XOR U14808 ( .A(DB[2336]), .B(DB[2305]), .Z(n10951) );
  AND U14809 ( .A(n216), .B(n10952), .Z(n10950) );
  XOR U14810 ( .A(n10953), .B(n10954), .Z(n10952) );
  XOR U14811 ( .A(DB[2305]), .B(DB[2274]), .Z(n10954) );
  AND U14812 ( .A(n220), .B(n10955), .Z(n10953) );
  XOR U14813 ( .A(n10956), .B(n10957), .Z(n10955) );
  XOR U14814 ( .A(DB[2274]), .B(DB[2243]), .Z(n10957) );
  AND U14815 ( .A(n224), .B(n10958), .Z(n10956) );
  XOR U14816 ( .A(n10959), .B(n10960), .Z(n10958) );
  XOR U14817 ( .A(DB[2243]), .B(DB[2212]), .Z(n10960) );
  AND U14818 ( .A(n228), .B(n10961), .Z(n10959) );
  XOR U14819 ( .A(n10962), .B(n10963), .Z(n10961) );
  XOR U14820 ( .A(DB[2212]), .B(DB[2181]), .Z(n10963) );
  AND U14821 ( .A(n232), .B(n10964), .Z(n10962) );
  XOR U14822 ( .A(n10965), .B(n10966), .Z(n10964) );
  XOR U14823 ( .A(DB[2181]), .B(DB[2150]), .Z(n10966) );
  AND U14824 ( .A(n236), .B(n10967), .Z(n10965) );
  XOR U14825 ( .A(n10968), .B(n10969), .Z(n10967) );
  XOR U14826 ( .A(DB[2150]), .B(DB[2119]), .Z(n10969) );
  AND U14827 ( .A(n240), .B(n10970), .Z(n10968) );
  XOR U14828 ( .A(n10971), .B(n10972), .Z(n10970) );
  XOR U14829 ( .A(DB[2119]), .B(DB[2088]), .Z(n10972) );
  AND U14830 ( .A(n244), .B(n10973), .Z(n10971) );
  XOR U14831 ( .A(n10974), .B(n10975), .Z(n10973) );
  XOR U14832 ( .A(DB[2088]), .B(DB[2057]), .Z(n10975) );
  AND U14833 ( .A(n248), .B(n10976), .Z(n10974) );
  XOR U14834 ( .A(n10977), .B(n10978), .Z(n10976) );
  XOR U14835 ( .A(DB[2057]), .B(DB[2026]), .Z(n10978) );
  AND U14836 ( .A(n252), .B(n10979), .Z(n10977) );
  XOR U14837 ( .A(n10980), .B(n10981), .Z(n10979) );
  XOR U14838 ( .A(DB[2026]), .B(DB[1995]), .Z(n10981) );
  AND U14839 ( .A(n256), .B(n10982), .Z(n10980) );
  XOR U14840 ( .A(n10983), .B(n10984), .Z(n10982) );
  XOR U14841 ( .A(DB[1995]), .B(DB[1964]), .Z(n10984) );
  AND U14842 ( .A(n260), .B(n10985), .Z(n10983) );
  XOR U14843 ( .A(n10986), .B(n10987), .Z(n10985) );
  XOR U14844 ( .A(DB[1964]), .B(DB[1933]), .Z(n10987) );
  AND U14845 ( .A(n264), .B(n10988), .Z(n10986) );
  XOR U14846 ( .A(n10989), .B(n10990), .Z(n10988) );
  XOR U14847 ( .A(DB[1933]), .B(DB[1902]), .Z(n10990) );
  AND U14848 ( .A(n268), .B(n10991), .Z(n10989) );
  XOR U14849 ( .A(n10992), .B(n10993), .Z(n10991) );
  XOR U14850 ( .A(DB[1902]), .B(DB[1871]), .Z(n10993) );
  AND U14851 ( .A(n272), .B(n10994), .Z(n10992) );
  XOR U14852 ( .A(n10995), .B(n10996), .Z(n10994) );
  XOR U14853 ( .A(DB[1871]), .B(DB[1840]), .Z(n10996) );
  AND U14854 ( .A(n276), .B(n10997), .Z(n10995) );
  XOR U14855 ( .A(n10998), .B(n10999), .Z(n10997) );
  XOR U14856 ( .A(DB[1840]), .B(DB[1809]), .Z(n10999) );
  AND U14857 ( .A(n280), .B(n11000), .Z(n10998) );
  XOR U14858 ( .A(n11001), .B(n11002), .Z(n11000) );
  XOR U14859 ( .A(DB[1809]), .B(DB[1778]), .Z(n11002) );
  AND U14860 ( .A(n284), .B(n11003), .Z(n11001) );
  XOR U14861 ( .A(n11004), .B(n11005), .Z(n11003) );
  XOR U14862 ( .A(DB[1778]), .B(DB[1747]), .Z(n11005) );
  AND U14863 ( .A(n288), .B(n11006), .Z(n11004) );
  XOR U14864 ( .A(n11007), .B(n11008), .Z(n11006) );
  XOR U14865 ( .A(DB[1747]), .B(DB[1716]), .Z(n11008) );
  AND U14866 ( .A(n292), .B(n11009), .Z(n11007) );
  XOR U14867 ( .A(n11010), .B(n11011), .Z(n11009) );
  XOR U14868 ( .A(DB[1716]), .B(DB[1685]), .Z(n11011) );
  AND U14869 ( .A(n296), .B(n11012), .Z(n11010) );
  XOR U14870 ( .A(n11013), .B(n11014), .Z(n11012) );
  XOR U14871 ( .A(DB[1685]), .B(DB[1654]), .Z(n11014) );
  AND U14872 ( .A(n300), .B(n11015), .Z(n11013) );
  XOR U14873 ( .A(n11016), .B(n11017), .Z(n11015) );
  XOR U14874 ( .A(DB[1654]), .B(DB[1623]), .Z(n11017) );
  AND U14875 ( .A(n304), .B(n11018), .Z(n11016) );
  XOR U14876 ( .A(n11019), .B(n11020), .Z(n11018) );
  XOR U14877 ( .A(DB[1623]), .B(DB[1592]), .Z(n11020) );
  AND U14878 ( .A(n308), .B(n11021), .Z(n11019) );
  XOR U14879 ( .A(n11022), .B(n11023), .Z(n11021) );
  XOR U14880 ( .A(DB[1592]), .B(DB[1561]), .Z(n11023) );
  AND U14881 ( .A(n312), .B(n11024), .Z(n11022) );
  XOR U14882 ( .A(n11025), .B(n11026), .Z(n11024) );
  XOR U14883 ( .A(DB[1561]), .B(DB[1530]), .Z(n11026) );
  AND U14884 ( .A(n316), .B(n11027), .Z(n11025) );
  XOR U14885 ( .A(n11028), .B(n11029), .Z(n11027) );
  XOR U14886 ( .A(DB[1530]), .B(DB[1499]), .Z(n11029) );
  AND U14887 ( .A(n320), .B(n11030), .Z(n11028) );
  XOR U14888 ( .A(n11031), .B(n11032), .Z(n11030) );
  XOR U14889 ( .A(DB[1499]), .B(DB[1468]), .Z(n11032) );
  AND U14890 ( .A(n324), .B(n11033), .Z(n11031) );
  XOR U14891 ( .A(n11034), .B(n11035), .Z(n11033) );
  XOR U14892 ( .A(DB[1468]), .B(DB[1437]), .Z(n11035) );
  AND U14893 ( .A(n328), .B(n11036), .Z(n11034) );
  XOR U14894 ( .A(n11037), .B(n11038), .Z(n11036) );
  XOR U14895 ( .A(DB[1437]), .B(DB[1406]), .Z(n11038) );
  AND U14896 ( .A(n332), .B(n11039), .Z(n11037) );
  XOR U14897 ( .A(n11040), .B(n11041), .Z(n11039) );
  XOR U14898 ( .A(DB[1406]), .B(DB[1375]), .Z(n11041) );
  AND U14899 ( .A(n336), .B(n11042), .Z(n11040) );
  XOR U14900 ( .A(n11043), .B(n11044), .Z(n11042) );
  XOR U14901 ( .A(DB[1375]), .B(DB[1344]), .Z(n11044) );
  AND U14902 ( .A(n340), .B(n11045), .Z(n11043) );
  XOR U14903 ( .A(n11046), .B(n11047), .Z(n11045) );
  XOR U14904 ( .A(DB[1344]), .B(DB[1313]), .Z(n11047) );
  AND U14905 ( .A(n344), .B(n11048), .Z(n11046) );
  XOR U14906 ( .A(n11049), .B(n11050), .Z(n11048) );
  XOR U14907 ( .A(DB[1313]), .B(DB[1282]), .Z(n11050) );
  AND U14908 ( .A(n348), .B(n11051), .Z(n11049) );
  XOR U14909 ( .A(n11052), .B(n11053), .Z(n11051) );
  XOR U14910 ( .A(DB[1282]), .B(DB[1251]), .Z(n11053) );
  AND U14911 ( .A(n352), .B(n11054), .Z(n11052) );
  XOR U14912 ( .A(n11055), .B(n11056), .Z(n11054) );
  XOR U14913 ( .A(DB[1251]), .B(DB[1220]), .Z(n11056) );
  AND U14914 ( .A(n356), .B(n11057), .Z(n11055) );
  XOR U14915 ( .A(n11058), .B(n11059), .Z(n11057) );
  XOR U14916 ( .A(DB[1220]), .B(DB[1189]), .Z(n11059) );
  AND U14917 ( .A(n360), .B(n11060), .Z(n11058) );
  XOR U14918 ( .A(n11061), .B(n11062), .Z(n11060) );
  XOR U14919 ( .A(DB[1189]), .B(DB[1158]), .Z(n11062) );
  AND U14920 ( .A(n364), .B(n11063), .Z(n11061) );
  XOR U14921 ( .A(n11064), .B(n11065), .Z(n11063) );
  XOR U14922 ( .A(DB[1158]), .B(DB[1127]), .Z(n11065) );
  AND U14923 ( .A(n368), .B(n11066), .Z(n11064) );
  XOR U14924 ( .A(n11067), .B(n11068), .Z(n11066) );
  XOR U14925 ( .A(DB[1127]), .B(DB[1096]), .Z(n11068) );
  AND U14926 ( .A(n372), .B(n11069), .Z(n11067) );
  XOR U14927 ( .A(n11070), .B(n11071), .Z(n11069) );
  XOR U14928 ( .A(DB[1096]), .B(DB[1065]), .Z(n11071) );
  AND U14929 ( .A(n376), .B(n11072), .Z(n11070) );
  XOR U14930 ( .A(n11073), .B(n11074), .Z(n11072) );
  XOR U14931 ( .A(DB[1065]), .B(DB[1034]), .Z(n11074) );
  AND U14932 ( .A(n380), .B(n11075), .Z(n11073) );
  XOR U14933 ( .A(n11076), .B(n11077), .Z(n11075) );
  XOR U14934 ( .A(DB[1034]), .B(DB[1003]), .Z(n11077) );
  AND U14935 ( .A(n384), .B(n11078), .Z(n11076) );
  XOR U14936 ( .A(n11079), .B(n11080), .Z(n11078) );
  XOR U14937 ( .A(DB[972]), .B(DB[1003]), .Z(n11080) );
  AND U14938 ( .A(n388), .B(n11081), .Z(n11079) );
  XOR U14939 ( .A(n11082), .B(n11083), .Z(n11081) );
  XOR U14940 ( .A(DB[972]), .B(DB[941]), .Z(n11083) );
  AND U14941 ( .A(n392), .B(n11084), .Z(n11082) );
  XOR U14942 ( .A(n11085), .B(n11086), .Z(n11084) );
  XOR U14943 ( .A(DB[941]), .B(DB[910]), .Z(n11086) );
  AND U14944 ( .A(n396), .B(n11087), .Z(n11085) );
  XOR U14945 ( .A(n11088), .B(n11089), .Z(n11087) );
  XOR U14946 ( .A(DB[910]), .B(DB[879]), .Z(n11089) );
  AND U14947 ( .A(n400), .B(n11090), .Z(n11088) );
  XOR U14948 ( .A(n11091), .B(n11092), .Z(n11090) );
  XOR U14949 ( .A(DB[879]), .B(DB[848]), .Z(n11092) );
  AND U14950 ( .A(n404), .B(n11093), .Z(n11091) );
  XOR U14951 ( .A(n11094), .B(n11095), .Z(n11093) );
  XOR U14952 ( .A(DB[848]), .B(DB[817]), .Z(n11095) );
  AND U14953 ( .A(n408), .B(n11096), .Z(n11094) );
  XOR U14954 ( .A(n11097), .B(n11098), .Z(n11096) );
  XOR U14955 ( .A(DB[817]), .B(DB[786]), .Z(n11098) );
  AND U14956 ( .A(n412), .B(n11099), .Z(n11097) );
  XOR U14957 ( .A(n11100), .B(n11101), .Z(n11099) );
  XOR U14958 ( .A(DB[786]), .B(DB[755]), .Z(n11101) );
  AND U14959 ( .A(n416), .B(n11102), .Z(n11100) );
  XOR U14960 ( .A(n11103), .B(n11104), .Z(n11102) );
  XOR U14961 ( .A(DB[755]), .B(DB[724]), .Z(n11104) );
  AND U14962 ( .A(n420), .B(n11105), .Z(n11103) );
  XOR U14963 ( .A(n11106), .B(n11107), .Z(n11105) );
  XOR U14964 ( .A(DB[724]), .B(DB[693]), .Z(n11107) );
  AND U14965 ( .A(n424), .B(n11108), .Z(n11106) );
  XOR U14966 ( .A(n11109), .B(n11110), .Z(n11108) );
  XOR U14967 ( .A(DB[693]), .B(DB[662]), .Z(n11110) );
  AND U14968 ( .A(n428), .B(n11111), .Z(n11109) );
  XOR U14969 ( .A(n11112), .B(n11113), .Z(n11111) );
  XOR U14970 ( .A(DB[662]), .B(DB[631]), .Z(n11113) );
  AND U14971 ( .A(n432), .B(n11114), .Z(n11112) );
  XOR U14972 ( .A(n11115), .B(n11116), .Z(n11114) );
  XOR U14973 ( .A(DB[631]), .B(DB[600]), .Z(n11116) );
  AND U14974 ( .A(n436), .B(n11117), .Z(n11115) );
  XOR U14975 ( .A(n11118), .B(n11119), .Z(n11117) );
  XOR U14976 ( .A(DB[600]), .B(DB[569]), .Z(n11119) );
  AND U14977 ( .A(n440), .B(n11120), .Z(n11118) );
  XOR U14978 ( .A(n11121), .B(n11122), .Z(n11120) );
  XOR U14979 ( .A(DB[569]), .B(DB[538]), .Z(n11122) );
  AND U14980 ( .A(n444), .B(n11123), .Z(n11121) );
  XOR U14981 ( .A(n11124), .B(n11125), .Z(n11123) );
  XOR U14982 ( .A(DB[538]), .B(DB[507]), .Z(n11125) );
  AND U14983 ( .A(n448), .B(n11126), .Z(n11124) );
  XOR U14984 ( .A(n11127), .B(n11128), .Z(n11126) );
  XOR U14985 ( .A(DB[507]), .B(DB[476]), .Z(n11128) );
  AND U14986 ( .A(n452), .B(n11129), .Z(n11127) );
  XOR U14987 ( .A(n11130), .B(n11131), .Z(n11129) );
  XOR U14988 ( .A(DB[476]), .B(DB[445]), .Z(n11131) );
  AND U14989 ( .A(n456), .B(n11132), .Z(n11130) );
  XOR U14990 ( .A(n11133), .B(n11134), .Z(n11132) );
  XOR U14991 ( .A(DB[445]), .B(DB[414]), .Z(n11134) );
  AND U14992 ( .A(n460), .B(n11135), .Z(n11133) );
  XOR U14993 ( .A(n11136), .B(n11137), .Z(n11135) );
  XOR U14994 ( .A(DB[414]), .B(DB[383]), .Z(n11137) );
  AND U14995 ( .A(n464), .B(n11138), .Z(n11136) );
  XOR U14996 ( .A(n11139), .B(n11140), .Z(n11138) );
  XOR U14997 ( .A(DB[383]), .B(DB[352]), .Z(n11140) );
  AND U14998 ( .A(n468), .B(n11141), .Z(n11139) );
  XOR U14999 ( .A(n11142), .B(n11143), .Z(n11141) );
  XOR U15000 ( .A(DB[352]), .B(DB[321]), .Z(n11143) );
  AND U15001 ( .A(n472), .B(n11144), .Z(n11142) );
  XOR U15002 ( .A(n11145), .B(n11146), .Z(n11144) );
  XOR U15003 ( .A(DB[321]), .B(DB[290]), .Z(n11146) );
  AND U15004 ( .A(n476), .B(n11147), .Z(n11145) );
  XOR U15005 ( .A(n11148), .B(n11149), .Z(n11147) );
  XOR U15006 ( .A(DB[290]), .B(DB[259]), .Z(n11149) );
  AND U15007 ( .A(n480), .B(n11150), .Z(n11148) );
  XOR U15008 ( .A(n11151), .B(n11152), .Z(n11150) );
  XOR U15009 ( .A(DB[259]), .B(DB[228]), .Z(n11152) );
  AND U15010 ( .A(n484), .B(n11153), .Z(n11151) );
  XOR U15011 ( .A(n11154), .B(n11155), .Z(n11153) );
  XOR U15012 ( .A(DB[228]), .B(DB[197]), .Z(n11155) );
  AND U15013 ( .A(n488), .B(n11156), .Z(n11154) );
  XOR U15014 ( .A(n11157), .B(n11158), .Z(n11156) );
  XOR U15015 ( .A(DB[197]), .B(DB[166]), .Z(n11158) );
  AND U15016 ( .A(n492), .B(n11159), .Z(n11157) );
  XOR U15017 ( .A(n11160), .B(n11161), .Z(n11159) );
  XOR U15018 ( .A(DB[166]), .B(DB[135]), .Z(n11161) );
  AND U15019 ( .A(n496), .B(n11162), .Z(n11160) );
  XOR U15020 ( .A(n11163), .B(n11164), .Z(n11162) );
  XOR U15021 ( .A(DB[135]), .B(DB[104]), .Z(n11164) );
  AND U15022 ( .A(n500), .B(n11165), .Z(n11163) );
  XOR U15023 ( .A(n11166), .B(n11167), .Z(n11165) );
  XOR U15024 ( .A(DB[73]), .B(DB[104]), .Z(n11167) );
  AND U15025 ( .A(n504), .B(n11168), .Z(n11166) );
  XOR U15026 ( .A(n11169), .B(n11170), .Z(n11168) );
  XOR U15027 ( .A(DB[73]), .B(DB[42]), .Z(n11170) );
  AND U15028 ( .A(n508), .B(n11171), .Z(n11169) );
  XOR U15029 ( .A(DB[42]), .B(DB[11]), .Z(n11171) );
  XOR U15030 ( .A(DB[3947]), .B(n11172), .Z(min_val_out[10]) );
  AND U15031 ( .A(n2), .B(n11173), .Z(n11172) );
  XOR U15032 ( .A(n11174), .B(n11175), .Z(n11173) );
  XOR U15033 ( .A(n11176), .B(n11177), .Z(n11175) );
  IV U15034 ( .A(DB[3947]), .Z(n11176) );
  AND U15035 ( .A(n8), .B(n11178), .Z(n11174) );
  XOR U15036 ( .A(n11179), .B(n11180), .Z(n11178) );
  XOR U15037 ( .A(DB[3916]), .B(DB[3885]), .Z(n11180) );
  AND U15038 ( .A(n12), .B(n11181), .Z(n11179) );
  XOR U15039 ( .A(n11182), .B(n11183), .Z(n11181) );
  XOR U15040 ( .A(DB[3885]), .B(DB[3854]), .Z(n11183) );
  AND U15041 ( .A(n16), .B(n11184), .Z(n11182) );
  XOR U15042 ( .A(n11185), .B(n11186), .Z(n11184) );
  XOR U15043 ( .A(DB[3854]), .B(DB[3823]), .Z(n11186) );
  AND U15044 ( .A(n20), .B(n11187), .Z(n11185) );
  XOR U15045 ( .A(n11188), .B(n11189), .Z(n11187) );
  XOR U15046 ( .A(DB[3823]), .B(DB[3792]), .Z(n11189) );
  AND U15047 ( .A(n24), .B(n11190), .Z(n11188) );
  XOR U15048 ( .A(n11191), .B(n11192), .Z(n11190) );
  XOR U15049 ( .A(DB[3792]), .B(DB[3761]), .Z(n11192) );
  AND U15050 ( .A(n28), .B(n11193), .Z(n11191) );
  XOR U15051 ( .A(n11194), .B(n11195), .Z(n11193) );
  XOR U15052 ( .A(DB[3761]), .B(DB[3730]), .Z(n11195) );
  AND U15053 ( .A(n32), .B(n11196), .Z(n11194) );
  XOR U15054 ( .A(n11197), .B(n11198), .Z(n11196) );
  XOR U15055 ( .A(DB[3730]), .B(DB[3699]), .Z(n11198) );
  AND U15056 ( .A(n36), .B(n11199), .Z(n11197) );
  XOR U15057 ( .A(n11200), .B(n11201), .Z(n11199) );
  XOR U15058 ( .A(DB[3699]), .B(DB[3668]), .Z(n11201) );
  AND U15059 ( .A(n40), .B(n11202), .Z(n11200) );
  XOR U15060 ( .A(n11203), .B(n11204), .Z(n11202) );
  XOR U15061 ( .A(DB[3668]), .B(DB[3637]), .Z(n11204) );
  AND U15062 ( .A(n44), .B(n11205), .Z(n11203) );
  XOR U15063 ( .A(n11206), .B(n11207), .Z(n11205) );
  XOR U15064 ( .A(DB[3637]), .B(DB[3606]), .Z(n11207) );
  AND U15065 ( .A(n48), .B(n11208), .Z(n11206) );
  XOR U15066 ( .A(n11209), .B(n11210), .Z(n11208) );
  XOR U15067 ( .A(DB[3606]), .B(DB[3575]), .Z(n11210) );
  AND U15068 ( .A(n52), .B(n11211), .Z(n11209) );
  XOR U15069 ( .A(n11212), .B(n11213), .Z(n11211) );
  XOR U15070 ( .A(DB[3575]), .B(DB[3544]), .Z(n11213) );
  AND U15071 ( .A(n56), .B(n11214), .Z(n11212) );
  XOR U15072 ( .A(n11215), .B(n11216), .Z(n11214) );
  XOR U15073 ( .A(DB[3544]), .B(DB[3513]), .Z(n11216) );
  AND U15074 ( .A(n60), .B(n11217), .Z(n11215) );
  XOR U15075 ( .A(n11218), .B(n11219), .Z(n11217) );
  XOR U15076 ( .A(DB[3513]), .B(DB[3482]), .Z(n11219) );
  AND U15077 ( .A(n64), .B(n11220), .Z(n11218) );
  XOR U15078 ( .A(n11221), .B(n11222), .Z(n11220) );
  XOR U15079 ( .A(DB[3482]), .B(DB[3451]), .Z(n11222) );
  AND U15080 ( .A(n68), .B(n11223), .Z(n11221) );
  XOR U15081 ( .A(n11224), .B(n11225), .Z(n11223) );
  XOR U15082 ( .A(DB[3451]), .B(DB[3420]), .Z(n11225) );
  AND U15083 ( .A(n72), .B(n11226), .Z(n11224) );
  XOR U15084 ( .A(n11227), .B(n11228), .Z(n11226) );
  XOR U15085 ( .A(DB[3420]), .B(DB[3389]), .Z(n11228) );
  AND U15086 ( .A(n76), .B(n11229), .Z(n11227) );
  XOR U15087 ( .A(n11230), .B(n11231), .Z(n11229) );
  XOR U15088 ( .A(DB[3389]), .B(DB[3358]), .Z(n11231) );
  AND U15089 ( .A(n80), .B(n11232), .Z(n11230) );
  XOR U15090 ( .A(n11233), .B(n11234), .Z(n11232) );
  XOR U15091 ( .A(DB[3358]), .B(DB[3327]), .Z(n11234) );
  AND U15092 ( .A(n84), .B(n11235), .Z(n11233) );
  XOR U15093 ( .A(n11236), .B(n11237), .Z(n11235) );
  XOR U15094 ( .A(DB[3327]), .B(DB[3296]), .Z(n11237) );
  AND U15095 ( .A(n88), .B(n11238), .Z(n11236) );
  XOR U15096 ( .A(n11239), .B(n11240), .Z(n11238) );
  XOR U15097 ( .A(DB[3296]), .B(DB[3265]), .Z(n11240) );
  AND U15098 ( .A(n92), .B(n11241), .Z(n11239) );
  XOR U15099 ( .A(n11242), .B(n11243), .Z(n11241) );
  XOR U15100 ( .A(DB[3265]), .B(DB[3234]), .Z(n11243) );
  AND U15101 ( .A(n96), .B(n11244), .Z(n11242) );
  XOR U15102 ( .A(n11245), .B(n11246), .Z(n11244) );
  XOR U15103 ( .A(DB[3234]), .B(DB[3203]), .Z(n11246) );
  AND U15104 ( .A(n100), .B(n11247), .Z(n11245) );
  XOR U15105 ( .A(n11248), .B(n11249), .Z(n11247) );
  XOR U15106 ( .A(DB[3203]), .B(DB[3172]), .Z(n11249) );
  AND U15107 ( .A(n104), .B(n11250), .Z(n11248) );
  XOR U15108 ( .A(n11251), .B(n11252), .Z(n11250) );
  XOR U15109 ( .A(DB[3172]), .B(DB[3141]), .Z(n11252) );
  AND U15110 ( .A(n108), .B(n11253), .Z(n11251) );
  XOR U15111 ( .A(n11254), .B(n11255), .Z(n11253) );
  XOR U15112 ( .A(DB[3141]), .B(DB[3110]), .Z(n11255) );
  AND U15113 ( .A(n112), .B(n11256), .Z(n11254) );
  XOR U15114 ( .A(n11257), .B(n11258), .Z(n11256) );
  XOR U15115 ( .A(DB[3110]), .B(DB[3079]), .Z(n11258) );
  AND U15116 ( .A(n116), .B(n11259), .Z(n11257) );
  XOR U15117 ( .A(n11260), .B(n11261), .Z(n11259) );
  XOR U15118 ( .A(DB[3079]), .B(DB[3048]), .Z(n11261) );
  AND U15119 ( .A(n120), .B(n11262), .Z(n11260) );
  XOR U15120 ( .A(n11263), .B(n11264), .Z(n11262) );
  XOR U15121 ( .A(DB[3048]), .B(DB[3017]), .Z(n11264) );
  AND U15122 ( .A(n124), .B(n11265), .Z(n11263) );
  XOR U15123 ( .A(n11266), .B(n11267), .Z(n11265) );
  XOR U15124 ( .A(DB[3017]), .B(DB[2986]), .Z(n11267) );
  AND U15125 ( .A(n128), .B(n11268), .Z(n11266) );
  XOR U15126 ( .A(n11269), .B(n11270), .Z(n11268) );
  XOR U15127 ( .A(DB[2986]), .B(DB[2955]), .Z(n11270) );
  AND U15128 ( .A(n132), .B(n11271), .Z(n11269) );
  XOR U15129 ( .A(n11272), .B(n11273), .Z(n11271) );
  XOR U15130 ( .A(DB[2955]), .B(DB[2924]), .Z(n11273) );
  AND U15131 ( .A(n136), .B(n11274), .Z(n11272) );
  XOR U15132 ( .A(n11275), .B(n11276), .Z(n11274) );
  XOR U15133 ( .A(DB[2924]), .B(DB[2893]), .Z(n11276) );
  AND U15134 ( .A(n140), .B(n11277), .Z(n11275) );
  XOR U15135 ( .A(n11278), .B(n11279), .Z(n11277) );
  XOR U15136 ( .A(DB[2893]), .B(DB[2862]), .Z(n11279) );
  AND U15137 ( .A(n144), .B(n11280), .Z(n11278) );
  XOR U15138 ( .A(n11281), .B(n11282), .Z(n11280) );
  XOR U15139 ( .A(DB[2862]), .B(DB[2831]), .Z(n11282) );
  AND U15140 ( .A(n148), .B(n11283), .Z(n11281) );
  XOR U15141 ( .A(n11284), .B(n11285), .Z(n11283) );
  XOR U15142 ( .A(DB[2831]), .B(DB[2800]), .Z(n11285) );
  AND U15143 ( .A(n152), .B(n11286), .Z(n11284) );
  XOR U15144 ( .A(n11287), .B(n11288), .Z(n11286) );
  XOR U15145 ( .A(DB[2800]), .B(DB[2769]), .Z(n11288) );
  AND U15146 ( .A(n156), .B(n11289), .Z(n11287) );
  XOR U15147 ( .A(n11290), .B(n11291), .Z(n11289) );
  XOR U15148 ( .A(DB[2769]), .B(DB[2738]), .Z(n11291) );
  AND U15149 ( .A(n160), .B(n11292), .Z(n11290) );
  XOR U15150 ( .A(n11293), .B(n11294), .Z(n11292) );
  XOR U15151 ( .A(DB[2738]), .B(DB[2707]), .Z(n11294) );
  AND U15152 ( .A(n164), .B(n11295), .Z(n11293) );
  XOR U15153 ( .A(n11296), .B(n11297), .Z(n11295) );
  XOR U15154 ( .A(DB[2707]), .B(DB[2676]), .Z(n11297) );
  AND U15155 ( .A(n168), .B(n11298), .Z(n11296) );
  XOR U15156 ( .A(n11299), .B(n11300), .Z(n11298) );
  XOR U15157 ( .A(DB[2676]), .B(DB[2645]), .Z(n11300) );
  AND U15158 ( .A(n172), .B(n11301), .Z(n11299) );
  XOR U15159 ( .A(n11302), .B(n11303), .Z(n11301) );
  XOR U15160 ( .A(DB[2645]), .B(DB[2614]), .Z(n11303) );
  AND U15161 ( .A(n176), .B(n11304), .Z(n11302) );
  XOR U15162 ( .A(n11305), .B(n11306), .Z(n11304) );
  XOR U15163 ( .A(DB[2614]), .B(DB[2583]), .Z(n11306) );
  AND U15164 ( .A(n180), .B(n11307), .Z(n11305) );
  XOR U15165 ( .A(n11308), .B(n11309), .Z(n11307) );
  XOR U15166 ( .A(DB[2583]), .B(DB[2552]), .Z(n11309) );
  AND U15167 ( .A(n184), .B(n11310), .Z(n11308) );
  XOR U15168 ( .A(n11311), .B(n11312), .Z(n11310) );
  XOR U15169 ( .A(DB[2552]), .B(DB[2521]), .Z(n11312) );
  AND U15170 ( .A(n188), .B(n11313), .Z(n11311) );
  XOR U15171 ( .A(n11314), .B(n11315), .Z(n11313) );
  XOR U15172 ( .A(DB[2521]), .B(DB[2490]), .Z(n11315) );
  AND U15173 ( .A(n192), .B(n11316), .Z(n11314) );
  XOR U15174 ( .A(n11317), .B(n11318), .Z(n11316) );
  XOR U15175 ( .A(DB[2490]), .B(DB[2459]), .Z(n11318) );
  AND U15176 ( .A(n196), .B(n11319), .Z(n11317) );
  XOR U15177 ( .A(n11320), .B(n11321), .Z(n11319) );
  XOR U15178 ( .A(DB[2459]), .B(DB[2428]), .Z(n11321) );
  AND U15179 ( .A(n200), .B(n11322), .Z(n11320) );
  XOR U15180 ( .A(n11323), .B(n11324), .Z(n11322) );
  XOR U15181 ( .A(DB[2428]), .B(DB[2397]), .Z(n11324) );
  AND U15182 ( .A(n204), .B(n11325), .Z(n11323) );
  XOR U15183 ( .A(n11326), .B(n11327), .Z(n11325) );
  XOR U15184 ( .A(DB[2397]), .B(DB[2366]), .Z(n11327) );
  AND U15185 ( .A(n208), .B(n11328), .Z(n11326) );
  XOR U15186 ( .A(n11329), .B(n11330), .Z(n11328) );
  XOR U15187 ( .A(DB[2366]), .B(DB[2335]), .Z(n11330) );
  AND U15188 ( .A(n212), .B(n11331), .Z(n11329) );
  XOR U15189 ( .A(n11332), .B(n11333), .Z(n11331) );
  XOR U15190 ( .A(DB[2335]), .B(DB[2304]), .Z(n11333) );
  AND U15191 ( .A(n216), .B(n11334), .Z(n11332) );
  XOR U15192 ( .A(n11335), .B(n11336), .Z(n11334) );
  XOR U15193 ( .A(DB[2304]), .B(DB[2273]), .Z(n11336) );
  AND U15194 ( .A(n220), .B(n11337), .Z(n11335) );
  XOR U15195 ( .A(n11338), .B(n11339), .Z(n11337) );
  XOR U15196 ( .A(DB[2273]), .B(DB[2242]), .Z(n11339) );
  AND U15197 ( .A(n224), .B(n11340), .Z(n11338) );
  XOR U15198 ( .A(n11341), .B(n11342), .Z(n11340) );
  XOR U15199 ( .A(DB[2242]), .B(DB[2211]), .Z(n11342) );
  AND U15200 ( .A(n228), .B(n11343), .Z(n11341) );
  XOR U15201 ( .A(n11344), .B(n11345), .Z(n11343) );
  XOR U15202 ( .A(DB[2211]), .B(DB[2180]), .Z(n11345) );
  AND U15203 ( .A(n232), .B(n11346), .Z(n11344) );
  XOR U15204 ( .A(n11347), .B(n11348), .Z(n11346) );
  XOR U15205 ( .A(DB[2180]), .B(DB[2149]), .Z(n11348) );
  AND U15206 ( .A(n236), .B(n11349), .Z(n11347) );
  XOR U15207 ( .A(n11350), .B(n11351), .Z(n11349) );
  XOR U15208 ( .A(DB[2149]), .B(DB[2118]), .Z(n11351) );
  AND U15209 ( .A(n240), .B(n11352), .Z(n11350) );
  XOR U15210 ( .A(n11353), .B(n11354), .Z(n11352) );
  XOR U15211 ( .A(DB[2118]), .B(DB[2087]), .Z(n11354) );
  AND U15212 ( .A(n244), .B(n11355), .Z(n11353) );
  XOR U15213 ( .A(n11356), .B(n11357), .Z(n11355) );
  XOR U15214 ( .A(DB[2087]), .B(DB[2056]), .Z(n11357) );
  AND U15215 ( .A(n248), .B(n11358), .Z(n11356) );
  XOR U15216 ( .A(n11359), .B(n11360), .Z(n11358) );
  XOR U15217 ( .A(DB[2056]), .B(DB[2025]), .Z(n11360) );
  AND U15218 ( .A(n252), .B(n11361), .Z(n11359) );
  XOR U15219 ( .A(n11362), .B(n11363), .Z(n11361) );
  XOR U15220 ( .A(DB[2025]), .B(DB[1994]), .Z(n11363) );
  AND U15221 ( .A(n256), .B(n11364), .Z(n11362) );
  XOR U15222 ( .A(n11365), .B(n11366), .Z(n11364) );
  XOR U15223 ( .A(DB[1994]), .B(DB[1963]), .Z(n11366) );
  AND U15224 ( .A(n260), .B(n11367), .Z(n11365) );
  XOR U15225 ( .A(n11368), .B(n11369), .Z(n11367) );
  XOR U15226 ( .A(DB[1963]), .B(DB[1932]), .Z(n11369) );
  AND U15227 ( .A(n264), .B(n11370), .Z(n11368) );
  XOR U15228 ( .A(n11371), .B(n11372), .Z(n11370) );
  XOR U15229 ( .A(DB[1932]), .B(DB[1901]), .Z(n11372) );
  AND U15230 ( .A(n268), .B(n11373), .Z(n11371) );
  XOR U15231 ( .A(n11374), .B(n11375), .Z(n11373) );
  XOR U15232 ( .A(DB[1901]), .B(DB[1870]), .Z(n11375) );
  AND U15233 ( .A(n272), .B(n11376), .Z(n11374) );
  XOR U15234 ( .A(n11377), .B(n11378), .Z(n11376) );
  XOR U15235 ( .A(DB[1870]), .B(DB[1839]), .Z(n11378) );
  AND U15236 ( .A(n276), .B(n11379), .Z(n11377) );
  XOR U15237 ( .A(n11380), .B(n11381), .Z(n11379) );
  XOR U15238 ( .A(DB[1839]), .B(DB[1808]), .Z(n11381) );
  AND U15239 ( .A(n280), .B(n11382), .Z(n11380) );
  XOR U15240 ( .A(n11383), .B(n11384), .Z(n11382) );
  XOR U15241 ( .A(DB[1808]), .B(DB[1777]), .Z(n11384) );
  AND U15242 ( .A(n284), .B(n11385), .Z(n11383) );
  XOR U15243 ( .A(n11386), .B(n11387), .Z(n11385) );
  XOR U15244 ( .A(DB[1777]), .B(DB[1746]), .Z(n11387) );
  AND U15245 ( .A(n288), .B(n11388), .Z(n11386) );
  XOR U15246 ( .A(n11389), .B(n11390), .Z(n11388) );
  XOR U15247 ( .A(DB[1746]), .B(DB[1715]), .Z(n11390) );
  AND U15248 ( .A(n292), .B(n11391), .Z(n11389) );
  XOR U15249 ( .A(n11392), .B(n11393), .Z(n11391) );
  XOR U15250 ( .A(DB[1715]), .B(DB[1684]), .Z(n11393) );
  AND U15251 ( .A(n296), .B(n11394), .Z(n11392) );
  XOR U15252 ( .A(n11395), .B(n11396), .Z(n11394) );
  XOR U15253 ( .A(DB[1684]), .B(DB[1653]), .Z(n11396) );
  AND U15254 ( .A(n300), .B(n11397), .Z(n11395) );
  XOR U15255 ( .A(n11398), .B(n11399), .Z(n11397) );
  XOR U15256 ( .A(DB[1653]), .B(DB[1622]), .Z(n11399) );
  AND U15257 ( .A(n304), .B(n11400), .Z(n11398) );
  XOR U15258 ( .A(n11401), .B(n11402), .Z(n11400) );
  XOR U15259 ( .A(DB[1622]), .B(DB[1591]), .Z(n11402) );
  AND U15260 ( .A(n308), .B(n11403), .Z(n11401) );
  XOR U15261 ( .A(n11404), .B(n11405), .Z(n11403) );
  XOR U15262 ( .A(DB[1591]), .B(DB[1560]), .Z(n11405) );
  AND U15263 ( .A(n312), .B(n11406), .Z(n11404) );
  XOR U15264 ( .A(n11407), .B(n11408), .Z(n11406) );
  XOR U15265 ( .A(DB[1560]), .B(DB[1529]), .Z(n11408) );
  AND U15266 ( .A(n316), .B(n11409), .Z(n11407) );
  XOR U15267 ( .A(n11410), .B(n11411), .Z(n11409) );
  XOR U15268 ( .A(DB[1529]), .B(DB[1498]), .Z(n11411) );
  AND U15269 ( .A(n320), .B(n11412), .Z(n11410) );
  XOR U15270 ( .A(n11413), .B(n11414), .Z(n11412) );
  XOR U15271 ( .A(DB[1498]), .B(DB[1467]), .Z(n11414) );
  AND U15272 ( .A(n324), .B(n11415), .Z(n11413) );
  XOR U15273 ( .A(n11416), .B(n11417), .Z(n11415) );
  XOR U15274 ( .A(DB[1467]), .B(DB[1436]), .Z(n11417) );
  AND U15275 ( .A(n328), .B(n11418), .Z(n11416) );
  XOR U15276 ( .A(n11419), .B(n11420), .Z(n11418) );
  XOR U15277 ( .A(DB[1436]), .B(DB[1405]), .Z(n11420) );
  AND U15278 ( .A(n332), .B(n11421), .Z(n11419) );
  XOR U15279 ( .A(n11422), .B(n11423), .Z(n11421) );
  XOR U15280 ( .A(DB[1405]), .B(DB[1374]), .Z(n11423) );
  AND U15281 ( .A(n336), .B(n11424), .Z(n11422) );
  XOR U15282 ( .A(n11425), .B(n11426), .Z(n11424) );
  XOR U15283 ( .A(DB[1374]), .B(DB[1343]), .Z(n11426) );
  AND U15284 ( .A(n340), .B(n11427), .Z(n11425) );
  XOR U15285 ( .A(n11428), .B(n11429), .Z(n11427) );
  XOR U15286 ( .A(DB[1343]), .B(DB[1312]), .Z(n11429) );
  AND U15287 ( .A(n344), .B(n11430), .Z(n11428) );
  XOR U15288 ( .A(n11431), .B(n11432), .Z(n11430) );
  XOR U15289 ( .A(DB[1312]), .B(DB[1281]), .Z(n11432) );
  AND U15290 ( .A(n348), .B(n11433), .Z(n11431) );
  XOR U15291 ( .A(n11434), .B(n11435), .Z(n11433) );
  XOR U15292 ( .A(DB[1281]), .B(DB[1250]), .Z(n11435) );
  AND U15293 ( .A(n352), .B(n11436), .Z(n11434) );
  XOR U15294 ( .A(n11437), .B(n11438), .Z(n11436) );
  XOR U15295 ( .A(DB[1250]), .B(DB[1219]), .Z(n11438) );
  AND U15296 ( .A(n356), .B(n11439), .Z(n11437) );
  XOR U15297 ( .A(n11440), .B(n11441), .Z(n11439) );
  XOR U15298 ( .A(DB[1219]), .B(DB[1188]), .Z(n11441) );
  AND U15299 ( .A(n360), .B(n11442), .Z(n11440) );
  XOR U15300 ( .A(n11443), .B(n11444), .Z(n11442) );
  XOR U15301 ( .A(DB[1188]), .B(DB[1157]), .Z(n11444) );
  AND U15302 ( .A(n364), .B(n11445), .Z(n11443) );
  XOR U15303 ( .A(n11446), .B(n11447), .Z(n11445) );
  XOR U15304 ( .A(DB[1157]), .B(DB[1126]), .Z(n11447) );
  AND U15305 ( .A(n368), .B(n11448), .Z(n11446) );
  XOR U15306 ( .A(n11449), .B(n11450), .Z(n11448) );
  XOR U15307 ( .A(DB[1126]), .B(DB[1095]), .Z(n11450) );
  AND U15308 ( .A(n372), .B(n11451), .Z(n11449) );
  XOR U15309 ( .A(n11452), .B(n11453), .Z(n11451) );
  XOR U15310 ( .A(DB[1095]), .B(DB[1064]), .Z(n11453) );
  AND U15311 ( .A(n376), .B(n11454), .Z(n11452) );
  XOR U15312 ( .A(n11455), .B(n11456), .Z(n11454) );
  XOR U15313 ( .A(DB[1064]), .B(DB[1033]), .Z(n11456) );
  AND U15314 ( .A(n380), .B(n11457), .Z(n11455) );
  XOR U15315 ( .A(n11458), .B(n11459), .Z(n11457) );
  XOR U15316 ( .A(DB[1033]), .B(DB[1002]), .Z(n11459) );
  AND U15317 ( .A(n384), .B(n11460), .Z(n11458) );
  XOR U15318 ( .A(n11461), .B(n11462), .Z(n11460) );
  XOR U15319 ( .A(DB[971]), .B(DB[1002]), .Z(n11462) );
  AND U15320 ( .A(n388), .B(n11463), .Z(n11461) );
  XOR U15321 ( .A(n11464), .B(n11465), .Z(n11463) );
  XOR U15322 ( .A(DB[971]), .B(DB[940]), .Z(n11465) );
  AND U15323 ( .A(n392), .B(n11466), .Z(n11464) );
  XOR U15324 ( .A(n11467), .B(n11468), .Z(n11466) );
  XOR U15325 ( .A(DB[940]), .B(DB[909]), .Z(n11468) );
  AND U15326 ( .A(n396), .B(n11469), .Z(n11467) );
  XOR U15327 ( .A(n11470), .B(n11471), .Z(n11469) );
  XOR U15328 ( .A(DB[909]), .B(DB[878]), .Z(n11471) );
  AND U15329 ( .A(n400), .B(n11472), .Z(n11470) );
  XOR U15330 ( .A(n11473), .B(n11474), .Z(n11472) );
  XOR U15331 ( .A(DB[878]), .B(DB[847]), .Z(n11474) );
  AND U15332 ( .A(n404), .B(n11475), .Z(n11473) );
  XOR U15333 ( .A(n11476), .B(n11477), .Z(n11475) );
  XOR U15334 ( .A(DB[847]), .B(DB[816]), .Z(n11477) );
  AND U15335 ( .A(n408), .B(n11478), .Z(n11476) );
  XOR U15336 ( .A(n11479), .B(n11480), .Z(n11478) );
  XOR U15337 ( .A(DB[816]), .B(DB[785]), .Z(n11480) );
  AND U15338 ( .A(n412), .B(n11481), .Z(n11479) );
  XOR U15339 ( .A(n11482), .B(n11483), .Z(n11481) );
  XOR U15340 ( .A(DB[785]), .B(DB[754]), .Z(n11483) );
  AND U15341 ( .A(n416), .B(n11484), .Z(n11482) );
  XOR U15342 ( .A(n11485), .B(n11486), .Z(n11484) );
  XOR U15343 ( .A(DB[754]), .B(DB[723]), .Z(n11486) );
  AND U15344 ( .A(n420), .B(n11487), .Z(n11485) );
  XOR U15345 ( .A(n11488), .B(n11489), .Z(n11487) );
  XOR U15346 ( .A(DB[723]), .B(DB[692]), .Z(n11489) );
  AND U15347 ( .A(n424), .B(n11490), .Z(n11488) );
  XOR U15348 ( .A(n11491), .B(n11492), .Z(n11490) );
  XOR U15349 ( .A(DB[692]), .B(DB[661]), .Z(n11492) );
  AND U15350 ( .A(n428), .B(n11493), .Z(n11491) );
  XOR U15351 ( .A(n11494), .B(n11495), .Z(n11493) );
  XOR U15352 ( .A(DB[661]), .B(DB[630]), .Z(n11495) );
  AND U15353 ( .A(n432), .B(n11496), .Z(n11494) );
  XOR U15354 ( .A(n11497), .B(n11498), .Z(n11496) );
  XOR U15355 ( .A(DB[630]), .B(DB[599]), .Z(n11498) );
  AND U15356 ( .A(n436), .B(n11499), .Z(n11497) );
  XOR U15357 ( .A(n11500), .B(n11501), .Z(n11499) );
  XOR U15358 ( .A(DB[599]), .B(DB[568]), .Z(n11501) );
  AND U15359 ( .A(n440), .B(n11502), .Z(n11500) );
  XOR U15360 ( .A(n11503), .B(n11504), .Z(n11502) );
  XOR U15361 ( .A(DB[568]), .B(DB[537]), .Z(n11504) );
  AND U15362 ( .A(n444), .B(n11505), .Z(n11503) );
  XOR U15363 ( .A(n11506), .B(n11507), .Z(n11505) );
  XOR U15364 ( .A(DB[537]), .B(DB[506]), .Z(n11507) );
  AND U15365 ( .A(n448), .B(n11508), .Z(n11506) );
  XOR U15366 ( .A(n11509), .B(n11510), .Z(n11508) );
  XOR U15367 ( .A(DB[506]), .B(DB[475]), .Z(n11510) );
  AND U15368 ( .A(n452), .B(n11511), .Z(n11509) );
  XOR U15369 ( .A(n11512), .B(n11513), .Z(n11511) );
  XOR U15370 ( .A(DB[475]), .B(DB[444]), .Z(n11513) );
  AND U15371 ( .A(n456), .B(n11514), .Z(n11512) );
  XOR U15372 ( .A(n11515), .B(n11516), .Z(n11514) );
  XOR U15373 ( .A(DB[444]), .B(DB[413]), .Z(n11516) );
  AND U15374 ( .A(n460), .B(n11517), .Z(n11515) );
  XOR U15375 ( .A(n11518), .B(n11519), .Z(n11517) );
  XOR U15376 ( .A(DB[413]), .B(DB[382]), .Z(n11519) );
  AND U15377 ( .A(n464), .B(n11520), .Z(n11518) );
  XOR U15378 ( .A(n11521), .B(n11522), .Z(n11520) );
  XOR U15379 ( .A(DB[382]), .B(DB[351]), .Z(n11522) );
  AND U15380 ( .A(n468), .B(n11523), .Z(n11521) );
  XOR U15381 ( .A(n11524), .B(n11525), .Z(n11523) );
  XOR U15382 ( .A(DB[351]), .B(DB[320]), .Z(n11525) );
  AND U15383 ( .A(n472), .B(n11526), .Z(n11524) );
  XOR U15384 ( .A(n11527), .B(n11528), .Z(n11526) );
  XOR U15385 ( .A(DB[320]), .B(DB[289]), .Z(n11528) );
  AND U15386 ( .A(n476), .B(n11529), .Z(n11527) );
  XOR U15387 ( .A(n11530), .B(n11531), .Z(n11529) );
  XOR U15388 ( .A(DB[289]), .B(DB[258]), .Z(n11531) );
  AND U15389 ( .A(n480), .B(n11532), .Z(n11530) );
  XOR U15390 ( .A(n11533), .B(n11534), .Z(n11532) );
  XOR U15391 ( .A(DB[258]), .B(DB[227]), .Z(n11534) );
  AND U15392 ( .A(n484), .B(n11535), .Z(n11533) );
  XOR U15393 ( .A(n11536), .B(n11537), .Z(n11535) );
  XOR U15394 ( .A(DB[227]), .B(DB[196]), .Z(n11537) );
  AND U15395 ( .A(n488), .B(n11538), .Z(n11536) );
  XOR U15396 ( .A(n11539), .B(n11540), .Z(n11538) );
  XOR U15397 ( .A(DB[196]), .B(DB[165]), .Z(n11540) );
  AND U15398 ( .A(n492), .B(n11541), .Z(n11539) );
  XOR U15399 ( .A(n11542), .B(n11543), .Z(n11541) );
  XOR U15400 ( .A(DB[165]), .B(DB[134]), .Z(n11543) );
  AND U15401 ( .A(n496), .B(n11544), .Z(n11542) );
  XOR U15402 ( .A(n11545), .B(n11546), .Z(n11544) );
  XOR U15403 ( .A(DB[134]), .B(DB[103]), .Z(n11546) );
  AND U15404 ( .A(n500), .B(n11547), .Z(n11545) );
  XOR U15405 ( .A(n11548), .B(n11549), .Z(n11547) );
  XOR U15406 ( .A(DB[72]), .B(DB[103]), .Z(n11549) );
  AND U15407 ( .A(n504), .B(n11550), .Z(n11548) );
  XOR U15408 ( .A(n11551), .B(n11552), .Z(n11550) );
  XOR U15409 ( .A(DB[72]), .B(DB[41]), .Z(n11552) );
  AND U15410 ( .A(n508), .B(n11553), .Z(n11551) );
  XOR U15411 ( .A(DB[41]), .B(DB[10]), .Z(n11553) );
  XOR U15412 ( .A(DB[3937]), .B(n11554), .Z(min_val_out[0]) );
  AND U15413 ( .A(n2), .B(n11555), .Z(n11554) );
  XOR U15414 ( .A(n11556), .B(n11557), .Z(n11555) );
  XOR U15415 ( .A(DB[3937]), .B(DB[3906]), .Z(n11557) );
  AND U15416 ( .A(n8), .B(n11558), .Z(n11556) );
  XOR U15417 ( .A(n11559), .B(n11560), .Z(n11558) );
  XOR U15418 ( .A(DB[3906]), .B(DB[3875]), .Z(n11560) );
  AND U15419 ( .A(n12), .B(n11561), .Z(n11559) );
  XOR U15420 ( .A(n11562), .B(n11563), .Z(n11561) );
  XOR U15421 ( .A(DB[3875]), .B(DB[3844]), .Z(n11563) );
  AND U15422 ( .A(n16), .B(n11564), .Z(n11562) );
  XOR U15423 ( .A(n11565), .B(n11566), .Z(n11564) );
  XOR U15424 ( .A(DB[3844]), .B(DB[3813]), .Z(n11566) );
  AND U15425 ( .A(n20), .B(n11567), .Z(n11565) );
  XOR U15426 ( .A(n11568), .B(n11569), .Z(n11567) );
  XOR U15427 ( .A(DB[3813]), .B(DB[3782]), .Z(n11569) );
  AND U15428 ( .A(n24), .B(n11570), .Z(n11568) );
  XOR U15429 ( .A(n11571), .B(n11572), .Z(n11570) );
  XOR U15430 ( .A(DB[3782]), .B(DB[3751]), .Z(n11572) );
  AND U15431 ( .A(n28), .B(n11573), .Z(n11571) );
  XOR U15432 ( .A(n11574), .B(n11575), .Z(n11573) );
  XOR U15433 ( .A(DB[3751]), .B(DB[3720]), .Z(n11575) );
  AND U15434 ( .A(n32), .B(n11576), .Z(n11574) );
  XOR U15435 ( .A(n11577), .B(n11578), .Z(n11576) );
  XOR U15436 ( .A(DB[3720]), .B(DB[3689]), .Z(n11578) );
  AND U15437 ( .A(n36), .B(n11579), .Z(n11577) );
  XOR U15438 ( .A(n11580), .B(n11581), .Z(n11579) );
  XOR U15439 ( .A(DB[3689]), .B(DB[3658]), .Z(n11581) );
  AND U15440 ( .A(n40), .B(n11582), .Z(n11580) );
  XOR U15441 ( .A(n11583), .B(n11584), .Z(n11582) );
  XOR U15442 ( .A(DB[3658]), .B(DB[3627]), .Z(n11584) );
  AND U15443 ( .A(n44), .B(n11585), .Z(n11583) );
  XOR U15444 ( .A(n11586), .B(n11587), .Z(n11585) );
  XOR U15445 ( .A(DB[3627]), .B(DB[3596]), .Z(n11587) );
  AND U15446 ( .A(n48), .B(n11588), .Z(n11586) );
  XOR U15447 ( .A(n11589), .B(n11590), .Z(n11588) );
  XOR U15448 ( .A(DB[3596]), .B(DB[3565]), .Z(n11590) );
  AND U15449 ( .A(n52), .B(n11591), .Z(n11589) );
  XOR U15450 ( .A(n11592), .B(n11593), .Z(n11591) );
  XOR U15451 ( .A(DB[3565]), .B(DB[3534]), .Z(n11593) );
  AND U15452 ( .A(n56), .B(n11594), .Z(n11592) );
  XOR U15453 ( .A(n11595), .B(n11596), .Z(n11594) );
  XOR U15454 ( .A(DB[3534]), .B(DB[3503]), .Z(n11596) );
  AND U15455 ( .A(n60), .B(n11597), .Z(n11595) );
  XOR U15456 ( .A(n11598), .B(n11599), .Z(n11597) );
  XOR U15457 ( .A(DB[3503]), .B(DB[3472]), .Z(n11599) );
  AND U15458 ( .A(n64), .B(n11600), .Z(n11598) );
  XOR U15459 ( .A(n11601), .B(n11602), .Z(n11600) );
  XOR U15460 ( .A(DB[3472]), .B(DB[3441]), .Z(n11602) );
  AND U15461 ( .A(n68), .B(n11603), .Z(n11601) );
  XOR U15462 ( .A(n11604), .B(n11605), .Z(n11603) );
  XOR U15463 ( .A(DB[3441]), .B(DB[3410]), .Z(n11605) );
  AND U15464 ( .A(n72), .B(n11606), .Z(n11604) );
  XOR U15465 ( .A(n11607), .B(n11608), .Z(n11606) );
  XOR U15466 ( .A(DB[3410]), .B(DB[3379]), .Z(n11608) );
  AND U15467 ( .A(n76), .B(n11609), .Z(n11607) );
  XOR U15468 ( .A(n11610), .B(n11611), .Z(n11609) );
  XOR U15469 ( .A(DB[3379]), .B(DB[3348]), .Z(n11611) );
  AND U15470 ( .A(n80), .B(n11612), .Z(n11610) );
  XOR U15471 ( .A(n11613), .B(n11614), .Z(n11612) );
  XOR U15472 ( .A(DB[3348]), .B(DB[3317]), .Z(n11614) );
  AND U15473 ( .A(n84), .B(n11615), .Z(n11613) );
  XOR U15474 ( .A(n11616), .B(n11617), .Z(n11615) );
  XOR U15475 ( .A(DB[3317]), .B(DB[3286]), .Z(n11617) );
  AND U15476 ( .A(n88), .B(n11618), .Z(n11616) );
  XOR U15477 ( .A(n11619), .B(n11620), .Z(n11618) );
  XOR U15478 ( .A(DB[3286]), .B(DB[3255]), .Z(n11620) );
  AND U15479 ( .A(n92), .B(n11621), .Z(n11619) );
  XOR U15480 ( .A(n11622), .B(n11623), .Z(n11621) );
  XOR U15481 ( .A(DB[3255]), .B(DB[3224]), .Z(n11623) );
  AND U15482 ( .A(n96), .B(n11624), .Z(n11622) );
  XOR U15483 ( .A(n11625), .B(n11626), .Z(n11624) );
  XOR U15484 ( .A(DB[3224]), .B(DB[3193]), .Z(n11626) );
  AND U15485 ( .A(n100), .B(n11627), .Z(n11625) );
  XOR U15486 ( .A(n11628), .B(n11629), .Z(n11627) );
  XOR U15487 ( .A(DB[3193]), .B(DB[3162]), .Z(n11629) );
  AND U15488 ( .A(n104), .B(n11630), .Z(n11628) );
  XOR U15489 ( .A(n11631), .B(n11632), .Z(n11630) );
  XOR U15490 ( .A(DB[3162]), .B(DB[3131]), .Z(n11632) );
  AND U15491 ( .A(n108), .B(n11633), .Z(n11631) );
  XOR U15492 ( .A(n11634), .B(n11635), .Z(n11633) );
  XOR U15493 ( .A(DB[3131]), .B(DB[3100]), .Z(n11635) );
  AND U15494 ( .A(n112), .B(n11636), .Z(n11634) );
  XOR U15495 ( .A(n11637), .B(n11638), .Z(n11636) );
  XOR U15496 ( .A(DB[3100]), .B(DB[3069]), .Z(n11638) );
  AND U15497 ( .A(n116), .B(n11639), .Z(n11637) );
  XOR U15498 ( .A(n11640), .B(n11641), .Z(n11639) );
  XOR U15499 ( .A(DB[3069]), .B(DB[3038]), .Z(n11641) );
  AND U15500 ( .A(n120), .B(n11642), .Z(n11640) );
  XOR U15501 ( .A(n11643), .B(n11644), .Z(n11642) );
  XOR U15502 ( .A(DB[3038]), .B(DB[3007]), .Z(n11644) );
  AND U15503 ( .A(n124), .B(n11645), .Z(n11643) );
  XOR U15504 ( .A(n11646), .B(n11647), .Z(n11645) );
  XOR U15505 ( .A(DB[3007]), .B(DB[2976]), .Z(n11647) );
  AND U15506 ( .A(n128), .B(n11648), .Z(n11646) );
  XOR U15507 ( .A(n11649), .B(n11650), .Z(n11648) );
  XOR U15508 ( .A(DB[2976]), .B(DB[2945]), .Z(n11650) );
  AND U15509 ( .A(n132), .B(n11651), .Z(n11649) );
  XOR U15510 ( .A(n11652), .B(n11653), .Z(n11651) );
  XOR U15511 ( .A(DB[2945]), .B(DB[2914]), .Z(n11653) );
  AND U15512 ( .A(n136), .B(n11654), .Z(n11652) );
  XOR U15513 ( .A(n11655), .B(n11656), .Z(n11654) );
  XOR U15514 ( .A(DB[2914]), .B(DB[2883]), .Z(n11656) );
  AND U15515 ( .A(n140), .B(n11657), .Z(n11655) );
  XOR U15516 ( .A(n11658), .B(n11659), .Z(n11657) );
  XOR U15517 ( .A(DB[2883]), .B(DB[2852]), .Z(n11659) );
  AND U15518 ( .A(n144), .B(n11660), .Z(n11658) );
  XOR U15519 ( .A(n11661), .B(n11662), .Z(n11660) );
  XOR U15520 ( .A(DB[2852]), .B(DB[2821]), .Z(n11662) );
  AND U15521 ( .A(n148), .B(n11663), .Z(n11661) );
  XOR U15522 ( .A(n11664), .B(n11665), .Z(n11663) );
  XOR U15523 ( .A(DB[2821]), .B(DB[2790]), .Z(n11665) );
  AND U15524 ( .A(n152), .B(n11666), .Z(n11664) );
  XOR U15525 ( .A(n11667), .B(n11668), .Z(n11666) );
  XOR U15526 ( .A(DB[2790]), .B(DB[2759]), .Z(n11668) );
  AND U15527 ( .A(n156), .B(n11669), .Z(n11667) );
  XOR U15528 ( .A(n11670), .B(n11671), .Z(n11669) );
  XOR U15529 ( .A(DB[2759]), .B(DB[2728]), .Z(n11671) );
  AND U15530 ( .A(n160), .B(n11672), .Z(n11670) );
  XOR U15531 ( .A(n11673), .B(n11674), .Z(n11672) );
  XOR U15532 ( .A(DB[2728]), .B(DB[2697]), .Z(n11674) );
  AND U15533 ( .A(n164), .B(n11675), .Z(n11673) );
  XOR U15534 ( .A(n11676), .B(n11677), .Z(n11675) );
  XOR U15535 ( .A(DB[2697]), .B(DB[2666]), .Z(n11677) );
  AND U15536 ( .A(n168), .B(n11678), .Z(n11676) );
  XOR U15537 ( .A(n11679), .B(n11680), .Z(n11678) );
  XOR U15538 ( .A(DB[2666]), .B(DB[2635]), .Z(n11680) );
  AND U15539 ( .A(n172), .B(n11681), .Z(n11679) );
  XOR U15540 ( .A(n11682), .B(n11683), .Z(n11681) );
  XOR U15541 ( .A(DB[2635]), .B(DB[2604]), .Z(n11683) );
  AND U15542 ( .A(n176), .B(n11684), .Z(n11682) );
  XOR U15543 ( .A(n11685), .B(n11686), .Z(n11684) );
  XOR U15544 ( .A(DB[2604]), .B(DB[2573]), .Z(n11686) );
  AND U15545 ( .A(n180), .B(n11687), .Z(n11685) );
  XOR U15546 ( .A(n11688), .B(n11689), .Z(n11687) );
  XOR U15547 ( .A(DB[2573]), .B(DB[2542]), .Z(n11689) );
  AND U15548 ( .A(n184), .B(n11690), .Z(n11688) );
  XOR U15549 ( .A(n11691), .B(n11692), .Z(n11690) );
  XOR U15550 ( .A(DB[2542]), .B(DB[2511]), .Z(n11692) );
  AND U15551 ( .A(n188), .B(n11693), .Z(n11691) );
  XOR U15552 ( .A(n11694), .B(n11695), .Z(n11693) );
  XOR U15553 ( .A(DB[2511]), .B(DB[2480]), .Z(n11695) );
  AND U15554 ( .A(n192), .B(n11696), .Z(n11694) );
  XOR U15555 ( .A(n11697), .B(n11698), .Z(n11696) );
  XOR U15556 ( .A(DB[2480]), .B(DB[2449]), .Z(n11698) );
  AND U15557 ( .A(n196), .B(n11699), .Z(n11697) );
  XOR U15558 ( .A(n11700), .B(n11701), .Z(n11699) );
  XOR U15559 ( .A(DB[2449]), .B(DB[2418]), .Z(n11701) );
  AND U15560 ( .A(n200), .B(n11702), .Z(n11700) );
  XOR U15561 ( .A(n11703), .B(n11704), .Z(n11702) );
  XOR U15562 ( .A(DB[2418]), .B(DB[2387]), .Z(n11704) );
  AND U15563 ( .A(n204), .B(n11705), .Z(n11703) );
  XOR U15564 ( .A(n11706), .B(n11707), .Z(n11705) );
  XOR U15565 ( .A(DB[2387]), .B(DB[2356]), .Z(n11707) );
  AND U15566 ( .A(n208), .B(n11708), .Z(n11706) );
  XOR U15567 ( .A(n11709), .B(n11710), .Z(n11708) );
  XOR U15568 ( .A(DB[2356]), .B(DB[2325]), .Z(n11710) );
  AND U15569 ( .A(n212), .B(n11711), .Z(n11709) );
  XOR U15570 ( .A(n11712), .B(n11713), .Z(n11711) );
  XOR U15571 ( .A(DB[2325]), .B(DB[2294]), .Z(n11713) );
  AND U15572 ( .A(n216), .B(n11714), .Z(n11712) );
  XOR U15573 ( .A(n11715), .B(n11716), .Z(n11714) );
  XOR U15574 ( .A(DB[2294]), .B(DB[2263]), .Z(n11716) );
  AND U15575 ( .A(n220), .B(n11717), .Z(n11715) );
  XOR U15576 ( .A(n11718), .B(n11719), .Z(n11717) );
  XOR U15577 ( .A(DB[2263]), .B(DB[2232]), .Z(n11719) );
  AND U15578 ( .A(n224), .B(n11720), .Z(n11718) );
  XOR U15579 ( .A(n11721), .B(n11722), .Z(n11720) );
  XOR U15580 ( .A(DB[2232]), .B(DB[2201]), .Z(n11722) );
  AND U15581 ( .A(n228), .B(n11723), .Z(n11721) );
  XOR U15582 ( .A(n11724), .B(n11725), .Z(n11723) );
  XOR U15583 ( .A(DB[2201]), .B(DB[2170]), .Z(n11725) );
  AND U15584 ( .A(n232), .B(n11726), .Z(n11724) );
  XOR U15585 ( .A(n11727), .B(n11728), .Z(n11726) );
  XOR U15586 ( .A(DB[2170]), .B(DB[2139]), .Z(n11728) );
  AND U15587 ( .A(n236), .B(n11729), .Z(n11727) );
  XOR U15588 ( .A(n11730), .B(n11731), .Z(n11729) );
  XOR U15589 ( .A(DB[2139]), .B(DB[2108]), .Z(n11731) );
  AND U15590 ( .A(n240), .B(n11732), .Z(n11730) );
  XOR U15591 ( .A(n11733), .B(n11734), .Z(n11732) );
  XOR U15592 ( .A(DB[2108]), .B(DB[2077]), .Z(n11734) );
  AND U15593 ( .A(n244), .B(n11735), .Z(n11733) );
  XOR U15594 ( .A(n11736), .B(n11737), .Z(n11735) );
  XOR U15595 ( .A(DB[2077]), .B(DB[2046]), .Z(n11737) );
  AND U15596 ( .A(n248), .B(n11738), .Z(n11736) );
  XOR U15597 ( .A(n11739), .B(n11740), .Z(n11738) );
  XOR U15598 ( .A(DB[2046]), .B(DB[2015]), .Z(n11740) );
  AND U15599 ( .A(n252), .B(n11741), .Z(n11739) );
  XOR U15600 ( .A(n11742), .B(n11743), .Z(n11741) );
  XOR U15601 ( .A(DB[2015]), .B(DB[1984]), .Z(n11743) );
  AND U15602 ( .A(n256), .B(n11744), .Z(n11742) );
  XOR U15603 ( .A(n11745), .B(n11746), .Z(n11744) );
  XOR U15604 ( .A(DB[1984]), .B(DB[1953]), .Z(n11746) );
  AND U15605 ( .A(n260), .B(n11747), .Z(n11745) );
  XOR U15606 ( .A(n11748), .B(n11749), .Z(n11747) );
  XOR U15607 ( .A(DB[1953]), .B(DB[1922]), .Z(n11749) );
  AND U15608 ( .A(n264), .B(n11750), .Z(n11748) );
  XOR U15609 ( .A(n11751), .B(n11752), .Z(n11750) );
  XOR U15610 ( .A(DB[1922]), .B(DB[1891]), .Z(n11752) );
  AND U15611 ( .A(n268), .B(n11753), .Z(n11751) );
  XOR U15612 ( .A(n11754), .B(n11755), .Z(n11753) );
  XOR U15613 ( .A(DB[1891]), .B(DB[1860]), .Z(n11755) );
  AND U15614 ( .A(n272), .B(n11756), .Z(n11754) );
  XOR U15615 ( .A(n11757), .B(n11758), .Z(n11756) );
  XOR U15616 ( .A(DB[1860]), .B(DB[1829]), .Z(n11758) );
  AND U15617 ( .A(n276), .B(n11759), .Z(n11757) );
  XOR U15618 ( .A(n11760), .B(n11761), .Z(n11759) );
  XOR U15619 ( .A(DB[1829]), .B(DB[1798]), .Z(n11761) );
  AND U15620 ( .A(n280), .B(n11762), .Z(n11760) );
  XOR U15621 ( .A(n11763), .B(n11764), .Z(n11762) );
  XOR U15622 ( .A(DB[1798]), .B(DB[1767]), .Z(n11764) );
  AND U15623 ( .A(n284), .B(n11765), .Z(n11763) );
  XOR U15624 ( .A(n11766), .B(n11767), .Z(n11765) );
  XOR U15625 ( .A(DB[1767]), .B(DB[1736]), .Z(n11767) );
  AND U15626 ( .A(n288), .B(n11768), .Z(n11766) );
  XOR U15627 ( .A(n11769), .B(n11770), .Z(n11768) );
  XOR U15628 ( .A(DB[1736]), .B(DB[1705]), .Z(n11770) );
  AND U15629 ( .A(n292), .B(n11771), .Z(n11769) );
  XOR U15630 ( .A(n11772), .B(n11773), .Z(n11771) );
  XOR U15631 ( .A(DB[1705]), .B(DB[1674]), .Z(n11773) );
  AND U15632 ( .A(n296), .B(n11774), .Z(n11772) );
  XOR U15633 ( .A(n11775), .B(n11776), .Z(n11774) );
  XOR U15634 ( .A(DB[1674]), .B(DB[1643]), .Z(n11776) );
  AND U15635 ( .A(n300), .B(n11777), .Z(n11775) );
  XOR U15636 ( .A(n11778), .B(n11779), .Z(n11777) );
  XOR U15637 ( .A(DB[1643]), .B(DB[1612]), .Z(n11779) );
  AND U15638 ( .A(n304), .B(n11780), .Z(n11778) );
  XOR U15639 ( .A(n11781), .B(n11782), .Z(n11780) );
  XOR U15640 ( .A(DB[1612]), .B(DB[1581]), .Z(n11782) );
  AND U15641 ( .A(n308), .B(n11783), .Z(n11781) );
  XOR U15642 ( .A(n11784), .B(n11785), .Z(n11783) );
  XOR U15643 ( .A(DB[1581]), .B(DB[1550]), .Z(n11785) );
  AND U15644 ( .A(n312), .B(n11786), .Z(n11784) );
  XOR U15645 ( .A(n11787), .B(n11788), .Z(n11786) );
  XOR U15646 ( .A(DB[1550]), .B(DB[1519]), .Z(n11788) );
  AND U15647 ( .A(n316), .B(n11789), .Z(n11787) );
  XOR U15648 ( .A(n11790), .B(n11791), .Z(n11789) );
  XOR U15649 ( .A(DB[1519]), .B(DB[1488]), .Z(n11791) );
  AND U15650 ( .A(n320), .B(n11792), .Z(n11790) );
  XOR U15651 ( .A(n11793), .B(n11794), .Z(n11792) );
  XOR U15652 ( .A(DB[1488]), .B(DB[1457]), .Z(n11794) );
  AND U15653 ( .A(n324), .B(n11795), .Z(n11793) );
  XOR U15654 ( .A(n11796), .B(n11797), .Z(n11795) );
  XOR U15655 ( .A(DB[1457]), .B(DB[1426]), .Z(n11797) );
  AND U15656 ( .A(n328), .B(n11798), .Z(n11796) );
  XOR U15657 ( .A(n11799), .B(n11800), .Z(n11798) );
  XOR U15658 ( .A(DB[1426]), .B(DB[1395]), .Z(n11800) );
  AND U15659 ( .A(n332), .B(n11801), .Z(n11799) );
  XOR U15660 ( .A(n11802), .B(n11803), .Z(n11801) );
  XOR U15661 ( .A(DB[1395]), .B(DB[1364]), .Z(n11803) );
  AND U15662 ( .A(n336), .B(n11804), .Z(n11802) );
  XOR U15663 ( .A(n11805), .B(n11806), .Z(n11804) );
  XOR U15664 ( .A(DB[1364]), .B(DB[1333]), .Z(n11806) );
  AND U15665 ( .A(n340), .B(n11807), .Z(n11805) );
  XOR U15666 ( .A(n11808), .B(n11809), .Z(n11807) );
  XOR U15667 ( .A(DB[1333]), .B(DB[1302]), .Z(n11809) );
  AND U15668 ( .A(n344), .B(n11810), .Z(n11808) );
  XOR U15669 ( .A(n11811), .B(n11812), .Z(n11810) );
  XOR U15670 ( .A(DB[1302]), .B(DB[1271]), .Z(n11812) );
  AND U15671 ( .A(n348), .B(n11813), .Z(n11811) );
  XOR U15672 ( .A(n11814), .B(n11815), .Z(n11813) );
  XOR U15673 ( .A(DB[1271]), .B(DB[1240]), .Z(n11815) );
  AND U15674 ( .A(n352), .B(n11816), .Z(n11814) );
  XOR U15675 ( .A(n11817), .B(n11818), .Z(n11816) );
  XOR U15676 ( .A(DB[1240]), .B(DB[1209]), .Z(n11818) );
  AND U15677 ( .A(n356), .B(n11819), .Z(n11817) );
  XOR U15678 ( .A(n11820), .B(n11821), .Z(n11819) );
  XOR U15679 ( .A(DB[1209]), .B(DB[1178]), .Z(n11821) );
  AND U15680 ( .A(n360), .B(n11822), .Z(n11820) );
  XOR U15681 ( .A(n11823), .B(n11824), .Z(n11822) );
  XOR U15682 ( .A(DB[1178]), .B(DB[1147]), .Z(n11824) );
  AND U15683 ( .A(n364), .B(n11825), .Z(n11823) );
  XOR U15684 ( .A(n11826), .B(n11827), .Z(n11825) );
  XOR U15685 ( .A(DB[1147]), .B(DB[1116]), .Z(n11827) );
  AND U15686 ( .A(n368), .B(n11828), .Z(n11826) );
  XOR U15687 ( .A(n11829), .B(n11830), .Z(n11828) );
  XOR U15688 ( .A(DB[1116]), .B(DB[1085]), .Z(n11830) );
  AND U15689 ( .A(n372), .B(n11831), .Z(n11829) );
  XOR U15690 ( .A(n11832), .B(n11833), .Z(n11831) );
  XOR U15691 ( .A(DB[1085]), .B(DB[1054]), .Z(n11833) );
  AND U15692 ( .A(n376), .B(n11834), .Z(n11832) );
  XOR U15693 ( .A(n11835), .B(n11836), .Z(n11834) );
  XOR U15694 ( .A(DB[1054]), .B(DB[1023]), .Z(n11836) );
  AND U15695 ( .A(n380), .B(n11837), .Z(n11835) );
  XOR U15696 ( .A(n11838), .B(n11839), .Z(n11837) );
  XOR U15697 ( .A(DB[992]), .B(DB[1023]), .Z(n11839) );
  AND U15698 ( .A(n384), .B(n11840), .Z(n11838) );
  XOR U15699 ( .A(n11841), .B(n11842), .Z(n11840) );
  XOR U15700 ( .A(DB[992]), .B(DB[961]), .Z(n11842) );
  AND U15701 ( .A(n388), .B(n11843), .Z(n11841) );
  XOR U15702 ( .A(n11844), .B(n11845), .Z(n11843) );
  XOR U15703 ( .A(DB[961]), .B(DB[930]), .Z(n11845) );
  AND U15704 ( .A(n392), .B(n11846), .Z(n11844) );
  XOR U15705 ( .A(n11847), .B(n11848), .Z(n11846) );
  XOR U15706 ( .A(DB[930]), .B(DB[899]), .Z(n11848) );
  AND U15707 ( .A(n396), .B(n11849), .Z(n11847) );
  XOR U15708 ( .A(n11850), .B(n11851), .Z(n11849) );
  XOR U15709 ( .A(DB[899]), .B(DB[868]), .Z(n11851) );
  AND U15710 ( .A(n400), .B(n11852), .Z(n11850) );
  XOR U15711 ( .A(n11853), .B(n11854), .Z(n11852) );
  XOR U15712 ( .A(DB[868]), .B(DB[837]), .Z(n11854) );
  AND U15713 ( .A(n404), .B(n11855), .Z(n11853) );
  XOR U15714 ( .A(n11856), .B(n11857), .Z(n11855) );
  XOR U15715 ( .A(DB[837]), .B(DB[806]), .Z(n11857) );
  AND U15716 ( .A(n408), .B(n11858), .Z(n11856) );
  XOR U15717 ( .A(n11859), .B(n11860), .Z(n11858) );
  XOR U15718 ( .A(DB[806]), .B(DB[775]), .Z(n11860) );
  AND U15719 ( .A(n412), .B(n11861), .Z(n11859) );
  XOR U15720 ( .A(n11862), .B(n11863), .Z(n11861) );
  XOR U15721 ( .A(DB[775]), .B(DB[744]), .Z(n11863) );
  AND U15722 ( .A(n416), .B(n11864), .Z(n11862) );
  XOR U15723 ( .A(n11865), .B(n11866), .Z(n11864) );
  XOR U15724 ( .A(DB[744]), .B(DB[713]), .Z(n11866) );
  AND U15725 ( .A(n420), .B(n11867), .Z(n11865) );
  XOR U15726 ( .A(n11868), .B(n11869), .Z(n11867) );
  XOR U15727 ( .A(DB[713]), .B(DB[682]), .Z(n11869) );
  AND U15728 ( .A(n424), .B(n11870), .Z(n11868) );
  XOR U15729 ( .A(n11871), .B(n11872), .Z(n11870) );
  XOR U15730 ( .A(DB[682]), .B(DB[651]), .Z(n11872) );
  AND U15731 ( .A(n428), .B(n11873), .Z(n11871) );
  XOR U15732 ( .A(n11874), .B(n11875), .Z(n11873) );
  XOR U15733 ( .A(DB[651]), .B(DB[620]), .Z(n11875) );
  AND U15734 ( .A(n432), .B(n11876), .Z(n11874) );
  XOR U15735 ( .A(n11877), .B(n11878), .Z(n11876) );
  XOR U15736 ( .A(DB[620]), .B(DB[589]), .Z(n11878) );
  AND U15737 ( .A(n436), .B(n11879), .Z(n11877) );
  XOR U15738 ( .A(n11880), .B(n11881), .Z(n11879) );
  XOR U15739 ( .A(DB[589]), .B(DB[558]), .Z(n11881) );
  AND U15740 ( .A(n440), .B(n11882), .Z(n11880) );
  XOR U15741 ( .A(n11883), .B(n11884), .Z(n11882) );
  XOR U15742 ( .A(DB[558]), .B(DB[527]), .Z(n11884) );
  AND U15743 ( .A(n444), .B(n11885), .Z(n11883) );
  XOR U15744 ( .A(n11886), .B(n11887), .Z(n11885) );
  XOR U15745 ( .A(DB[527]), .B(DB[496]), .Z(n11887) );
  AND U15746 ( .A(n448), .B(n11888), .Z(n11886) );
  XOR U15747 ( .A(n11889), .B(n11890), .Z(n11888) );
  XOR U15748 ( .A(DB[496]), .B(DB[465]), .Z(n11890) );
  AND U15749 ( .A(n452), .B(n11891), .Z(n11889) );
  XOR U15750 ( .A(n11892), .B(n11893), .Z(n11891) );
  XOR U15751 ( .A(DB[465]), .B(DB[434]), .Z(n11893) );
  AND U15752 ( .A(n456), .B(n11894), .Z(n11892) );
  XOR U15753 ( .A(n11895), .B(n11896), .Z(n11894) );
  XOR U15754 ( .A(DB[434]), .B(DB[403]), .Z(n11896) );
  AND U15755 ( .A(n460), .B(n11897), .Z(n11895) );
  XOR U15756 ( .A(n11898), .B(n11899), .Z(n11897) );
  XOR U15757 ( .A(DB[403]), .B(DB[372]), .Z(n11899) );
  AND U15758 ( .A(n464), .B(n11900), .Z(n11898) );
  XOR U15759 ( .A(n11901), .B(n11902), .Z(n11900) );
  XOR U15760 ( .A(DB[372]), .B(DB[341]), .Z(n11902) );
  AND U15761 ( .A(n468), .B(n11903), .Z(n11901) );
  XOR U15762 ( .A(n11904), .B(n11905), .Z(n11903) );
  XOR U15763 ( .A(DB[341]), .B(DB[310]), .Z(n11905) );
  AND U15764 ( .A(n472), .B(n11906), .Z(n11904) );
  XOR U15765 ( .A(n11907), .B(n11908), .Z(n11906) );
  XOR U15766 ( .A(DB[310]), .B(DB[279]), .Z(n11908) );
  AND U15767 ( .A(n476), .B(n11909), .Z(n11907) );
  XOR U15768 ( .A(n11910), .B(n11911), .Z(n11909) );
  XOR U15769 ( .A(DB[279]), .B(DB[248]), .Z(n11911) );
  AND U15770 ( .A(n480), .B(n11912), .Z(n11910) );
  XOR U15771 ( .A(n11913), .B(n11914), .Z(n11912) );
  XOR U15772 ( .A(DB[248]), .B(DB[217]), .Z(n11914) );
  AND U15773 ( .A(n484), .B(n11915), .Z(n11913) );
  XOR U15774 ( .A(n11916), .B(n11917), .Z(n11915) );
  XOR U15775 ( .A(DB[217]), .B(DB[186]), .Z(n11917) );
  AND U15776 ( .A(n488), .B(n11918), .Z(n11916) );
  XOR U15777 ( .A(n11919), .B(n11920), .Z(n11918) );
  XOR U15778 ( .A(DB[186]), .B(DB[155]), .Z(n11920) );
  AND U15779 ( .A(n492), .B(n11921), .Z(n11919) );
  XOR U15780 ( .A(n11922), .B(n11923), .Z(n11921) );
  XOR U15781 ( .A(DB[155]), .B(DB[124]), .Z(n11923) );
  AND U15782 ( .A(n496), .B(n11924), .Z(n11922) );
  XOR U15783 ( .A(n11925), .B(n11926), .Z(n11924) );
  XOR U15784 ( .A(DB[93]), .B(DB[124]), .Z(n11926) );
  AND U15785 ( .A(n500), .B(n11927), .Z(n11925) );
  XOR U15786 ( .A(n11928), .B(n11929), .Z(n11927) );
  XOR U15787 ( .A(DB[93]), .B(DB[62]), .Z(n11929) );
  AND U15788 ( .A(n504), .B(n11930), .Z(n11928) );
  XOR U15789 ( .A(n11931), .B(n11932), .Z(n11930) );
  XOR U15790 ( .A(DB[62]), .B(DB[31]), .Z(n11932) );
  AND U15791 ( .A(n508), .B(n11933), .Z(n11931) );
  XOR U15792 ( .A(DB[31]), .B(DB[0]), .Z(n11933) );
  XNOR U15793 ( .A(n11934), .B(n11935), .Z(n2) );
  AND U15794 ( .A(n11936), .B(n11937), .Z(n11934) );
  XOR U15795 ( .A(n11935), .B(n11938), .Z(n11937) );
  XOR U15796 ( .A(n11939), .B(n11940), .Z(n11938) );
  AND U15797 ( .A(n11941), .B(n11942), .Z(n11939) );
  XNOR U15798 ( .A(n11943), .B(n11944), .Z(n11942) );
  XOR U15799 ( .A(n11935), .B(n11945), .Z(n11936) );
  XNOR U15800 ( .A(n11946), .B(n11947), .Z(n11945) );
  AND U15801 ( .A(n8), .B(n11948), .Z(n11946) );
  XOR U15802 ( .A(n11949), .B(n11947), .Z(n11948) );
  XOR U15803 ( .A(n11950), .B(n11951), .Z(n11935) );
  AND U15804 ( .A(n11952), .B(n11953), .Z(n11950) );
  XOR U15805 ( .A(n11941), .B(n11954), .Z(n11953) );
  XOR U15806 ( .A(n11951), .B(n11943), .Z(n11954) );
  XNOR U15807 ( .A(n11955), .B(n11956), .Z(n11943) );
  ANDN U15808 ( .B(n11957), .A(n11958), .Z(n11955) );
  XOR U15809 ( .A(n11956), .B(n11959), .Z(n11957) );
  XNOR U15810 ( .A(n11940), .B(n11960), .Z(n11941) );
  XNOR U15811 ( .A(n11961), .B(n11962), .Z(n11960) );
  ANDN U15812 ( .B(n11963), .A(n11964), .Z(n11961) );
  XNOR U15813 ( .A(n11965), .B(n11966), .Z(n11963) );
  IV U15814 ( .A(n11944), .Z(n11940) );
  XOR U15815 ( .A(n11967), .B(n11968), .Z(n11944) );
  AND U15816 ( .A(n11969), .B(n11970), .Z(n11967) );
  XOR U15817 ( .A(n11971), .B(n11968), .Z(n11970) );
  XOR U15818 ( .A(n11951), .B(n11972), .Z(n11952) );
  XOR U15819 ( .A(n11973), .B(n11974), .Z(n11972) );
  AND U15820 ( .A(n8), .B(n11975), .Z(n11973) );
  XNOR U15821 ( .A(n11976), .B(n11974), .Z(n11975) );
  XNOR U15822 ( .A(n11977), .B(n11978), .Z(n11951) );
  AND U15823 ( .A(n11979), .B(n11980), .Z(n11977) );
  XOR U15824 ( .A(n11969), .B(n11981), .Z(n11980) );
  XOR U15825 ( .A(n11978), .B(n11971), .Z(n11981) );
  XOR U15826 ( .A(n11982), .B(n11959), .Z(n11971) );
  XNOR U15827 ( .A(n11983), .B(n11984), .Z(n11959) );
  ANDN U15828 ( .B(n11985), .A(n11986), .Z(n11983) );
  XOR U15829 ( .A(n11987), .B(n11988), .Z(n11985) );
  IV U15830 ( .A(n11958), .Z(n11982) );
  XOR U15831 ( .A(n11989), .B(n11990), .Z(n11958) );
  XNOR U15832 ( .A(n11991), .B(n11992), .Z(n11990) );
  ANDN U15833 ( .B(n11993), .A(n11994), .Z(n11991) );
  XNOR U15834 ( .A(n11995), .B(n11996), .Z(n11993) );
  IV U15835 ( .A(n11956), .Z(n11989) );
  XOR U15836 ( .A(n11997), .B(n11998), .Z(n11956) );
  ANDN U15837 ( .B(n11999), .A(n12000), .Z(n11997) );
  XOR U15838 ( .A(n11998), .B(n12001), .Z(n11999) );
  XNOR U15839 ( .A(n12002), .B(n12003), .Z(n11969) );
  XNOR U15840 ( .A(n11965), .B(n12004), .Z(n12003) );
  IV U15841 ( .A(n11968), .Z(n12004) );
  XOR U15842 ( .A(n12005), .B(n12006), .Z(n11968) );
  AND U15843 ( .A(n12007), .B(n12008), .Z(n12005) );
  XOR U15844 ( .A(n12009), .B(n12006), .Z(n12008) );
  XNOR U15845 ( .A(n12010), .B(n12011), .Z(n11965) );
  ANDN U15846 ( .B(n12012), .A(n12013), .Z(n12010) );
  XOR U15847 ( .A(n12011), .B(n12014), .Z(n12012) );
  IV U15848 ( .A(n11964), .Z(n12002) );
  XOR U15849 ( .A(n11962), .B(n12015), .Z(n11964) );
  XNOR U15850 ( .A(n12016), .B(n12017), .Z(n12015) );
  ANDN U15851 ( .B(n12018), .A(n12019), .Z(n12016) );
  XNOR U15852 ( .A(n12020), .B(n12021), .Z(n12018) );
  IV U15853 ( .A(n11966), .Z(n11962) );
  XOR U15854 ( .A(n12022), .B(n12023), .Z(n11966) );
  ANDN U15855 ( .B(n12024), .A(n12025), .Z(n12022) );
  XOR U15856 ( .A(n12026), .B(n12023), .Z(n12024) );
  XNOR U15857 ( .A(n11978), .B(n12027), .Z(n11979) );
  XOR U15858 ( .A(n12028), .B(n12029), .Z(n12027) );
  AND U15859 ( .A(n8), .B(n12030), .Z(n12028) );
  XNOR U15860 ( .A(n12031), .B(n12029), .Z(n12030) );
  XNOR U15861 ( .A(n12032), .B(n12033), .Z(n11978) );
  NAND U15862 ( .A(n12034), .B(n12035), .Z(n12033) );
  XOR U15863 ( .A(n12007), .B(n12036), .Z(n12035) );
  XOR U15864 ( .A(n12032), .B(n12009), .Z(n12036) );
  XOR U15865 ( .A(n12037), .B(n12001), .Z(n12009) );
  XOR U15866 ( .A(n12038), .B(n11988), .Z(n12001) );
  XNOR U15867 ( .A(n12039), .B(n12040), .Z(n11988) );
  ANDN U15868 ( .B(n12041), .A(n12042), .Z(n12039) );
  XNOR U15869 ( .A(n12040), .B(n12043), .Z(n12041) );
  IV U15870 ( .A(n11986), .Z(n12038) );
  XOR U15871 ( .A(n11984), .B(n12044), .Z(n11986) );
  XNOR U15872 ( .A(n12045), .B(n12046), .Z(n12044) );
  ANDN U15873 ( .B(n12047), .A(n12048), .Z(n12045) );
  XNOR U15874 ( .A(n12049), .B(n12050), .Z(n12047) );
  IV U15875 ( .A(n12046), .Z(n12050) );
  IV U15876 ( .A(n11987), .Z(n11984) );
  XNOR U15877 ( .A(n12051), .B(n12052), .Z(n11987) );
  ANDN U15878 ( .B(n12053), .A(n12054), .Z(n12051) );
  XNOR U15879 ( .A(n12052), .B(n12055), .Z(n12053) );
  IV U15880 ( .A(n12000), .Z(n12037) );
  XOR U15881 ( .A(n12056), .B(n12057), .Z(n12000) );
  XNOR U15882 ( .A(n11995), .B(n12058), .Z(n12057) );
  IV U15883 ( .A(n11998), .Z(n12058) );
  XNOR U15884 ( .A(n12059), .B(n12060), .Z(n11998) );
  ANDN U15885 ( .B(n12061), .A(n12062), .Z(n12059) );
  XNOR U15886 ( .A(n12060), .B(n12063), .Z(n12061) );
  XOR U15887 ( .A(n12064), .B(n12065), .Z(n11995) );
  ANDN U15888 ( .B(n12066), .A(n12067), .Z(n12064) );
  XNOR U15889 ( .A(n12065), .B(n12068), .Z(n12066) );
  IV U15890 ( .A(n11994), .Z(n12056) );
  XOR U15891 ( .A(n11992), .B(n12069), .Z(n11994) );
  XNOR U15892 ( .A(n12070), .B(n12071), .Z(n12069) );
  ANDN U15893 ( .B(n12072), .A(n12073), .Z(n12070) );
  XNOR U15894 ( .A(n12074), .B(n12075), .Z(n12072) );
  IV U15895 ( .A(n12071), .Z(n12075) );
  IV U15896 ( .A(n11996), .Z(n11992) );
  XNOR U15897 ( .A(n12076), .B(n12077), .Z(n11996) );
  ANDN U15898 ( .B(n12078), .A(n12079), .Z(n12076) );
  XNOR U15899 ( .A(n12080), .B(n12077), .Z(n12078) );
  XNOR U15900 ( .A(n12081), .B(n12082), .Z(n12007) );
  XOR U15901 ( .A(n12026), .B(n12083), .Z(n12082) );
  IV U15902 ( .A(n12006), .Z(n12083) );
  XNOR U15903 ( .A(n12084), .B(n12085), .Z(n12006) );
  AND U15904 ( .A(n12086), .B(n12087), .Z(n12084) );
  XNOR U15905 ( .A(n12085), .B(n12088), .Z(n12087) );
  XOR U15906 ( .A(n12089), .B(n12014), .Z(n12026) );
  XNOR U15907 ( .A(n12090), .B(n12091), .Z(n12014) );
  ANDN U15908 ( .B(n12092), .A(n12093), .Z(n12090) );
  XNOR U15909 ( .A(n12091), .B(n12094), .Z(n12092) );
  IV U15910 ( .A(n12013), .Z(n12089) );
  XOR U15911 ( .A(n12095), .B(n12096), .Z(n12013) );
  XNOR U15912 ( .A(n12097), .B(n12098), .Z(n12096) );
  ANDN U15913 ( .B(n12099), .A(n12100), .Z(n12097) );
  XNOR U15914 ( .A(n12101), .B(n12102), .Z(n12099) );
  IV U15915 ( .A(n12098), .Z(n12102) );
  IV U15916 ( .A(n12011), .Z(n12095) );
  XNOR U15917 ( .A(n12103), .B(n12104), .Z(n12011) );
  ANDN U15918 ( .B(n12105), .A(n12106), .Z(n12103) );
  XNOR U15919 ( .A(n12104), .B(n12107), .Z(n12105) );
  IV U15920 ( .A(n12025), .Z(n12081) );
  XOR U15921 ( .A(n12108), .B(n12109), .Z(n12025) );
  XNOR U15922 ( .A(n12020), .B(n12110), .Z(n12109) );
  IV U15923 ( .A(n12023), .Z(n12110) );
  XNOR U15924 ( .A(n12111), .B(n12112), .Z(n12023) );
  ANDN U15925 ( .B(n12113), .A(n12114), .Z(n12111) );
  XNOR U15926 ( .A(n12115), .B(n12112), .Z(n12113) );
  XOR U15927 ( .A(n12116), .B(n12117), .Z(n12020) );
  ANDN U15928 ( .B(n12118), .A(n12119), .Z(n12116) );
  XNOR U15929 ( .A(n12117), .B(n12120), .Z(n12118) );
  IV U15930 ( .A(n12019), .Z(n12108) );
  XOR U15931 ( .A(n12017), .B(n12121), .Z(n12019) );
  XNOR U15932 ( .A(n12122), .B(n12123), .Z(n12121) );
  ANDN U15933 ( .B(n12124), .A(n12125), .Z(n12122) );
  XNOR U15934 ( .A(n12126), .B(n12127), .Z(n12124) );
  IV U15935 ( .A(n12123), .Z(n12127) );
  IV U15936 ( .A(n12021), .Z(n12017) );
  XNOR U15937 ( .A(n12128), .B(n12129), .Z(n12021) );
  ANDN U15938 ( .B(n12130), .A(n12131), .Z(n12128) );
  XNOR U15939 ( .A(n12132), .B(n12129), .Z(n12130) );
  XOR U15940 ( .A(n12133), .B(n12134), .Z(n12034) );
  XNOR U15941 ( .A(n12032), .B(n12135), .Z(n12134) );
  NAND U15942 ( .A(n12136), .B(n8), .Z(n12135) );
  XOR U15943 ( .A(n12137), .B(n12133), .Z(n12136) );
  NAND U15944 ( .A(n12138), .B(n12139), .Z(n12032) );
  XNOR U15945 ( .A(n12086), .B(n12088), .Z(n12139) );
  XOR U15946 ( .A(n12140), .B(n12063), .Z(n12088) );
  XOR U15947 ( .A(n12141), .B(n12055), .Z(n12063) );
  XOR U15948 ( .A(n12142), .B(n12043), .Z(n12055) );
  XNOR U15949 ( .A(q[30]), .B(DB[3967]), .Z(n12043) );
  IV U15950 ( .A(n12042), .Z(n12142) );
  XOR U15951 ( .A(n12040), .B(n12143), .Z(n12042) );
  XNOR U15952 ( .A(q[29]), .B(DB[3966]), .Z(n12143) );
  XOR U15953 ( .A(q[28]), .B(DB[3965]), .Z(n12040) );
  IV U15954 ( .A(n12054), .Z(n12141) );
  XOR U15955 ( .A(n12144), .B(n12145), .Z(n12054) );
  XNOR U15956 ( .A(n12049), .B(n12052), .Z(n12145) );
  XOR U15957 ( .A(q[24]), .B(DB[3961]), .Z(n12052) );
  XOR U15958 ( .A(q[27]), .B(DB[3964]), .Z(n12049) );
  IV U15959 ( .A(n12048), .Z(n12144) );
  XOR U15960 ( .A(n12046), .B(n12146), .Z(n12048) );
  XNOR U15961 ( .A(q[26]), .B(DB[3963]), .Z(n12146) );
  XOR U15962 ( .A(q[25]), .B(DB[3962]), .Z(n12046) );
  IV U15963 ( .A(n12062), .Z(n12140) );
  XOR U15964 ( .A(n12147), .B(n12148), .Z(n12062) );
  XOR U15965 ( .A(n12080), .B(n12060), .Z(n12148) );
  XOR U15966 ( .A(q[16]), .B(DB[3953]), .Z(n12060) );
  XOR U15967 ( .A(n12149), .B(n12068), .Z(n12080) );
  XNOR U15968 ( .A(q[23]), .B(DB[3960]), .Z(n12068) );
  IV U15969 ( .A(n12067), .Z(n12149) );
  XOR U15970 ( .A(n12065), .B(n12150), .Z(n12067) );
  XNOR U15971 ( .A(q[22]), .B(DB[3959]), .Z(n12150) );
  XOR U15972 ( .A(q[21]), .B(DB[3958]), .Z(n12065) );
  IV U15973 ( .A(n12079), .Z(n12147) );
  XOR U15974 ( .A(n12151), .B(n12152), .Z(n12079) );
  XNOR U15975 ( .A(n12074), .B(n12077), .Z(n12152) );
  XOR U15976 ( .A(q[17]), .B(DB[3954]), .Z(n12077) );
  XOR U15977 ( .A(q[20]), .B(DB[3957]), .Z(n12074) );
  IV U15978 ( .A(n12073), .Z(n12151) );
  XOR U15979 ( .A(n12071), .B(n12153), .Z(n12073) );
  XNOR U15980 ( .A(q[19]), .B(DB[3956]), .Z(n12153) );
  XOR U15981 ( .A(q[18]), .B(DB[3955]), .Z(n12071) );
  XNOR U15982 ( .A(n12154), .B(n12155), .Z(n12086) );
  XOR U15983 ( .A(n12115), .B(n12085), .Z(n12155) );
  XOR U15984 ( .A(q[0]), .B(DB[3937]), .Z(n12085) );
  XOR U15985 ( .A(n12156), .B(n12107), .Z(n12115) );
  XOR U15986 ( .A(n12157), .B(n12094), .Z(n12107) );
  XNOR U15987 ( .A(q[15]), .B(DB[3952]), .Z(n12094) );
  IV U15988 ( .A(n12093), .Z(n12157) );
  XOR U15989 ( .A(n12091), .B(n12158), .Z(n12093) );
  XNOR U15990 ( .A(q[14]), .B(DB[3951]), .Z(n12158) );
  XOR U15991 ( .A(q[13]), .B(DB[3950]), .Z(n12091) );
  IV U15992 ( .A(n12106), .Z(n12156) );
  XOR U15993 ( .A(n12159), .B(n12160), .Z(n12106) );
  XNOR U15994 ( .A(n12101), .B(n12104), .Z(n12160) );
  XOR U15995 ( .A(q[9]), .B(DB[3946]), .Z(n12104) );
  XOR U15996 ( .A(q[12]), .B(DB[3949]), .Z(n12101) );
  IV U15997 ( .A(n12100), .Z(n12159) );
  XOR U15998 ( .A(n12098), .B(n12161), .Z(n12100) );
  XNOR U15999 ( .A(q[11]), .B(DB[3948]), .Z(n12161) );
  XOR U16000 ( .A(q[10]), .B(DB[3947]), .Z(n12098) );
  IV U16001 ( .A(n12114), .Z(n12154) );
  XOR U16002 ( .A(n12162), .B(n12163), .Z(n12114) );
  XOR U16003 ( .A(n12132), .B(n12112), .Z(n12163) );
  XOR U16004 ( .A(q[1]), .B(DB[3938]), .Z(n12112) );
  XOR U16005 ( .A(n12164), .B(n12120), .Z(n12132) );
  XNOR U16006 ( .A(q[8]), .B(DB[3945]), .Z(n12120) );
  IV U16007 ( .A(n12119), .Z(n12164) );
  XOR U16008 ( .A(n12117), .B(n12165), .Z(n12119) );
  XNOR U16009 ( .A(q[7]), .B(DB[3944]), .Z(n12165) );
  XOR U16010 ( .A(q[6]), .B(DB[3943]), .Z(n12117) );
  IV U16011 ( .A(n12131), .Z(n12162) );
  XOR U16012 ( .A(n12166), .B(n12167), .Z(n12131) );
  XNOR U16013 ( .A(n12126), .B(n12129), .Z(n12167) );
  XOR U16014 ( .A(q[2]), .B(DB[3939]), .Z(n12129) );
  XOR U16015 ( .A(q[5]), .B(DB[3942]), .Z(n12126) );
  IV U16016 ( .A(n12125), .Z(n12166) );
  XOR U16017 ( .A(n12123), .B(n12168), .Z(n12125) );
  XNOR U16018 ( .A(q[4]), .B(DB[3941]), .Z(n12168) );
  XOR U16019 ( .A(q[3]), .B(DB[3940]), .Z(n12123) );
  XOR U16020 ( .A(n12169), .B(n12170), .Z(n12138) );
  AND U16021 ( .A(n8), .B(n12171), .Z(n12169) );
  XOR U16022 ( .A(n12170), .B(n12172), .Z(n12171) );
  XNOR U16023 ( .A(n12173), .B(n12174), .Z(n8) );
  AND U16024 ( .A(n12175), .B(n12176), .Z(n12173) );
  XOR U16025 ( .A(n12174), .B(n11947), .Z(n12176) );
  XNOR U16026 ( .A(n12177), .B(n12178), .Z(n11947) );
  ANDN U16027 ( .B(n12179), .A(n12180), .Z(n12177) );
  XOR U16028 ( .A(n12178), .B(n12181), .Z(n12179) );
  XNOR U16029 ( .A(n12174), .B(n11949), .Z(n12175) );
  XOR U16030 ( .A(n12182), .B(n12183), .Z(n11949) );
  AND U16031 ( .A(n12), .B(n12184), .Z(n12182) );
  XOR U16032 ( .A(n12185), .B(n12183), .Z(n12184) );
  XOR U16033 ( .A(n12186), .B(n12187), .Z(n12174) );
  AND U16034 ( .A(n12188), .B(n12189), .Z(n12186) );
  XNOR U16035 ( .A(n12187), .B(n11974), .Z(n12189) );
  XOR U16036 ( .A(n12190), .B(n12181), .Z(n11974) );
  XNOR U16037 ( .A(n12191), .B(n12192), .Z(n12181) );
  ANDN U16038 ( .B(n12193), .A(n12194), .Z(n12191) );
  XOR U16039 ( .A(n12195), .B(n12196), .Z(n12193) );
  IV U16040 ( .A(n12180), .Z(n12190) );
  XOR U16041 ( .A(n12197), .B(n12198), .Z(n12180) );
  XNOR U16042 ( .A(n12199), .B(n12200), .Z(n12198) );
  ANDN U16043 ( .B(n12201), .A(n12202), .Z(n12199) );
  XNOR U16044 ( .A(n12203), .B(n12204), .Z(n12201) );
  IV U16045 ( .A(n12178), .Z(n12197) );
  XOR U16046 ( .A(n12205), .B(n12206), .Z(n12178) );
  ANDN U16047 ( .B(n12207), .A(n12208), .Z(n12205) );
  XOR U16048 ( .A(n12206), .B(n12209), .Z(n12207) );
  XNOR U16049 ( .A(n12187), .B(n11976), .Z(n12188) );
  XOR U16050 ( .A(n12210), .B(n12211), .Z(n11976) );
  AND U16051 ( .A(n12), .B(n12212), .Z(n12210) );
  XOR U16052 ( .A(n12213), .B(n12211), .Z(n12212) );
  XNOR U16053 ( .A(n12214), .B(n12215), .Z(n12187) );
  AND U16054 ( .A(n12216), .B(n12217), .Z(n12214) );
  XOR U16055 ( .A(n12215), .B(n12029), .Z(n12217) );
  XOR U16056 ( .A(n12218), .B(n12209), .Z(n12029) );
  XOR U16057 ( .A(n12219), .B(n12196), .Z(n12209) );
  XNOR U16058 ( .A(n12220), .B(n12221), .Z(n12196) );
  ANDN U16059 ( .B(n12222), .A(n12223), .Z(n12220) );
  XOR U16060 ( .A(n12224), .B(n12225), .Z(n12222) );
  IV U16061 ( .A(n12194), .Z(n12219) );
  XOR U16062 ( .A(n12192), .B(n12226), .Z(n12194) );
  XNOR U16063 ( .A(n12227), .B(n12228), .Z(n12226) );
  ANDN U16064 ( .B(n12229), .A(n12230), .Z(n12227) );
  XNOR U16065 ( .A(n12231), .B(n12232), .Z(n12229) );
  IV U16066 ( .A(n12195), .Z(n12192) );
  XOR U16067 ( .A(n12233), .B(n12234), .Z(n12195) );
  ANDN U16068 ( .B(n12235), .A(n12236), .Z(n12233) );
  XOR U16069 ( .A(n12234), .B(n12237), .Z(n12235) );
  IV U16070 ( .A(n12208), .Z(n12218) );
  XOR U16071 ( .A(n12238), .B(n12239), .Z(n12208) );
  XNOR U16072 ( .A(n12203), .B(n12240), .Z(n12239) );
  IV U16073 ( .A(n12206), .Z(n12240) );
  XOR U16074 ( .A(n12241), .B(n12242), .Z(n12206) );
  ANDN U16075 ( .B(n12243), .A(n12244), .Z(n12241) );
  XOR U16076 ( .A(n12242), .B(n12245), .Z(n12243) );
  XNOR U16077 ( .A(n12246), .B(n12247), .Z(n12203) );
  ANDN U16078 ( .B(n12248), .A(n12249), .Z(n12246) );
  XOR U16079 ( .A(n12247), .B(n12250), .Z(n12248) );
  IV U16080 ( .A(n12202), .Z(n12238) );
  XOR U16081 ( .A(n12200), .B(n12251), .Z(n12202) );
  XNOR U16082 ( .A(n12252), .B(n12253), .Z(n12251) );
  ANDN U16083 ( .B(n12254), .A(n12255), .Z(n12252) );
  XNOR U16084 ( .A(n12256), .B(n12257), .Z(n12254) );
  IV U16085 ( .A(n12204), .Z(n12200) );
  XOR U16086 ( .A(n12258), .B(n12259), .Z(n12204) );
  ANDN U16087 ( .B(n12260), .A(n12261), .Z(n12258) );
  XOR U16088 ( .A(n12262), .B(n12259), .Z(n12260) );
  XOR U16089 ( .A(n12215), .B(n12031), .Z(n12216) );
  XOR U16090 ( .A(n12263), .B(n12264), .Z(n12031) );
  AND U16091 ( .A(n12), .B(n12265), .Z(n12263) );
  XOR U16092 ( .A(n12266), .B(n12264), .Z(n12265) );
  XNOR U16093 ( .A(n12267), .B(n12268), .Z(n12215) );
  NAND U16094 ( .A(n12269), .B(n12270), .Z(n12268) );
  XOR U16095 ( .A(n12271), .B(n12133), .Z(n12270) );
  XNOR U16096 ( .A(n12272), .B(n12245), .Z(n12133) );
  XOR U16097 ( .A(n12273), .B(n12237), .Z(n12245) );
  XOR U16098 ( .A(n12274), .B(n12225), .Z(n12237) );
  XOR U16099 ( .A(n12275), .B(n12276), .Z(n12225) );
  ANDN U16100 ( .B(n12277), .A(n12278), .Z(n12275) );
  XOR U16101 ( .A(n12276), .B(n12279), .Z(n12277) );
  IV U16102 ( .A(n12223), .Z(n12274) );
  XOR U16103 ( .A(n12221), .B(n12280), .Z(n12223) );
  XOR U16104 ( .A(n12281), .B(n12282), .Z(n12280) );
  ANDN U16105 ( .B(n12283), .A(n12284), .Z(n12281) );
  XOR U16106 ( .A(n12285), .B(n12282), .Z(n12283) );
  IV U16107 ( .A(n12224), .Z(n12221) );
  XOR U16108 ( .A(n12286), .B(n12287), .Z(n12224) );
  ANDN U16109 ( .B(n12288), .A(n12289), .Z(n12286) );
  XOR U16110 ( .A(n12287), .B(n12290), .Z(n12288) );
  IV U16111 ( .A(n12236), .Z(n12273) );
  XOR U16112 ( .A(n12291), .B(n12292), .Z(n12236) );
  XNOR U16113 ( .A(n12231), .B(n12293), .Z(n12292) );
  IV U16114 ( .A(n12234), .Z(n12293) );
  XOR U16115 ( .A(n12294), .B(n12295), .Z(n12234) );
  ANDN U16116 ( .B(n12296), .A(n12297), .Z(n12294) );
  XOR U16117 ( .A(n12295), .B(n12298), .Z(n12296) );
  XNOR U16118 ( .A(n12299), .B(n12300), .Z(n12231) );
  ANDN U16119 ( .B(n12301), .A(n12302), .Z(n12299) );
  XOR U16120 ( .A(n12300), .B(n12303), .Z(n12301) );
  IV U16121 ( .A(n12230), .Z(n12291) );
  XOR U16122 ( .A(n12228), .B(n12304), .Z(n12230) );
  XOR U16123 ( .A(n12305), .B(n12306), .Z(n12304) );
  ANDN U16124 ( .B(n12307), .A(n12308), .Z(n12305) );
  XOR U16125 ( .A(n12309), .B(n12306), .Z(n12307) );
  IV U16126 ( .A(n12232), .Z(n12228) );
  XOR U16127 ( .A(n12310), .B(n12311), .Z(n12232) );
  ANDN U16128 ( .B(n12312), .A(n12313), .Z(n12310) );
  XOR U16129 ( .A(n12314), .B(n12311), .Z(n12312) );
  IV U16130 ( .A(n12244), .Z(n12272) );
  XOR U16131 ( .A(n12315), .B(n12316), .Z(n12244) );
  XOR U16132 ( .A(n12262), .B(n12317), .Z(n12316) );
  IV U16133 ( .A(n12242), .Z(n12317) );
  XOR U16134 ( .A(n12318), .B(n12319), .Z(n12242) );
  ANDN U16135 ( .B(n12320), .A(n12321), .Z(n12318) );
  XOR U16136 ( .A(n12319), .B(n12322), .Z(n12320) );
  XOR U16137 ( .A(n12323), .B(n12250), .Z(n12262) );
  XOR U16138 ( .A(n12324), .B(n12325), .Z(n12250) );
  ANDN U16139 ( .B(n12326), .A(n12327), .Z(n12324) );
  XOR U16140 ( .A(n12325), .B(n12328), .Z(n12326) );
  IV U16141 ( .A(n12249), .Z(n12323) );
  XOR U16142 ( .A(n12329), .B(n12330), .Z(n12249) );
  XOR U16143 ( .A(n12331), .B(n12332), .Z(n12330) );
  ANDN U16144 ( .B(n12333), .A(n12334), .Z(n12331) );
  XOR U16145 ( .A(n12335), .B(n12332), .Z(n12333) );
  IV U16146 ( .A(n12247), .Z(n12329) );
  XOR U16147 ( .A(n12336), .B(n12337), .Z(n12247) );
  ANDN U16148 ( .B(n12338), .A(n12339), .Z(n12336) );
  XOR U16149 ( .A(n12337), .B(n12340), .Z(n12338) );
  IV U16150 ( .A(n12261), .Z(n12315) );
  XOR U16151 ( .A(n12341), .B(n12342), .Z(n12261) );
  XNOR U16152 ( .A(n12256), .B(n12343), .Z(n12342) );
  IV U16153 ( .A(n12259), .Z(n12343) );
  XOR U16154 ( .A(n12344), .B(n12345), .Z(n12259) );
  ANDN U16155 ( .B(n12346), .A(n12347), .Z(n12344) );
  XOR U16156 ( .A(n12348), .B(n12345), .Z(n12346) );
  XNOR U16157 ( .A(n12349), .B(n12350), .Z(n12256) );
  ANDN U16158 ( .B(n12351), .A(n12352), .Z(n12349) );
  XOR U16159 ( .A(n12350), .B(n12353), .Z(n12351) );
  IV U16160 ( .A(n12255), .Z(n12341) );
  XOR U16161 ( .A(n12253), .B(n12354), .Z(n12255) );
  XOR U16162 ( .A(n12355), .B(n12356), .Z(n12354) );
  ANDN U16163 ( .B(n12357), .A(n12358), .Z(n12355) );
  XOR U16164 ( .A(n12359), .B(n12356), .Z(n12357) );
  IV U16165 ( .A(n12257), .Z(n12253) );
  XOR U16166 ( .A(n12360), .B(n12361), .Z(n12257) );
  ANDN U16167 ( .B(n12362), .A(n12363), .Z(n12360) );
  XOR U16168 ( .A(n12364), .B(n12361), .Z(n12362) );
  IV U16169 ( .A(n12267), .Z(n12271) );
  XOR U16170 ( .A(n12267), .B(n12137), .Z(n12269) );
  XOR U16171 ( .A(n12365), .B(n12366), .Z(n12137) );
  AND U16172 ( .A(n12), .B(n12367), .Z(n12365) );
  XOR U16173 ( .A(n12368), .B(n12366), .Z(n12367) );
  NANDN U16174 ( .A(n12170), .B(n12172), .Z(n12267) );
  XOR U16175 ( .A(n12369), .B(n12370), .Z(n12172) );
  AND U16176 ( .A(n12), .B(n12371), .Z(n12369) );
  XOR U16177 ( .A(n12370), .B(n12372), .Z(n12371) );
  XNOR U16178 ( .A(n12373), .B(n12374), .Z(n12) );
  AND U16179 ( .A(n12375), .B(n12376), .Z(n12373) );
  XOR U16180 ( .A(n12374), .B(n12183), .Z(n12376) );
  XNOR U16181 ( .A(n12377), .B(n12378), .Z(n12183) );
  ANDN U16182 ( .B(n12379), .A(n12380), .Z(n12377) );
  XOR U16183 ( .A(n12378), .B(n12381), .Z(n12379) );
  XNOR U16184 ( .A(n12374), .B(n12185), .Z(n12375) );
  XOR U16185 ( .A(n12382), .B(n12383), .Z(n12185) );
  AND U16186 ( .A(n16), .B(n12384), .Z(n12382) );
  XOR U16187 ( .A(n12385), .B(n12383), .Z(n12384) );
  XOR U16188 ( .A(n12386), .B(n12387), .Z(n12374) );
  AND U16189 ( .A(n12388), .B(n12389), .Z(n12386) );
  XOR U16190 ( .A(n12387), .B(n12211), .Z(n12389) );
  XOR U16191 ( .A(n12380), .B(n12381), .Z(n12211) );
  XNOR U16192 ( .A(n12390), .B(n12391), .Z(n12381) );
  ANDN U16193 ( .B(n12392), .A(n12393), .Z(n12390) );
  XOR U16194 ( .A(n12394), .B(n12395), .Z(n12392) );
  XOR U16195 ( .A(n12396), .B(n12397), .Z(n12380) );
  XNOR U16196 ( .A(n12398), .B(n12399), .Z(n12397) );
  ANDN U16197 ( .B(n12400), .A(n12401), .Z(n12398) );
  XNOR U16198 ( .A(n12402), .B(n12403), .Z(n12400) );
  IV U16199 ( .A(n12378), .Z(n12396) );
  XOR U16200 ( .A(n12404), .B(n12405), .Z(n12378) );
  ANDN U16201 ( .B(n12406), .A(n12407), .Z(n12404) );
  XOR U16202 ( .A(n12405), .B(n12408), .Z(n12406) );
  XNOR U16203 ( .A(n12387), .B(n12213), .Z(n12388) );
  XOR U16204 ( .A(n12409), .B(n12410), .Z(n12213) );
  AND U16205 ( .A(n16), .B(n12411), .Z(n12409) );
  XOR U16206 ( .A(n12412), .B(n12410), .Z(n12411) );
  XNOR U16207 ( .A(n12413), .B(n12414), .Z(n12387) );
  AND U16208 ( .A(n12415), .B(n12416), .Z(n12413) );
  XNOR U16209 ( .A(n12414), .B(n12264), .Z(n12416) );
  XOR U16210 ( .A(n12407), .B(n12408), .Z(n12264) );
  XOR U16211 ( .A(n12417), .B(n12395), .Z(n12408) );
  XNOR U16212 ( .A(n12418), .B(n12419), .Z(n12395) );
  ANDN U16213 ( .B(n12420), .A(n12421), .Z(n12418) );
  XOR U16214 ( .A(n12422), .B(n12423), .Z(n12420) );
  IV U16215 ( .A(n12393), .Z(n12417) );
  XOR U16216 ( .A(n12391), .B(n12424), .Z(n12393) );
  XNOR U16217 ( .A(n12425), .B(n12426), .Z(n12424) );
  ANDN U16218 ( .B(n12427), .A(n12428), .Z(n12425) );
  XNOR U16219 ( .A(n12429), .B(n12430), .Z(n12427) );
  IV U16220 ( .A(n12394), .Z(n12391) );
  XOR U16221 ( .A(n12431), .B(n12432), .Z(n12394) );
  ANDN U16222 ( .B(n12433), .A(n12434), .Z(n12431) );
  XOR U16223 ( .A(n12432), .B(n12435), .Z(n12433) );
  XOR U16224 ( .A(n12436), .B(n12437), .Z(n12407) );
  XNOR U16225 ( .A(n12402), .B(n12438), .Z(n12437) );
  IV U16226 ( .A(n12405), .Z(n12438) );
  XOR U16227 ( .A(n12439), .B(n12440), .Z(n12405) );
  ANDN U16228 ( .B(n12441), .A(n12442), .Z(n12439) );
  XOR U16229 ( .A(n12440), .B(n12443), .Z(n12441) );
  XNOR U16230 ( .A(n12444), .B(n12445), .Z(n12402) );
  ANDN U16231 ( .B(n12446), .A(n12447), .Z(n12444) );
  XOR U16232 ( .A(n12445), .B(n12448), .Z(n12446) );
  IV U16233 ( .A(n12401), .Z(n12436) );
  XOR U16234 ( .A(n12399), .B(n12449), .Z(n12401) );
  XNOR U16235 ( .A(n12450), .B(n12451), .Z(n12449) );
  ANDN U16236 ( .B(n12452), .A(n12453), .Z(n12450) );
  XNOR U16237 ( .A(n12454), .B(n12455), .Z(n12452) );
  IV U16238 ( .A(n12403), .Z(n12399) );
  XOR U16239 ( .A(n12456), .B(n12457), .Z(n12403) );
  ANDN U16240 ( .B(n12458), .A(n12459), .Z(n12456) );
  XOR U16241 ( .A(n12460), .B(n12457), .Z(n12458) );
  XOR U16242 ( .A(n12414), .B(n12266), .Z(n12415) );
  XOR U16243 ( .A(n12461), .B(n12462), .Z(n12266) );
  AND U16244 ( .A(n16), .B(n12463), .Z(n12461) );
  XOR U16245 ( .A(n12464), .B(n12462), .Z(n12463) );
  XNOR U16246 ( .A(n12465), .B(n12466), .Z(n12414) );
  NAND U16247 ( .A(n12467), .B(n12468), .Z(n12466) );
  XOR U16248 ( .A(n12469), .B(n12366), .Z(n12468) );
  XOR U16249 ( .A(n12442), .B(n12443), .Z(n12366) );
  XOR U16250 ( .A(n12470), .B(n12435), .Z(n12443) );
  XOR U16251 ( .A(n12471), .B(n12423), .Z(n12435) );
  XOR U16252 ( .A(n12472), .B(n12473), .Z(n12423) );
  ANDN U16253 ( .B(n12474), .A(n12475), .Z(n12472) );
  XOR U16254 ( .A(n12473), .B(n12476), .Z(n12474) );
  IV U16255 ( .A(n12421), .Z(n12471) );
  XOR U16256 ( .A(n12419), .B(n12477), .Z(n12421) );
  XOR U16257 ( .A(n12478), .B(n12479), .Z(n12477) );
  ANDN U16258 ( .B(n12480), .A(n12481), .Z(n12478) );
  XOR U16259 ( .A(n12482), .B(n12479), .Z(n12480) );
  IV U16260 ( .A(n12422), .Z(n12419) );
  XOR U16261 ( .A(n12483), .B(n12484), .Z(n12422) );
  ANDN U16262 ( .B(n12485), .A(n12486), .Z(n12483) );
  XOR U16263 ( .A(n12484), .B(n12487), .Z(n12485) );
  IV U16264 ( .A(n12434), .Z(n12470) );
  XOR U16265 ( .A(n12488), .B(n12489), .Z(n12434) );
  XNOR U16266 ( .A(n12429), .B(n12490), .Z(n12489) );
  IV U16267 ( .A(n12432), .Z(n12490) );
  XOR U16268 ( .A(n12491), .B(n12492), .Z(n12432) );
  ANDN U16269 ( .B(n12493), .A(n12494), .Z(n12491) );
  XOR U16270 ( .A(n12492), .B(n12495), .Z(n12493) );
  XNOR U16271 ( .A(n12496), .B(n12497), .Z(n12429) );
  ANDN U16272 ( .B(n12498), .A(n12499), .Z(n12496) );
  XOR U16273 ( .A(n12497), .B(n12500), .Z(n12498) );
  IV U16274 ( .A(n12428), .Z(n12488) );
  XOR U16275 ( .A(n12426), .B(n12501), .Z(n12428) );
  XOR U16276 ( .A(n12502), .B(n12503), .Z(n12501) );
  ANDN U16277 ( .B(n12504), .A(n12505), .Z(n12502) );
  XOR U16278 ( .A(n12506), .B(n12503), .Z(n12504) );
  IV U16279 ( .A(n12430), .Z(n12426) );
  XOR U16280 ( .A(n12507), .B(n12508), .Z(n12430) );
  ANDN U16281 ( .B(n12509), .A(n12510), .Z(n12507) );
  XOR U16282 ( .A(n12511), .B(n12508), .Z(n12509) );
  XOR U16283 ( .A(n12512), .B(n12513), .Z(n12442) );
  XOR U16284 ( .A(n12460), .B(n12514), .Z(n12513) );
  IV U16285 ( .A(n12440), .Z(n12514) );
  XOR U16286 ( .A(n12515), .B(n12516), .Z(n12440) );
  ANDN U16287 ( .B(n12517), .A(n12518), .Z(n12515) );
  XOR U16288 ( .A(n12516), .B(n12519), .Z(n12517) );
  XOR U16289 ( .A(n12520), .B(n12448), .Z(n12460) );
  XOR U16290 ( .A(n12521), .B(n12522), .Z(n12448) );
  ANDN U16291 ( .B(n12523), .A(n12524), .Z(n12521) );
  XOR U16292 ( .A(n12522), .B(n12525), .Z(n12523) );
  IV U16293 ( .A(n12447), .Z(n12520) );
  XOR U16294 ( .A(n12526), .B(n12527), .Z(n12447) );
  XOR U16295 ( .A(n12528), .B(n12529), .Z(n12527) );
  ANDN U16296 ( .B(n12530), .A(n12531), .Z(n12528) );
  XOR U16297 ( .A(n12532), .B(n12529), .Z(n12530) );
  IV U16298 ( .A(n12445), .Z(n12526) );
  XOR U16299 ( .A(n12533), .B(n12534), .Z(n12445) );
  ANDN U16300 ( .B(n12535), .A(n12536), .Z(n12533) );
  XOR U16301 ( .A(n12534), .B(n12537), .Z(n12535) );
  IV U16302 ( .A(n12459), .Z(n12512) );
  XOR U16303 ( .A(n12538), .B(n12539), .Z(n12459) );
  XNOR U16304 ( .A(n12454), .B(n12540), .Z(n12539) );
  IV U16305 ( .A(n12457), .Z(n12540) );
  XOR U16306 ( .A(n12541), .B(n12542), .Z(n12457) );
  ANDN U16307 ( .B(n12543), .A(n12544), .Z(n12541) );
  XOR U16308 ( .A(n12545), .B(n12542), .Z(n12543) );
  XNOR U16309 ( .A(n12546), .B(n12547), .Z(n12454) );
  ANDN U16310 ( .B(n12548), .A(n12549), .Z(n12546) );
  XOR U16311 ( .A(n12547), .B(n12550), .Z(n12548) );
  IV U16312 ( .A(n12453), .Z(n12538) );
  XOR U16313 ( .A(n12451), .B(n12551), .Z(n12453) );
  XOR U16314 ( .A(n12552), .B(n12553), .Z(n12551) );
  ANDN U16315 ( .B(n12554), .A(n12555), .Z(n12552) );
  XOR U16316 ( .A(n12556), .B(n12553), .Z(n12554) );
  IV U16317 ( .A(n12455), .Z(n12451) );
  XOR U16318 ( .A(n12557), .B(n12558), .Z(n12455) );
  ANDN U16319 ( .B(n12559), .A(n12560), .Z(n12557) );
  XOR U16320 ( .A(n12561), .B(n12558), .Z(n12559) );
  IV U16321 ( .A(n12465), .Z(n12469) );
  XOR U16322 ( .A(n12465), .B(n12368), .Z(n12467) );
  XOR U16323 ( .A(n12562), .B(n12563), .Z(n12368) );
  AND U16324 ( .A(n16), .B(n12564), .Z(n12562) );
  XOR U16325 ( .A(n12565), .B(n12563), .Z(n12564) );
  NANDN U16326 ( .A(n12370), .B(n12372), .Z(n12465) );
  XOR U16327 ( .A(n12566), .B(n12567), .Z(n12372) );
  AND U16328 ( .A(n16), .B(n12568), .Z(n12566) );
  XOR U16329 ( .A(n12567), .B(n12569), .Z(n12568) );
  XNOR U16330 ( .A(n12570), .B(n12571), .Z(n16) );
  AND U16331 ( .A(n12572), .B(n12573), .Z(n12570) );
  XOR U16332 ( .A(n12571), .B(n12383), .Z(n12573) );
  XNOR U16333 ( .A(n12574), .B(n12575), .Z(n12383) );
  ANDN U16334 ( .B(n12576), .A(n12577), .Z(n12574) );
  XOR U16335 ( .A(n12575), .B(n12578), .Z(n12576) );
  XNOR U16336 ( .A(n12571), .B(n12385), .Z(n12572) );
  XOR U16337 ( .A(n12579), .B(n12580), .Z(n12385) );
  AND U16338 ( .A(n20), .B(n12581), .Z(n12579) );
  XOR U16339 ( .A(n12582), .B(n12580), .Z(n12581) );
  XOR U16340 ( .A(n12583), .B(n12584), .Z(n12571) );
  AND U16341 ( .A(n12585), .B(n12586), .Z(n12583) );
  XOR U16342 ( .A(n12584), .B(n12410), .Z(n12586) );
  XOR U16343 ( .A(n12577), .B(n12578), .Z(n12410) );
  XNOR U16344 ( .A(n12587), .B(n12588), .Z(n12578) );
  ANDN U16345 ( .B(n12589), .A(n12590), .Z(n12587) );
  XOR U16346 ( .A(n12591), .B(n12592), .Z(n12589) );
  XOR U16347 ( .A(n12593), .B(n12594), .Z(n12577) );
  XNOR U16348 ( .A(n12595), .B(n12596), .Z(n12594) );
  ANDN U16349 ( .B(n12597), .A(n12598), .Z(n12595) );
  XNOR U16350 ( .A(n12599), .B(n12600), .Z(n12597) );
  IV U16351 ( .A(n12575), .Z(n12593) );
  XOR U16352 ( .A(n12601), .B(n12602), .Z(n12575) );
  ANDN U16353 ( .B(n12603), .A(n12604), .Z(n12601) );
  XOR U16354 ( .A(n12602), .B(n12605), .Z(n12603) );
  XNOR U16355 ( .A(n12584), .B(n12412), .Z(n12585) );
  XOR U16356 ( .A(n12606), .B(n12607), .Z(n12412) );
  AND U16357 ( .A(n20), .B(n12608), .Z(n12606) );
  XOR U16358 ( .A(n12609), .B(n12607), .Z(n12608) );
  XNOR U16359 ( .A(n12610), .B(n12611), .Z(n12584) );
  AND U16360 ( .A(n12612), .B(n12613), .Z(n12610) );
  XNOR U16361 ( .A(n12611), .B(n12462), .Z(n12613) );
  XOR U16362 ( .A(n12604), .B(n12605), .Z(n12462) );
  XOR U16363 ( .A(n12614), .B(n12592), .Z(n12605) );
  XNOR U16364 ( .A(n12615), .B(n12616), .Z(n12592) );
  ANDN U16365 ( .B(n12617), .A(n12618), .Z(n12615) );
  XOR U16366 ( .A(n12619), .B(n12620), .Z(n12617) );
  IV U16367 ( .A(n12590), .Z(n12614) );
  XOR U16368 ( .A(n12588), .B(n12621), .Z(n12590) );
  XNOR U16369 ( .A(n12622), .B(n12623), .Z(n12621) );
  ANDN U16370 ( .B(n12624), .A(n12625), .Z(n12622) );
  XNOR U16371 ( .A(n12626), .B(n12627), .Z(n12624) );
  IV U16372 ( .A(n12591), .Z(n12588) );
  XOR U16373 ( .A(n12628), .B(n12629), .Z(n12591) );
  ANDN U16374 ( .B(n12630), .A(n12631), .Z(n12628) );
  XOR U16375 ( .A(n12629), .B(n12632), .Z(n12630) );
  XOR U16376 ( .A(n12633), .B(n12634), .Z(n12604) );
  XNOR U16377 ( .A(n12599), .B(n12635), .Z(n12634) );
  IV U16378 ( .A(n12602), .Z(n12635) );
  XOR U16379 ( .A(n12636), .B(n12637), .Z(n12602) );
  ANDN U16380 ( .B(n12638), .A(n12639), .Z(n12636) );
  XOR U16381 ( .A(n12637), .B(n12640), .Z(n12638) );
  XNOR U16382 ( .A(n12641), .B(n12642), .Z(n12599) );
  ANDN U16383 ( .B(n12643), .A(n12644), .Z(n12641) );
  XOR U16384 ( .A(n12642), .B(n12645), .Z(n12643) );
  IV U16385 ( .A(n12598), .Z(n12633) );
  XOR U16386 ( .A(n12596), .B(n12646), .Z(n12598) );
  XNOR U16387 ( .A(n12647), .B(n12648), .Z(n12646) );
  ANDN U16388 ( .B(n12649), .A(n12650), .Z(n12647) );
  XNOR U16389 ( .A(n12651), .B(n12652), .Z(n12649) );
  IV U16390 ( .A(n12600), .Z(n12596) );
  XOR U16391 ( .A(n12653), .B(n12654), .Z(n12600) );
  ANDN U16392 ( .B(n12655), .A(n12656), .Z(n12653) );
  XOR U16393 ( .A(n12657), .B(n12654), .Z(n12655) );
  XOR U16394 ( .A(n12611), .B(n12464), .Z(n12612) );
  XOR U16395 ( .A(n12658), .B(n12659), .Z(n12464) );
  AND U16396 ( .A(n20), .B(n12660), .Z(n12658) );
  XOR U16397 ( .A(n12661), .B(n12659), .Z(n12660) );
  XNOR U16398 ( .A(n12662), .B(n12663), .Z(n12611) );
  NAND U16399 ( .A(n12664), .B(n12665), .Z(n12663) );
  XOR U16400 ( .A(n12666), .B(n12563), .Z(n12665) );
  XOR U16401 ( .A(n12639), .B(n12640), .Z(n12563) );
  XOR U16402 ( .A(n12667), .B(n12632), .Z(n12640) );
  XOR U16403 ( .A(n12668), .B(n12620), .Z(n12632) );
  XOR U16404 ( .A(n12669), .B(n12670), .Z(n12620) );
  ANDN U16405 ( .B(n12671), .A(n12672), .Z(n12669) );
  XOR U16406 ( .A(n12670), .B(n12673), .Z(n12671) );
  IV U16407 ( .A(n12618), .Z(n12668) );
  XOR U16408 ( .A(n12616), .B(n12674), .Z(n12618) );
  XOR U16409 ( .A(n12675), .B(n12676), .Z(n12674) );
  ANDN U16410 ( .B(n12677), .A(n12678), .Z(n12675) );
  XOR U16411 ( .A(n12679), .B(n12676), .Z(n12677) );
  IV U16412 ( .A(n12619), .Z(n12616) );
  XOR U16413 ( .A(n12680), .B(n12681), .Z(n12619) );
  ANDN U16414 ( .B(n12682), .A(n12683), .Z(n12680) );
  XOR U16415 ( .A(n12681), .B(n12684), .Z(n12682) );
  IV U16416 ( .A(n12631), .Z(n12667) );
  XOR U16417 ( .A(n12685), .B(n12686), .Z(n12631) );
  XNOR U16418 ( .A(n12626), .B(n12687), .Z(n12686) );
  IV U16419 ( .A(n12629), .Z(n12687) );
  XOR U16420 ( .A(n12688), .B(n12689), .Z(n12629) );
  ANDN U16421 ( .B(n12690), .A(n12691), .Z(n12688) );
  XOR U16422 ( .A(n12689), .B(n12692), .Z(n12690) );
  XNOR U16423 ( .A(n12693), .B(n12694), .Z(n12626) );
  ANDN U16424 ( .B(n12695), .A(n12696), .Z(n12693) );
  XOR U16425 ( .A(n12694), .B(n12697), .Z(n12695) );
  IV U16426 ( .A(n12625), .Z(n12685) );
  XOR U16427 ( .A(n12623), .B(n12698), .Z(n12625) );
  XOR U16428 ( .A(n12699), .B(n12700), .Z(n12698) );
  ANDN U16429 ( .B(n12701), .A(n12702), .Z(n12699) );
  XOR U16430 ( .A(n12703), .B(n12700), .Z(n12701) );
  IV U16431 ( .A(n12627), .Z(n12623) );
  XOR U16432 ( .A(n12704), .B(n12705), .Z(n12627) );
  ANDN U16433 ( .B(n12706), .A(n12707), .Z(n12704) );
  XOR U16434 ( .A(n12708), .B(n12705), .Z(n12706) );
  XOR U16435 ( .A(n12709), .B(n12710), .Z(n12639) );
  XOR U16436 ( .A(n12657), .B(n12711), .Z(n12710) );
  IV U16437 ( .A(n12637), .Z(n12711) );
  XOR U16438 ( .A(n12712), .B(n12713), .Z(n12637) );
  ANDN U16439 ( .B(n12714), .A(n12715), .Z(n12712) );
  XOR U16440 ( .A(n12713), .B(n12716), .Z(n12714) );
  XOR U16441 ( .A(n12717), .B(n12645), .Z(n12657) );
  XOR U16442 ( .A(n12718), .B(n12719), .Z(n12645) );
  ANDN U16443 ( .B(n12720), .A(n12721), .Z(n12718) );
  XOR U16444 ( .A(n12719), .B(n12722), .Z(n12720) );
  IV U16445 ( .A(n12644), .Z(n12717) );
  XOR U16446 ( .A(n12723), .B(n12724), .Z(n12644) );
  XOR U16447 ( .A(n12725), .B(n12726), .Z(n12724) );
  ANDN U16448 ( .B(n12727), .A(n12728), .Z(n12725) );
  XOR U16449 ( .A(n12729), .B(n12726), .Z(n12727) );
  IV U16450 ( .A(n12642), .Z(n12723) );
  XOR U16451 ( .A(n12730), .B(n12731), .Z(n12642) );
  ANDN U16452 ( .B(n12732), .A(n12733), .Z(n12730) );
  XOR U16453 ( .A(n12731), .B(n12734), .Z(n12732) );
  IV U16454 ( .A(n12656), .Z(n12709) );
  XOR U16455 ( .A(n12735), .B(n12736), .Z(n12656) );
  XNOR U16456 ( .A(n12651), .B(n12737), .Z(n12736) );
  IV U16457 ( .A(n12654), .Z(n12737) );
  XOR U16458 ( .A(n12738), .B(n12739), .Z(n12654) );
  ANDN U16459 ( .B(n12740), .A(n12741), .Z(n12738) );
  XOR U16460 ( .A(n12742), .B(n12739), .Z(n12740) );
  XNOR U16461 ( .A(n12743), .B(n12744), .Z(n12651) );
  ANDN U16462 ( .B(n12745), .A(n12746), .Z(n12743) );
  XOR U16463 ( .A(n12744), .B(n12747), .Z(n12745) );
  IV U16464 ( .A(n12650), .Z(n12735) );
  XOR U16465 ( .A(n12648), .B(n12748), .Z(n12650) );
  XOR U16466 ( .A(n12749), .B(n12750), .Z(n12748) );
  ANDN U16467 ( .B(n12751), .A(n12752), .Z(n12749) );
  XOR U16468 ( .A(n12753), .B(n12750), .Z(n12751) );
  IV U16469 ( .A(n12652), .Z(n12648) );
  XOR U16470 ( .A(n12754), .B(n12755), .Z(n12652) );
  ANDN U16471 ( .B(n12756), .A(n12757), .Z(n12754) );
  XOR U16472 ( .A(n12758), .B(n12755), .Z(n12756) );
  IV U16473 ( .A(n12662), .Z(n12666) );
  XOR U16474 ( .A(n12662), .B(n12565), .Z(n12664) );
  XOR U16475 ( .A(n12759), .B(n12760), .Z(n12565) );
  AND U16476 ( .A(n20), .B(n12761), .Z(n12759) );
  XOR U16477 ( .A(n12762), .B(n12760), .Z(n12761) );
  NANDN U16478 ( .A(n12567), .B(n12569), .Z(n12662) );
  XOR U16479 ( .A(n12763), .B(n12764), .Z(n12569) );
  AND U16480 ( .A(n20), .B(n12765), .Z(n12763) );
  XOR U16481 ( .A(n12764), .B(n12766), .Z(n12765) );
  XNOR U16482 ( .A(n12767), .B(n12768), .Z(n20) );
  AND U16483 ( .A(n12769), .B(n12770), .Z(n12767) );
  XOR U16484 ( .A(n12768), .B(n12580), .Z(n12770) );
  XNOR U16485 ( .A(n12771), .B(n12772), .Z(n12580) );
  ANDN U16486 ( .B(n12773), .A(n12774), .Z(n12771) );
  XOR U16487 ( .A(n12772), .B(n12775), .Z(n12773) );
  XNOR U16488 ( .A(n12768), .B(n12582), .Z(n12769) );
  XOR U16489 ( .A(n12776), .B(n12777), .Z(n12582) );
  AND U16490 ( .A(n24), .B(n12778), .Z(n12776) );
  XOR U16491 ( .A(n12779), .B(n12777), .Z(n12778) );
  XOR U16492 ( .A(n12780), .B(n12781), .Z(n12768) );
  AND U16493 ( .A(n12782), .B(n12783), .Z(n12780) );
  XOR U16494 ( .A(n12781), .B(n12607), .Z(n12783) );
  XOR U16495 ( .A(n12774), .B(n12775), .Z(n12607) );
  XNOR U16496 ( .A(n12784), .B(n12785), .Z(n12775) );
  ANDN U16497 ( .B(n12786), .A(n12787), .Z(n12784) );
  XOR U16498 ( .A(n12788), .B(n12789), .Z(n12786) );
  XOR U16499 ( .A(n12790), .B(n12791), .Z(n12774) );
  XNOR U16500 ( .A(n12792), .B(n12793), .Z(n12791) );
  ANDN U16501 ( .B(n12794), .A(n12795), .Z(n12792) );
  XNOR U16502 ( .A(n12796), .B(n12797), .Z(n12794) );
  IV U16503 ( .A(n12772), .Z(n12790) );
  XOR U16504 ( .A(n12798), .B(n12799), .Z(n12772) );
  ANDN U16505 ( .B(n12800), .A(n12801), .Z(n12798) );
  XOR U16506 ( .A(n12799), .B(n12802), .Z(n12800) );
  XNOR U16507 ( .A(n12781), .B(n12609), .Z(n12782) );
  XOR U16508 ( .A(n12803), .B(n12804), .Z(n12609) );
  AND U16509 ( .A(n24), .B(n12805), .Z(n12803) );
  XOR U16510 ( .A(n12806), .B(n12804), .Z(n12805) );
  XNOR U16511 ( .A(n12807), .B(n12808), .Z(n12781) );
  AND U16512 ( .A(n12809), .B(n12810), .Z(n12807) );
  XNOR U16513 ( .A(n12808), .B(n12659), .Z(n12810) );
  XOR U16514 ( .A(n12801), .B(n12802), .Z(n12659) );
  XOR U16515 ( .A(n12811), .B(n12789), .Z(n12802) );
  XNOR U16516 ( .A(n12812), .B(n12813), .Z(n12789) );
  ANDN U16517 ( .B(n12814), .A(n12815), .Z(n12812) );
  XOR U16518 ( .A(n12816), .B(n12817), .Z(n12814) );
  IV U16519 ( .A(n12787), .Z(n12811) );
  XOR U16520 ( .A(n12785), .B(n12818), .Z(n12787) );
  XNOR U16521 ( .A(n12819), .B(n12820), .Z(n12818) );
  ANDN U16522 ( .B(n12821), .A(n12822), .Z(n12819) );
  XNOR U16523 ( .A(n12823), .B(n12824), .Z(n12821) );
  IV U16524 ( .A(n12788), .Z(n12785) );
  XOR U16525 ( .A(n12825), .B(n12826), .Z(n12788) );
  ANDN U16526 ( .B(n12827), .A(n12828), .Z(n12825) );
  XOR U16527 ( .A(n12826), .B(n12829), .Z(n12827) );
  XOR U16528 ( .A(n12830), .B(n12831), .Z(n12801) );
  XNOR U16529 ( .A(n12796), .B(n12832), .Z(n12831) );
  IV U16530 ( .A(n12799), .Z(n12832) );
  XOR U16531 ( .A(n12833), .B(n12834), .Z(n12799) );
  ANDN U16532 ( .B(n12835), .A(n12836), .Z(n12833) );
  XOR U16533 ( .A(n12834), .B(n12837), .Z(n12835) );
  XNOR U16534 ( .A(n12838), .B(n12839), .Z(n12796) );
  ANDN U16535 ( .B(n12840), .A(n12841), .Z(n12838) );
  XOR U16536 ( .A(n12839), .B(n12842), .Z(n12840) );
  IV U16537 ( .A(n12795), .Z(n12830) );
  XOR U16538 ( .A(n12793), .B(n12843), .Z(n12795) );
  XNOR U16539 ( .A(n12844), .B(n12845), .Z(n12843) );
  ANDN U16540 ( .B(n12846), .A(n12847), .Z(n12844) );
  XNOR U16541 ( .A(n12848), .B(n12849), .Z(n12846) );
  IV U16542 ( .A(n12797), .Z(n12793) );
  XOR U16543 ( .A(n12850), .B(n12851), .Z(n12797) );
  ANDN U16544 ( .B(n12852), .A(n12853), .Z(n12850) );
  XOR U16545 ( .A(n12854), .B(n12851), .Z(n12852) );
  XOR U16546 ( .A(n12808), .B(n12661), .Z(n12809) );
  XOR U16547 ( .A(n12855), .B(n12856), .Z(n12661) );
  AND U16548 ( .A(n24), .B(n12857), .Z(n12855) );
  XOR U16549 ( .A(n12858), .B(n12856), .Z(n12857) );
  XNOR U16550 ( .A(n12859), .B(n12860), .Z(n12808) );
  NAND U16551 ( .A(n12861), .B(n12862), .Z(n12860) );
  XOR U16552 ( .A(n12863), .B(n12760), .Z(n12862) );
  XOR U16553 ( .A(n12836), .B(n12837), .Z(n12760) );
  XOR U16554 ( .A(n12864), .B(n12829), .Z(n12837) );
  XOR U16555 ( .A(n12865), .B(n12817), .Z(n12829) );
  XOR U16556 ( .A(n12866), .B(n12867), .Z(n12817) );
  ANDN U16557 ( .B(n12868), .A(n12869), .Z(n12866) );
  XOR U16558 ( .A(n12867), .B(n12870), .Z(n12868) );
  IV U16559 ( .A(n12815), .Z(n12865) );
  XOR U16560 ( .A(n12813), .B(n12871), .Z(n12815) );
  XOR U16561 ( .A(n12872), .B(n12873), .Z(n12871) );
  ANDN U16562 ( .B(n12874), .A(n12875), .Z(n12872) );
  XOR U16563 ( .A(n12876), .B(n12873), .Z(n12874) );
  IV U16564 ( .A(n12816), .Z(n12813) );
  XOR U16565 ( .A(n12877), .B(n12878), .Z(n12816) );
  ANDN U16566 ( .B(n12879), .A(n12880), .Z(n12877) );
  XOR U16567 ( .A(n12878), .B(n12881), .Z(n12879) );
  IV U16568 ( .A(n12828), .Z(n12864) );
  XOR U16569 ( .A(n12882), .B(n12883), .Z(n12828) );
  XNOR U16570 ( .A(n12823), .B(n12884), .Z(n12883) );
  IV U16571 ( .A(n12826), .Z(n12884) );
  XOR U16572 ( .A(n12885), .B(n12886), .Z(n12826) );
  ANDN U16573 ( .B(n12887), .A(n12888), .Z(n12885) );
  XOR U16574 ( .A(n12886), .B(n12889), .Z(n12887) );
  XNOR U16575 ( .A(n12890), .B(n12891), .Z(n12823) );
  ANDN U16576 ( .B(n12892), .A(n12893), .Z(n12890) );
  XOR U16577 ( .A(n12891), .B(n12894), .Z(n12892) );
  IV U16578 ( .A(n12822), .Z(n12882) );
  XOR U16579 ( .A(n12820), .B(n12895), .Z(n12822) );
  XOR U16580 ( .A(n12896), .B(n12897), .Z(n12895) );
  ANDN U16581 ( .B(n12898), .A(n12899), .Z(n12896) );
  XOR U16582 ( .A(n12900), .B(n12897), .Z(n12898) );
  IV U16583 ( .A(n12824), .Z(n12820) );
  XOR U16584 ( .A(n12901), .B(n12902), .Z(n12824) );
  ANDN U16585 ( .B(n12903), .A(n12904), .Z(n12901) );
  XOR U16586 ( .A(n12905), .B(n12902), .Z(n12903) );
  XOR U16587 ( .A(n12906), .B(n12907), .Z(n12836) );
  XOR U16588 ( .A(n12854), .B(n12908), .Z(n12907) );
  IV U16589 ( .A(n12834), .Z(n12908) );
  XOR U16590 ( .A(n12909), .B(n12910), .Z(n12834) );
  ANDN U16591 ( .B(n12911), .A(n12912), .Z(n12909) );
  XOR U16592 ( .A(n12910), .B(n12913), .Z(n12911) );
  XOR U16593 ( .A(n12914), .B(n12842), .Z(n12854) );
  XOR U16594 ( .A(n12915), .B(n12916), .Z(n12842) );
  ANDN U16595 ( .B(n12917), .A(n12918), .Z(n12915) );
  XOR U16596 ( .A(n12916), .B(n12919), .Z(n12917) );
  IV U16597 ( .A(n12841), .Z(n12914) );
  XOR U16598 ( .A(n12920), .B(n12921), .Z(n12841) );
  XOR U16599 ( .A(n12922), .B(n12923), .Z(n12921) );
  ANDN U16600 ( .B(n12924), .A(n12925), .Z(n12922) );
  XOR U16601 ( .A(n12926), .B(n12923), .Z(n12924) );
  IV U16602 ( .A(n12839), .Z(n12920) );
  XOR U16603 ( .A(n12927), .B(n12928), .Z(n12839) );
  ANDN U16604 ( .B(n12929), .A(n12930), .Z(n12927) );
  XOR U16605 ( .A(n12928), .B(n12931), .Z(n12929) );
  IV U16606 ( .A(n12853), .Z(n12906) );
  XOR U16607 ( .A(n12932), .B(n12933), .Z(n12853) );
  XNOR U16608 ( .A(n12848), .B(n12934), .Z(n12933) );
  IV U16609 ( .A(n12851), .Z(n12934) );
  XOR U16610 ( .A(n12935), .B(n12936), .Z(n12851) );
  ANDN U16611 ( .B(n12937), .A(n12938), .Z(n12935) );
  XOR U16612 ( .A(n12939), .B(n12936), .Z(n12937) );
  XNOR U16613 ( .A(n12940), .B(n12941), .Z(n12848) );
  ANDN U16614 ( .B(n12942), .A(n12943), .Z(n12940) );
  XOR U16615 ( .A(n12941), .B(n12944), .Z(n12942) );
  IV U16616 ( .A(n12847), .Z(n12932) );
  XOR U16617 ( .A(n12845), .B(n12945), .Z(n12847) );
  XOR U16618 ( .A(n12946), .B(n12947), .Z(n12945) );
  ANDN U16619 ( .B(n12948), .A(n12949), .Z(n12946) );
  XOR U16620 ( .A(n12950), .B(n12947), .Z(n12948) );
  IV U16621 ( .A(n12849), .Z(n12845) );
  XOR U16622 ( .A(n12951), .B(n12952), .Z(n12849) );
  ANDN U16623 ( .B(n12953), .A(n12954), .Z(n12951) );
  XOR U16624 ( .A(n12955), .B(n12952), .Z(n12953) );
  IV U16625 ( .A(n12859), .Z(n12863) );
  XOR U16626 ( .A(n12859), .B(n12762), .Z(n12861) );
  XOR U16627 ( .A(n12956), .B(n12957), .Z(n12762) );
  AND U16628 ( .A(n24), .B(n12958), .Z(n12956) );
  XOR U16629 ( .A(n12959), .B(n12957), .Z(n12958) );
  NANDN U16630 ( .A(n12764), .B(n12766), .Z(n12859) );
  XOR U16631 ( .A(n12960), .B(n12961), .Z(n12766) );
  AND U16632 ( .A(n24), .B(n12962), .Z(n12960) );
  XOR U16633 ( .A(n12961), .B(n12963), .Z(n12962) );
  XNOR U16634 ( .A(n12964), .B(n12965), .Z(n24) );
  AND U16635 ( .A(n12966), .B(n12967), .Z(n12964) );
  XOR U16636 ( .A(n12965), .B(n12777), .Z(n12967) );
  XNOR U16637 ( .A(n12968), .B(n12969), .Z(n12777) );
  ANDN U16638 ( .B(n12970), .A(n12971), .Z(n12968) );
  XOR U16639 ( .A(n12969), .B(n12972), .Z(n12970) );
  XNOR U16640 ( .A(n12965), .B(n12779), .Z(n12966) );
  XOR U16641 ( .A(n12973), .B(n12974), .Z(n12779) );
  AND U16642 ( .A(n28), .B(n12975), .Z(n12973) );
  XOR U16643 ( .A(n12976), .B(n12974), .Z(n12975) );
  XOR U16644 ( .A(n12977), .B(n12978), .Z(n12965) );
  AND U16645 ( .A(n12979), .B(n12980), .Z(n12977) );
  XOR U16646 ( .A(n12978), .B(n12804), .Z(n12980) );
  XOR U16647 ( .A(n12971), .B(n12972), .Z(n12804) );
  XNOR U16648 ( .A(n12981), .B(n12982), .Z(n12972) );
  ANDN U16649 ( .B(n12983), .A(n12984), .Z(n12981) );
  XOR U16650 ( .A(n12985), .B(n12986), .Z(n12983) );
  XOR U16651 ( .A(n12987), .B(n12988), .Z(n12971) );
  XNOR U16652 ( .A(n12989), .B(n12990), .Z(n12988) );
  ANDN U16653 ( .B(n12991), .A(n12992), .Z(n12989) );
  XNOR U16654 ( .A(n12993), .B(n12994), .Z(n12991) );
  IV U16655 ( .A(n12969), .Z(n12987) );
  XOR U16656 ( .A(n12995), .B(n12996), .Z(n12969) );
  ANDN U16657 ( .B(n12997), .A(n12998), .Z(n12995) );
  XOR U16658 ( .A(n12996), .B(n12999), .Z(n12997) );
  XNOR U16659 ( .A(n12978), .B(n12806), .Z(n12979) );
  XOR U16660 ( .A(n13000), .B(n13001), .Z(n12806) );
  AND U16661 ( .A(n28), .B(n13002), .Z(n13000) );
  XOR U16662 ( .A(n13003), .B(n13001), .Z(n13002) );
  XNOR U16663 ( .A(n13004), .B(n13005), .Z(n12978) );
  AND U16664 ( .A(n13006), .B(n13007), .Z(n13004) );
  XNOR U16665 ( .A(n13005), .B(n12856), .Z(n13007) );
  XOR U16666 ( .A(n12998), .B(n12999), .Z(n12856) );
  XOR U16667 ( .A(n13008), .B(n12986), .Z(n12999) );
  XNOR U16668 ( .A(n13009), .B(n13010), .Z(n12986) );
  ANDN U16669 ( .B(n13011), .A(n13012), .Z(n13009) );
  XOR U16670 ( .A(n13013), .B(n13014), .Z(n13011) );
  IV U16671 ( .A(n12984), .Z(n13008) );
  XOR U16672 ( .A(n12982), .B(n13015), .Z(n12984) );
  XNOR U16673 ( .A(n13016), .B(n13017), .Z(n13015) );
  ANDN U16674 ( .B(n13018), .A(n13019), .Z(n13016) );
  XNOR U16675 ( .A(n13020), .B(n13021), .Z(n13018) );
  IV U16676 ( .A(n12985), .Z(n12982) );
  XOR U16677 ( .A(n13022), .B(n13023), .Z(n12985) );
  ANDN U16678 ( .B(n13024), .A(n13025), .Z(n13022) );
  XOR U16679 ( .A(n13023), .B(n13026), .Z(n13024) );
  XOR U16680 ( .A(n13027), .B(n13028), .Z(n12998) );
  XNOR U16681 ( .A(n12993), .B(n13029), .Z(n13028) );
  IV U16682 ( .A(n12996), .Z(n13029) );
  XOR U16683 ( .A(n13030), .B(n13031), .Z(n12996) );
  ANDN U16684 ( .B(n13032), .A(n13033), .Z(n13030) );
  XOR U16685 ( .A(n13031), .B(n13034), .Z(n13032) );
  XNOR U16686 ( .A(n13035), .B(n13036), .Z(n12993) );
  ANDN U16687 ( .B(n13037), .A(n13038), .Z(n13035) );
  XOR U16688 ( .A(n13036), .B(n13039), .Z(n13037) );
  IV U16689 ( .A(n12992), .Z(n13027) );
  XOR U16690 ( .A(n12990), .B(n13040), .Z(n12992) );
  XNOR U16691 ( .A(n13041), .B(n13042), .Z(n13040) );
  ANDN U16692 ( .B(n13043), .A(n13044), .Z(n13041) );
  XNOR U16693 ( .A(n13045), .B(n13046), .Z(n13043) );
  IV U16694 ( .A(n12994), .Z(n12990) );
  XOR U16695 ( .A(n13047), .B(n13048), .Z(n12994) );
  ANDN U16696 ( .B(n13049), .A(n13050), .Z(n13047) );
  XOR U16697 ( .A(n13051), .B(n13048), .Z(n13049) );
  XOR U16698 ( .A(n13005), .B(n12858), .Z(n13006) );
  XOR U16699 ( .A(n13052), .B(n13053), .Z(n12858) );
  AND U16700 ( .A(n28), .B(n13054), .Z(n13052) );
  XOR U16701 ( .A(n13055), .B(n13053), .Z(n13054) );
  XNOR U16702 ( .A(n13056), .B(n13057), .Z(n13005) );
  NAND U16703 ( .A(n13058), .B(n13059), .Z(n13057) );
  XOR U16704 ( .A(n13060), .B(n12957), .Z(n13059) );
  XOR U16705 ( .A(n13033), .B(n13034), .Z(n12957) );
  XOR U16706 ( .A(n13061), .B(n13026), .Z(n13034) );
  XOR U16707 ( .A(n13062), .B(n13014), .Z(n13026) );
  XOR U16708 ( .A(n13063), .B(n13064), .Z(n13014) );
  ANDN U16709 ( .B(n13065), .A(n13066), .Z(n13063) );
  XOR U16710 ( .A(n13064), .B(n13067), .Z(n13065) );
  IV U16711 ( .A(n13012), .Z(n13062) );
  XOR U16712 ( .A(n13010), .B(n13068), .Z(n13012) );
  XOR U16713 ( .A(n13069), .B(n13070), .Z(n13068) );
  ANDN U16714 ( .B(n13071), .A(n13072), .Z(n13069) );
  XOR U16715 ( .A(n13073), .B(n13070), .Z(n13071) );
  IV U16716 ( .A(n13013), .Z(n13010) );
  XOR U16717 ( .A(n13074), .B(n13075), .Z(n13013) );
  ANDN U16718 ( .B(n13076), .A(n13077), .Z(n13074) );
  XOR U16719 ( .A(n13075), .B(n13078), .Z(n13076) );
  IV U16720 ( .A(n13025), .Z(n13061) );
  XOR U16721 ( .A(n13079), .B(n13080), .Z(n13025) );
  XNOR U16722 ( .A(n13020), .B(n13081), .Z(n13080) );
  IV U16723 ( .A(n13023), .Z(n13081) );
  XOR U16724 ( .A(n13082), .B(n13083), .Z(n13023) );
  ANDN U16725 ( .B(n13084), .A(n13085), .Z(n13082) );
  XOR U16726 ( .A(n13083), .B(n13086), .Z(n13084) );
  XNOR U16727 ( .A(n13087), .B(n13088), .Z(n13020) );
  ANDN U16728 ( .B(n13089), .A(n13090), .Z(n13087) );
  XOR U16729 ( .A(n13088), .B(n13091), .Z(n13089) );
  IV U16730 ( .A(n13019), .Z(n13079) );
  XOR U16731 ( .A(n13017), .B(n13092), .Z(n13019) );
  XOR U16732 ( .A(n13093), .B(n13094), .Z(n13092) );
  ANDN U16733 ( .B(n13095), .A(n13096), .Z(n13093) );
  XOR U16734 ( .A(n13097), .B(n13094), .Z(n13095) );
  IV U16735 ( .A(n13021), .Z(n13017) );
  XOR U16736 ( .A(n13098), .B(n13099), .Z(n13021) );
  ANDN U16737 ( .B(n13100), .A(n13101), .Z(n13098) );
  XOR U16738 ( .A(n13102), .B(n13099), .Z(n13100) );
  XOR U16739 ( .A(n13103), .B(n13104), .Z(n13033) );
  XOR U16740 ( .A(n13051), .B(n13105), .Z(n13104) );
  IV U16741 ( .A(n13031), .Z(n13105) );
  XOR U16742 ( .A(n13106), .B(n13107), .Z(n13031) );
  ANDN U16743 ( .B(n13108), .A(n13109), .Z(n13106) );
  XOR U16744 ( .A(n13107), .B(n13110), .Z(n13108) );
  XOR U16745 ( .A(n13111), .B(n13039), .Z(n13051) );
  XOR U16746 ( .A(n13112), .B(n13113), .Z(n13039) );
  ANDN U16747 ( .B(n13114), .A(n13115), .Z(n13112) );
  XOR U16748 ( .A(n13113), .B(n13116), .Z(n13114) );
  IV U16749 ( .A(n13038), .Z(n13111) );
  XOR U16750 ( .A(n13117), .B(n13118), .Z(n13038) );
  XOR U16751 ( .A(n13119), .B(n13120), .Z(n13118) );
  ANDN U16752 ( .B(n13121), .A(n13122), .Z(n13119) );
  XOR U16753 ( .A(n13123), .B(n13120), .Z(n13121) );
  IV U16754 ( .A(n13036), .Z(n13117) );
  XOR U16755 ( .A(n13124), .B(n13125), .Z(n13036) );
  ANDN U16756 ( .B(n13126), .A(n13127), .Z(n13124) );
  XOR U16757 ( .A(n13125), .B(n13128), .Z(n13126) );
  IV U16758 ( .A(n13050), .Z(n13103) );
  XOR U16759 ( .A(n13129), .B(n13130), .Z(n13050) );
  XNOR U16760 ( .A(n13045), .B(n13131), .Z(n13130) );
  IV U16761 ( .A(n13048), .Z(n13131) );
  XOR U16762 ( .A(n13132), .B(n13133), .Z(n13048) );
  ANDN U16763 ( .B(n13134), .A(n13135), .Z(n13132) );
  XOR U16764 ( .A(n13136), .B(n13133), .Z(n13134) );
  XNOR U16765 ( .A(n13137), .B(n13138), .Z(n13045) );
  ANDN U16766 ( .B(n13139), .A(n13140), .Z(n13137) );
  XOR U16767 ( .A(n13138), .B(n13141), .Z(n13139) );
  IV U16768 ( .A(n13044), .Z(n13129) );
  XOR U16769 ( .A(n13042), .B(n13142), .Z(n13044) );
  XOR U16770 ( .A(n13143), .B(n13144), .Z(n13142) );
  ANDN U16771 ( .B(n13145), .A(n13146), .Z(n13143) );
  XOR U16772 ( .A(n13147), .B(n13144), .Z(n13145) );
  IV U16773 ( .A(n13046), .Z(n13042) );
  XOR U16774 ( .A(n13148), .B(n13149), .Z(n13046) );
  ANDN U16775 ( .B(n13150), .A(n13151), .Z(n13148) );
  XOR U16776 ( .A(n13152), .B(n13149), .Z(n13150) );
  IV U16777 ( .A(n13056), .Z(n13060) );
  XOR U16778 ( .A(n13056), .B(n12959), .Z(n13058) );
  XOR U16779 ( .A(n13153), .B(n13154), .Z(n12959) );
  AND U16780 ( .A(n28), .B(n13155), .Z(n13153) );
  XOR U16781 ( .A(n13156), .B(n13154), .Z(n13155) );
  NANDN U16782 ( .A(n12961), .B(n12963), .Z(n13056) );
  XOR U16783 ( .A(n13157), .B(n13158), .Z(n12963) );
  AND U16784 ( .A(n28), .B(n13159), .Z(n13157) );
  XOR U16785 ( .A(n13158), .B(n13160), .Z(n13159) );
  XNOR U16786 ( .A(n13161), .B(n13162), .Z(n28) );
  AND U16787 ( .A(n13163), .B(n13164), .Z(n13161) );
  XOR U16788 ( .A(n13162), .B(n12974), .Z(n13164) );
  XNOR U16789 ( .A(n13165), .B(n13166), .Z(n12974) );
  ANDN U16790 ( .B(n13167), .A(n13168), .Z(n13165) );
  XOR U16791 ( .A(n13166), .B(n13169), .Z(n13167) );
  XNOR U16792 ( .A(n13162), .B(n12976), .Z(n13163) );
  XOR U16793 ( .A(n13170), .B(n13171), .Z(n12976) );
  AND U16794 ( .A(n32), .B(n13172), .Z(n13170) );
  XOR U16795 ( .A(n13173), .B(n13171), .Z(n13172) );
  XOR U16796 ( .A(n13174), .B(n13175), .Z(n13162) );
  AND U16797 ( .A(n13176), .B(n13177), .Z(n13174) );
  XOR U16798 ( .A(n13175), .B(n13001), .Z(n13177) );
  XOR U16799 ( .A(n13168), .B(n13169), .Z(n13001) );
  XNOR U16800 ( .A(n13178), .B(n13179), .Z(n13169) );
  ANDN U16801 ( .B(n13180), .A(n13181), .Z(n13178) );
  XOR U16802 ( .A(n13182), .B(n13183), .Z(n13180) );
  XOR U16803 ( .A(n13184), .B(n13185), .Z(n13168) );
  XNOR U16804 ( .A(n13186), .B(n13187), .Z(n13185) );
  ANDN U16805 ( .B(n13188), .A(n13189), .Z(n13186) );
  XNOR U16806 ( .A(n13190), .B(n13191), .Z(n13188) );
  IV U16807 ( .A(n13166), .Z(n13184) );
  XOR U16808 ( .A(n13192), .B(n13193), .Z(n13166) );
  ANDN U16809 ( .B(n13194), .A(n13195), .Z(n13192) );
  XOR U16810 ( .A(n13193), .B(n13196), .Z(n13194) );
  XNOR U16811 ( .A(n13175), .B(n13003), .Z(n13176) );
  XOR U16812 ( .A(n13197), .B(n13198), .Z(n13003) );
  AND U16813 ( .A(n32), .B(n13199), .Z(n13197) );
  XOR U16814 ( .A(n13200), .B(n13198), .Z(n13199) );
  XNOR U16815 ( .A(n13201), .B(n13202), .Z(n13175) );
  AND U16816 ( .A(n13203), .B(n13204), .Z(n13201) );
  XNOR U16817 ( .A(n13202), .B(n13053), .Z(n13204) );
  XOR U16818 ( .A(n13195), .B(n13196), .Z(n13053) );
  XOR U16819 ( .A(n13205), .B(n13183), .Z(n13196) );
  XNOR U16820 ( .A(n13206), .B(n13207), .Z(n13183) );
  ANDN U16821 ( .B(n13208), .A(n13209), .Z(n13206) );
  XOR U16822 ( .A(n13210), .B(n13211), .Z(n13208) );
  IV U16823 ( .A(n13181), .Z(n13205) );
  XOR U16824 ( .A(n13179), .B(n13212), .Z(n13181) );
  XNOR U16825 ( .A(n13213), .B(n13214), .Z(n13212) );
  ANDN U16826 ( .B(n13215), .A(n13216), .Z(n13213) );
  XNOR U16827 ( .A(n13217), .B(n13218), .Z(n13215) );
  IV U16828 ( .A(n13182), .Z(n13179) );
  XOR U16829 ( .A(n13219), .B(n13220), .Z(n13182) );
  ANDN U16830 ( .B(n13221), .A(n13222), .Z(n13219) );
  XOR U16831 ( .A(n13220), .B(n13223), .Z(n13221) );
  XOR U16832 ( .A(n13224), .B(n13225), .Z(n13195) );
  XNOR U16833 ( .A(n13190), .B(n13226), .Z(n13225) );
  IV U16834 ( .A(n13193), .Z(n13226) );
  XOR U16835 ( .A(n13227), .B(n13228), .Z(n13193) );
  ANDN U16836 ( .B(n13229), .A(n13230), .Z(n13227) );
  XOR U16837 ( .A(n13228), .B(n13231), .Z(n13229) );
  XNOR U16838 ( .A(n13232), .B(n13233), .Z(n13190) );
  ANDN U16839 ( .B(n13234), .A(n13235), .Z(n13232) );
  XOR U16840 ( .A(n13233), .B(n13236), .Z(n13234) );
  IV U16841 ( .A(n13189), .Z(n13224) );
  XOR U16842 ( .A(n13187), .B(n13237), .Z(n13189) );
  XNOR U16843 ( .A(n13238), .B(n13239), .Z(n13237) );
  ANDN U16844 ( .B(n13240), .A(n13241), .Z(n13238) );
  XNOR U16845 ( .A(n13242), .B(n13243), .Z(n13240) );
  IV U16846 ( .A(n13191), .Z(n13187) );
  XOR U16847 ( .A(n13244), .B(n13245), .Z(n13191) );
  ANDN U16848 ( .B(n13246), .A(n13247), .Z(n13244) );
  XOR U16849 ( .A(n13248), .B(n13245), .Z(n13246) );
  XOR U16850 ( .A(n13202), .B(n13055), .Z(n13203) );
  XOR U16851 ( .A(n13249), .B(n13250), .Z(n13055) );
  AND U16852 ( .A(n32), .B(n13251), .Z(n13249) );
  XOR U16853 ( .A(n13252), .B(n13250), .Z(n13251) );
  XNOR U16854 ( .A(n13253), .B(n13254), .Z(n13202) );
  NAND U16855 ( .A(n13255), .B(n13256), .Z(n13254) );
  XOR U16856 ( .A(n13257), .B(n13154), .Z(n13256) );
  XOR U16857 ( .A(n13230), .B(n13231), .Z(n13154) );
  XOR U16858 ( .A(n13258), .B(n13223), .Z(n13231) );
  XOR U16859 ( .A(n13259), .B(n13211), .Z(n13223) );
  XOR U16860 ( .A(n13260), .B(n13261), .Z(n13211) );
  ANDN U16861 ( .B(n13262), .A(n13263), .Z(n13260) );
  XOR U16862 ( .A(n13261), .B(n13264), .Z(n13262) );
  IV U16863 ( .A(n13209), .Z(n13259) );
  XOR U16864 ( .A(n13207), .B(n13265), .Z(n13209) );
  XOR U16865 ( .A(n13266), .B(n13267), .Z(n13265) );
  ANDN U16866 ( .B(n13268), .A(n13269), .Z(n13266) );
  XOR U16867 ( .A(n13270), .B(n13267), .Z(n13268) );
  IV U16868 ( .A(n13210), .Z(n13207) );
  XOR U16869 ( .A(n13271), .B(n13272), .Z(n13210) );
  ANDN U16870 ( .B(n13273), .A(n13274), .Z(n13271) );
  XOR U16871 ( .A(n13272), .B(n13275), .Z(n13273) );
  IV U16872 ( .A(n13222), .Z(n13258) );
  XOR U16873 ( .A(n13276), .B(n13277), .Z(n13222) );
  XNOR U16874 ( .A(n13217), .B(n13278), .Z(n13277) );
  IV U16875 ( .A(n13220), .Z(n13278) );
  XOR U16876 ( .A(n13279), .B(n13280), .Z(n13220) );
  ANDN U16877 ( .B(n13281), .A(n13282), .Z(n13279) );
  XOR U16878 ( .A(n13280), .B(n13283), .Z(n13281) );
  XNOR U16879 ( .A(n13284), .B(n13285), .Z(n13217) );
  ANDN U16880 ( .B(n13286), .A(n13287), .Z(n13284) );
  XOR U16881 ( .A(n13285), .B(n13288), .Z(n13286) );
  IV U16882 ( .A(n13216), .Z(n13276) );
  XOR U16883 ( .A(n13214), .B(n13289), .Z(n13216) );
  XOR U16884 ( .A(n13290), .B(n13291), .Z(n13289) );
  ANDN U16885 ( .B(n13292), .A(n13293), .Z(n13290) );
  XOR U16886 ( .A(n13294), .B(n13291), .Z(n13292) );
  IV U16887 ( .A(n13218), .Z(n13214) );
  XOR U16888 ( .A(n13295), .B(n13296), .Z(n13218) );
  ANDN U16889 ( .B(n13297), .A(n13298), .Z(n13295) );
  XOR U16890 ( .A(n13299), .B(n13296), .Z(n13297) );
  XOR U16891 ( .A(n13300), .B(n13301), .Z(n13230) );
  XOR U16892 ( .A(n13248), .B(n13302), .Z(n13301) );
  IV U16893 ( .A(n13228), .Z(n13302) );
  XOR U16894 ( .A(n13303), .B(n13304), .Z(n13228) );
  ANDN U16895 ( .B(n13305), .A(n13306), .Z(n13303) );
  XOR U16896 ( .A(n13304), .B(n13307), .Z(n13305) );
  XOR U16897 ( .A(n13308), .B(n13236), .Z(n13248) );
  XOR U16898 ( .A(n13309), .B(n13310), .Z(n13236) );
  ANDN U16899 ( .B(n13311), .A(n13312), .Z(n13309) );
  XOR U16900 ( .A(n13310), .B(n13313), .Z(n13311) );
  IV U16901 ( .A(n13235), .Z(n13308) );
  XOR U16902 ( .A(n13314), .B(n13315), .Z(n13235) );
  XOR U16903 ( .A(n13316), .B(n13317), .Z(n13315) );
  ANDN U16904 ( .B(n13318), .A(n13319), .Z(n13316) );
  XOR U16905 ( .A(n13320), .B(n13317), .Z(n13318) );
  IV U16906 ( .A(n13233), .Z(n13314) );
  XOR U16907 ( .A(n13321), .B(n13322), .Z(n13233) );
  ANDN U16908 ( .B(n13323), .A(n13324), .Z(n13321) );
  XOR U16909 ( .A(n13322), .B(n13325), .Z(n13323) );
  IV U16910 ( .A(n13247), .Z(n13300) );
  XOR U16911 ( .A(n13326), .B(n13327), .Z(n13247) );
  XNOR U16912 ( .A(n13242), .B(n13328), .Z(n13327) );
  IV U16913 ( .A(n13245), .Z(n13328) );
  XOR U16914 ( .A(n13329), .B(n13330), .Z(n13245) );
  ANDN U16915 ( .B(n13331), .A(n13332), .Z(n13329) );
  XOR U16916 ( .A(n13333), .B(n13330), .Z(n13331) );
  XNOR U16917 ( .A(n13334), .B(n13335), .Z(n13242) );
  ANDN U16918 ( .B(n13336), .A(n13337), .Z(n13334) );
  XOR U16919 ( .A(n13335), .B(n13338), .Z(n13336) );
  IV U16920 ( .A(n13241), .Z(n13326) );
  XOR U16921 ( .A(n13239), .B(n13339), .Z(n13241) );
  XOR U16922 ( .A(n13340), .B(n13341), .Z(n13339) );
  ANDN U16923 ( .B(n13342), .A(n13343), .Z(n13340) );
  XOR U16924 ( .A(n13344), .B(n13341), .Z(n13342) );
  IV U16925 ( .A(n13243), .Z(n13239) );
  XOR U16926 ( .A(n13345), .B(n13346), .Z(n13243) );
  ANDN U16927 ( .B(n13347), .A(n13348), .Z(n13345) );
  XOR U16928 ( .A(n13349), .B(n13346), .Z(n13347) );
  IV U16929 ( .A(n13253), .Z(n13257) );
  XOR U16930 ( .A(n13253), .B(n13156), .Z(n13255) );
  XOR U16931 ( .A(n13350), .B(n13351), .Z(n13156) );
  AND U16932 ( .A(n32), .B(n13352), .Z(n13350) );
  XOR U16933 ( .A(n13353), .B(n13351), .Z(n13352) );
  NANDN U16934 ( .A(n13158), .B(n13160), .Z(n13253) );
  XOR U16935 ( .A(n13354), .B(n13355), .Z(n13160) );
  AND U16936 ( .A(n32), .B(n13356), .Z(n13354) );
  XOR U16937 ( .A(n13355), .B(n13357), .Z(n13356) );
  XNOR U16938 ( .A(n13358), .B(n13359), .Z(n32) );
  AND U16939 ( .A(n13360), .B(n13361), .Z(n13358) );
  XOR U16940 ( .A(n13359), .B(n13171), .Z(n13361) );
  XNOR U16941 ( .A(n13362), .B(n13363), .Z(n13171) );
  ANDN U16942 ( .B(n13364), .A(n13365), .Z(n13362) );
  XOR U16943 ( .A(n13363), .B(n13366), .Z(n13364) );
  XNOR U16944 ( .A(n13359), .B(n13173), .Z(n13360) );
  XOR U16945 ( .A(n13367), .B(n13368), .Z(n13173) );
  AND U16946 ( .A(n36), .B(n13369), .Z(n13367) );
  XOR U16947 ( .A(n13370), .B(n13368), .Z(n13369) );
  XOR U16948 ( .A(n13371), .B(n13372), .Z(n13359) );
  AND U16949 ( .A(n13373), .B(n13374), .Z(n13371) );
  XOR U16950 ( .A(n13372), .B(n13198), .Z(n13374) );
  XOR U16951 ( .A(n13365), .B(n13366), .Z(n13198) );
  XNOR U16952 ( .A(n13375), .B(n13376), .Z(n13366) );
  ANDN U16953 ( .B(n13377), .A(n13378), .Z(n13375) );
  XOR U16954 ( .A(n13379), .B(n13380), .Z(n13377) );
  XOR U16955 ( .A(n13381), .B(n13382), .Z(n13365) );
  XNOR U16956 ( .A(n13383), .B(n13384), .Z(n13382) );
  ANDN U16957 ( .B(n13385), .A(n13386), .Z(n13383) );
  XNOR U16958 ( .A(n13387), .B(n13388), .Z(n13385) );
  IV U16959 ( .A(n13363), .Z(n13381) );
  XOR U16960 ( .A(n13389), .B(n13390), .Z(n13363) );
  ANDN U16961 ( .B(n13391), .A(n13392), .Z(n13389) );
  XOR U16962 ( .A(n13390), .B(n13393), .Z(n13391) );
  XNOR U16963 ( .A(n13372), .B(n13200), .Z(n13373) );
  XOR U16964 ( .A(n13394), .B(n13395), .Z(n13200) );
  AND U16965 ( .A(n36), .B(n13396), .Z(n13394) );
  XOR U16966 ( .A(n13397), .B(n13395), .Z(n13396) );
  XNOR U16967 ( .A(n13398), .B(n13399), .Z(n13372) );
  AND U16968 ( .A(n13400), .B(n13401), .Z(n13398) );
  XNOR U16969 ( .A(n13399), .B(n13250), .Z(n13401) );
  XOR U16970 ( .A(n13392), .B(n13393), .Z(n13250) );
  XOR U16971 ( .A(n13402), .B(n13380), .Z(n13393) );
  XNOR U16972 ( .A(n13403), .B(n13404), .Z(n13380) );
  ANDN U16973 ( .B(n13405), .A(n13406), .Z(n13403) );
  XOR U16974 ( .A(n13407), .B(n13408), .Z(n13405) );
  IV U16975 ( .A(n13378), .Z(n13402) );
  XOR U16976 ( .A(n13376), .B(n13409), .Z(n13378) );
  XNOR U16977 ( .A(n13410), .B(n13411), .Z(n13409) );
  ANDN U16978 ( .B(n13412), .A(n13413), .Z(n13410) );
  XNOR U16979 ( .A(n13414), .B(n13415), .Z(n13412) );
  IV U16980 ( .A(n13379), .Z(n13376) );
  XOR U16981 ( .A(n13416), .B(n13417), .Z(n13379) );
  ANDN U16982 ( .B(n13418), .A(n13419), .Z(n13416) );
  XOR U16983 ( .A(n13417), .B(n13420), .Z(n13418) );
  XOR U16984 ( .A(n13421), .B(n13422), .Z(n13392) );
  XNOR U16985 ( .A(n13387), .B(n13423), .Z(n13422) );
  IV U16986 ( .A(n13390), .Z(n13423) );
  XOR U16987 ( .A(n13424), .B(n13425), .Z(n13390) );
  ANDN U16988 ( .B(n13426), .A(n13427), .Z(n13424) );
  XOR U16989 ( .A(n13425), .B(n13428), .Z(n13426) );
  XNOR U16990 ( .A(n13429), .B(n13430), .Z(n13387) );
  ANDN U16991 ( .B(n13431), .A(n13432), .Z(n13429) );
  XOR U16992 ( .A(n13430), .B(n13433), .Z(n13431) );
  IV U16993 ( .A(n13386), .Z(n13421) );
  XOR U16994 ( .A(n13384), .B(n13434), .Z(n13386) );
  XNOR U16995 ( .A(n13435), .B(n13436), .Z(n13434) );
  ANDN U16996 ( .B(n13437), .A(n13438), .Z(n13435) );
  XNOR U16997 ( .A(n13439), .B(n13440), .Z(n13437) );
  IV U16998 ( .A(n13388), .Z(n13384) );
  XOR U16999 ( .A(n13441), .B(n13442), .Z(n13388) );
  ANDN U17000 ( .B(n13443), .A(n13444), .Z(n13441) );
  XOR U17001 ( .A(n13445), .B(n13442), .Z(n13443) );
  XOR U17002 ( .A(n13399), .B(n13252), .Z(n13400) );
  XOR U17003 ( .A(n13446), .B(n13447), .Z(n13252) );
  AND U17004 ( .A(n36), .B(n13448), .Z(n13446) );
  XOR U17005 ( .A(n13449), .B(n13447), .Z(n13448) );
  XNOR U17006 ( .A(n13450), .B(n13451), .Z(n13399) );
  NAND U17007 ( .A(n13452), .B(n13453), .Z(n13451) );
  XOR U17008 ( .A(n13454), .B(n13351), .Z(n13453) );
  XOR U17009 ( .A(n13427), .B(n13428), .Z(n13351) );
  XOR U17010 ( .A(n13455), .B(n13420), .Z(n13428) );
  XOR U17011 ( .A(n13456), .B(n13408), .Z(n13420) );
  XOR U17012 ( .A(n13457), .B(n13458), .Z(n13408) );
  ANDN U17013 ( .B(n13459), .A(n13460), .Z(n13457) );
  XOR U17014 ( .A(n13458), .B(n13461), .Z(n13459) );
  IV U17015 ( .A(n13406), .Z(n13456) );
  XOR U17016 ( .A(n13404), .B(n13462), .Z(n13406) );
  XOR U17017 ( .A(n13463), .B(n13464), .Z(n13462) );
  ANDN U17018 ( .B(n13465), .A(n13466), .Z(n13463) );
  XOR U17019 ( .A(n13467), .B(n13464), .Z(n13465) );
  IV U17020 ( .A(n13407), .Z(n13404) );
  XOR U17021 ( .A(n13468), .B(n13469), .Z(n13407) );
  ANDN U17022 ( .B(n13470), .A(n13471), .Z(n13468) );
  XOR U17023 ( .A(n13469), .B(n13472), .Z(n13470) );
  IV U17024 ( .A(n13419), .Z(n13455) );
  XOR U17025 ( .A(n13473), .B(n13474), .Z(n13419) );
  XNOR U17026 ( .A(n13414), .B(n13475), .Z(n13474) );
  IV U17027 ( .A(n13417), .Z(n13475) );
  XOR U17028 ( .A(n13476), .B(n13477), .Z(n13417) );
  ANDN U17029 ( .B(n13478), .A(n13479), .Z(n13476) );
  XOR U17030 ( .A(n13477), .B(n13480), .Z(n13478) );
  XNOR U17031 ( .A(n13481), .B(n13482), .Z(n13414) );
  ANDN U17032 ( .B(n13483), .A(n13484), .Z(n13481) );
  XOR U17033 ( .A(n13482), .B(n13485), .Z(n13483) );
  IV U17034 ( .A(n13413), .Z(n13473) );
  XOR U17035 ( .A(n13411), .B(n13486), .Z(n13413) );
  XOR U17036 ( .A(n13487), .B(n13488), .Z(n13486) );
  ANDN U17037 ( .B(n13489), .A(n13490), .Z(n13487) );
  XOR U17038 ( .A(n13491), .B(n13488), .Z(n13489) );
  IV U17039 ( .A(n13415), .Z(n13411) );
  XOR U17040 ( .A(n13492), .B(n13493), .Z(n13415) );
  ANDN U17041 ( .B(n13494), .A(n13495), .Z(n13492) );
  XOR U17042 ( .A(n13496), .B(n13493), .Z(n13494) );
  XOR U17043 ( .A(n13497), .B(n13498), .Z(n13427) );
  XOR U17044 ( .A(n13445), .B(n13499), .Z(n13498) );
  IV U17045 ( .A(n13425), .Z(n13499) );
  XOR U17046 ( .A(n13500), .B(n13501), .Z(n13425) );
  ANDN U17047 ( .B(n13502), .A(n13503), .Z(n13500) );
  XOR U17048 ( .A(n13501), .B(n13504), .Z(n13502) );
  XOR U17049 ( .A(n13505), .B(n13433), .Z(n13445) );
  XOR U17050 ( .A(n13506), .B(n13507), .Z(n13433) );
  ANDN U17051 ( .B(n13508), .A(n13509), .Z(n13506) );
  XOR U17052 ( .A(n13507), .B(n13510), .Z(n13508) );
  IV U17053 ( .A(n13432), .Z(n13505) );
  XOR U17054 ( .A(n13511), .B(n13512), .Z(n13432) );
  XOR U17055 ( .A(n13513), .B(n13514), .Z(n13512) );
  ANDN U17056 ( .B(n13515), .A(n13516), .Z(n13513) );
  XOR U17057 ( .A(n13517), .B(n13514), .Z(n13515) );
  IV U17058 ( .A(n13430), .Z(n13511) );
  XOR U17059 ( .A(n13518), .B(n13519), .Z(n13430) );
  ANDN U17060 ( .B(n13520), .A(n13521), .Z(n13518) );
  XOR U17061 ( .A(n13519), .B(n13522), .Z(n13520) );
  IV U17062 ( .A(n13444), .Z(n13497) );
  XOR U17063 ( .A(n13523), .B(n13524), .Z(n13444) );
  XNOR U17064 ( .A(n13439), .B(n13525), .Z(n13524) );
  IV U17065 ( .A(n13442), .Z(n13525) );
  XOR U17066 ( .A(n13526), .B(n13527), .Z(n13442) );
  ANDN U17067 ( .B(n13528), .A(n13529), .Z(n13526) );
  XOR U17068 ( .A(n13530), .B(n13527), .Z(n13528) );
  XNOR U17069 ( .A(n13531), .B(n13532), .Z(n13439) );
  ANDN U17070 ( .B(n13533), .A(n13534), .Z(n13531) );
  XOR U17071 ( .A(n13532), .B(n13535), .Z(n13533) );
  IV U17072 ( .A(n13438), .Z(n13523) );
  XOR U17073 ( .A(n13436), .B(n13536), .Z(n13438) );
  XOR U17074 ( .A(n13537), .B(n13538), .Z(n13536) );
  ANDN U17075 ( .B(n13539), .A(n13540), .Z(n13537) );
  XOR U17076 ( .A(n13541), .B(n13538), .Z(n13539) );
  IV U17077 ( .A(n13440), .Z(n13436) );
  XOR U17078 ( .A(n13542), .B(n13543), .Z(n13440) );
  ANDN U17079 ( .B(n13544), .A(n13545), .Z(n13542) );
  XOR U17080 ( .A(n13546), .B(n13543), .Z(n13544) );
  IV U17081 ( .A(n13450), .Z(n13454) );
  XOR U17082 ( .A(n13450), .B(n13353), .Z(n13452) );
  XOR U17083 ( .A(n13547), .B(n13548), .Z(n13353) );
  AND U17084 ( .A(n36), .B(n13549), .Z(n13547) );
  XOR U17085 ( .A(n13550), .B(n13548), .Z(n13549) );
  NANDN U17086 ( .A(n13355), .B(n13357), .Z(n13450) );
  XOR U17087 ( .A(n13551), .B(n13552), .Z(n13357) );
  AND U17088 ( .A(n36), .B(n13553), .Z(n13551) );
  XOR U17089 ( .A(n13552), .B(n13554), .Z(n13553) );
  XNOR U17090 ( .A(n13555), .B(n13556), .Z(n36) );
  AND U17091 ( .A(n13557), .B(n13558), .Z(n13555) );
  XOR U17092 ( .A(n13556), .B(n13368), .Z(n13558) );
  XNOR U17093 ( .A(n13559), .B(n13560), .Z(n13368) );
  ANDN U17094 ( .B(n13561), .A(n13562), .Z(n13559) );
  XOR U17095 ( .A(n13560), .B(n13563), .Z(n13561) );
  XNOR U17096 ( .A(n13556), .B(n13370), .Z(n13557) );
  XOR U17097 ( .A(n13564), .B(n13565), .Z(n13370) );
  AND U17098 ( .A(n40), .B(n13566), .Z(n13564) );
  XOR U17099 ( .A(n13567), .B(n13565), .Z(n13566) );
  XOR U17100 ( .A(n13568), .B(n13569), .Z(n13556) );
  AND U17101 ( .A(n13570), .B(n13571), .Z(n13568) );
  XOR U17102 ( .A(n13569), .B(n13395), .Z(n13571) );
  XOR U17103 ( .A(n13562), .B(n13563), .Z(n13395) );
  XNOR U17104 ( .A(n13572), .B(n13573), .Z(n13563) );
  ANDN U17105 ( .B(n13574), .A(n13575), .Z(n13572) );
  XOR U17106 ( .A(n13576), .B(n13577), .Z(n13574) );
  XOR U17107 ( .A(n13578), .B(n13579), .Z(n13562) );
  XNOR U17108 ( .A(n13580), .B(n13581), .Z(n13579) );
  ANDN U17109 ( .B(n13582), .A(n13583), .Z(n13580) );
  XNOR U17110 ( .A(n13584), .B(n13585), .Z(n13582) );
  IV U17111 ( .A(n13560), .Z(n13578) );
  XOR U17112 ( .A(n13586), .B(n13587), .Z(n13560) );
  ANDN U17113 ( .B(n13588), .A(n13589), .Z(n13586) );
  XOR U17114 ( .A(n13587), .B(n13590), .Z(n13588) );
  XNOR U17115 ( .A(n13569), .B(n13397), .Z(n13570) );
  XOR U17116 ( .A(n13591), .B(n13592), .Z(n13397) );
  AND U17117 ( .A(n40), .B(n13593), .Z(n13591) );
  XOR U17118 ( .A(n13594), .B(n13592), .Z(n13593) );
  XNOR U17119 ( .A(n13595), .B(n13596), .Z(n13569) );
  AND U17120 ( .A(n13597), .B(n13598), .Z(n13595) );
  XNOR U17121 ( .A(n13596), .B(n13447), .Z(n13598) );
  XOR U17122 ( .A(n13589), .B(n13590), .Z(n13447) );
  XOR U17123 ( .A(n13599), .B(n13577), .Z(n13590) );
  XNOR U17124 ( .A(n13600), .B(n13601), .Z(n13577) );
  ANDN U17125 ( .B(n13602), .A(n13603), .Z(n13600) );
  XOR U17126 ( .A(n13604), .B(n13605), .Z(n13602) );
  IV U17127 ( .A(n13575), .Z(n13599) );
  XOR U17128 ( .A(n13573), .B(n13606), .Z(n13575) );
  XNOR U17129 ( .A(n13607), .B(n13608), .Z(n13606) );
  ANDN U17130 ( .B(n13609), .A(n13610), .Z(n13607) );
  XNOR U17131 ( .A(n13611), .B(n13612), .Z(n13609) );
  IV U17132 ( .A(n13576), .Z(n13573) );
  XOR U17133 ( .A(n13613), .B(n13614), .Z(n13576) );
  ANDN U17134 ( .B(n13615), .A(n13616), .Z(n13613) );
  XOR U17135 ( .A(n13614), .B(n13617), .Z(n13615) );
  XOR U17136 ( .A(n13618), .B(n13619), .Z(n13589) );
  XNOR U17137 ( .A(n13584), .B(n13620), .Z(n13619) );
  IV U17138 ( .A(n13587), .Z(n13620) );
  XOR U17139 ( .A(n13621), .B(n13622), .Z(n13587) );
  ANDN U17140 ( .B(n13623), .A(n13624), .Z(n13621) );
  XOR U17141 ( .A(n13622), .B(n13625), .Z(n13623) );
  XNOR U17142 ( .A(n13626), .B(n13627), .Z(n13584) );
  ANDN U17143 ( .B(n13628), .A(n13629), .Z(n13626) );
  XOR U17144 ( .A(n13627), .B(n13630), .Z(n13628) );
  IV U17145 ( .A(n13583), .Z(n13618) );
  XOR U17146 ( .A(n13581), .B(n13631), .Z(n13583) );
  XNOR U17147 ( .A(n13632), .B(n13633), .Z(n13631) );
  ANDN U17148 ( .B(n13634), .A(n13635), .Z(n13632) );
  XNOR U17149 ( .A(n13636), .B(n13637), .Z(n13634) );
  IV U17150 ( .A(n13585), .Z(n13581) );
  XOR U17151 ( .A(n13638), .B(n13639), .Z(n13585) );
  ANDN U17152 ( .B(n13640), .A(n13641), .Z(n13638) );
  XOR U17153 ( .A(n13642), .B(n13639), .Z(n13640) );
  XOR U17154 ( .A(n13596), .B(n13449), .Z(n13597) );
  XOR U17155 ( .A(n13643), .B(n13644), .Z(n13449) );
  AND U17156 ( .A(n40), .B(n13645), .Z(n13643) );
  XOR U17157 ( .A(n13646), .B(n13644), .Z(n13645) );
  XNOR U17158 ( .A(n13647), .B(n13648), .Z(n13596) );
  NAND U17159 ( .A(n13649), .B(n13650), .Z(n13648) );
  XOR U17160 ( .A(n13651), .B(n13548), .Z(n13650) );
  XOR U17161 ( .A(n13624), .B(n13625), .Z(n13548) );
  XOR U17162 ( .A(n13652), .B(n13617), .Z(n13625) );
  XOR U17163 ( .A(n13653), .B(n13605), .Z(n13617) );
  XOR U17164 ( .A(n13654), .B(n13655), .Z(n13605) );
  ANDN U17165 ( .B(n13656), .A(n13657), .Z(n13654) );
  XOR U17166 ( .A(n13655), .B(n13658), .Z(n13656) );
  IV U17167 ( .A(n13603), .Z(n13653) );
  XOR U17168 ( .A(n13601), .B(n13659), .Z(n13603) );
  XOR U17169 ( .A(n13660), .B(n13661), .Z(n13659) );
  ANDN U17170 ( .B(n13662), .A(n13663), .Z(n13660) );
  XOR U17171 ( .A(n13664), .B(n13661), .Z(n13662) );
  IV U17172 ( .A(n13604), .Z(n13601) );
  XOR U17173 ( .A(n13665), .B(n13666), .Z(n13604) );
  ANDN U17174 ( .B(n13667), .A(n13668), .Z(n13665) );
  XOR U17175 ( .A(n13666), .B(n13669), .Z(n13667) );
  IV U17176 ( .A(n13616), .Z(n13652) );
  XOR U17177 ( .A(n13670), .B(n13671), .Z(n13616) );
  XNOR U17178 ( .A(n13611), .B(n13672), .Z(n13671) );
  IV U17179 ( .A(n13614), .Z(n13672) );
  XOR U17180 ( .A(n13673), .B(n13674), .Z(n13614) );
  ANDN U17181 ( .B(n13675), .A(n13676), .Z(n13673) );
  XOR U17182 ( .A(n13674), .B(n13677), .Z(n13675) );
  XNOR U17183 ( .A(n13678), .B(n13679), .Z(n13611) );
  ANDN U17184 ( .B(n13680), .A(n13681), .Z(n13678) );
  XOR U17185 ( .A(n13679), .B(n13682), .Z(n13680) );
  IV U17186 ( .A(n13610), .Z(n13670) );
  XOR U17187 ( .A(n13608), .B(n13683), .Z(n13610) );
  XOR U17188 ( .A(n13684), .B(n13685), .Z(n13683) );
  ANDN U17189 ( .B(n13686), .A(n13687), .Z(n13684) );
  XOR U17190 ( .A(n13688), .B(n13685), .Z(n13686) );
  IV U17191 ( .A(n13612), .Z(n13608) );
  XOR U17192 ( .A(n13689), .B(n13690), .Z(n13612) );
  ANDN U17193 ( .B(n13691), .A(n13692), .Z(n13689) );
  XOR U17194 ( .A(n13693), .B(n13690), .Z(n13691) );
  XOR U17195 ( .A(n13694), .B(n13695), .Z(n13624) );
  XOR U17196 ( .A(n13642), .B(n13696), .Z(n13695) );
  IV U17197 ( .A(n13622), .Z(n13696) );
  XOR U17198 ( .A(n13697), .B(n13698), .Z(n13622) );
  ANDN U17199 ( .B(n13699), .A(n13700), .Z(n13697) );
  XOR U17200 ( .A(n13698), .B(n13701), .Z(n13699) );
  XOR U17201 ( .A(n13702), .B(n13630), .Z(n13642) );
  XOR U17202 ( .A(n13703), .B(n13704), .Z(n13630) );
  ANDN U17203 ( .B(n13705), .A(n13706), .Z(n13703) );
  XOR U17204 ( .A(n13704), .B(n13707), .Z(n13705) );
  IV U17205 ( .A(n13629), .Z(n13702) );
  XOR U17206 ( .A(n13708), .B(n13709), .Z(n13629) );
  XOR U17207 ( .A(n13710), .B(n13711), .Z(n13709) );
  ANDN U17208 ( .B(n13712), .A(n13713), .Z(n13710) );
  XOR U17209 ( .A(n13714), .B(n13711), .Z(n13712) );
  IV U17210 ( .A(n13627), .Z(n13708) );
  XOR U17211 ( .A(n13715), .B(n13716), .Z(n13627) );
  ANDN U17212 ( .B(n13717), .A(n13718), .Z(n13715) );
  XOR U17213 ( .A(n13716), .B(n13719), .Z(n13717) );
  IV U17214 ( .A(n13641), .Z(n13694) );
  XOR U17215 ( .A(n13720), .B(n13721), .Z(n13641) );
  XNOR U17216 ( .A(n13636), .B(n13722), .Z(n13721) );
  IV U17217 ( .A(n13639), .Z(n13722) );
  XOR U17218 ( .A(n13723), .B(n13724), .Z(n13639) );
  ANDN U17219 ( .B(n13725), .A(n13726), .Z(n13723) );
  XOR U17220 ( .A(n13727), .B(n13724), .Z(n13725) );
  XNOR U17221 ( .A(n13728), .B(n13729), .Z(n13636) );
  ANDN U17222 ( .B(n13730), .A(n13731), .Z(n13728) );
  XOR U17223 ( .A(n13729), .B(n13732), .Z(n13730) );
  IV U17224 ( .A(n13635), .Z(n13720) );
  XOR U17225 ( .A(n13633), .B(n13733), .Z(n13635) );
  XOR U17226 ( .A(n13734), .B(n13735), .Z(n13733) );
  ANDN U17227 ( .B(n13736), .A(n13737), .Z(n13734) );
  XOR U17228 ( .A(n13738), .B(n13735), .Z(n13736) );
  IV U17229 ( .A(n13637), .Z(n13633) );
  XOR U17230 ( .A(n13739), .B(n13740), .Z(n13637) );
  ANDN U17231 ( .B(n13741), .A(n13742), .Z(n13739) );
  XOR U17232 ( .A(n13743), .B(n13740), .Z(n13741) );
  IV U17233 ( .A(n13647), .Z(n13651) );
  XOR U17234 ( .A(n13647), .B(n13550), .Z(n13649) );
  XOR U17235 ( .A(n13744), .B(n13745), .Z(n13550) );
  AND U17236 ( .A(n40), .B(n13746), .Z(n13744) );
  XOR U17237 ( .A(n13747), .B(n13745), .Z(n13746) );
  NANDN U17238 ( .A(n13552), .B(n13554), .Z(n13647) );
  XOR U17239 ( .A(n13748), .B(n13749), .Z(n13554) );
  AND U17240 ( .A(n40), .B(n13750), .Z(n13748) );
  XOR U17241 ( .A(n13749), .B(n13751), .Z(n13750) );
  XNOR U17242 ( .A(n13752), .B(n13753), .Z(n40) );
  AND U17243 ( .A(n13754), .B(n13755), .Z(n13752) );
  XOR U17244 ( .A(n13753), .B(n13565), .Z(n13755) );
  XNOR U17245 ( .A(n13756), .B(n13757), .Z(n13565) );
  ANDN U17246 ( .B(n13758), .A(n13759), .Z(n13756) );
  XOR U17247 ( .A(n13757), .B(n13760), .Z(n13758) );
  XNOR U17248 ( .A(n13753), .B(n13567), .Z(n13754) );
  XOR U17249 ( .A(n13761), .B(n13762), .Z(n13567) );
  AND U17250 ( .A(n44), .B(n13763), .Z(n13761) );
  XOR U17251 ( .A(n13764), .B(n13762), .Z(n13763) );
  XOR U17252 ( .A(n13765), .B(n13766), .Z(n13753) );
  AND U17253 ( .A(n13767), .B(n13768), .Z(n13765) );
  XOR U17254 ( .A(n13766), .B(n13592), .Z(n13768) );
  XOR U17255 ( .A(n13759), .B(n13760), .Z(n13592) );
  XNOR U17256 ( .A(n13769), .B(n13770), .Z(n13760) );
  ANDN U17257 ( .B(n13771), .A(n13772), .Z(n13769) );
  XOR U17258 ( .A(n13773), .B(n13774), .Z(n13771) );
  XOR U17259 ( .A(n13775), .B(n13776), .Z(n13759) );
  XNOR U17260 ( .A(n13777), .B(n13778), .Z(n13776) );
  ANDN U17261 ( .B(n13779), .A(n13780), .Z(n13777) );
  XNOR U17262 ( .A(n13781), .B(n13782), .Z(n13779) );
  IV U17263 ( .A(n13757), .Z(n13775) );
  XOR U17264 ( .A(n13783), .B(n13784), .Z(n13757) );
  ANDN U17265 ( .B(n13785), .A(n13786), .Z(n13783) );
  XOR U17266 ( .A(n13784), .B(n13787), .Z(n13785) );
  XNOR U17267 ( .A(n13766), .B(n13594), .Z(n13767) );
  XOR U17268 ( .A(n13788), .B(n13789), .Z(n13594) );
  AND U17269 ( .A(n44), .B(n13790), .Z(n13788) );
  XOR U17270 ( .A(n13791), .B(n13789), .Z(n13790) );
  XNOR U17271 ( .A(n13792), .B(n13793), .Z(n13766) );
  AND U17272 ( .A(n13794), .B(n13795), .Z(n13792) );
  XNOR U17273 ( .A(n13793), .B(n13644), .Z(n13795) );
  XOR U17274 ( .A(n13786), .B(n13787), .Z(n13644) );
  XOR U17275 ( .A(n13796), .B(n13774), .Z(n13787) );
  XNOR U17276 ( .A(n13797), .B(n13798), .Z(n13774) );
  ANDN U17277 ( .B(n13799), .A(n13800), .Z(n13797) );
  XOR U17278 ( .A(n13801), .B(n13802), .Z(n13799) );
  IV U17279 ( .A(n13772), .Z(n13796) );
  XOR U17280 ( .A(n13770), .B(n13803), .Z(n13772) );
  XNOR U17281 ( .A(n13804), .B(n13805), .Z(n13803) );
  ANDN U17282 ( .B(n13806), .A(n13807), .Z(n13804) );
  XNOR U17283 ( .A(n13808), .B(n13809), .Z(n13806) );
  IV U17284 ( .A(n13773), .Z(n13770) );
  XOR U17285 ( .A(n13810), .B(n13811), .Z(n13773) );
  ANDN U17286 ( .B(n13812), .A(n13813), .Z(n13810) );
  XOR U17287 ( .A(n13811), .B(n13814), .Z(n13812) );
  XOR U17288 ( .A(n13815), .B(n13816), .Z(n13786) );
  XNOR U17289 ( .A(n13781), .B(n13817), .Z(n13816) );
  IV U17290 ( .A(n13784), .Z(n13817) );
  XOR U17291 ( .A(n13818), .B(n13819), .Z(n13784) );
  ANDN U17292 ( .B(n13820), .A(n13821), .Z(n13818) );
  XOR U17293 ( .A(n13819), .B(n13822), .Z(n13820) );
  XNOR U17294 ( .A(n13823), .B(n13824), .Z(n13781) );
  ANDN U17295 ( .B(n13825), .A(n13826), .Z(n13823) );
  XOR U17296 ( .A(n13824), .B(n13827), .Z(n13825) );
  IV U17297 ( .A(n13780), .Z(n13815) );
  XOR U17298 ( .A(n13778), .B(n13828), .Z(n13780) );
  XNOR U17299 ( .A(n13829), .B(n13830), .Z(n13828) );
  ANDN U17300 ( .B(n13831), .A(n13832), .Z(n13829) );
  XNOR U17301 ( .A(n13833), .B(n13834), .Z(n13831) );
  IV U17302 ( .A(n13782), .Z(n13778) );
  XOR U17303 ( .A(n13835), .B(n13836), .Z(n13782) );
  ANDN U17304 ( .B(n13837), .A(n13838), .Z(n13835) );
  XOR U17305 ( .A(n13839), .B(n13836), .Z(n13837) );
  XOR U17306 ( .A(n13793), .B(n13646), .Z(n13794) );
  XOR U17307 ( .A(n13840), .B(n13841), .Z(n13646) );
  AND U17308 ( .A(n44), .B(n13842), .Z(n13840) );
  XOR U17309 ( .A(n13843), .B(n13841), .Z(n13842) );
  XNOR U17310 ( .A(n13844), .B(n13845), .Z(n13793) );
  NAND U17311 ( .A(n13846), .B(n13847), .Z(n13845) );
  XOR U17312 ( .A(n13848), .B(n13745), .Z(n13847) );
  XOR U17313 ( .A(n13821), .B(n13822), .Z(n13745) );
  XOR U17314 ( .A(n13849), .B(n13814), .Z(n13822) );
  XOR U17315 ( .A(n13850), .B(n13802), .Z(n13814) );
  XOR U17316 ( .A(n13851), .B(n13852), .Z(n13802) );
  ANDN U17317 ( .B(n13853), .A(n13854), .Z(n13851) );
  XOR U17318 ( .A(n13852), .B(n13855), .Z(n13853) );
  IV U17319 ( .A(n13800), .Z(n13850) );
  XOR U17320 ( .A(n13798), .B(n13856), .Z(n13800) );
  XOR U17321 ( .A(n13857), .B(n13858), .Z(n13856) );
  ANDN U17322 ( .B(n13859), .A(n13860), .Z(n13857) );
  XOR U17323 ( .A(n13861), .B(n13858), .Z(n13859) );
  IV U17324 ( .A(n13801), .Z(n13798) );
  XOR U17325 ( .A(n13862), .B(n13863), .Z(n13801) );
  ANDN U17326 ( .B(n13864), .A(n13865), .Z(n13862) );
  XOR U17327 ( .A(n13863), .B(n13866), .Z(n13864) );
  IV U17328 ( .A(n13813), .Z(n13849) );
  XOR U17329 ( .A(n13867), .B(n13868), .Z(n13813) );
  XNOR U17330 ( .A(n13808), .B(n13869), .Z(n13868) );
  IV U17331 ( .A(n13811), .Z(n13869) );
  XOR U17332 ( .A(n13870), .B(n13871), .Z(n13811) );
  ANDN U17333 ( .B(n13872), .A(n13873), .Z(n13870) );
  XOR U17334 ( .A(n13871), .B(n13874), .Z(n13872) );
  XNOR U17335 ( .A(n13875), .B(n13876), .Z(n13808) );
  ANDN U17336 ( .B(n13877), .A(n13878), .Z(n13875) );
  XOR U17337 ( .A(n13876), .B(n13879), .Z(n13877) );
  IV U17338 ( .A(n13807), .Z(n13867) );
  XOR U17339 ( .A(n13805), .B(n13880), .Z(n13807) );
  XOR U17340 ( .A(n13881), .B(n13882), .Z(n13880) );
  ANDN U17341 ( .B(n13883), .A(n13884), .Z(n13881) );
  XOR U17342 ( .A(n13885), .B(n13882), .Z(n13883) );
  IV U17343 ( .A(n13809), .Z(n13805) );
  XOR U17344 ( .A(n13886), .B(n13887), .Z(n13809) );
  ANDN U17345 ( .B(n13888), .A(n13889), .Z(n13886) );
  XOR U17346 ( .A(n13890), .B(n13887), .Z(n13888) );
  XOR U17347 ( .A(n13891), .B(n13892), .Z(n13821) );
  XOR U17348 ( .A(n13839), .B(n13893), .Z(n13892) );
  IV U17349 ( .A(n13819), .Z(n13893) );
  XOR U17350 ( .A(n13894), .B(n13895), .Z(n13819) );
  ANDN U17351 ( .B(n13896), .A(n13897), .Z(n13894) );
  XOR U17352 ( .A(n13895), .B(n13898), .Z(n13896) );
  XOR U17353 ( .A(n13899), .B(n13827), .Z(n13839) );
  XOR U17354 ( .A(n13900), .B(n13901), .Z(n13827) );
  ANDN U17355 ( .B(n13902), .A(n13903), .Z(n13900) );
  XOR U17356 ( .A(n13901), .B(n13904), .Z(n13902) );
  IV U17357 ( .A(n13826), .Z(n13899) );
  XOR U17358 ( .A(n13905), .B(n13906), .Z(n13826) );
  XOR U17359 ( .A(n13907), .B(n13908), .Z(n13906) );
  ANDN U17360 ( .B(n13909), .A(n13910), .Z(n13907) );
  XOR U17361 ( .A(n13911), .B(n13908), .Z(n13909) );
  IV U17362 ( .A(n13824), .Z(n13905) );
  XOR U17363 ( .A(n13912), .B(n13913), .Z(n13824) );
  ANDN U17364 ( .B(n13914), .A(n13915), .Z(n13912) );
  XOR U17365 ( .A(n13913), .B(n13916), .Z(n13914) );
  IV U17366 ( .A(n13838), .Z(n13891) );
  XOR U17367 ( .A(n13917), .B(n13918), .Z(n13838) );
  XNOR U17368 ( .A(n13833), .B(n13919), .Z(n13918) );
  IV U17369 ( .A(n13836), .Z(n13919) );
  XOR U17370 ( .A(n13920), .B(n13921), .Z(n13836) );
  ANDN U17371 ( .B(n13922), .A(n13923), .Z(n13920) );
  XOR U17372 ( .A(n13924), .B(n13921), .Z(n13922) );
  XNOR U17373 ( .A(n13925), .B(n13926), .Z(n13833) );
  ANDN U17374 ( .B(n13927), .A(n13928), .Z(n13925) );
  XOR U17375 ( .A(n13926), .B(n13929), .Z(n13927) );
  IV U17376 ( .A(n13832), .Z(n13917) );
  XOR U17377 ( .A(n13830), .B(n13930), .Z(n13832) );
  XOR U17378 ( .A(n13931), .B(n13932), .Z(n13930) );
  ANDN U17379 ( .B(n13933), .A(n13934), .Z(n13931) );
  XOR U17380 ( .A(n13935), .B(n13932), .Z(n13933) );
  IV U17381 ( .A(n13834), .Z(n13830) );
  XOR U17382 ( .A(n13936), .B(n13937), .Z(n13834) );
  ANDN U17383 ( .B(n13938), .A(n13939), .Z(n13936) );
  XOR U17384 ( .A(n13940), .B(n13937), .Z(n13938) );
  IV U17385 ( .A(n13844), .Z(n13848) );
  XOR U17386 ( .A(n13844), .B(n13747), .Z(n13846) );
  XOR U17387 ( .A(n13941), .B(n13942), .Z(n13747) );
  AND U17388 ( .A(n44), .B(n13943), .Z(n13941) );
  XOR U17389 ( .A(n13944), .B(n13942), .Z(n13943) );
  NANDN U17390 ( .A(n13749), .B(n13751), .Z(n13844) );
  XOR U17391 ( .A(n13945), .B(n13946), .Z(n13751) );
  AND U17392 ( .A(n44), .B(n13947), .Z(n13945) );
  XOR U17393 ( .A(n13946), .B(n13948), .Z(n13947) );
  XNOR U17394 ( .A(n13949), .B(n13950), .Z(n44) );
  AND U17395 ( .A(n13951), .B(n13952), .Z(n13949) );
  XOR U17396 ( .A(n13950), .B(n13762), .Z(n13952) );
  XNOR U17397 ( .A(n13953), .B(n13954), .Z(n13762) );
  ANDN U17398 ( .B(n13955), .A(n13956), .Z(n13953) );
  XOR U17399 ( .A(n13954), .B(n13957), .Z(n13955) );
  XNOR U17400 ( .A(n13950), .B(n13764), .Z(n13951) );
  XOR U17401 ( .A(n13958), .B(n13959), .Z(n13764) );
  AND U17402 ( .A(n48), .B(n13960), .Z(n13958) );
  XOR U17403 ( .A(n13961), .B(n13959), .Z(n13960) );
  XOR U17404 ( .A(n13962), .B(n13963), .Z(n13950) );
  AND U17405 ( .A(n13964), .B(n13965), .Z(n13962) );
  XOR U17406 ( .A(n13963), .B(n13789), .Z(n13965) );
  XOR U17407 ( .A(n13956), .B(n13957), .Z(n13789) );
  XNOR U17408 ( .A(n13966), .B(n13967), .Z(n13957) );
  ANDN U17409 ( .B(n13968), .A(n13969), .Z(n13966) );
  XOR U17410 ( .A(n13970), .B(n13971), .Z(n13968) );
  XOR U17411 ( .A(n13972), .B(n13973), .Z(n13956) );
  XNOR U17412 ( .A(n13974), .B(n13975), .Z(n13973) );
  ANDN U17413 ( .B(n13976), .A(n13977), .Z(n13974) );
  XNOR U17414 ( .A(n13978), .B(n13979), .Z(n13976) );
  IV U17415 ( .A(n13954), .Z(n13972) );
  XOR U17416 ( .A(n13980), .B(n13981), .Z(n13954) );
  ANDN U17417 ( .B(n13982), .A(n13983), .Z(n13980) );
  XOR U17418 ( .A(n13981), .B(n13984), .Z(n13982) );
  XNOR U17419 ( .A(n13963), .B(n13791), .Z(n13964) );
  XOR U17420 ( .A(n13985), .B(n13986), .Z(n13791) );
  AND U17421 ( .A(n48), .B(n13987), .Z(n13985) );
  XOR U17422 ( .A(n13988), .B(n13986), .Z(n13987) );
  XNOR U17423 ( .A(n13989), .B(n13990), .Z(n13963) );
  AND U17424 ( .A(n13991), .B(n13992), .Z(n13989) );
  XNOR U17425 ( .A(n13990), .B(n13841), .Z(n13992) );
  XOR U17426 ( .A(n13983), .B(n13984), .Z(n13841) );
  XOR U17427 ( .A(n13993), .B(n13971), .Z(n13984) );
  XNOR U17428 ( .A(n13994), .B(n13995), .Z(n13971) );
  ANDN U17429 ( .B(n13996), .A(n13997), .Z(n13994) );
  XOR U17430 ( .A(n13998), .B(n13999), .Z(n13996) );
  IV U17431 ( .A(n13969), .Z(n13993) );
  XOR U17432 ( .A(n13967), .B(n14000), .Z(n13969) );
  XNOR U17433 ( .A(n14001), .B(n14002), .Z(n14000) );
  ANDN U17434 ( .B(n14003), .A(n14004), .Z(n14001) );
  XNOR U17435 ( .A(n14005), .B(n14006), .Z(n14003) );
  IV U17436 ( .A(n13970), .Z(n13967) );
  XOR U17437 ( .A(n14007), .B(n14008), .Z(n13970) );
  ANDN U17438 ( .B(n14009), .A(n14010), .Z(n14007) );
  XOR U17439 ( .A(n14008), .B(n14011), .Z(n14009) );
  XOR U17440 ( .A(n14012), .B(n14013), .Z(n13983) );
  XNOR U17441 ( .A(n13978), .B(n14014), .Z(n14013) );
  IV U17442 ( .A(n13981), .Z(n14014) );
  XOR U17443 ( .A(n14015), .B(n14016), .Z(n13981) );
  ANDN U17444 ( .B(n14017), .A(n14018), .Z(n14015) );
  XOR U17445 ( .A(n14016), .B(n14019), .Z(n14017) );
  XNOR U17446 ( .A(n14020), .B(n14021), .Z(n13978) );
  ANDN U17447 ( .B(n14022), .A(n14023), .Z(n14020) );
  XOR U17448 ( .A(n14021), .B(n14024), .Z(n14022) );
  IV U17449 ( .A(n13977), .Z(n14012) );
  XOR U17450 ( .A(n13975), .B(n14025), .Z(n13977) );
  XNOR U17451 ( .A(n14026), .B(n14027), .Z(n14025) );
  ANDN U17452 ( .B(n14028), .A(n14029), .Z(n14026) );
  XNOR U17453 ( .A(n14030), .B(n14031), .Z(n14028) );
  IV U17454 ( .A(n13979), .Z(n13975) );
  XOR U17455 ( .A(n14032), .B(n14033), .Z(n13979) );
  ANDN U17456 ( .B(n14034), .A(n14035), .Z(n14032) );
  XOR U17457 ( .A(n14036), .B(n14033), .Z(n14034) );
  XOR U17458 ( .A(n13990), .B(n13843), .Z(n13991) );
  XOR U17459 ( .A(n14037), .B(n14038), .Z(n13843) );
  AND U17460 ( .A(n48), .B(n14039), .Z(n14037) );
  XOR U17461 ( .A(n14040), .B(n14038), .Z(n14039) );
  XNOR U17462 ( .A(n14041), .B(n14042), .Z(n13990) );
  NAND U17463 ( .A(n14043), .B(n14044), .Z(n14042) );
  XOR U17464 ( .A(n14045), .B(n13942), .Z(n14044) );
  XOR U17465 ( .A(n14018), .B(n14019), .Z(n13942) );
  XOR U17466 ( .A(n14046), .B(n14011), .Z(n14019) );
  XOR U17467 ( .A(n14047), .B(n13999), .Z(n14011) );
  XOR U17468 ( .A(n14048), .B(n14049), .Z(n13999) );
  ANDN U17469 ( .B(n14050), .A(n14051), .Z(n14048) );
  XOR U17470 ( .A(n14049), .B(n14052), .Z(n14050) );
  IV U17471 ( .A(n13997), .Z(n14047) );
  XOR U17472 ( .A(n13995), .B(n14053), .Z(n13997) );
  XOR U17473 ( .A(n14054), .B(n14055), .Z(n14053) );
  ANDN U17474 ( .B(n14056), .A(n14057), .Z(n14054) );
  XOR U17475 ( .A(n14058), .B(n14055), .Z(n14056) );
  IV U17476 ( .A(n13998), .Z(n13995) );
  XOR U17477 ( .A(n14059), .B(n14060), .Z(n13998) );
  ANDN U17478 ( .B(n14061), .A(n14062), .Z(n14059) );
  XOR U17479 ( .A(n14060), .B(n14063), .Z(n14061) );
  IV U17480 ( .A(n14010), .Z(n14046) );
  XOR U17481 ( .A(n14064), .B(n14065), .Z(n14010) );
  XNOR U17482 ( .A(n14005), .B(n14066), .Z(n14065) );
  IV U17483 ( .A(n14008), .Z(n14066) );
  XOR U17484 ( .A(n14067), .B(n14068), .Z(n14008) );
  ANDN U17485 ( .B(n14069), .A(n14070), .Z(n14067) );
  XOR U17486 ( .A(n14068), .B(n14071), .Z(n14069) );
  XNOR U17487 ( .A(n14072), .B(n14073), .Z(n14005) );
  ANDN U17488 ( .B(n14074), .A(n14075), .Z(n14072) );
  XOR U17489 ( .A(n14073), .B(n14076), .Z(n14074) );
  IV U17490 ( .A(n14004), .Z(n14064) );
  XOR U17491 ( .A(n14002), .B(n14077), .Z(n14004) );
  XOR U17492 ( .A(n14078), .B(n14079), .Z(n14077) );
  ANDN U17493 ( .B(n14080), .A(n14081), .Z(n14078) );
  XOR U17494 ( .A(n14082), .B(n14079), .Z(n14080) );
  IV U17495 ( .A(n14006), .Z(n14002) );
  XOR U17496 ( .A(n14083), .B(n14084), .Z(n14006) );
  ANDN U17497 ( .B(n14085), .A(n14086), .Z(n14083) );
  XOR U17498 ( .A(n14087), .B(n14084), .Z(n14085) );
  XOR U17499 ( .A(n14088), .B(n14089), .Z(n14018) );
  XOR U17500 ( .A(n14036), .B(n14090), .Z(n14089) );
  IV U17501 ( .A(n14016), .Z(n14090) );
  XOR U17502 ( .A(n14091), .B(n14092), .Z(n14016) );
  ANDN U17503 ( .B(n14093), .A(n14094), .Z(n14091) );
  XOR U17504 ( .A(n14092), .B(n14095), .Z(n14093) );
  XOR U17505 ( .A(n14096), .B(n14024), .Z(n14036) );
  XOR U17506 ( .A(n14097), .B(n14098), .Z(n14024) );
  ANDN U17507 ( .B(n14099), .A(n14100), .Z(n14097) );
  XOR U17508 ( .A(n14098), .B(n14101), .Z(n14099) );
  IV U17509 ( .A(n14023), .Z(n14096) );
  XOR U17510 ( .A(n14102), .B(n14103), .Z(n14023) );
  XOR U17511 ( .A(n14104), .B(n14105), .Z(n14103) );
  ANDN U17512 ( .B(n14106), .A(n14107), .Z(n14104) );
  XOR U17513 ( .A(n14108), .B(n14105), .Z(n14106) );
  IV U17514 ( .A(n14021), .Z(n14102) );
  XOR U17515 ( .A(n14109), .B(n14110), .Z(n14021) );
  ANDN U17516 ( .B(n14111), .A(n14112), .Z(n14109) );
  XOR U17517 ( .A(n14110), .B(n14113), .Z(n14111) );
  IV U17518 ( .A(n14035), .Z(n14088) );
  XOR U17519 ( .A(n14114), .B(n14115), .Z(n14035) );
  XNOR U17520 ( .A(n14030), .B(n14116), .Z(n14115) );
  IV U17521 ( .A(n14033), .Z(n14116) );
  XOR U17522 ( .A(n14117), .B(n14118), .Z(n14033) );
  ANDN U17523 ( .B(n14119), .A(n14120), .Z(n14117) );
  XOR U17524 ( .A(n14121), .B(n14118), .Z(n14119) );
  XNOR U17525 ( .A(n14122), .B(n14123), .Z(n14030) );
  ANDN U17526 ( .B(n14124), .A(n14125), .Z(n14122) );
  XOR U17527 ( .A(n14123), .B(n14126), .Z(n14124) );
  IV U17528 ( .A(n14029), .Z(n14114) );
  XOR U17529 ( .A(n14027), .B(n14127), .Z(n14029) );
  XOR U17530 ( .A(n14128), .B(n14129), .Z(n14127) );
  ANDN U17531 ( .B(n14130), .A(n14131), .Z(n14128) );
  XOR U17532 ( .A(n14132), .B(n14129), .Z(n14130) );
  IV U17533 ( .A(n14031), .Z(n14027) );
  XOR U17534 ( .A(n14133), .B(n14134), .Z(n14031) );
  ANDN U17535 ( .B(n14135), .A(n14136), .Z(n14133) );
  XOR U17536 ( .A(n14137), .B(n14134), .Z(n14135) );
  IV U17537 ( .A(n14041), .Z(n14045) );
  XOR U17538 ( .A(n14041), .B(n13944), .Z(n14043) );
  XOR U17539 ( .A(n14138), .B(n14139), .Z(n13944) );
  AND U17540 ( .A(n48), .B(n14140), .Z(n14138) );
  XOR U17541 ( .A(n14141), .B(n14139), .Z(n14140) );
  NANDN U17542 ( .A(n13946), .B(n13948), .Z(n14041) );
  XOR U17543 ( .A(n14142), .B(n14143), .Z(n13948) );
  AND U17544 ( .A(n48), .B(n14144), .Z(n14142) );
  XOR U17545 ( .A(n14143), .B(n14145), .Z(n14144) );
  XNOR U17546 ( .A(n14146), .B(n14147), .Z(n48) );
  AND U17547 ( .A(n14148), .B(n14149), .Z(n14146) );
  XOR U17548 ( .A(n14147), .B(n13959), .Z(n14149) );
  XNOR U17549 ( .A(n14150), .B(n14151), .Z(n13959) );
  ANDN U17550 ( .B(n14152), .A(n14153), .Z(n14150) );
  XOR U17551 ( .A(n14151), .B(n14154), .Z(n14152) );
  XNOR U17552 ( .A(n14147), .B(n13961), .Z(n14148) );
  XOR U17553 ( .A(n14155), .B(n14156), .Z(n13961) );
  AND U17554 ( .A(n52), .B(n14157), .Z(n14155) );
  XOR U17555 ( .A(n14158), .B(n14156), .Z(n14157) );
  XOR U17556 ( .A(n14159), .B(n14160), .Z(n14147) );
  AND U17557 ( .A(n14161), .B(n14162), .Z(n14159) );
  XOR U17558 ( .A(n14160), .B(n13986), .Z(n14162) );
  XOR U17559 ( .A(n14153), .B(n14154), .Z(n13986) );
  XNOR U17560 ( .A(n14163), .B(n14164), .Z(n14154) );
  ANDN U17561 ( .B(n14165), .A(n14166), .Z(n14163) );
  XOR U17562 ( .A(n14167), .B(n14168), .Z(n14165) );
  XOR U17563 ( .A(n14169), .B(n14170), .Z(n14153) );
  XNOR U17564 ( .A(n14171), .B(n14172), .Z(n14170) );
  ANDN U17565 ( .B(n14173), .A(n14174), .Z(n14171) );
  XNOR U17566 ( .A(n14175), .B(n14176), .Z(n14173) );
  IV U17567 ( .A(n14151), .Z(n14169) );
  XOR U17568 ( .A(n14177), .B(n14178), .Z(n14151) );
  ANDN U17569 ( .B(n14179), .A(n14180), .Z(n14177) );
  XOR U17570 ( .A(n14178), .B(n14181), .Z(n14179) );
  XNOR U17571 ( .A(n14160), .B(n13988), .Z(n14161) );
  XOR U17572 ( .A(n14182), .B(n14183), .Z(n13988) );
  AND U17573 ( .A(n52), .B(n14184), .Z(n14182) );
  XOR U17574 ( .A(n14185), .B(n14183), .Z(n14184) );
  XNOR U17575 ( .A(n14186), .B(n14187), .Z(n14160) );
  AND U17576 ( .A(n14188), .B(n14189), .Z(n14186) );
  XNOR U17577 ( .A(n14187), .B(n14038), .Z(n14189) );
  XOR U17578 ( .A(n14180), .B(n14181), .Z(n14038) );
  XOR U17579 ( .A(n14190), .B(n14168), .Z(n14181) );
  XNOR U17580 ( .A(n14191), .B(n14192), .Z(n14168) );
  ANDN U17581 ( .B(n14193), .A(n14194), .Z(n14191) );
  XOR U17582 ( .A(n14195), .B(n14196), .Z(n14193) );
  IV U17583 ( .A(n14166), .Z(n14190) );
  XOR U17584 ( .A(n14164), .B(n14197), .Z(n14166) );
  XNOR U17585 ( .A(n14198), .B(n14199), .Z(n14197) );
  ANDN U17586 ( .B(n14200), .A(n14201), .Z(n14198) );
  XNOR U17587 ( .A(n14202), .B(n14203), .Z(n14200) );
  IV U17588 ( .A(n14167), .Z(n14164) );
  XOR U17589 ( .A(n14204), .B(n14205), .Z(n14167) );
  ANDN U17590 ( .B(n14206), .A(n14207), .Z(n14204) );
  XOR U17591 ( .A(n14205), .B(n14208), .Z(n14206) );
  XOR U17592 ( .A(n14209), .B(n14210), .Z(n14180) );
  XNOR U17593 ( .A(n14175), .B(n14211), .Z(n14210) );
  IV U17594 ( .A(n14178), .Z(n14211) );
  XOR U17595 ( .A(n14212), .B(n14213), .Z(n14178) );
  ANDN U17596 ( .B(n14214), .A(n14215), .Z(n14212) );
  XOR U17597 ( .A(n14213), .B(n14216), .Z(n14214) );
  XNOR U17598 ( .A(n14217), .B(n14218), .Z(n14175) );
  ANDN U17599 ( .B(n14219), .A(n14220), .Z(n14217) );
  XOR U17600 ( .A(n14218), .B(n14221), .Z(n14219) );
  IV U17601 ( .A(n14174), .Z(n14209) );
  XOR U17602 ( .A(n14172), .B(n14222), .Z(n14174) );
  XNOR U17603 ( .A(n14223), .B(n14224), .Z(n14222) );
  ANDN U17604 ( .B(n14225), .A(n14226), .Z(n14223) );
  XNOR U17605 ( .A(n14227), .B(n14228), .Z(n14225) );
  IV U17606 ( .A(n14176), .Z(n14172) );
  XOR U17607 ( .A(n14229), .B(n14230), .Z(n14176) );
  ANDN U17608 ( .B(n14231), .A(n14232), .Z(n14229) );
  XOR U17609 ( .A(n14233), .B(n14230), .Z(n14231) );
  XOR U17610 ( .A(n14187), .B(n14040), .Z(n14188) );
  XOR U17611 ( .A(n14234), .B(n14235), .Z(n14040) );
  AND U17612 ( .A(n52), .B(n14236), .Z(n14234) );
  XOR U17613 ( .A(n14237), .B(n14235), .Z(n14236) );
  XNOR U17614 ( .A(n14238), .B(n14239), .Z(n14187) );
  NAND U17615 ( .A(n14240), .B(n14241), .Z(n14239) );
  XOR U17616 ( .A(n14242), .B(n14139), .Z(n14241) );
  XOR U17617 ( .A(n14215), .B(n14216), .Z(n14139) );
  XOR U17618 ( .A(n14243), .B(n14208), .Z(n14216) );
  XOR U17619 ( .A(n14244), .B(n14196), .Z(n14208) );
  XOR U17620 ( .A(n14245), .B(n14246), .Z(n14196) );
  ANDN U17621 ( .B(n14247), .A(n14248), .Z(n14245) );
  XOR U17622 ( .A(n14246), .B(n14249), .Z(n14247) );
  IV U17623 ( .A(n14194), .Z(n14244) );
  XOR U17624 ( .A(n14192), .B(n14250), .Z(n14194) );
  XOR U17625 ( .A(n14251), .B(n14252), .Z(n14250) );
  ANDN U17626 ( .B(n14253), .A(n14254), .Z(n14251) );
  XOR U17627 ( .A(n14255), .B(n14252), .Z(n14253) );
  IV U17628 ( .A(n14195), .Z(n14192) );
  XOR U17629 ( .A(n14256), .B(n14257), .Z(n14195) );
  ANDN U17630 ( .B(n14258), .A(n14259), .Z(n14256) );
  XOR U17631 ( .A(n14257), .B(n14260), .Z(n14258) );
  IV U17632 ( .A(n14207), .Z(n14243) );
  XOR U17633 ( .A(n14261), .B(n14262), .Z(n14207) );
  XNOR U17634 ( .A(n14202), .B(n14263), .Z(n14262) );
  IV U17635 ( .A(n14205), .Z(n14263) );
  XOR U17636 ( .A(n14264), .B(n14265), .Z(n14205) );
  ANDN U17637 ( .B(n14266), .A(n14267), .Z(n14264) );
  XOR U17638 ( .A(n14265), .B(n14268), .Z(n14266) );
  XNOR U17639 ( .A(n14269), .B(n14270), .Z(n14202) );
  ANDN U17640 ( .B(n14271), .A(n14272), .Z(n14269) );
  XOR U17641 ( .A(n14270), .B(n14273), .Z(n14271) );
  IV U17642 ( .A(n14201), .Z(n14261) );
  XOR U17643 ( .A(n14199), .B(n14274), .Z(n14201) );
  XOR U17644 ( .A(n14275), .B(n14276), .Z(n14274) );
  ANDN U17645 ( .B(n14277), .A(n14278), .Z(n14275) );
  XOR U17646 ( .A(n14279), .B(n14276), .Z(n14277) );
  IV U17647 ( .A(n14203), .Z(n14199) );
  XOR U17648 ( .A(n14280), .B(n14281), .Z(n14203) );
  ANDN U17649 ( .B(n14282), .A(n14283), .Z(n14280) );
  XOR U17650 ( .A(n14284), .B(n14281), .Z(n14282) );
  XOR U17651 ( .A(n14285), .B(n14286), .Z(n14215) );
  XOR U17652 ( .A(n14233), .B(n14287), .Z(n14286) );
  IV U17653 ( .A(n14213), .Z(n14287) );
  XOR U17654 ( .A(n14288), .B(n14289), .Z(n14213) );
  ANDN U17655 ( .B(n14290), .A(n14291), .Z(n14288) );
  XOR U17656 ( .A(n14289), .B(n14292), .Z(n14290) );
  XOR U17657 ( .A(n14293), .B(n14221), .Z(n14233) );
  XOR U17658 ( .A(n14294), .B(n14295), .Z(n14221) );
  ANDN U17659 ( .B(n14296), .A(n14297), .Z(n14294) );
  XOR U17660 ( .A(n14295), .B(n14298), .Z(n14296) );
  IV U17661 ( .A(n14220), .Z(n14293) );
  XOR U17662 ( .A(n14299), .B(n14300), .Z(n14220) );
  XOR U17663 ( .A(n14301), .B(n14302), .Z(n14300) );
  ANDN U17664 ( .B(n14303), .A(n14304), .Z(n14301) );
  XOR U17665 ( .A(n14305), .B(n14302), .Z(n14303) );
  IV U17666 ( .A(n14218), .Z(n14299) );
  XOR U17667 ( .A(n14306), .B(n14307), .Z(n14218) );
  ANDN U17668 ( .B(n14308), .A(n14309), .Z(n14306) );
  XOR U17669 ( .A(n14307), .B(n14310), .Z(n14308) );
  IV U17670 ( .A(n14232), .Z(n14285) );
  XOR U17671 ( .A(n14311), .B(n14312), .Z(n14232) );
  XNOR U17672 ( .A(n14227), .B(n14313), .Z(n14312) );
  IV U17673 ( .A(n14230), .Z(n14313) );
  XOR U17674 ( .A(n14314), .B(n14315), .Z(n14230) );
  ANDN U17675 ( .B(n14316), .A(n14317), .Z(n14314) );
  XOR U17676 ( .A(n14318), .B(n14315), .Z(n14316) );
  XNOR U17677 ( .A(n14319), .B(n14320), .Z(n14227) );
  ANDN U17678 ( .B(n14321), .A(n14322), .Z(n14319) );
  XOR U17679 ( .A(n14320), .B(n14323), .Z(n14321) );
  IV U17680 ( .A(n14226), .Z(n14311) );
  XOR U17681 ( .A(n14224), .B(n14324), .Z(n14226) );
  XOR U17682 ( .A(n14325), .B(n14326), .Z(n14324) );
  ANDN U17683 ( .B(n14327), .A(n14328), .Z(n14325) );
  XOR U17684 ( .A(n14329), .B(n14326), .Z(n14327) );
  IV U17685 ( .A(n14228), .Z(n14224) );
  XOR U17686 ( .A(n14330), .B(n14331), .Z(n14228) );
  ANDN U17687 ( .B(n14332), .A(n14333), .Z(n14330) );
  XOR U17688 ( .A(n14334), .B(n14331), .Z(n14332) );
  IV U17689 ( .A(n14238), .Z(n14242) );
  XOR U17690 ( .A(n14238), .B(n14141), .Z(n14240) );
  XOR U17691 ( .A(n14335), .B(n14336), .Z(n14141) );
  AND U17692 ( .A(n52), .B(n14337), .Z(n14335) );
  XOR U17693 ( .A(n14338), .B(n14336), .Z(n14337) );
  NANDN U17694 ( .A(n14143), .B(n14145), .Z(n14238) );
  XOR U17695 ( .A(n14339), .B(n14340), .Z(n14145) );
  AND U17696 ( .A(n52), .B(n14341), .Z(n14339) );
  XOR U17697 ( .A(n14340), .B(n14342), .Z(n14341) );
  XNOR U17698 ( .A(n14343), .B(n14344), .Z(n52) );
  AND U17699 ( .A(n14345), .B(n14346), .Z(n14343) );
  XOR U17700 ( .A(n14344), .B(n14156), .Z(n14346) );
  XNOR U17701 ( .A(n14347), .B(n14348), .Z(n14156) );
  ANDN U17702 ( .B(n14349), .A(n14350), .Z(n14347) );
  XOR U17703 ( .A(n14348), .B(n14351), .Z(n14349) );
  XNOR U17704 ( .A(n14344), .B(n14158), .Z(n14345) );
  XOR U17705 ( .A(n14352), .B(n14353), .Z(n14158) );
  AND U17706 ( .A(n56), .B(n14354), .Z(n14352) );
  XOR U17707 ( .A(n14355), .B(n14353), .Z(n14354) );
  XOR U17708 ( .A(n14356), .B(n14357), .Z(n14344) );
  AND U17709 ( .A(n14358), .B(n14359), .Z(n14356) );
  XOR U17710 ( .A(n14357), .B(n14183), .Z(n14359) );
  XOR U17711 ( .A(n14350), .B(n14351), .Z(n14183) );
  XNOR U17712 ( .A(n14360), .B(n14361), .Z(n14351) );
  ANDN U17713 ( .B(n14362), .A(n14363), .Z(n14360) );
  XOR U17714 ( .A(n14364), .B(n14365), .Z(n14362) );
  XOR U17715 ( .A(n14366), .B(n14367), .Z(n14350) );
  XNOR U17716 ( .A(n14368), .B(n14369), .Z(n14367) );
  ANDN U17717 ( .B(n14370), .A(n14371), .Z(n14368) );
  XNOR U17718 ( .A(n14372), .B(n14373), .Z(n14370) );
  IV U17719 ( .A(n14348), .Z(n14366) );
  XOR U17720 ( .A(n14374), .B(n14375), .Z(n14348) );
  ANDN U17721 ( .B(n14376), .A(n14377), .Z(n14374) );
  XOR U17722 ( .A(n14375), .B(n14378), .Z(n14376) );
  XNOR U17723 ( .A(n14357), .B(n14185), .Z(n14358) );
  XOR U17724 ( .A(n14379), .B(n14380), .Z(n14185) );
  AND U17725 ( .A(n56), .B(n14381), .Z(n14379) );
  XOR U17726 ( .A(n14382), .B(n14380), .Z(n14381) );
  XNOR U17727 ( .A(n14383), .B(n14384), .Z(n14357) );
  AND U17728 ( .A(n14385), .B(n14386), .Z(n14383) );
  XNOR U17729 ( .A(n14384), .B(n14235), .Z(n14386) );
  XOR U17730 ( .A(n14377), .B(n14378), .Z(n14235) );
  XOR U17731 ( .A(n14387), .B(n14365), .Z(n14378) );
  XNOR U17732 ( .A(n14388), .B(n14389), .Z(n14365) );
  ANDN U17733 ( .B(n14390), .A(n14391), .Z(n14388) );
  XOR U17734 ( .A(n14392), .B(n14393), .Z(n14390) );
  IV U17735 ( .A(n14363), .Z(n14387) );
  XOR U17736 ( .A(n14361), .B(n14394), .Z(n14363) );
  XNOR U17737 ( .A(n14395), .B(n14396), .Z(n14394) );
  ANDN U17738 ( .B(n14397), .A(n14398), .Z(n14395) );
  XNOR U17739 ( .A(n14399), .B(n14400), .Z(n14397) );
  IV U17740 ( .A(n14364), .Z(n14361) );
  XOR U17741 ( .A(n14401), .B(n14402), .Z(n14364) );
  ANDN U17742 ( .B(n14403), .A(n14404), .Z(n14401) );
  XOR U17743 ( .A(n14402), .B(n14405), .Z(n14403) );
  XOR U17744 ( .A(n14406), .B(n14407), .Z(n14377) );
  XNOR U17745 ( .A(n14372), .B(n14408), .Z(n14407) );
  IV U17746 ( .A(n14375), .Z(n14408) );
  XOR U17747 ( .A(n14409), .B(n14410), .Z(n14375) );
  ANDN U17748 ( .B(n14411), .A(n14412), .Z(n14409) );
  XOR U17749 ( .A(n14410), .B(n14413), .Z(n14411) );
  XNOR U17750 ( .A(n14414), .B(n14415), .Z(n14372) );
  ANDN U17751 ( .B(n14416), .A(n14417), .Z(n14414) );
  XOR U17752 ( .A(n14415), .B(n14418), .Z(n14416) );
  IV U17753 ( .A(n14371), .Z(n14406) );
  XOR U17754 ( .A(n14369), .B(n14419), .Z(n14371) );
  XNOR U17755 ( .A(n14420), .B(n14421), .Z(n14419) );
  ANDN U17756 ( .B(n14422), .A(n14423), .Z(n14420) );
  XNOR U17757 ( .A(n14424), .B(n14425), .Z(n14422) );
  IV U17758 ( .A(n14373), .Z(n14369) );
  XOR U17759 ( .A(n14426), .B(n14427), .Z(n14373) );
  ANDN U17760 ( .B(n14428), .A(n14429), .Z(n14426) );
  XOR U17761 ( .A(n14430), .B(n14427), .Z(n14428) );
  XOR U17762 ( .A(n14384), .B(n14237), .Z(n14385) );
  XOR U17763 ( .A(n14431), .B(n14432), .Z(n14237) );
  AND U17764 ( .A(n56), .B(n14433), .Z(n14431) );
  XOR U17765 ( .A(n14434), .B(n14432), .Z(n14433) );
  XNOR U17766 ( .A(n14435), .B(n14436), .Z(n14384) );
  NAND U17767 ( .A(n14437), .B(n14438), .Z(n14436) );
  XOR U17768 ( .A(n14439), .B(n14336), .Z(n14438) );
  XOR U17769 ( .A(n14412), .B(n14413), .Z(n14336) );
  XOR U17770 ( .A(n14440), .B(n14405), .Z(n14413) );
  XOR U17771 ( .A(n14441), .B(n14393), .Z(n14405) );
  XOR U17772 ( .A(n14442), .B(n14443), .Z(n14393) );
  ANDN U17773 ( .B(n14444), .A(n14445), .Z(n14442) );
  XOR U17774 ( .A(n14443), .B(n14446), .Z(n14444) );
  IV U17775 ( .A(n14391), .Z(n14441) );
  XOR U17776 ( .A(n14389), .B(n14447), .Z(n14391) );
  XOR U17777 ( .A(n14448), .B(n14449), .Z(n14447) );
  ANDN U17778 ( .B(n14450), .A(n14451), .Z(n14448) );
  XOR U17779 ( .A(n14452), .B(n14449), .Z(n14450) );
  IV U17780 ( .A(n14392), .Z(n14389) );
  XOR U17781 ( .A(n14453), .B(n14454), .Z(n14392) );
  ANDN U17782 ( .B(n14455), .A(n14456), .Z(n14453) );
  XOR U17783 ( .A(n14454), .B(n14457), .Z(n14455) );
  IV U17784 ( .A(n14404), .Z(n14440) );
  XOR U17785 ( .A(n14458), .B(n14459), .Z(n14404) );
  XNOR U17786 ( .A(n14399), .B(n14460), .Z(n14459) );
  IV U17787 ( .A(n14402), .Z(n14460) );
  XOR U17788 ( .A(n14461), .B(n14462), .Z(n14402) );
  ANDN U17789 ( .B(n14463), .A(n14464), .Z(n14461) );
  XOR U17790 ( .A(n14462), .B(n14465), .Z(n14463) );
  XNOR U17791 ( .A(n14466), .B(n14467), .Z(n14399) );
  ANDN U17792 ( .B(n14468), .A(n14469), .Z(n14466) );
  XOR U17793 ( .A(n14467), .B(n14470), .Z(n14468) );
  IV U17794 ( .A(n14398), .Z(n14458) );
  XOR U17795 ( .A(n14396), .B(n14471), .Z(n14398) );
  XOR U17796 ( .A(n14472), .B(n14473), .Z(n14471) );
  ANDN U17797 ( .B(n14474), .A(n14475), .Z(n14472) );
  XOR U17798 ( .A(n14476), .B(n14473), .Z(n14474) );
  IV U17799 ( .A(n14400), .Z(n14396) );
  XOR U17800 ( .A(n14477), .B(n14478), .Z(n14400) );
  ANDN U17801 ( .B(n14479), .A(n14480), .Z(n14477) );
  XOR U17802 ( .A(n14481), .B(n14478), .Z(n14479) );
  XOR U17803 ( .A(n14482), .B(n14483), .Z(n14412) );
  XOR U17804 ( .A(n14430), .B(n14484), .Z(n14483) );
  IV U17805 ( .A(n14410), .Z(n14484) );
  XOR U17806 ( .A(n14485), .B(n14486), .Z(n14410) );
  ANDN U17807 ( .B(n14487), .A(n14488), .Z(n14485) );
  XOR U17808 ( .A(n14486), .B(n14489), .Z(n14487) );
  XOR U17809 ( .A(n14490), .B(n14418), .Z(n14430) );
  XOR U17810 ( .A(n14491), .B(n14492), .Z(n14418) );
  ANDN U17811 ( .B(n14493), .A(n14494), .Z(n14491) );
  XOR U17812 ( .A(n14492), .B(n14495), .Z(n14493) );
  IV U17813 ( .A(n14417), .Z(n14490) );
  XOR U17814 ( .A(n14496), .B(n14497), .Z(n14417) );
  XOR U17815 ( .A(n14498), .B(n14499), .Z(n14497) );
  ANDN U17816 ( .B(n14500), .A(n14501), .Z(n14498) );
  XOR U17817 ( .A(n14502), .B(n14499), .Z(n14500) );
  IV U17818 ( .A(n14415), .Z(n14496) );
  XOR U17819 ( .A(n14503), .B(n14504), .Z(n14415) );
  ANDN U17820 ( .B(n14505), .A(n14506), .Z(n14503) );
  XOR U17821 ( .A(n14504), .B(n14507), .Z(n14505) );
  IV U17822 ( .A(n14429), .Z(n14482) );
  XOR U17823 ( .A(n14508), .B(n14509), .Z(n14429) );
  XNOR U17824 ( .A(n14424), .B(n14510), .Z(n14509) );
  IV U17825 ( .A(n14427), .Z(n14510) );
  XOR U17826 ( .A(n14511), .B(n14512), .Z(n14427) );
  ANDN U17827 ( .B(n14513), .A(n14514), .Z(n14511) );
  XOR U17828 ( .A(n14515), .B(n14512), .Z(n14513) );
  XNOR U17829 ( .A(n14516), .B(n14517), .Z(n14424) );
  ANDN U17830 ( .B(n14518), .A(n14519), .Z(n14516) );
  XOR U17831 ( .A(n14517), .B(n14520), .Z(n14518) );
  IV U17832 ( .A(n14423), .Z(n14508) );
  XOR U17833 ( .A(n14421), .B(n14521), .Z(n14423) );
  XOR U17834 ( .A(n14522), .B(n14523), .Z(n14521) );
  ANDN U17835 ( .B(n14524), .A(n14525), .Z(n14522) );
  XOR U17836 ( .A(n14526), .B(n14523), .Z(n14524) );
  IV U17837 ( .A(n14425), .Z(n14421) );
  XOR U17838 ( .A(n14527), .B(n14528), .Z(n14425) );
  ANDN U17839 ( .B(n14529), .A(n14530), .Z(n14527) );
  XOR U17840 ( .A(n14531), .B(n14528), .Z(n14529) );
  IV U17841 ( .A(n14435), .Z(n14439) );
  XOR U17842 ( .A(n14435), .B(n14338), .Z(n14437) );
  XOR U17843 ( .A(n14532), .B(n14533), .Z(n14338) );
  AND U17844 ( .A(n56), .B(n14534), .Z(n14532) );
  XOR U17845 ( .A(n14535), .B(n14533), .Z(n14534) );
  NANDN U17846 ( .A(n14340), .B(n14342), .Z(n14435) );
  XOR U17847 ( .A(n14536), .B(n14537), .Z(n14342) );
  AND U17848 ( .A(n56), .B(n14538), .Z(n14536) );
  XOR U17849 ( .A(n14537), .B(n14539), .Z(n14538) );
  XNOR U17850 ( .A(n14540), .B(n14541), .Z(n56) );
  AND U17851 ( .A(n14542), .B(n14543), .Z(n14540) );
  XOR U17852 ( .A(n14541), .B(n14353), .Z(n14543) );
  XNOR U17853 ( .A(n14544), .B(n14545), .Z(n14353) );
  ANDN U17854 ( .B(n14546), .A(n14547), .Z(n14544) );
  XOR U17855 ( .A(n14545), .B(n14548), .Z(n14546) );
  XNOR U17856 ( .A(n14541), .B(n14355), .Z(n14542) );
  XOR U17857 ( .A(n14549), .B(n14550), .Z(n14355) );
  AND U17858 ( .A(n60), .B(n14551), .Z(n14549) );
  XOR U17859 ( .A(n14552), .B(n14550), .Z(n14551) );
  XOR U17860 ( .A(n14553), .B(n14554), .Z(n14541) );
  AND U17861 ( .A(n14555), .B(n14556), .Z(n14553) );
  XOR U17862 ( .A(n14554), .B(n14380), .Z(n14556) );
  XOR U17863 ( .A(n14547), .B(n14548), .Z(n14380) );
  XNOR U17864 ( .A(n14557), .B(n14558), .Z(n14548) );
  ANDN U17865 ( .B(n14559), .A(n14560), .Z(n14557) );
  XOR U17866 ( .A(n14561), .B(n14562), .Z(n14559) );
  XOR U17867 ( .A(n14563), .B(n14564), .Z(n14547) );
  XNOR U17868 ( .A(n14565), .B(n14566), .Z(n14564) );
  ANDN U17869 ( .B(n14567), .A(n14568), .Z(n14565) );
  XNOR U17870 ( .A(n14569), .B(n14570), .Z(n14567) );
  IV U17871 ( .A(n14545), .Z(n14563) );
  XOR U17872 ( .A(n14571), .B(n14572), .Z(n14545) );
  ANDN U17873 ( .B(n14573), .A(n14574), .Z(n14571) );
  XOR U17874 ( .A(n14572), .B(n14575), .Z(n14573) );
  XNOR U17875 ( .A(n14554), .B(n14382), .Z(n14555) );
  XOR U17876 ( .A(n14576), .B(n14577), .Z(n14382) );
  AND U17877 ( .A(n60), .B(n14578), .Z(n14576) );
  XOR U17878 ( .A(n14579), .B(n14577), .Z(n14578) );
  XNOR U17879 ( .A(n14580), .B(n14581), .Z(n14554) );
  AND U17880 ( .A(n14582), .B(n14583), .Z(n14580) );
  XNOR U17881 ( .A(n14581), .B(n14432), .Z(n14583) );
  XOR U17882 ( .A(n14574), .B(n14575), .Z(n14432) );
  XOR U17883 ( .A(n14584), .B(n14562), .Z(n14575) );
  XNOR U17884 ( .A(n14585), .B(n14586), .Z(n14562) );
  ANDN U17885 ( .B(n14587), .A(n14588), .Z(n14585) );
  XOR U17886 ( .A(n14589), .B(n14590), .Z(n14587) );
  IV U17887 ( .A(n14560), .Z(n14584) );
  XOR U17888 ( .A(n14558), .B(n14591), .Z(n14560) );
  XNOR U17889 ( .A(n14592), .B(n14593), .Z(n14591) );
  ANDN U17890 ( .B(n14594), .A(n14595), .Z(n14592) );
  XNOR U17891 ( .A(n14596), .B(n14597), .Z(n14594) );
  IV U17892 ( .A(n14561), .Z(n14558) );
  XOR U17893 ( .A(n14598), .B(n14599), .Z(n14561) );
  ANDN U17894 ( .B(n14600), .A(n14601), .Z(n14598) );
  XOR U17895 ( .A(n14599), .B(n14602), .Z(n14600) );
  XOR U17896 ( .A(n14603), .B(n14604), .Z(n14574) );
  XNOR U17897 ( .A(n14569), .B(n14605), .Z(n14604) );
  IV U17898 ( .A(n14572), .Z(n14605) );
  XOR U17899 ( .A(n14606), .B(n14607), .Z(n14572) );
  ANDN U17900 ( .B(n14608), .A(n14609), .Z(n14606) );
  XOR U17901 ( .A(n14607), .B(n14610), .Z(n14608) );
  XNOR U17902 ( .A(n14611), .B(n14612), .Z(n14569) );
  ANDN U17903 ( .B(n14613), .A(n14614), .Z(n14611) );
  XOR U17904 ( .A(n14612), .B(n14615), .Z(n14613) );
  IV U17905 ( .A(n14568), .Z(n14603) );
  XOR U17906 ( .A(n14566), .B(n14616), .Z(n14568) );
  XNOR U17907 ( .A(n14617), .B(n14618), .Z(n14616) );
  ANDN U17908 ( .B(n14619), .A(n14620), .Z(n14617) );
  XNOR U17909 ( .A(n14621), .B(n14622), .Z(n14619) );
  IV U17910 ( .A(n14570), .Z(n14566) );
  XOR U17911 ( .A(n14623), .B(n14624), .Z(n14570) );
  ANDN U17912 ( .B(n14625), .A(n14626), .Z(n14623) );
  XOR U17913 ( .A(n14627), .B(n14624), .Z(n14625) );
  XOR U17914 ( .A(n14581), .B(n14434), .Z(n14582) );
  XOR U17915 ( .A(n14628), .B(n14629), .Z(n14434) );
  AND U17916 ( .A(n60), .B(n14630), .Z(n14628) );
  XOR U17917 ( .A(n14631), .B(n14629), .Z(n14630) );
  XNOR U17918 ( .A(n14632), .B(n14633), .Z(n14581) );
  NAND U17919 ( .A(n14634), .B(n14635), .Z(n14633) );
  XOR U17920 ( .A(n14636), .B(n14533), .Z(n14635) );
  XOR U17921 ( .A(n14609), .B(n14610), .Z(n14533) );
  XOR U17922 ( .A(n14637), .B(n14602), .Z(n14610) );
  XOR U17923 ( .A(n14638), .B(n14590), .Z(n14602) );
  XOR U17924 ( .A(n14639), .B(n14640), .Z(n14590) );
  ANDN U17925 ( .B(n14641), .A(n14642), .Z(n14639) );
  XOR U17926 ( .A(n14640), .B(n14643), .Z(n14641) );
  IV U17927 ( .A(n14588), .Z(n14638) );
  XOR U17928 ( .A(n14586), .B(n14644), .Z(n14588) );
  XOR U17929 ( .A(n14645), .B(n14646), .Z(n14644) );
  ANDN U17930 ( .B(n14647), .A(n14648), .Z(n14645) );
  XOR U17931 ( .A(n14649), .B(n14646), .Z(n14647) );
  IV U17932 ( .A(n14589), .Z(n14586) );
  XOR U17933 ( .A(n14650), .B(n14651), .Z(n14589) );
  ANDN U17934 ( .B(n14652), .A(n14653), .Z(n14650) );
  XOR U17935 ( .A(n14651), .B(n14654), .Z(n14652) );
  IV U17936 ( .A(n14601), .Z(n14637) );
  XOR U17937 ( .A(n14655), .B(n14656), .Z(n14601) );
  XNOR U17938 ( .A(n14596), .B(n14657), .Z(n14656) );
  IV U17939 ( .A(n14599), .Z(n14657) );
  XOR U17940 ( .A(n14658), .B(n14659), .Z(n14599) );
  ANDN U17941 ( .B(n14660), .A(n14661), .Z(n14658) );
  XOR U17942 ( .A(n14659), .B(n14662), .Z(n14660) );
  XNOR U17943 ( .A(n14663), .B(n14664), .Z(n14596) );
  ANDN U17944 ( .B(n14665), .A(n14666), .Z(n14663) );
  XOR U17945 ( .A(n14664), .B(n14667), .Z(n14665) );
  IV U17946 ( .A(n14595), .Z(n14655) );
  XOR U17947 ( .A(n14593), .B(n14668), .Z(n14595) );
  XOR U17948 ( .A(n14669), .B(n14670), .Z(n14668) );
  ANDN U17949 ( .B(n14671), .A(n14672), .Z(n14669) );
  XOR U17950 ( .A(n14673), .B(n14670), .Z(n14671) );
  IV U17951 ( .A(n14597), .Z(n14593) );
  XOR U17952 ( .A(n14674), .B(n14675), .Z(n14597) );
  ANDN U17953 ( .B(n14676), .A(n14677), .Z(n14674) );
  XOR U17954 ( .A(n14678), .B(n14675), .Z(n14676) );
  XOR U17955 ( .A(n14679), .B(n14680), .Z(n14609) );
  XOR U17956 ( .A(n14627), .B(n14681), .Z(n14680) );
  IV U17957 ( .A(n14607), .Z(n14681) );
  XOR U17958 ( .A(n14682), .B(n14683), .Z(n14607) );
  ANDN U17959 ( .B(n14684), .A(n14685), .Z(n14682) );
  XOR U17960 ( .A(n14683), .B(n14686), .Z(n14684) );
  XOR U17961 ( .A(n14687), .B(n14615), .Z(n14627) );
  XOR U17962 ( .A(n14688), .B(n14689), .Z(n14615) );
  ANDN U17963 ( .B(n14690), .A(n14691), .Z(n14688) );
  XOR U17964 ( .A(n14689), .B(n14692), .Z(n14690) );
  IV U17965 ( .A(n14614), .Z(n14687) );
  XOR U17966 ( .A(n14693), .B(n14694), .Z(n14614) );
  XOR U17967 ( .A(n14695), .B(n14696), .Z(n14694) );
  ANDN U17968 ( .B(n14697), .A(n14698), .Z(n14695) );
  XOR U17969 ( .A(n14699), .B(n14696), .Z(n14697) );
  IV U17970 ( .A(n14612), .Z(n14693) );
  XOR U17971 ( .A(n14700), .B(n14701), .Z(n14612) );
  ANDN U17972 ( .B(n14702), .A(n14703), .Z(n14700) );
  XOR U17973 ( .A(n14701), .B(n14704), .Z(n14702) );
  IV U17974 ( .A(n14626), .Z(n14679) );
  XOR U17975 ( .A(n14705), .B(n14706), .Z(n14626) );
  XNOR U17976 ( .A(n14621), .B(n14707), .Z(n14706) );
  IV U17977 ( .A(n14624), .Z(n14707) );
  XOR U17978 ( .A(n14708), .B(n14709), .Z(n14624) );
  ANDN U17979 ( .B(n14710), .A(n14711), .Z(n14708) );
  XOR U17980 ( .A(n14712), .B(n14709), .Z(n14710) );
  XNOR U17981 ( .A(n14713), .B(n14714), .Z(n14621) );
  ANDN U17982 ( .B(n14715), .A(n14716), .Z(n14713) );
  XOR U17983 ( .A(n14714), .B(n14717), .Z(n14715) );
  IV U17984 ( .A(n14620), .Z(n14705) );
  XOR U17985 ( .A(n14618), .B(n14718), .Z(n14620) );
  XOR U17986 ( .A(n14719), .B(n14720), .Z(n14718) );
  ANDN U17987 ( .B(n14721), .A(n14722), .Z(n14719) );
  XOR U17988 ( .A(n14723), .B(n14720), .Z(n14721) );
  IV U17989 ( .A(n14622), .Z(n14618) );
  XOR U17990 ( .A(n14724), .B(n14725), .Z(n14622) );
  ANDN U17991 ( .B(n14726), .A(n14727), .Z(n14724) );
  XOR U17992 ( .A(n14728), .B(n14725), .Z(n14726) );
  IV U17993 ( .A(n14632), .Z(n14636) );
  XOR U17994 ( .A(n14632), .B(n14535), .Z(n14634) );
  XOR U17995 ( .A(n14729), .B(n14730), .Z(n14535) );
  AND U17996 ( .A(n60), .B(n14731), .Z(n14729) );
  XOR U17997 ( .A(n14732), .B(n14730), .Z(n14731) );
  NANDN U17998 ( .A(n14537), .B(n14539), .Z(n14632) );
  XOR U17999 ( .A(n14733), .B(n14734), .Z(n14539) );
  AND U18000 ( .A(n60), .B(n14735), .Z(n14733) );
  XOR U18001 ( .A(n14734), .B(n14736), .Z(n14735) );
  XNOR U18002 ( .A(n14737), .B(n14738), .Z(n60) );
  AND U18003 ( .A(n14739), .B(n14740), .Z(n14737) );
  XOR U18004 ( .A(n14738), .B(n14550), .Z(n14740) );
  XNOR U18005 ( .A(n14741), .B(n14742), .Z(n14550) );
  ANDN U18006 ( .B(n14743), .A(n14744), .Z(n14741) );
  XOR U18007 ( .A(n14742), .B(n14745), .Z(n14743) );
  XNOR U18008 ( .A(n14738), .B(n14552), .Z(n14739) );
  XOR U18009 ( .A(n14746), .B(n14747), .Z(n14552) );
  AND U18010 ( .A(n64), .B(n14748), .Z(n14746) );
  XOR U18011 ( .A(n14749), .B(n14747), .Z(n14748) );
  XOR U18012 ( .A(n14750), .B(n14751), .Z(n14738) );
  AND U18013 ( .A(n14752), .B(n14753), .Z(n14750) );
  XOR U18014 ( .A(n14751), .B(n14577), .Z(n14753) );
  XOR U18015 ( .A(n14744), .B(n14745), .Z(n14577) );
  XNOR U18016 ( .A(n14754), .B(n14755), .Z(n14745) );
  ANDN U18017 ( .B(n14756), .A(n14757), .Z(n14754) );
  XOR U18018 ( .A(n14758), .B(n14759), .Z(n14756) );
  XOR U18019 ( .A(n14760), .B(n14761), .Z(n14744) );
  XNOR U18020 ( .A(n14762), .B(n14763), .Z(n14761) );
  ANDN U18021 ( .B(n14764), .A(n14765), .Z(n14762) );
  XNOR U18022 ( .A(n14766), .B(n14767), .Z(n14764) );
  IV U18023 ( .A(n14742), .Z(n14760) );
  XOR U18024 ( .A(n14768), .B(n14769), .Z(n14742) );
  ANDN U18025 ( .B(n14770), .A(n14771), .Z(n14768) );
  XOR U18026 ( .A(n14769), .B(n14772), .Z(n14770) );
  XNOR U18027 ( .A(n14751), .B(n14579), .Z(n14752) );
  XOR U18028 ( .A(n14773), .B(n14774), .Z(n14579) );
  AND U18029 ( .A(n64), .B(n14775), .Z(n14773) );
  XOR U18030 ( .A(n14776), .B(n14774), .Z(n14775) );
  XNOR U18031 ( .A(n14777), .B(n14778), .Z(n14751) );
  AND U18032 ( .A(n14779), .B(n14780), .Z(n14777) );
  XNOR U18033 ( .A(n14778), .B(n14629), .Z(n14780) );
  XOR U18034 ( .A(n14771), .B(n14772), .Z(n14629) );
  XOR U18035 ( .A(n14781), .B(n14759), .Z(n14772) );
  XNOR U18036 ( .A(n14782), .B(n14783), .Z(n14759) );
  ANDN U18037 ( .B(n14784), .A(n14785), .Z(n14782) );
  XOR U18038 ( .A(n14786), .B(n14787), .Z(n14784) );
  IV U18039 ( .A(n14757), .Z(n14781) );
  XOR U18040 ( .A(n14755), .B(n14788), .Z(n14757) );
  XNOR U18041 ( .A(n14789), .B(n14790), .Z(n14788) );
  ANDN U18042 ( .B(n14791), .A(n14792), .Z(n14789) );
  XNOR U18043 ( .A(n14793), .B(n14794), .Z(n14791) );
  IV U18044 ( .A(n14758), .Z(n14755) );
  XOR U18045 ( .A(n14795), .B(n14796), .Z(n14758) );
  ANDN U18046 ( .B(n14797), .A(n14798), .Z(n14795) );
  XOR U18047 ( .A(n14796), .B(n14799), .Z(n14797) );
  XOR U18048 ( .A(n14800), .B(n14801), .Z(n14771) );
  XNOR U18049 ( .A(n14766), .B(n14802), .Z(n14801) );
  IV U18050 ( .A(n14769), .Z(n14802) );
  XOR U18051 ( .A(n14803), .B(n14804), .Z(n14769) );
  ANDN U18052 ( .B(n14805), .A(n14806), .Z(n14803) );
  XOR U18053 ( .A(n14804), .B(n14807), .Z(n14805) );
  XNOR U18054 ( .A(n14808), .B(n14809), .Z(n14766) );
  ANDN U18055 ( .B(n14810), .A(n14811), .Z(n14808) );
  XOR U18056 ( .A(n14809), .B(n14812), .Z(n14810) );
  IV U18057 ( .A(n14765), .Z(n14800) );
  XOR U18058 ( .A(n14763), .B(n14813), .Z(n14765) );
  XNOR U18059 ( .A(n14814), .B(n14815), .Z(n14813) );
  ANDN U18060 ( .B(n14816), .A(n14817), .Z(n14814) );
  XNOR U18061 ( .A(n14818), .B(n14819), .Z(n14816) );
  IV U18062 ( .A(n14767), .Z(n14763) );
  XOR U18063 ( .A(n14820), .B(n14821), .Z(n14767) );
  ANDN U18064 ( .B(n14822), .A(n14823), .Z(n14820) );
  XOR U18065 ( .A(n14824), .B(n14821), .Z(n14822) );
  XOR U18066 ( .A(n14778), .B(n14631), .Z(n14779) );
  XOR U18067 ( .A(n14825), .B(n14826), .Z(n14631) );
  AND U18068 ( .A(n64), .B(n14827), .Z(n14825) );
  XOR U18069 ( .A(n14828), .B(n14826), .Z(n14827) );
  XNOR U18070 ( .A(n14829), .B(n14830), .Z(n14778) );
  NAND U18071 ( .A(n14831), .B(n14832), .Z(n14830) );
  XOR U18072 ( .A(n14833), .B(n14730), .Z(n14832) );
  XOR U18073 ( .A(n14806), .B(n14807), .Z(n14730) );
  XOR U18074 ( .A(n14834), .B(n14799), .Z(n14807) );
  XOR U18075 ( .A(n14835), .B(n14787), .Z(n14799) );
  XOR U18076 ( .A(n14836), .B(n14837), .Z(n14787) );
  ANDN U18077 ( .B(n14838), .A(n14839), .Z(n14836) );
  XOR U18078 ( .A(n14837), .B(n14840), .Z(n14838) );
  IV U18079 ( .A(n14785), .Z(n14835) );
  XOR U18080 ( .A(n14783), .B(n14841), .Z(n14785) );
  XOR U18081 ( .A(n14842), .B(n14843), .Z(n14841) );
  ANDN U18082 ( .B(n14844), .A(n14845), .Z(n14842) );
  XOR U18083 ( .A(n14846), .B(n14843), .Z(n14844) );
  IV U18084 ( .A(n14786), .Z(n14783) );
  XOR U18085 ( .A(n14847), .B(n14848), .Z(n14786) );
  ANDN U18086 ( .B(n14849), .A(n14850), .Z(n14847) );
  XOR U18087 ( .A(n14848), .B(n14851), .Z(n14849) );
  IV U18088 ( .A(n14798), .Z(n14834) );
  XOR U18089 ( .A(n14852), .B(n14853), .Z(n14798) );
  XNOR U18090 ( .A(n14793), .B(n14854), .Z(n14853) );
  IV U18091 ( .A(n14796), .Z(n14854) );
  XOR U18092 ( .A(n14855), .B(n14856), .Z(n14796) );
  ANDN U18093 ( .B(n14857), .A(n14858), .Z(n14855) );
  XOR U18094 ( .A(n14856), .B(n14859), .Z(n14857) );
  XNOR U18095 ( .A(n14860), .B(n14861), .Z(n14793) );
  ANDN U18096 ( .B(n14862), .A(n14863), .Z(n14860) );
  XOR U18097 ( .A(n14861), .B(n14864), .Z(n14862) );
  IV U18098 ( .A(n14792), .Z(n14852) );
  XOR U18099 ( .A(n14790), .B(n14865), .Z(n14792) );
  XOR U18100 ( .A(n14866), .B(n14867), .Z(n14865) );
  ANDN U18101 ( .B(n14868), .A(n14869), .Z(n14866) );
  XOR U18102 ( .A(n14870), .B(n14867), .Z(n14868) );
  IV U18103 ( .A(n14794), .Z(n14790) );
  XOR U18104 ( .A(n14871), .B(n14872), .Z(n14794) );
  ANDN U18105 ( .B(n14873), .A(n14874), .Z(n14871) );
  XOR U18106 ( .A(n14875), .B(n14872), .Z(n14873) );
  XOR U18107 ( .A(n14876), .B(n14877), .Z(n14806) );
  XOR U18108 ( .A(n14824), .B(n14878), .Z(n14877) );
  IV U18109 ( .A(n14804), .Z(n14878) );
  XOR U18110 ( .A(n14879), .B(n14880), .Z(n14804) );
  ANDN U18111 ( .B(n14881), .A(n14882), .Z(n14879) );
  XOR U18112 ( .A(n14880), .B(n14883), .Z(n14881) );
  XOR U18113 ( .A(n14884), .B(n14812), .Z(n14824) );
  XOR U18114 ( .A(n14885), .B(n14886), .Z(n14812) );
  ANDN U18115 ( .B(n14887), .A(n14888), .Z(n14885) );
  XOR U18116 ( .A(n14886), .B(n14889), .Z(n14887) );
  IV U18117 ( .A(n14811), .Z(n14884) );
  XOR U18118 ( .A(n14890), .B(n14891), .Z(n14811) );
  XOR U18119 ( .A(n14892), .B(n14893), .Z(n14891) );
  ANDN U18120 ( .B(n14894), .A(n14895), .Z(n14892) );
  XOR U18121 ( .A(n14896), .B(n14893), .Z(n14894) );
  IV U18122 ( .A(n14809), .Z(n14890) );
  XOR U18123 ( .A(n14897), .B(n14898), .Z(n14809) );
  ANDN U18124 ( .B(n14899), .A(n14900), .Z(n14897) );
  XOR U18125 ( .A(n14898), .B(n14901), .Z(n14899) );
  IV U18126 ( .A(n14823), .Z(n14876) );
  XOR U18127 ( .A(n14902), .B(n14903), .Z(n14823) );
  XNOR U18128 ( .A(n14818), .B(n14904), .Z(n14903) );
  IV U18129 ( .A(n14821), .Z(n14904) );
  XOR U18130 ( .A(n14905), .B(n14906), .Z(n14821) );
  ANDN U18131 ( .B(n14907), .A(n14908), .Z(n14905) );
  XOR U18132 ( .A(n14909), .B(n14906), .Z(n14907) );
  XNOR U18133 ( .A(n14910), .B(n14911), .Z(n14818) );
  ANDN U18134 ( .B(n14912), .A(n14913), .Z(n14910) );
  XOR U18135 ( .A(n14911), .B(n14914), .Z(n14912) );
  IV U18136 ( .A(n14817), .Z(n14902) );
  XOR U18137 ( .A(n14815), .B(n14915), .Z(n14817) );
  XOR U18138 ( .A(n14916), .B(n14917), .Z(n14915) );
  ANDN U18139 ( .B(n14918), .A(n14919), .Z(n14916) );
  XOR U18140 ( .A(n14920), .B(n14917), .Z(n14918) );
  IV U18141 ( .A(n14819), .Z(n14815) );
  XOR U18142 ( .A(n14921), .B(n14922), .Z(n14819) );
  ANDN U18143 ( .B(n14923), .A(n14924), .Z(n14921) );
  XOR U18144 ( .A(n14925), .B(n14922), .Z(n14923) );
  IV U18145 ( .A(n14829), .Z(n14833) );
  XOR U18146 ( .A(n14829), .B(n14732), .Z(n14831) );
  XOR U18147 ( .A(n14926), .B(n14927), .Z(n14732) );
  AND U18148 ( .A(n64), .B(n14928), .Z(n14926) );
  XOR U18149 ( .A(n14929), .B(n14927), .Z(n14928) );
  NANDN U18150 ( .A(n14734), .B(n14736), .Z(n14829) );
  XOR U18151 ( .A(n14930), .B(n14931), .Z(n14736) );
  AND U18152 ( .A(n64), .B(n14932), .Z(n14930) );
  XOR U18153 ( .A(n14931), .B(n14933), .Z(n14932) );
  XNOR U18154 ( .A(n14934), .B(n14935), .Z(n64) );
  AND U18155 ( .A(n14936), .B(n14937), .Z(n14934) );
  XOR U18156 ( .A(n14935), .B(n14747), .Z(n14937) );
  XNOR U18157 ( .A(n14938), .B(n14939), .Z(n14747) );
  ANDN U18158 ( .B(n14940), .A(n14941), .Z(n14938) );
  XOR U18159 ( .A(n14939), .B(n14942), .Z(n14940) );
  XNOR U18160 ( .A(n14935), .B(n14749), .Z(n14936) );
  XOR U18161 ( .A(n14943), .B(n14944), .Z(n14749) );
  AND U18162 ( .A(n68), .B(n14945), .Z(n14943) );
  XOR U18163 ( .A(n14946), .B(n14944), .Z(n14945) );
  XOR U18164 ( .A(n14947), .B(n14948), .Z(n14935) );
  AND U18165 ( .A(n14949), .B(n14950), .Z(n14947) );
  XOR U18166 ( .A(n14948), .B(n14774), .Z(n14950) );
  XOR U18167 ( .A(n14941), .B(n14942), .Z(n14774) );
  XNOR U18168 ( .A(n14951), .B(n14952), .Z(n14942) );
  ANDN U18169 ( .B(n14953), .A(n14954), .Z(n14951) );
  XOR U18170 ( .A(n14955), .B(n14956), .Z(n14953) );
  XOR U18171 ( .A(n14957), .B(n14958), .Z(n14941) );
  XNOR U18172 ( .A(n14959), .B(n14960), .Z(n14958) );
  ANDN U18173 ( .B(n14961), .A(n14962), .Z(n14959) );
  XNOR U18174 ( .A(n14963), .B(n14964), .Z(n14961) );
  IV U18175 ( .A(n14939), .Z(n14957) );
  XOR U18176 ( .A(n14965), .B(n14966), .Z(n14939) );
  ANDN U18177 ( .B(n14967), .A(n14968), .Z(n14965) );
  XOR U18178 ( .A(n14966), .B(n14969), .Z(n14967) );
  XNOR U18179 ( .A(n14948), .B(n14776), .Z(n14949) );
  XOR U18180 ( .A(n14970), .B(n14971), .Z(n14776) );
  AND U18181 ( .A(n68), .B(n14972), .Z(n14970) );
  XOR U18182 ( .A(n14973), .B(n14971), .Z(n14972) );
  XNOR U18183 ( .A(n14974), .B(n14975), .Z(n14948) );
  AND U18184 ( .A(n14976), .B(n14977), .Z(n14974) );
  XNOR U18185 ( .A(n14975), .B(n14826), .Z(n14977) );
  XOR U18186 ( .A(n14968), .B(n14969), .Z(n14826) );
  XOR U18187 ( .A(n14978), .B(n14956), .Z(n14969) );
  XNOR U18188 ( .A(n14979), .B(n14980), .Z(n14956) );
  ANDN U18189 ( .B(n14981), .A(n14982), .Z(n14979) );
  XOR U18190 ( .A(n14983), .B(n14984), .Z(n14981) );
  IV U18191 ( .A(n14954), .Z(n14978) );
  XOR U18192 ( .A(n14952), .B(n14985), .Z(n14954) );
  XNOR U18193 ( .A(n14986), .B(n14987), .Z(n14985) );
  ANDN U18194 ( .B(n14988), .A(n14989), .Z(n14986) );
  XNOR U18195 ( .A(n14990), .B(n14991), .Z(n14988) );
  IV U18196 ( .A(n14955), .Z(n14952) );
  XOR U18197 ( .A(n14992), .B(n14993), .Z(n14955) );
  ANDN U18198 ( .B(n14994), .A(n14995), .Z(n14992) );
  XOR U18199 ( .A(n14993), .B(n14996), .Z(n14994) );
  XOR U18200 ( .A(n14997), .B(n14998), .Z(n14968) );
  XNOR U18201 ( .A(n14963), .B(n14999), .Z(n14998) );
  IV U18202 ( .A(n14966), .Z(n14999) );
  XOR U18203 ( .A(n15000), .B(n15001), .Z(n14966) );
  ANDN U18204 ( .B(n15002), .A(n15003), .Z(n15000) );
  XOR U18205 ( .A(n15001), .B(n15004), .Z(n15002) );
  XNOR U18206 ( .A(n15005), .B(n15006), .Z(n14963) );
  ANDN U18207 ( .B(n15007), .A(n15008), .Z(n15005) );
  XOR U18208 ( .A(n15006), .B(n15009), .Z(n15007) );
  IV U18209 ( .A(n14962), .Z(n14997) );
  XOR U18210 ( .A(n14960), .B(n15010), .Z(n14962) );
  XNOR U18211 ( .A(n15011), .B(n15012), .Z(n15010) );
  ANDN U18212 ( .B(n15013), .A(n15014), .Z(n15011) );
  XNOR U18213 ( .A(n15015), .B(n15016), .Z(n15013) );
  IV U18214 ( .A(n14964), .Z(n14960) );
  XOR U18215 ( .A(n15017), .B(n15018), .Z(n14964) );
  ANDN U18216 ( .B(n15019), .A(n15020), .Z(n15017) );
  XOR U18217 ( .A(n15021), .B(n15018), .Z(n15019) );
  XOR U18218 ( .A(n14975), .B(n14828), .Z(n14976) );
  XOR U18219 ( .A(n15022), .B(n15023), .Z(n14828) );
  AND U18220 ( .A(n68), .B(n15024), .Z(n15022) );
  XOR U18221 ( .A(n15025), .B(n15023), .Z(n15024) );
  XNOR U18222 ( .A(n15026), .B(n15027), .Z(n14975) );
  NAND U18223 ( .A(n15028), .B(n15029), .Z(n15027) );
  XOR U18224 ( .A(n15030), .B(n14927), .Z(n15029) );
  XOR U18225 ( .A(n15003), .B(n15004), .Z(n14927) );
  XOR U18226 ( .A(n15031), .B(n14996), .Z(n15004) );
  XOR U18227 ( .A(n15032), .B(n14984), .Z(n14996) );
  XOR U18228 ( .A(n15033), .B(n15034), .Z(n14984) );
  ANDN U18229 ( .B(n15035), .A(n15036), .Z(n15033) );
  XOR U18230 ( .A(n15034), .B(n15037), .Z(n15035) );
  IV U18231 ( .A(n14982), .Z(n15032) );
  XOR U18232 ( .A(n14980), .B(n15038), .Z(n14982) );
  XOR U18233 ( .A(n15039), .B(n15040), .Z(n15038) );
  ANDN U18234 ( .B(n15041), .A(n15042), .Z(n15039) );
  XOR U18235 ( .A(n15043), .B(n15040), .Z(n15041) );
  IV U18236 ( .A(n14983), .Z(n14980) );
  XOR U18237 ( .A(n15044), .B(n15045), .Z(n14983) );
  ANDN U18238 ( .B(n15046), .A(n15047), .Z(n15044) );
  XOR U18239 ( .A(n15045), .B(n15048), .Z(n15046) );
  IV U18240 ( .A(n14995), .Z(n15031) );
  XOR U18241 ( .A(n15049), .B(n15050), .Z(n14995) );
  XNOR U18242 ( .A(n14990), .B(n15051), .Z(n15050) );
  IV U18243 ( .A(n14993), .Z(n15051) );
  XOR U18244 ( .A(n15052), .B(n15053), .Z(n14993) );
  ANDN U18245 ( .B(n15054), .A(n15055), .Z(n15052) );
  XOR U18246 ( .A(n15053), .B(n15056), .Z(n15054) );
  XNOR U18247 ( .A(n15057), .B(n15058), .Z(n14990) );
  ANDN U18248 ( .B(n15059), .A(n15060), .Z(n15057) );
  XOR U18249 ( .A(n15058), .B(n15061), .Z(n15059) );
  IV U18250 ( .A(n14989), .Z(n15049) );
  XOR U18251 ( .A(n14987), .B(n15062), .Z(n14989) );
  XOR U18252 ( .A(n15063), .B(n15064), .Z(n15062) );
  ANDN U18253 ( .B(n15065), .A(n15066), .Z(n15063) );
  XOR U18254 ( .A(n15067), .B(n15064), .Z(n15065) );
  IV U18255 ( .A(n14991), .Z(n14987) );
  XOR U18256 ( .A(n15068), .B(n15069), .Z(n14991) );
  ANDN U18257 ( .B(n15070), .A(n15071), .Z(n15068) );
  XOR U18258 ( .A(n15072), .B(n15069), .Z(n15070) );
  XOR U18259 ( .A(n15073), .B(n15074), .Z(n15003) );
  XOR U18260 ( .A(n15021), .B(n15075), .Z(n15074) );
  IV U18261 ( .A(n15001), .Z(n15075) );
  XOR U18262 ( .A(n15076), .B(n15077), .Z(n15001) );
  ANDN U18263 ( .B(n15078), .A(n15079), .Z(n15076) );
  XOR U18264 ( .A(n15077), .B(n15080), .Z(n15078) );
  XOR U18265 ( .A(n15081), .B(n15009), .Z(n15021) );
  XOR U18266 ( .A(n15082), .B(n15083), .Z(n15009) );
  ANDN U18267 ( .B(n15084), .A(n15085), .Z(n15082) );
  XOR U18268 ( .A(n15083), .B(n15086), .Z(n15084) );
  IV U18269 ( .A(n15008), .Z(n15081) );
  XOR U18270 ( .A(n15087), .B(n15088), .Z(n15008) );
  XOR U18271 ( .A(n15089), .B(n15090), .Z(n15088) );
  ANDN U18272 ( .B(n15091), .A(n15092), .Z(n15089) );
  XOR U18273 ( .A(n15093), .B(n15090), .Z(n15091) );
  IV U18274 ( .A(n15006), .Z(n15087) );
  XOR U18275 ( .A(n15094), .B(n15095), .Z(n15006) );
  ANDN U18276 ( .B(n15096), .A(n15097), .Z(n15094) );
  XOR U18277 ( .A(n15095), .B(n15098), .Z(n15096) );
  IV U18278 ( .A(n15020), .Z(n15073) );
  XOR U18279 ( .A(n15099), .B(n15100), .Z(n15020) );
  XNOR U18280 ( .A(n15015), .B(n15101), .Z(n15100) );
  IV U18281 ( .A(n15018), .Z(n15101) );
  XOR U18282 ( .A(n15102), .B(n15103), .Z(n15018) );
  ANDN U18283 ( .B(n15104), .A(n15105), .Z(n15102) );
  XOR U18284 ( .A(n15106), .B(n15103), .Z(n15104) );
  XNOR U18285 ( .A(n15107), .B(n15108), .Z(n15015) );
  ANDN U18286 ( .B(n15109), .A(n15110), .Z(n15107) );
  XOR U18287 ( .A(n15108), .B(n15111), .Z(n15109) );
  IV U18288 ( .A(n15014), .Z(n15099) );
  XOR U18289 ( .A(n15012), .B(n15112), .Z(n15014) );
  XOR U18290 ( .A(n15113), .B(n15114), .Z(n15112) );
  ANDN U18291 ( .B(n15115), .A(n15116), .Z(n15113) );
  XOR U18292 ( .A(n15117), .B(n15114), .Z(n15115) );
  IV U18293 ( .A(n15016), .Z(n15012) );
  XOR U18294 ( .A(n15118), .B(n15119), .Z(n15016) );
  ANDN U18295 ( .B(n15120), .A(n15121), .Z(n15118) );
  XOR U18296 ( .A(n15122), .B(n15119), .Z(n15120) );
  IV U18297 ( .A(n15026), .Z(n15030) );
  XOR U18298 ( .A(n15026), .B(n14929), .Z(n15028) );
  XOR U18299 ( .A(n15123), .B(n15124), .Z(n14929) );
  AND U18300 ( .A(n68), .B(n15125), .Z(n15123) );
  XOR U18301 ( .A(n15126), .B(n15124), .Z(n15125) );
  NANDN U18302 ( .A(n14931), .B(n14933), .Z(n15026) );
  XOR U18303 ( .A(n15127), .B(n15128), .Z(n14933) );
  AND U18304 ( .A(n68), .B(n15129), .Z(n15127) );
  XOR U18305 ( .A(n15128), .B(n15130), .Z(n15129) );
  XNOR U18306 ( .A(n15131), .B(n15132), .Z(n68) );
  AND U18307 ( .A(n15133), .B(n15134), .Z(n15131) );
  XOR U18308 ( .A(n15132), .B(n14944), .Z(n15134) );
  XNOR U18309 ( .A(n15135), .B(n15136), .Z(n14944) );
  ANDN U18310 ( .B(n15137), .A(n15138), .Z(n15135) );
  XOR U18311 ( .A(n15136), .B(n15139), .Z(n15137) );
  XNOR U18312 ( .A(n15132), .B(n14946), .Z(n15133) );
  XOR U18313 ( .A(n15140), .B(n15141), .Z(n14946) );
  AND U18314 ( .A(n72), .B(n15142), .Z(n15140) );
  XOR U18315 ( .A(n15143), .B(n15141), .Z(n15142) );
  XOR U18316 ( .A(n15144), .B(n15145), .Z(n15132) );
  AND U18317 ( .A(n15146), .B(n15147), .Z(n15144) );
  XOR U18318 ( .A(n15145), .B(n14971), .Z(n15147) );
  XOR U18319 ( .A(n15138), .B(n15139), .Z(n14971) );
  XNOR U18320 ( .A(n15148), .B(n15149), .Z(n15139) );
  ANDN U18321 ( .B(n15150), .A(n15151), .Z(n15148) );
  XOR U18322 ( .A(n15152), .B(n15153), .Z(n15150) );
  XOR U18323 ( .A(n15154), .B(n15155), .Z(n15138) );
  XNOR U18324 ( .A(n15156), .B(n15157), .Z(n15155) );
  ANDN U18325 ( .B(n15158), .A(n15159), .Z(n15156) );
  XNOR U18326 ( .A(n15160), .B(n15161), .Z(n15158) );
  IV U18327 ( .A(n15136), .Z(n15154) );
  XOR U18328 ( .A(n15162), .B(n15163), .Z(n15136) );
  ANDN U18329 ( .B(n15164), .A(n15165), .Z(n15162) );
  XOR U18330 ( .A(n15163), .B(n15166), .Z(n15164) );
  XNOR U18331 ( .A(n15145), .B(n14973), .Z(n15146) );
  XOR U18332 ( .A(n15167), .B(n15168), .Z(n14973) );
  AND U18333 ( .A(n72), .B(n15169), .Z(n15167) );
  XOR U18334 ( .A(n15170), .B(n15168), .Z(n15169) );
  XNOR U18335 ( .A(n15171), .B(n15172), .Z(n15145) );
  AND U18336 ( .A(n15173), .B(n15174), .Z(n15171) );
  XNOR U18337 ( .A(n15172), .B(n15023), .Z(n15174) );
  XOR U18338 ( .A(n15165), .B(n15166), .Z(n15023) );
  XOR U18339 ( .A(n15175), .B(n15153), .Z(n15166) );
  XNOR U18340 ( .A(n15176), .B(n15177), .Z(n15153) );
  ANDN U18341 ( .B(n15178), .A(n15179), .Z(n15176) );
  XOR U18342 ( .A(n15180), .B(n15181), .Z(n15178) );
  IV U18343 ( .A(n15151), .Z(n15175) );
  XOR U18344 ( .A(n15149), .B(n15182), .Z(n15151) );
  XNOR U18345 ( .A(n15183), .B(n15184), .Z(n15182) );
  ANDN U18346 ( .B(n15185), .A(n15186), .Z(n15183) );
  XNOR U18347 ( .A(n15187), .B(n15188), .Z(n15185) );
  IV U18348 ( .A(n15152), .Z(n15149) );
  XOR U18349 ( .A(n15189), .B(n15190), .Z(n15152) );
  ANDN U18350 ( .B(n15191), .A(n15192), .Z(n15189) );
  XOR U18351 ( .A(n15190), .B(n15193), .Z(n15191) );
  XOR U18352 ( .A(n15194), .B(n15195), .Z(n15165) );
  XNOR U18353 ( .A(n15160), .B(n15196), .Z(n15195) );
  IV U18354 ( .A(n15163), .Z(n15196) );
  XOR U18355 ( .A(n15197), .B(n15198), .Z(n15163) );
  ANDN U18356 ( .B(n15199), .A(n15200), .Z(n15197) );
  XOR U18357 ( .A(n15198), .B(n15201), .Z(n15199) );
  XNOR U18358 ( .A(n15202), .B(n15203), .Z(n15160) );
  ANDN U18359 ( .B(n15204), .A(n15205), .Z(n15202) );
  XOR U18360 ( .A(n15203), .B(n15206), .Z(n15204) );
  IV U18361 ( .A(n15159), .Z(n15194) );
  XOR U18362 ( .A(n15157), .B(n15207), .Z(n15159) );
  XNOR U18363 ( .A(n15208), .B(n15209), .Z(n15207) );
  ANDN U18364 ( .B(n15210), .A(n15211), .Z(n15208) );
  XNOR U18365 ( .A(n15212), .B(n15213), .Z(n15210) );
  IV U18366 ( .A(n15161), .Z(n15157) );
  XOR U18367 ( .A(n15214), .B(n15215), .Z(n15161) );
  ANDN U18368 ( .B(n15216), .A(n15217), .Z(n15214) );
  XOR U18369 ( .A(n15218), .B(n15215), .Z(n15216) );
  XOR U18370 ( .A(n15172), .B(n15025), .Z(n15173) );
  XOR U18371 ( .A(n15219), .B(n15220), .Z(n15025) );
  AND U18372 ( .A(n72), .B(n15221), .Z(n15219) );
  XOR U18373 ( .A(n15222), .B(n15220), .Z(n15221) );
  XNOR U18374 ( .A(n15223), .B(n15224), .Z(n15172) );
  NAND U18375 ( .A(n15225), .B(n15226), .Z(n15224) );
  XOR U18376 ( .A(n15227), .B(n15124), .Z(n15226) );
  XOR U18377 ( .A(n15200), .B(n15201), .Z(n15124) );
  XOR U18378 ( .A(n15228), .B(n15193), .Z(n15201) );
  XOR U18379 ( .A(n15229), .B(n15181), .Z(n15193) );
  XOR U18380 ( .A(n15230), .B(n15231), .Z(n15181) );
  ANDN U18381 ( .B(n15232), .A(n15233), .Z(n15230) );
  XOR U18382 ( .A(n15231), .B(n15234), .Z(n15232) );
  IV U18383 ( .A(n15179), .Z(n15229) );
  XOR U18384 ( .A(n15177), .B(n15235), .Z(n15179) );
  XOR U18385 ( .A(n15236), .B(n15237), .Z(n15235) );
  ANDN U18386 ( .B(n15238), .A(n15239), .Z(n15236) );
  XOR U18387 ( .A(n15240), .B(n15237), .Z(n15238) );
  IV U18388 ( .A(n15180), .Z(n15177) );
  XOR U18389 ( .A(n15241), .B(n15242), .Z(n15180) );
  ANDN U18390 ( .B(n15243), .A(n15244), .Z(n15241) );
  XOR U18391 ( .A(n15242), .B(n15245), .Z(n15243) );
  IV U18392 ( .A(n15192), .Z(n15228) );
  XOR U18393 ( .A(n15246), .B(n15247), .Z(n15192) );
  XNOR U18394 ( .A(n15187), .B(n15248), .Z(n15247) );
  IV U18395 ( .A(n15190), .Z(n15248) );
  XOR U18396 ( .A(n15249), .B(n15250), .Z(n15190) );
  ANDN U18397 ( .B(n15251), .A(n15252), .Z(n15249) );
  XOR U18398 ( .A(n15250), .B(n15253), .Z(n15251) );
  XNOR U18399 ( .A(n15254), .B(n15255), .Z(n15187) );
  ANDN U18400 ( .B(n15256), .A(n15257), .Z(n15254) );
  XOR U18401 ( .A(n15255), .B(n15258), .Z(n15256) );
  IV U18402 ( .A(n15186), .Z(n15246) );
  XOR U18403 ( .A(n15184), .B(n15259), .Z(n15186) );
  XOR U18404 ( .A(n15260), .B(n15261), .Z(n15259) );
  ANDN U18405 ( .B(n15262), .A(n15263), .Z(n15260) );
  XOR U18406 ( .A(n15264), .B(n15261), .Z(n15262) );
  IV U18407 ( .A(n15188), .Z(n15184) );
  XOR U18408 ( .A(n15265), .B(n15266), .Z(n15188) );
  ANDN U18409 ( .B(n15267), .A(n15268), .Z(n15265) );
  XOR U18410 ( .A(n15269), .B(n15266), .Z(n15267) );
  XOR U18411 ( .A(n15270), .B(n15271), .Z(n15200) );
  XOR U18412 ( .A(n15218), .B(n15272), .Z(n15271) );
  IV U18413 ( .A(n15198), .Z(n15272) );
  XOR U18414 ( .A(n15273), .B(n15274), .Z(n15198) );
  ANDN U18415 ( .B(n15275), .A(n15276), .Z(n15273) );
  XOR U18416 ( .A(n15274), .B(n15277), .Z(n15275) );
  XOR U18417 ( .A(n15278), .B(n15206), .Z(n15218) );
  XOR U18418 ( .A(n15279), .B(n15280), .Z(n15206) );
  ANDN U18419 ( .B(n15281), .A(n15282), .Z(n15279) );
  XOR U18420 ( .A(n15280), .B(n15283), .Z(n15281) );
  IV U18421 ( .A(n15205), .Z(n15278) );
  XOR U18422 ( .A(n15284), .B(n15285), .Z(n15205) );
  XOR U18423 ( .A(n15286), .B(n15287), .Z(n15285) );
  ANDN U18424 ( .B(n15288), .A(n15289), .Z(n15286) );
  XOR U18425 ( .A(n15290), .B(n15287), .Z(n15288) );
  IV U18426 ( .A(n15203), .Z(n15284) );
  XOR U18427 ( .A(n15291), .B(n15292), .Z(n15203) );
  ANDN U18428 ( .B(n15293), .A(n15294), .Z(n15291) );
  XOR U18429 ( .A(n15292), .B(n15295), .Z(n15293) );
  IV U18430 ( .A(n15217), .Z(n15270) );
  XOR U18431 ( .A(n15296), .B(n15297), .Z(n15217) );
  XNOR U18432 ( .A(n15212), .B(n15298), .Z(n15297) );
  IV U18433 ( .A(n15215), .Z(n15298) );
  XOR U18434 ( .A(n15299), .B(n15300), .Z(n15215) );
  ANDN U18435 ( .B(n15301), .A(n15302), .Z(n15299) );
  XOR U18436 ( .A(n15303), .B(n15300), .Z(n15301) );
  XNOR U18437 ( .A(n15304), .B(n15305), .Z(n15212) );
  ANDN U18438 ( .B(n15306), .A(n15307), .Z(n15304) );
  XOR U18439 ( .A(n15305), .B(n15308), .Z(n15306) );
  IV U18440 ( .A(n15211), .Z(n15296) );
  XOR U18441 ( .A(n15209), .B(n15309), .Z(n15211) );
  XOR U18442 ( .A(n15310), .B(n15311), .Z(n15309) );
  ANDN U18443 ( .B(n15312), .A(n15313), .Z(n15310) );
  XOR U18444 ( .A(n15314), .B(n15311), .Z(n15312) );
  IV U18445 ( .A(n15213), .Z(n15209) );
  XOR U18446 ( .A(n15315), .B(n15316), .Z(n15213) );
  ANDN U18447 ( .B(n15317), .A(n15318), .Z(n15315) );
  XOR U18448 ( .A(n15319), .B(n15316), .Z(n15317) );
  IV U18449 ( .A(n15223), .Z(n15227) );
  XOR U18450 ( .A(n15223), .B(n15126), .Z(n15225) );
  XOR U18451 ( .A(n15320), .B(n15321), .Z(n15126) );
  AND U18452 ( .A(n72), .B(n15322), .Z(n15320) );
  XOR U18453 ( .A(n15323), .B(n15321), .Z(n15322) );
  NANDN U18454 ( .A(n15128), .B(n15130), .Z(n15223) );
  XOR U18455 ( .A(n15324), .B(n15325), .Z(n15130) );
  AND U18456 ( .A(n72), .B(n15326), .Z(n15324) );
  XOR U18457 ( .A(n15325), .B(n15327), .Z(n15326) );
  XNOR U18458 ( .A(n15328), .B(n15329), .Z(n72) );
  AND U18459 ( .A(n15330), .B(n15331), .Z(n15328) );
  XOR U18460 ( .A(n15329), .B(n15141), .Z(n15331) );
  XNOR U18461 ( .A(n15332), .B(n15333), .Z(n15141) );
  ANDN U18462 ( .B(n15334), .A(n15335), .Z(n15332) );
  XOR U18463 ( .A(n15333), .B(n15336), .Z(n15334) );
  XNOR U18464 ( .A(n15329), .B(n15143), .Z(n15330) );
  XOR U18465 ( .A(n15337), .B(n15338), .Z(n15143) );
  AND U18466 ( .A(n76), .B(n15339), .Z(n15337) );
  XOR U18467 ( .A(n15340), .B(n15338), .Z(n15339) );
  XOR U18468 ( .A(n15341), .B(n15342), .Z(n15329) );
  AND U18469 ( .A(n15343), .B(n15344), .Z(n15341) );
  XOR U18470 ( .A(n15342), .B(n15168), .Z(n15344) );
  XOR U18471 ( .A(n15335), .B(n15336), .Z(n15168) );
  XNOR U18472 ( .A(n15345), .B(n15346), .Z(n15336) );
  ANDN U18473 ( .B(n15347), .A(n15348), .Z(n15345) );
  XOR U18474 ( .A(n15349), .B(n15350), .Z(n15347) );
  XOR U18475 ( .A(n15351), .B(n15352), .Z(n15335) );
  XNOR U18476 ( .A(n15353), .B(n15354), .Z(n15352) );
  ANDN U18477 ( .B(n15355), .A(n15356), .Z(n15353) );
  XNOR U18478 ( .A(n15357), .B(n15358), .Z(n15355) );
  IV U18479 ( .A(n15333), .Z(n15351) );
  XOR U18480 ( .A(n15359), .B(n15360), .Z(n15333) );
  ANDN U18481 ( .B(n15361), .A(n15362), .Z(n15359) );
  XOR U18482 ( .A(n15360), .B(n15363), .Z(n15361) );
  XNOR U18483 ( .A(n15342), .B(n15170), .Z(n15343) );
  XOR U18484 ( .A(n15364), .B(n15365), .Z(n15170) );
  AND U18485 ( .A(n76), .B(n15366), .Z(n15364) );
  XOR U18486 ( .A(n15367), .B(n15365), .Z(n15366) );
  XNOR U18487 ( .A(n15368), .B(n15369), .Z(n15342) );
  AND U18488 ( .A(n15370), .B(n15371), .Z(n15368) );
  XNOR U18489 ( .A(n15369), .B(n15220), .Z(n15371) );
  XOR U18490 ( .A(n15362), .B(n15363), .Z(n15220) );
  XOR U18491 ( .A(n15372), .B(n15350), .Z(n15363) );
  XNOR U18492 ( .A(n15373), .B(n15374), .Z(n15350) );
  ANDN U18493 ( .B(n15375), .A(n15376), .Z(n15373) );
  XOR U18494 ( .A(n15377), .B(n15378), .Z(n15375) );
  IV U18495 ( .A(n15348), .Z(n15372) );
  XOR U18496 ( .A(n15346), .B(n15379), .Z(n15348) );
  XNOR U18497 ( .A(n15380), .B(n15381), .Z(n15379) );
  ANDN U18498 ( .B(n15382), .A(n15383), .Z(n15380) );
  XNOR U18499 ( .A(n15384), .B(n15385), .Z(n15382) );
  IV U18500 ( .A(n15349), .Z(n15346) );
  XOR U18501 ( .A(n15386), .B(n15387), .Z(n15349) );
  ANDN U18502 ( .B(n15388), .A(n15389), .Z(n15386) );
  XOR U18503 ( .A(n15387), .B(n15390), .Z(n15388) );
  XOR U18504 ( .A(n15391), .B(n15392), .Z(n15362) );
  XNOR U18505 ( .A(n15357), .B(n15393), .Z(n15392) );
  IV U18506 ( .A(n15360), .Z(n15393) );
  XOR U18507 ( .A(n15394), .B(n15395), .Z(n15360) );
  ANDN U18508 ( .B(n15396), .A(n15397), .Z(n15394) );
  XOR U18509 ( .A(n15395), .B(n15398), .Z(n15396) );
  XNOR U18510 ( .A(n15399), .B(n15400), .Z(n15357) );
  ANDN U18511 ( .B(n15401), .A(n15402), .Z(n15399) );
  XOR U18512 ( .A(n15400), .B(n15403), .Z(n15401) );
  IV U18513 ( .A(n15356), .Z(n15391) );
  XOR U18514 ( .A(n15354), .B(n15404), .Z(n15356) );
  XNOR U18515 ( .A(n15405), .B(n15406), .Z(n15404) );
  ANDN U18516 ( .B(n15407), .A(n15408), .Z(n15405) );
  XNOR U18517 ( .A(n15409), .B(n15410), .Z(n15407) );
  IV U18518 ( .A(n15358), .Z(n15354) );
  XOR U18519 ( .A(n15411), .B(n15412), .Z(n15358) );
  ANDN U18520 ( .B(n15413), .A(n15414), .Z(n15411) );
  XOR U18521 ( .A(n15415), .B(n15412), .Z(n15413) );
  XOR U18522 ( .A(n15369), .B(n15222), .Z(n15370) );
  XOR U18523 ( .A(n15416), .B(n15417), .Z(n15222) );
  AND U18524 ( .A(n76), .B(n15418), .Z(n15416) );
  XOR U18525 ( .A(n15419), .B(n15417), .Z(n15418) );
  XNOR U18526 ( .A(n15420), .B(n15421), .Z(n15369) );
  NAND U18527 ( .A(n15422), .B(n15423), .Z(n15421) );
  XOR U18528 ( .A(n15424), .B(n15321), .Z(n15423) );
  XOR U18529 ( .A(n15397), .B(n15398), .Z(n15321) );
  XOR U18530 ( .A(n15425), .B(n15390), .Z(n15398) );
  XOR U18531 ( .A(n15426), .B(n15378), .Z(n15390) );
  XOR U18532 ( .A(n15427), .B(n15428), .Z(n15378) );
  ANDN U18533 ( .B(n15429), .A(n15430), .Z(n15427) );
  XOR U18534 ( .A(n15428), .B(n15431), .Z(n15429) );
  IV U18535 ( .A(n15376), .Z(n15426) );
  XOR U18536 ( .A(n15374), .B(n15432), .Z(n15376) );
  XOR U18537 ( .A(n15433), .B(n15434), .Z(n15432) );
  ANDN U18538 ( .B(n15435), .A(n15436), .Z(n15433) );
  XOR U18539 ( .A(n15437), .B(n15434), .Z(n15435) );
  IV U18540 ( .A(n15377), .Z(n15374) );
  XOR U18541 ( .A(n15438), .B(n15439), .Z(n15377) );
  ANDN U18542 ( .B(n15440), .A(n15441), .Z(n15438) );
  XOR U18543 ( .A(n15439), .B(n15442), .Z(n15440) );
  IV U18544 ( .A(n15389), .Z(n15425) );
  XOR U18545 ( .A(n15443), .B(n15444), .Z(n15389) );
  XNOR U18546 ( .A(n15384), .B(n15445), .Z(n15444) );
  IV U18547 ( .A(n15387), .Z(n15445) );
  XOR U18548 ( .A(n15446), .B(n15447), .Z(n15387) );
  ANDN U18549 ( .B(n15448), .A(n15449), .Z(n15446) );
  XOR U18550 ( .A(n15447), .B(n15450), .Z(n15448) );
  XNOR U18551 ( .A(n15451), .B(n15452), .Z(n15384) );
  ANDN U18552 ( .B(n15453), .A(n15454), .Z(n15451) );
  XOR U18553 ( .A(n15452), .B(n15455), .Z(n15453) );
  IV U18554 ( .A(n15383), .Z(n15443) );
  XOR U18555 ( .A(n15381), .B(n15456), .Z(n15383) );
  XOR U18556 ( .A(n15457), .B(n15458), .Z(n15456) );
  ANDN U18557 ( .B(n15459), .A(n15460), .Z(n15457) );
  XOR U18558 ( .A(n15461), .B(n15458), .Z(n15459) );
  IV U18559 ( .A(n15385), .Z(n15381) );
  XOR U18560 ( .A(n15462), .B(n15463), .Z(n15385) );
  ANDN U18561 ( .B(n15464), .A(n15465), .Z(n15462) );
  XOR U18562 ( .A(n15466), .B(n15463), .Z(n15464) );
  XOR U18563 ( .A(n15467), .B(n15468), .Z(n15397) );
  XOR U18564 ( .A(n15415), .B(n15469), .Z(n15468) );
  IV U18565 ( .A(n15395), .Z(n15469) );
  XOR U18566 ( .A(n15470), .B(n15471), .Z(n15395) );
  ANDN U18567 ( .B(n15472), .A(n15473), .Z(n15470) );
  XOR U18568 ( .A(n15471), .B(n15474), .Z(n15472) );
  XOR U18569 ( .A(n15475), .B(n15403), .Z(n15415) );
  XOR U18570 ( .A(n15476), .B(n15477), .Z(n15403) );
  ANDN U18571 ( .B(n15478), .A(n15479), .Z(n15476) );
  XOR U18572 ( .A(n15477), .B(n15480), .Z(n15478) );
  IV U18573 ( .A(n15402), .Z(n15475) );
  XOR U18574 ( .A(n15481), .B(n15482), .Z(n15402) );
  XOR U18575 ( .A(n15483), .B(n15484), .Z(n15482) );
  ANDN U18576 ( .B(n15485), .A(n15486), .Z(n15483) );
  XOR U18577 ( .A(n15487), .B(n15484), .Z(n15485) );
  IV U18578 ( .A(n15400), .Z(n15481) );
  XOR U18579 ( .A(n15488), .B(n15489), .Z(n15400) );
  ANDN U18580 ( .B(n15490), .A(n15491), .Z(n15488) );
  XOR U18581 ( .A(n15489), .B(n15492), .Z(n15490) );
  IV U18582 ( .A(n15414), .Z(n15467) );
  XOR U18583 ( .A(n15493), .B(n15494), .Z(n15414) );
  XNOR U18584 ( .A(n15409), .B(n15495), .Z(n15494) );
  IV U18585 ( .A(n15412), .Z(n15495) );
  XOR U18586 ( .A(n15496), .B(n15497), .Z(n15412) );
  ANDN U18587 ( .B(n15498), .A(n15499), .Z(n15496) );
  XOR U18588 ( .A(n15500), .B(n15497), .Z(n15498) );
  XNOR U18589 ( .A(n15501), .B(n15502), .Z(n15409) );
  ANDN U18590 ( .B(n15503), .A(n15504), .Z(n15501) );
  XOR U18591 ( .A(n15502), .B(n15505), .Z(n15503) );
  IV U18592 ( .A(n15408), .Z(n15493) );
  XOR U18593 ( .A(n15406), .B(n15506), .Z(n15408) );
  XOR U18594 ( .A(n15507), .B(n15508), .Z(n15506) );
  ANDN U18595 ( .B(n15509), .A(n15510), .Z(n15507) );
  XOR U18596 ( .A(n15511), .B(n15508), .Z(n15509) );
  IV U18597 ( .A(n15410), .Z(n15406) );
  XOR U18598 ( .A(n15512), .B(n15513), .Z(n15410) );
  ANDN U18599 ( .B(n15514), .A(n15515), .Z(n15512) );
  XOR U18600 ( .A(n15516), .B(n15513), .Z(n15514) );
  IV U18601 ( .A(n15420), .Z(n15424) );
  XOR U18602 ( .A(n15420), .B(n15323), .Z(n15422) );
  XOR U18603 ( .A(n15517), .B(n15518), .Z(n15323) );
  AND U18604 ( .A(n76), .B(n15519), .Z(n15517) );
  XOR U18605 ( .A(n15520), .B(n15518), .Z(n15519) );
  NANDN U18606 ( .A(n15325), .B(n15327), .Z(n15420) );
  XOR U18607 ( .A(n15521), .B(n15522), .Z(n15327) );
  AND U18608 ( .A(n76), .B(n15523), .Z(n15521) );
  XOR U18609 ( .A(n15522), .B(n15524), .Z(n15523) );
  XNOR U18610 ( .A(n15525), .B(n15526), .Z(n76) );
  AND U18611 ( .A(n15527), .B(n15528), .Z(n15525) );
  XOR U18612 ( .A(n15526), .B(n15338), .Z(n15528) );
  XNOR U18613 ( .A(n15529), .B(n15530), .Z(n15338) );
  ANDN U18614 ( .B(n15531), .A(n15532), .Z(n15529) );
  XOR U18615 ( .A(n15530), .B(n15533), .Z(n15531) );
  XNOR U18616 ( .A(n15526), .B(n15340), .Z(n15527) );
  XOR U18617 ( .A(n15534), .B(n15535), .Z(n15340) );
  AND U18618 ( .A(n80), .B(n15536), .Z(n15534) );
  XOR U18619 ( .A(n15537), .B(n15535), .Z(n15536) );
  XOR U18620 ( .A(n15538), .B(n15539), .Z(n15526) );
  AND U18621 ( .A(n15540), .B(n15541), .Z(n15538) );
  XOR U18622 ( .A(n15539), .B(n15365), .Z(n15541) );
  XOR U18623 ( .A(n15532), .B(n15533), .Z(n15365) );
  XNOR U18624 ( .A(n15542), .B(n15543), .Z(n15533) );
  ANDN U18625 ( .B(n15544), .A(n15545), .Z(n15542) );
  XOR U18626 ( .A(n15546), .B(n15547), .Z(n15544) );
  XOR U18627 ( .A(n15548), .B(n15549), .Z(n15532) );
  XNOR U18628 ( .A(n15550), .B(n15551), .Z(n15549) );
  ANDN U18629 ( .B(n15552), .A(n15553), .Z(n15550) );
  XNOR U18630 ( .A(n15554), .B(n15555), .Z(n15552) );
  IV U18631 ( .A(n15530), .Z(n15548) );
  XOR U18632 ( .A(n15556), .B(n15557), .Z(n15530) );
  ANDN U18633 ( .B(n15558), .A(n15559), .Z(n15556) );
  XOR U18634 ( .A(n15557), .B(n15560), .Z(n15558) );
  XNOR U18635 ( .A(n15539), .B(n15367), .Z(n15540) );
  XOR U18636 ( .A(n15561), .B(n15562), .Z(n15367) );
  AND U18637 ( .A(n80), .B(n15563), .Z(n15561) );
  XOR U18638 ( .A(n15564), .B(n15562), .Z(n15563) );
  XNOR U18639 ( .A(n15565), .B(n15566), .Z(n15539) );
  AND U18640 ( .A(n15567), .B(n15568), .Z(n15565) );
  XNOR U18641 ( .A(n15566), .B(n15417), .Z(n15568) );
  XOR U18642 ( .A(n15559), .B(n15560), .Z(n15417) );
  XOR U18643 ( .A(n15569), .B(n15547), .Z(n15560) );
  XNOR U18644 ( .A(n15570), .B(n15571), .Z(n15547) );
  ANDN U18645 ( .B(n15572), .A(n15573), .Z(n15570) );
  XOR U18646 ( .A(n15574), .B(n15575), .Z(n15572) );
  IV U18647 ( .A(n15545), .Z(n15569) );
  XOR U18648 ( .A(n15543), .B(n15576), .Z(n15545) );
  XNOR U18649 ( .A(n15577), .B(n15578), .Z(n15576) );
  ANDN U18650 ( .B(n15579), .A(n15580), .Z(n15577) );
  XNOR U18651 ( .A(n15581), .B(n15582), .Z(n15579) );
  IV U18652 ( .A(n15546), .Z(n15543) );
  XOR U18653 ( .A(n15583), .B(n15584), .Z(n15546) );
  ANDN U18654 ( .B(n15585), .A(n15586), .Z(n15583) );
  XOR U18655 ( .A(n15584), .B(n15587), .Z(n15585) );
  XOR U18656 ( .A(n15588), .B(n15589), .Z(n15559) );
  XNOR U18657 ( .A(n15554), .B(n15590), .Z(n15589) );
  IV U18658 ( .A(n15557), .Z(n15590) );
  XOR U18659 ( .A(n15591), .B(n15592), .Z(n15557) );
  ANDN U18660 ( .B(n15593), .A(n15594), .Z(n15591) );
  XOR U18661 ( .A(n15592), .B(n15595), .Z(n15593) );
  XNOR U18662 ( .A(n15596), .B(n15597), .Z(n15554) );
  ANDN U18663 ( .B(n15598), .A(n15599), .Z(n15596) );
  XOR U18664 ( .A(n15597), .B(n15600), .Z(n15598) );
  IV U18665 ( .A(n15553), .Z(n15588) );
  XOR U18666 ( .A(n15551), .B(n15601), .Z(n15553) );
  XNOR U18667 ( .A(n15602), .B(n15603), .Z(n15601) );
  ANDN U18668 ( .B(n15604), .A(n15605), .Z(n15602) );
  XNOR U18669 ( .A(n15606), .B(n15607), .Z(n15604) );
  IV U18670 ( .A(n15555), .Z(n15551) );
  XOR U18671 ( .A(n15608), .B(n15609), .Z(n15555) );
  ANDN U18672 ( .B(n15610), .A(n15611), .Z(n15608) );
  XOR U18673 ( .A(n15612), .B(n15609), .Z(n15610) );
  XOR U18674 ( .A(n15566), .B(n15419), .Z(n15567) );
  XOR U18675 ( .A(n15613), .B(n15614), .Z(n15419) );
  AND U18676 ( .A(n80), .B(n15615), .Z(n15613) );
  XOR U18677 ( .A(n15616), .B(n15614), .Z(n15615) );
  XNOR U18678 ( .A(n15617), .B(n15618), .Z(n15566) );
  NAND U18679 ( .A(n15619), .B(n15620), .Z(n15618) );
  XOR U18680 ( .A(n15621), .B(n15518), .Z(n15620) );
  XOR U18681 ( .A(n15594), .B(n15595), .Z(n15518) );
  XOR U18682 ( .A(n15622), .B(n15587), .Z(n15595) );
  XOR U18683 ( .A(n15623), .B(n15575), .Z(n15587) );
  XOR U18684 ( .A(n15624), .B(n15625), .Z(n15575) );
  ANDN U18685 ( .B(n15626), .A(n15627), .Z(n15624) );
  XOR U18686 ( .A(n15625), .B(n15628), .Z(n15626) );
  IV U18687 ( .A(n15573), .Z(n15623) );
  XOR U18688 ( .A(n15571), .B(n15629), .Z(n15573) );
  XOR U18689 ( .A(n15630), .B(n15631), .Z(n15629) );
  ANDN U18690 ( .B(n15632), .A(n15633), .Z(n15630) );
  XOR U18691 ( .A(n15634), .B(n15631), .Z(n15632) );
  IV U18692 ( .A(n15574), .Z(n15571) );
  XOR U18693 ( .A(n15635), .B(n15636), .Z(n15574) );
  ANDN U18694 ( .B(n15637), .A(n15638), .Z(n15635) );
  XOR U18695 ( .A(n15636), .B(n15639), .Z(n15637) );
  IV U18696 ( .A(n15586), .Z(n15622) );
  XOR U18697 ( .A(n15640), .B(n15641), .Z(n15586) );
  XNOR U18698 ( .A(n15581), .B(n15642), .Z(n15641) );
  IV U18699 ( .A(n15584), .Z(n15642) );
  XOR U18700 ( .A(n15643), .B(n15644), .Z(n15584) );
  ANDN U18701 ( .B(n15645), .A(n15646), .Z(n15643) );
  XOR U18702 ( .A(n15644), .B(n15647), .Z(n15645) );
  XNOR U18703 ( .A(n15648), .B(n15649), .Z(n15581) );
  ANDN U18704 ( .B(n15650), .A(n15651), .Z(n15648) );
  XOR U18705 ( .A(n15649), .B(n15652), .Z(n15650) );
  IV U18706 ( .A(n15580), .Z(n15640) );
  XOR U18707 ( .A(n15578), .B(n15653), .Z(n15580) );
  XOR U18708 ( .A(n15654), .B(n15655), .Z(n15653) );
  ANDN U18709 ( .B(n15656), .A(n15657), .Z(n15654) );
  XOR U18710 ( .A(n15658), .B(n15655), .Z(n15656) );
  IV U18711 ( .A(n15582), .Z(n15578) );
  XOR U18712 ( .A(n15659), .B(n15660), .Z(n15582) );
  ANDN U18713 ( .B(n15661), .A(n15662), .Z(n15659) );
  XOR U18714 ( .A(n15663), .B(n15660), .Z(n15661) );
  XOR U18715 ( .A(n15664), .B(n15665), .Z(n15594) );
  XOR U18716 ( .A(n15612), .B(n15666), .Z(n15665) );
  IV U18717 ( .A(n15592), .Z(n15666) );
  XOR U18718 ( .A(n15667), .B(n15668), .Z(n15592) );
  ANDN U18719 ( .B(n15669), .A(n15670), .Z(n15667) );
  XOR U18720 ( .A(n15668), .B(n15671), .Z(n15669) );
  XOR U18721 ( .A(n15672), .B(n15600), .Z(n15612) );
  XOR U18722 ( .A(n15673), .B(n15674), .Z(n15600) );
  ANDN U18723 ( .B(n15675), .A(n15676), .Z(n15673) );
  XOR U18724 ( .A(n15674), .B(n15677), .Z(n15675) );
  IV U18725 ( .A(n15599), .Z(n15672) );
  XOR U18726 ( .A(n15678), .B(n15679), .Z(n15599) );
  XOR U18727 ( .A(n15680), .B(n15681), .Z(n15679) );
  ANDN U18728 ( .B(n15682), .A(n15683), .Z(n15680) );
  XOR U18729 ( .A(n15684), .B(n15681), .Z(n15682) );
  IV U18730 ( .A(n15597), .Z(n15678) );
  XOR U18731 ( .A(n15685), .B(n15686), .Z(n15597) );
  ANDN U18732 ( .B(n15687), .A(n15688), .Z(n15685) );
  XOR U18733 ( .A(n15686), .B(n15689), .Z(n15687) );
  IV U18734 ( .A(n15611), .Z(n15664) );
  XOR U18735 ( .A(n15690), .B(n15691), .Z(n15611) );
  XNOR U18736 ( .A(n15606), .B(n15692), .Z(n15691) );
  IV U18737 ( .A(n15609), .Z(n15692) );
  XOR U18738 ( .A(n15693), .B(n15694), .Z(n15609) );
  ANDN U18739 ( .B(n15695), .A(n15696), .Z(n15693) );
  XOR U18740 ( .A(n15697), .B(n15694), .Z(n15695) );
  XNOR U18741 ( .A(n15698), .B(n15699), .Z(n15606) );
  ANDN U18742 ( .B(n15700), .A(n15701), .Z(n15698) );
  XOR U18743 ( .A(n15699), .B(n15702), .Z(n15700) );
  IV U18744 ( .A(n15605), .Z(n15690) );
  XOR U18745 ( .A(n15603), .B(n15703), .Z(n15605) );
  XOR U18746 ( .A(n15704), .B(n15705), .Z(n15703) );
  ANDN U18747 ( .B(n15706), .A(n15707), .Z(n15704) );
  XOR U18748 ( .A(n15708), .B(n15705), .Z(n15706) );
  IV U18749 ( .A(n15607), .Z(n15603) );
  XOR U18750 ( .A(n15709), .B(n15710), .Z(n15607) );
  ANDN U18751 ( .B(n15711), .A(n15712), .Z(n15709) );
  XOR U18752 ( .A(n15713), .B(n15710), .Z(n15711) );
  IV U18753 ( .A(n15617), .Z(n15621) );
  XOR U18754 ( .A(n15617), .B(n15520), .Z(n15619) );
  XOR U18755 ( .A(n15714), .B(n15715), .Z(n15520) );
  AND U18756 ( .A(n80), .B(n15716), .Z(n15714) );
  XOR U18757 ( .A(n15717), .B(n15715), .Z(n15716) );
  NANDN U18758 ( .A(n15522), .B(n15524), .Z(n15617) );
  XOR U18759 ( .A(n15718), .B(n15719), .Z(n15524) );
  AND U18760 ( .A(n80), .B(n15720), .Z(n15718) );
  XOR U18761 ( .A(n15719), .B(n15721), .Z(n15720) );
  XNOR U18762 ( .A(n15722), .B(n15723), .Z(n80) );
  AND U18763 ( .A(n15724), .B(n15725), .Z(n15722) );
  XOR U18764 ( .A(n15723), .B(n15535), .Z(n15725) );
  XNOR U18765 ( .A(n15726), .B(n15727), .Z(n15535) );
  ANDN U18766 ( .B(n15728), .A(n15729), .Z(n15726) );
  XOR U18767 ( .A(n15727), .B(n15730), .Z(n15728) );
  XNOR U18768 ( .A(n15723), .B(n15537), .Z(n15724) );
  XOR U18769 ( .A(n15731), .B(n15732), .Z(n15537) );
  AND U18770 ( .A(n84), .B(n15733), .Z(n15731) );
  XOR U18771 ( .A(n15734), .B(n15732), .Z(n15733) );
  XOR U18772 ( .A(n15735), .B(n15736), .Z(n15723) );
  AND U18773 ( .A(n15737), .B(n15738), .Z(n15735) );
  XOR U18774 ( .A(n15736), .B(n15562), .Z(n15738) );
  XOR U18775 ( .A(n15729), .B(n15730), .Z(n15562) );
  XNOR U18776 ( .A(n15739), .B(n15740), .Z(n15730) );
  ANDN U18777 ( .B(n15741), .A(n15742), .Z(n15739) );
  XOR U18778 ( .A(n15743), .B(n15744), .Z(n15741) );
  XOR U18779 ( .A(n15745), .B(n15746), .Z(n15729) );
  XNOR U18780 ( .A(n15747), .B(n15748), .Z(n15746) );
  ANDN U18781 ( .B(n15749), .A(n15750), .Z(n15747) );
  XNOR U18782 ( .A(n15751), .B(n15752), .Z(n15749) );
  IV U18783 ( .A(n15727), .Z(n15745) );
  XOR U18784 ( .A(n15753), .B(n15754), .Z(n15727) );
  ANDN U18785 ( .B(n15755), .A(n15756), .Z(n15753) );
  XOR U18786 ( .A(n15754), .B(n15757), .Z(n15755) );
  XNOR U18787 ( .A(n15736), .B(n15564), .Z(n15737) );
  XOR U18788 ( .A(n15758), .B(n15759), .Z(n15564) );
  AND U18789 ( .A(n84), .B(n15760), .Z(n15758) );
  XOR U18790 ( .A(n15761), .B(n15759), .Z(n15760) );
  XNOR U18791 ( .A(n15762), .B(n15763), .Z(n15736) );
  AND U18792 ( .A(n15764), .B(n15765), .Z(n15762) );
  XNOR U18793 ( .A(n15763), .B(n15614), .Z(n15765) );
  XOR U18794 ( .A(n15756), .B(n15757), .Z(n15614) );
  XOR U18795 ( .A(n15766), .B(n15744), .Z(n15757) );
  XNOR U18796 ( .A(n15767), .B(n15768), .Z(n15744) );
  ANDN U18797 ( .B(n15769), .A(n15770), .Z(n15767) );
  XOR U18798 ( .A(n15771), .B(n15772), .Z(n15769) );
  IV U18799 ( .A(n15742), .Z(n15766) );
  XOR U18800 ( .A(n15740), .B(n15773), .Z(n15742) );
  XNOR U18801 ( .A(n15774), .B(n15775), .Z(n15773) );
  ANDN U18802 ( .B(n15776), .A(n15777), .Z(n15774) );
  XNOR U18803 ( .A(n15778), .B(n15779), .Z(n15776) );
  IV U18804 ( .A(n15743), .Z(n15740) );
  XOR U18805 ( .A(n15780), .B(n15781), .Z(n15743) );
  ANDN U18806 ( .B(n15782), .A(n15783), .Z(n15780) );
  XOR U18807 ( .A(n15781), .B(n15784), .Z(n15782) );
  XOR U18808 ( .A(n15785), .B(n15786), .Z(n15756) );
  XNOR U18809 ( .A(n15751), .B(n15787), .Z(n15786) );
  IV U18810 ( .A(n15754), .Z(n15787) );
  XOR U18811 ( .A(n15788), .B(n15789), .Z(n15754) );
  ANDN U18812 ( .B(n15790), .A(n15791), .Z(n15788) );
  XOR U18813 ( .A(n15789), .B(n15792), .Z(n15790) );
  XNOR U18814 ( .A(n15793), .B(n15794), .Z(n15751) );
  ANDN U18815 ( .B(n15795), .A(n15796), .Z(n15793) );
  XOR U18816 ( .A(n15794), .B(n15797), .Z(n15795) );
  IV U18817 ( .A(n15750), .Z(n15785) );
  XOR U18818 ( .A(n15748), .B(n15798), .Z(n15750) );
  XNOR U18819 ( .A(n15799), .B(n15800), .Z(n15798) );
  ANDN U18820 ( .B(n15801), .A(n15802), .Z(n15799) );
  XNOR U18821 ( .A(n15803), .B(n15804), .Z(n15801) );
  IV U18822 ( .A(n15752), .Z(n15748) );
  XOR U18823 ( .A(n15805), .B(n15806), .Z(n15752) );
  ANDN U18824 ( .B(n15807), .A(n15808), .Z(n15805) );
  XOR U18825 ( .A(n15809), .B(n15806), .Z(n15807) );
  XOR U18826 ( .A(n15763), .B(n15616), .Z(n15764) );
  XOR U18827 ( .A(n15810), .B(n15811), .Z(n15616) );
  AND U18828 ( .A(n84), .B(n15812), .Z(n15810) );
  XOR U18829 ( .A(n15813), .B(n15811), .Z(n15812) );
  XNOR U18830 ( .A(n15814), .B(n15815), .Z(n15763) );
  NAND U18831 ( .A(n15816), .B(n15817), .Z(n15815) );
  XOR U18832 ( .A(n15818), .B(n15715), .Z(n15817) );
  XOR U18833 ( .A(n15791), .B(n15792), .Z(n15715) );
  XOR U18834 ( .A(n15819), .B(n15784), .Z(n15792) );
  XOR U18835 ( .A(n15820), .B(n15772), .Z(n15784) );
  XOR U18836 ( .A(n15821), .B(n15822), .Z(n15772) );
  ANDN U18837 ( .B(n15823), .A(n15824), .Z(n15821) );
  XOR U18838 ( .A(n15822), .B(n15825), .Z(n15823) );
  IV U18839 ( .A(n15770), .Z(n15820) );
  XOR U18840 ( .A(n15768), .B(n15826), .Z(n15770) );
  XOR U18841 ( .A(n15827), .B(n15828), .Z(n15826) );
  ANDN U18842 ( .B(n15829), .A(n15830), .Z(n15827) );
  XOR U18843 ( .A(n15831), .B(n15828), .Z(n15829) );
  IV U18844 ( .A(n15771), .Z(n15768) );
  XOR U18845 ( .A(n15832), .B(n15833), .Z(n15771) );
  ANDN U18846 ( .B(n15834), .A(n15835), .Z(n15832) );
  XOR U18847 ( .A(n15833), .B(n15836), .Z(n15834) );
  IV U18848 ( .A(n15783), .Z(n15819) );
  XOR U18849 ( .A(n15837), .B(n15838), .Z(n15783) );
  XNOR U18850 ( .A(n15778), .B(n15839), .Z(n15838) );
  IV U18851 ( .A(n15781), .Z(n15839) );
  XOR U18852 ( .A(n15840), .B(n15841), .Z(n15781) );
  ANDN U18853 ( .B(n15842), .A(n15843), .Z(n15840) );
  XOR U18854 ( .A(n15841), .B(n15844), .Z(n15842) );
  XNOR U18855 ( .A(n15845), .B(n15846), .Z(n15778) );
  ANDN U18856 ( .B(n15847), .A(n15848), .Z(n15845) );
  XOR U18857 ( .A(n15846), .B(n15849), .Z(n15847) );
  IV U18858 ( .A(n15777), .Z(n15837) );
  XOR U18859 ( .A(n15775), .B(n15850), .Z(n15777) );
  XOR U18860 ( .A(n15851), .B(n15852), .Z(n15850) );
  ANDN U18861 ( .B(n15853), .A(n15854), .Z(n15851) );
  XOR U18862 ( .A(n15855), .B(n15852), .Z(n15853) );
  IV U18863 ( .A(n15779), .Z(n15775) );
  XOR U18864 ( .A(n15856), .B(n15857), .Z(n15779) );
  ANDN U18865 ( .B(n15858), .A(n15859), .Z(n15856) );
  XOR U18866 ( .A(n15860), .B(n15857), .Z(n15858) );
  XOR U18867 ( .A(n15861), .B(n15862), .Z(n15791) );
  XOR U18868 ( .A(n15809), .B(n15863), .Z(n15862) );
  IV U18869 ( .A(n15789), .Z(n15863) );
  XOR U18870 ( .A(n15864), .B(n15865), .Z(n15789) );
  ANDN U18871 ( .B(n15866), .A(n15867), .Z(n15864) );
  XOR U18872 ( .A(n15865), .B(n15868), .Z(n15866) );
  XOR U18873 ( .A(n15869), .B(n15797), .Z(n15809) );
  XOR U18874 ( .A(n15870), .B(n15871), .Z(n15797) );
  ANDN U18875 ( .B(n15872), .A(n15873), .Z(n15870) );
  XOR U18876 ( .A(n15871), .B(n15874), .Z(n15872) );
  IV U18877 ( .A(n15796), .Z(n15869) );
  XOR U18878 ( .A(n15875), .B(n15876), .Z(n15796) );
  XOR U18879 ( .A(n15877), .B(n15878), .Z(n15876) );
  ANDN U18880 ( .B(n15879), .A(n15880), .Z(n15877) );
  XOR U18881 ( .A(n15881), .B(n15878), .Z(n15879) );
  IV U18882 ( .A(n15794), .Z(n15875) );
  XOR U18883 ( .A(n15882), .B(n15883), .Z(n15794) );
  ANDN U18884 ( .B(n15884), .A(n15885), .Z(n15882) );
  XOR U18885 ( .A(n15883), .B(n15886), .Z(n15884) );
  IV U18886 ( .A(n15808), .Z(n15861) );
  XOR U18887 ( .A(n15887), .B(n15888), .Z(n15808) );
  XNOR U18888 ( .A(n15803), .B(n15889), .Z(n15888) );
  IV U18889 ( .A(n15806), .Z(n15889) );
  XOR U18890 ( .A(n15890), .B(n15891), .Z(n15806) );
  ANDN U18891 ( .B(n15892), .A(n15893), .Z(n15890) );
  XOR U18892 ( .A(n15894), .B(n15891), .Z(n15892) );
  XNOR U18893 ( .A(n15895), .B(n15896), .Z(n15803) );
  ANDN U18894 ( .B(n15897), .A(n15898), .Z(n15895) );
  XOR U18895 ( .A(n15896), .B(n15899), .Z(n15897) );
  IV U18896 ( .A(n15802), .Z(n15887) );
  XOR U18897 ( .A(n15800), .B(n15900), .Z(n15802) );
  XOR U18898 ( .A(n15901), .B(n15902), .Z(n15900) );
  ANDN U18899 ( .B(n15903), .A(n15904), .Z(n15901) );
  XOR U18900 ( .A(n15905), .B(n15902), .Z(n15903) );
  IV U18901 ( .A(n15804), .Z(n15800) );
  XOR U18902 ( .A(n15906), .B(n15907), .Z(n15804) );
  ANDN U18903 ( .B(n15908), .A(n15909), .Z(n15906) );
  XOR U18904 ( .A(n15910), .B(n15907), .Z(n15908) );
  IV U18905 ( .A(n15814), .Z(n15818) );
  XOR U18906 ( .A(n15814), .B(n15717), .Z(n15816) );
  XOR U18907 ( .A(n15911), .B(n15912), .Z(n15717) );
  AND U18908 ( .A(n84), .B(n15913), .Z(n15911) );
  XOR U18909 ( .A(n15914), .B(n15912), .Z(n15913) );
  NANDN U18910 ( .A(n15719), .B(n15721), .Z(n15814) );
  XOR U18911 ( .A(n15915), .B(n15916), .Z(n15721) );
  AND U18912 ( .A(n84), .B(n15917), .Z(n15915) );
  XOR U18913 ( .A(n15916), .B(n15918), .Z(n15917) );
  XNOR U18914 ( .A(n15919), .B(n15920), .Z(n84) );
  AND U18915 ( .A(n15921), .B(n15922), .Z(n15919) );
  XOR U18916 ( .A(n15920), .B(n15732), .Z(n15922) );
  XNOR U18917 ( .A(n15923), .B(n15924), .Z(n15732) );
  ANDN U18918 ( .B(n15925), .A(n15926), .Z(n15923) );
  XOR U18919 ( .A(n15924), .B(n15927), .Z(n15925) );
  XNOR U18920 ( .A(n15920), .B(n15734), .Z(n15921) );
  XOR U18921 ( .A(n15928), .B(n15929), .Z(n15734) );
  AND U18922 ( .A(n88), .B(n15930), .Z(n15928) );
  XOR U18923 ( .A(n15931), .B(n15929), .Z(n15930) );
  XOR U18924 ( .A(n15932), .B(n15933), .Z(n15920) );
  AND U18925 ( .A(n15934), .B(n15935), .Z(n15932) );
  XOR U18926 ( .A(n15933), .B(n15759), .Z(n15935) );
  XOR U18927 ( .A(n15926), .B(n15927), .Z(n15759) );
  XNOR U18928 ( .A(n15936), .B(n15937), .Z(n15927) );
  ANDN U18929 ( .B(n15938), .A(n15939), .Z(n15936) );
  XOR U18930 ( .A(n15940), .B(n15941), .Z(n15938) );
  XOR U18931 ( .A(n15942), .B(n15943), .Z(n15926) );
  XNOR U18932 ( .A(n15944), .B(n15945), .Z(n15943) );
  ANDN U18933 ( .B(n15946), .A(n15947), .Z(n15944) );
  XNOR U18934 ( .A(n15948), .B(n15949), .Z(n15946) );
  IV U18935 ( .A(n15924), .Z(n15942) );
  XOR U18936 ( .A(n15950), .B(n15951), .Z(n15924) );
  ANDN U18937 ( .B(n15952), .A(n15953), .Z(n15950) );
  XOR U18938 ( .A(n15951), .B(n15954), .Z(n15952) );
  XNOR U18939 ( .A(n15933), .B(n15761), .Z(n15934) );
  XOR U18940 ( .A(n15955), .B(n15956), .Z(n15761) );
  AND U18941 ( .A(n88), .B(n15957), .Z(n15955) );
  XOR U18942 ( .A(n15958), .B(n15956), .Z(n15957) );
  XNOR U18943 ( .A(n15959), .B(n15960), .Z(n15933) );
  AND U18944 ( .A(n15961), .B(n15962), .Z(n15959) );
  XNOR U18945 ( .A(n15960), .B(n15811), .Z(n15962) );
  XOR U18946 ( .A(n15953), .B(n15954), .Z(n15811) );
  XOR U18947 ( .A(n15963), .B(n15941), .Z(n15954) );
  XNOR U18948 ( .A(n15964), .B(n15965), .Z(n15941) );
  ANDN U18949 ( .B(n15966), .A(n15967), .Z(n15964) );
  XOR U18950 ( .A(n15968), .B(n15969), .Z(n15966) );
  IV U18951 ( .A(n15939), .Z(n15963) );
  XOR U18952 ( .A(n15937), .B(n15970), .Z(n15939) );
  XNOR U18953 ( .A(n15971), .B(n15972), .Z(n15970) );
  ANDN U18954 ( .B(n15973), .A(n15974), .Z(n15971) );
  XNOR U18955 ( .A(n15975), .B(n15976), .Z(n15973) );
  IV U18956 ( .A(n15940), .Z(n15937) );
  XOR U18957 ( .A(n15977), .B(n15978), .Z(n15940) );
  ANDN U18958 ( .B(n15979), .A(n15980), .Z(n15977) );
  XOR U18959 ( .A(n15978), .B(n15981), .Z(n15979) );
  XOR U18960 ( .A(n15982), .B(n15983), .Z(n15953) );
  XNOR U18961 ( .A(n15948), .B(n15984), .Z(n15983) );
  IV U18962 ( .A(n15951), .Z(n15984) );
  XOR U18963 ( .A(n15985), .B(n15986), .Z(n15951) );
  ANDN U18964 ( .B(n15987), .A(n15988), .Z(n15985) );
  XOR U18965 ( .A(n15986), .B(n15989), .Z(n15987) );
  XNOR U18966 ( .A(n15990), .B(n15991), .Z(n15948) );
  ANDN U18967 ( .B(n15992), .A(n15993), .Z(n15990) );
  XOR U18968 ( .A(n15991), .B(n15994), .Z(n15992) );
  IV U18969 ( .A(n15947), .Z(n15982) );
  XOR U18970 ( .A(n15945), .B(n15995), .Z(n15947) );
  XNOR U18971 ( .A(n15996), .B(n15997), .Z(n15995) );
  ANDN U18972 ( .B(n15998), .A(n15999), .Z(n15996) );
  XNOR U18973 ( .A(n16000), .B(n16001), .Z(n15998) );
  IV U18974 ( .A(n15949), .Z(n15945) );
  XOR U18975 ( .A(n16002), .B(n16003), .Z(n15949) );
  ANDN U18976 ( .B(n16004), .A(n16005), .Z(n16002) );
  XOR U18977 ( .A(n16006), .B(n16003), .Z(n16004) );
  XOR U18978 ( .A(n15960), .B(n15813), .Z(n15961) );
  XOR U18979 ( .A(n16007), .B(n16008), .Z(n15813) );
  AND U18980 ( .A(n88), .B(n16009), .Z(n16007) );
  XOR U18981 ( .A(n16010), .B(n16008), .Z(n16009) );
  XNOR U18982 ( .A(n16011), .B(n16012), .Z(n15960) );
  NAND U18983 ( .A(n16013), .B(n16014), .Z(n16012) );
  XOR U18984 ( .A(n16015), .B(n15912), .Z(n16014) );
  XOR U18985 ( .A(n15988), .B(n15989), .Z(n15912) );
  XOR U18986 ( .A(n16016), .B(n15981), .Z(n15989) );
  XOR U18987 ( .A(n16017), .B(n15969), .Z(n15981) );
  XOR U18988 ( .A(n16018), .B(n16019), .Z(n15969) );
  ANDN U18989 ( .B(n16020), .A(n16021), .Z(n16018) );
  XOR U18990 ( .A(n16019), .B(n16022), .Z(n16020) );
  IV U18991 ( .A(n15967), .Z(n16017) );
  XOR U18992 ( .A(n15965), .B(n16023), .Z(n15967) );
  XOR U18993 ( .A(n16024), .B(n16025), .Z(n16023) );
  ANDN U18994 ( .B(n16026), .A(n16027), .Z(n16024) );
  XOR U18995 ( .A(n16028), .B(n16025), .Z(n16026) );
  IV U18996 ( .A(n15968), .Z(n15965) );
  XOR U18997 ( .A(n16029), .B(n16030), .Z(n15968) );
  ANDN U18998 ( .B(n16031), .A(n16032), .Z(n16029) );
  XOR U18999 ( .A(n16030), .B(n16033), .Z(n16031) );
  IV U19000 ( .A(n15980), .Z(n16016) );
  XOR U19001 ( .A(n16034), .B(n16035), .Z(n15980) );
  XNOR U19002 ( .A(n15975), .B(n16036), .Z(n16035) );
  IV U19003 ( .A(n15978), .Z(n16036) );
  XOR U19004 ( .A(n16037), .B(n16038), .Z(n15978) );
  ANDN U19005 ( .B(n16039), .A(n16040), .Z(n16037) );
  XOR U19006 ( .A(n16038), .B(n16041), .Z(n16039) );
  XNOR U19007 ( .A(n16042), .B(n16043), .Z(n15975) );
  ANDN U19008 ( .B(n16044), .A(n16045), .Z(n16042) );
  XOR U19009 ( .A(n16043), .B(n16046), .Z(n16044) );
  IV U19010 ( .A(n15974), .Z(n16034) );
  XOR U19011 ( .A(n15972), .B(n16047), .Z(n15974) );
  XOR U19012 ( .A(n16048), .B(n16049), .Z(n16047) );
  ANDN U19013 ( .B(n16050), .A(n16051), .Z(n16048) );
  XOR U19014 ( .A(n16052), .B(n16049), .Z(n16050) );
  IV U19015 ( .A(n15976), .Z(n15972) );
  XOR U19016 ( .A(n16053), .B(n16054), .Z(n15976) );
  ANDN U19017 ( .B(n16055), .A(n16056), .Z(n16053) );
  XOR U19018 ( .A(n16057), .B(n16054), .Z(n16055) );
  XOR U19019 ( .A(n16058), .B(n16059), .Z(n15988) );
  XOR U19020 ( .A(n16006), .B(n16060), .Z(n16059) );
  IV U19021 ( .A(n15986), .Z(n16060) );
  XOR U19022 ( .A(n16061), .B(n16062), .Z(n15986) );
  ANDN U19023 ( .B(n16063), .A(n16064), .Z(n16061) );
  XOR U19024 ( .A(n16062), .B(n16065), .Z(n16063) );
  XOR U19025 ( .A(n16066), .B(n15994), .Z(n16006) );
  XOR U19026 ( .A(n16067), .B(n16068), .Z(n15994) );
  ANDN U19027 ( .B(n16069), .A(n16070), .Z(n16067) );
  XOR U19028 ( .A(n16068), .B(n16071), .Z(n16069) );
  IV U19029 ( .A(n15993), .Z(n16066) );
  XOR U19030 ( .A(n16072), .B(n16073), .Z(n15993) );
  XOR U19031 ( .A(n16074), .B(n16075), .Z(n16073) );
  ANDN U19032 ( .B(n16076), .A(n16077), .Z(n16074) );
  XOR U19033 ( .A(n16078), .B(n16075), .Z(n16076) );
  IV U19034 ( .A(n15991), .Z(n16072) );
  XOR U19035 ( .A(n16079), .B(n16080), .Z(n15991) );
  ANDN U19036 ( .B(n16081), .A(n16082), .Z(n16079) );
  XOR U19037 ( .A(n16080), .B(n16083), .Z(n16081) );
  IV U19038 ( .A(n16005), .Z(n16058) );
  XOR U19039 ( .A(n16084), .B(n16085), .Z(n16005) );
  XNOR U19040 ( .A(n16000), .B(n16086), .Z(n16085) );
  IV U19041 ( .A(n16003), .Z(n16086) );
  XOR U19042 ( .A(n16087), .B(n16088), .Z(n16003) );
  ANDN U19043 ( .B(n16089), .A(n16090), .Z(n16087) );
  XOR U19044 ( .A(n16091), .B(n16088), .Z(n16089) );
  XNOR U19045 ( .A(n16092), .B(n16093), .Z(n16000) );
  ANDN U19046 ( .B(n16094), .A(n16095), .Z(n16092) );
  XOR U19047 ( .A(n16093), .B(n16096), .Z(n16094) );
  IV U19048 ( .A(n15999), .Z(n16084) );
  XOR U19049 ( .A(n15997), .B(n16097), .Z(n15999) );
  XOR U19050 ( .A(n16098), .B(n16099), .Z(n16097) );
  ANDN U19051 ( .B(n16100), .A(n16101), .Z(n16098) );
  XOR U19052 ( .A(n16102), .B(n16099), .Z(n16100) );
  IV U19053 ( .A(n16001), .Z(n15997) );
  XOR U19054 ( .A(n16103), .B(n16104), .Z(n16001) );
  ANDN U19055 ( .B(n16105), .A(n16106), .Z(n16103) );
  XOR U19056 ( .A(n16107), .B(n16104), .Z(n16105) );
  IV U19057 ( .A(n16011), .Z(n16015) );
  XOR U19058 ( .A(n16011), .B(n15914), .Z(n16013) );
  XOR U19059 ( .A(n16108), .B(n16109), .Z(n15914) );
  AND U19060 ( .A(n88), .B(n16110), .Z(n16108) );
  XOR U19061 ( .A(n16111), .B(n16109), .Z(n16110) );
  NANDN U19062 ( .A(n15916), .B(n15918), .Z(n16011) );
  XOR U19063 ( .A(n16112), .B(n16113), .Z(n15918) );
  AND U19064 ( .A(n88), .B(n16114), .Z(n16112) );
  XOR U19065 ( .A(n16113), .B(n16115), .Z(n16114) );
  XNOR U19066 ( .A(n16116), .B(n16117), .Z(n88) );
  AND U19067 ( .A(n16118), .B(n16119), .Z(n16116) );
  XOR U19068 ( .A(n16117), .B(n15929), .Z(n16119) );
  XNOR U19069 ( .A(n16120), .B(n16121), .Z(n15929) );
  ANDN U19070 ( .B(n16122), .A(n16123), .Z(n16120) );
  XOR U19071 ( .A(n16121), .B(n16124), .Z(n16122) );
  XNOR U19072 ( .A(n16117), .B(n15931), .Z(n16118) );
  XOR U19073 ( .A(n16125), .B(n16126), .Z(n15931) );
  AND U19074 ( .A(n92), .B(n16127), .Z(n16125) );
  XOR U19075 ( .A(n16128), .B(n16126), .Z(n16127) );
  XOR U19076 ( .A(n16129), .B(n16130), .Z(n16117) );
  AND U19077 ( .A(n16131), .B(n16132), .Z(n16129) );
  XOR U19078 ( .A(n16130), .B(n15956), .Z(n16132) );
  XOR U19079 ( .A(n16123), .B(n16124), .Z(n15956) );
  XNOR U19080 ( .A(n16133), .B(n16134), .Z(n16124) );
  ANDN U19081 ( .B(n16135), .A(n16136), .Z(n16133) );
  XOR U19082 ( .A(n16137), .B(n16138), .Z(n16135) );
  XOR U19083 ( .A(n16139), .B(n16140), .Z(n16123) );
  XNOR U19084 ( .A(n16141), .B(n16142), .Z(n16140) );
  ANDN U19085 ( .B(n16143), .A(n16144), .Z(n16141) );
  XNOR U19086 ( .A(n16145), .B(n16146), .Z(n16143) );
  IV U19087 ( .A(n16121), .Z(n16139) );
  XOR U19088 ( .A(n16147), .B(n16148), .Z(n16121) );
  ANDN U19089 ( .B(n16149), .A(n16150), .Z(n16147) );
  XOR U19090 ( .A(n16148), .B(n16151), .Z(n16149) );
  XNOR U19091 ( .A(n16130), .B(n15958), .Z(n16131) );
  XOR U19092 ( .A(n16152), .B(n16153), .Z(n15958) );
  AND U19093 ( .A(n92), .B(n16154), .Z(n16152) );
  XOR U19094 ( .A(n16155), .B(n16153), .Z(n16154) );
  XNOR U19095 ( .A(n16156), .B(n16157), .Z(n16130) );
  AND U19096 ( .A(n16158), .B(n16159), .Z(n16156) );
  XNOR U19097 ( .A(n16157), .B(n16008), .Z(n16159) );
  XOR U19098 ( .A(n16150), .B(n16151), .Z(n16008) );
  XOR U19099 ( .A(n16160), .B(n16138), .Z(n16151) );
  XNOR U19100 ( .A(n16161), .B(n16162), .Z(n16138) );
  ANDN U19101 ( .B(n16163), .A(n16164), .Z(n16161) );
  XOR U19102 ( .A(n16165), .B(n16166), .Z(n16163) );
  IV U19103 ( .A(n16136), .Z(n16160) );
  XOR U19104 ( .A(n16134), .B(n16167), .Z(n16136) );
  XNOR U19105 ( .A(n16168), .B(n16169), .Z(n16167) );
  ANDN U19106 ( .B(n16170), .A(n16171), .Z(n16168) );
  XNOR U19107 ( .A(n16172), .B(n16173), .Z(n16170) );
  IV U19108 ( .A(n16137), .Z(n16134) );
  XOR U19109 ( .A(n16174), .B(n16175), .Z(n16137) );
  ANDN U19110 ( .B(n16176), .A(n16177), .Z(n16174) );
  XOR U19111 ( .A(n16175), .B(n16178), .Z(n16176) );
  XOR U19112 ( .A(n16179), .B(n16180), .Z(n16150) );
  XNOR U19113 ( .A(n16145), .B(n16181), .Z(n16180) );
  IV U19114 ( .A(n16148), .Z(n16181) );
  XOR U19115 ( .A(n16182), .B(n16183), .Z(n16148) );
  ANDN U19116 ( .B(n16184), .A(n16185), .Z(n16182) );
  XOR U19117 ( .A(n16183), .B(n16186), .Z(n16184) );
  XNOR U19118 ( .A(n16187), .B(n16188), .Z(n16145) );
  ANDN U19119 ( .B(n16189), .A(n16190), .Z(n16187) );
  XOR U19120 ( .A(n16188), .B(n16191), .Z(n16189) );
  IV U19121 ( .A(n16144), .Z(n16179) );
  XOR U19122 ( .A(n16142), .B(n16192), .Z(n16144) );
  XNOR U19123 ( .A(n16193), .B(n16194), .Z(n16192) );
  ANDN U19124 ( .B(n16195), .A(n16196), .Z(n16193) );
  XNOR U19125 ( .A(n16197), .B(n16198), .Z(n16195) );
  IV U19126 ( .A(n16146), .Z(n16142) );
  XOR U19127 ( .A(n16199), .B(n16200), .Z(n16146) );
  ANDN U19128 ( .B(n16201), .A(n16202), .Z(n16199) );
  XOR U19129 ( .A(n16203), .B(n16200), .Z(n16201) );
  XOR U19130 ( .A(n16157), .B(n16010), .Z(n16158) );
  XOR U19131 ( .A(n16204), .B(n16205), .Z(n16010) );
  AND U19132 ( .A(n92), .B(n16206), .Z(n16204) );
  XOR U19133 ( .A(n16207), .B(n16205), .Z(n16206) );
  XNOR U19134 ( .A(n16208), .B(n16209), .Z(n16157) );
  NAND U19135 ( .A(n16210), .B(n16211), .Z(n16209) );
  XOR U19136 ( .A(n16212), .B(n16109), .Z(n16211) );
  XOR U19137 ( .A(n16185), .B(n16186), .Z(n16109) );
  XOR U19138 ( .A(n16213), .B(n16178), .Z(n16186) );
  XOR U19139 ( .A(n16214), .B(n16166), .Z(n16178) );
  XOR U19140 ( .A(n16215), .B(n16216), .Z(n16166) );
  ANDN U19141 ( .B(n16217), .A(n16218), .Z(n16215) );
  XOR U19142 ( .A(n16216), .B(n16219), .Z(n16217) );
  IV U19143 ( .A(n16164), .Z(n16214) );
  XOR U19144 ( .A(n16162), .B(n16220), .Z(n16164) );
  XOR U19145 ( .A(n16221), .B(n16222), .Z(n16220) );
  ANDN U19146 ( .B(n16223), .A(n16224), .Z(n16221) );
  XOR U19147 ( .A(n16225), .B(n16222), .Z(n16223) );
  IV U19148 ( .A(n16165), .Z(n16162) );
  XOR U19149 ( .A(n16226), .B(n16227), .Z(n16165) );
  ANDN U19150 ( .B(n16228), .A(n16229), .Z(n16226) );
  XOR U19151 ( .A(n16227), .B(n16230), .Z(n16228) );
  IV U19152 ( .A(n16177), .Z(n16213) );
  XOR U19153 ( .A(n16231), .B(n16232), .Z(n16177) );
  XNOR U19154 ( .A(n16172), .B(n16233), .Z(n16232) );
  IV U19155 ( .A(n16175), .Z(n16233) );
  XOR U19156 ( .A(n16234), .B(n16235), .Z(n16175) );
  ANDN U19157 ( .B(n16236), .A(n16237), .Z(n16234) );
  XOR U19158 ( .A(n16235), .B(n16238), .Z(n16236) );
  XNOR U19159 ( .A(n16239), .B(n16240), .Z(n16172) );
  ANDN U19160 ( .B(n16241), .A(n16242), .Z(n16239) );
  XOR U19161 ( .A(n16240), .B(n16243), .Z(n16241) );
  IV U19162 ( .A(n16171), .Z(n16231) );
  XOR U19163 ( .A(n16169), .B(n16244), .Z(n16171) );
  XOR U19164 ( .A(n16245), .B(n16246), .Z(n16244) );
  ANDN U19165 ( .B(n16247), .A(n16248), .Z(n16245) );
  XOR U19166 ( .A(n16249), .B(n16246), .Z(n16247) );
  IV U19167 ( .A(n16173), .Z(n16169) );
  XOR U19168 ( .A(n16250), .B(n16251), .Z(n16173) );
  ANDN U19169 ( .B(n16252), .A(n16253), .Z(n16250) );
  XOR U19170 ( .A(n16254), .B(n16251), .Z(n16252) );
  XOR U19171 ( .A(n16255), .B(n16256), .Z(n16185) );
  XOR U19172 ( .A(n16203), .B(n16257), .Z(n16256) );
  IV U19173 ( .A(n16183), .Z(n16257) );
  XOR U19174 ( .A(n16258), .B(n16259), .Z(n16183) );
  ANDN U19175 ( .B(n16260), .A(n16261), .Z(n16258) );
  XOR U19176 ( .A(n16259), .B(n16262), .Z(n16260) );
  XOR U19177 ( .A(n16263), .B(n16191), .Z(n16203) );
  XOR U19178 ( .A(n16264), .B(n16265), .Z(n16191) );
  ANDN U19179 ( .B(n16266), .A(n16267), .Z(n16264) );
  XOR U19180 ( .A(n16265), .B(n16268), .Z(n16266) );
  IV U19181 ( .A(n16190), .Z(n16263) );
  XOR U19182 ( .A(n16269), .B(n16270), .Z(n16190) );
  XOR U19183 ( .A(n16271), .B(n16272), .Z(n16270) );
  ANDN U19184 ( .B(n16273), .A(n16274), .Z(n16271) );
  XOR U19185 ( .A(n16275), .B(n16272), .Z(n16273) );
  IV U19186 ( .A(n16188), .Z(n16269) );
  XOR U19187 ( .A(n16276), .B(n16277), .Z(n16188) );
  ANDN U19188 ( .B(n16278), .A(n16279), .Z(n16276) );
  XOR U19189 ( .A(n16277), .B(n16280), .Z(n16278) );
  IV U19190 ( .A(n16202), .Z(n16255) );
  XOR U19191 ( .A(n16281), .B(n16282), .Z(n16202) );
  XNOR U19192 ( .A(n16197), .B(n16283), .Z(n16282) );
  IV U19193 ( .A(n16200), .Z(n16283) );
  XOR U19194 ( .A(n16284), .B(n16285), .Z(n16200) );
  ANDN U19195 ( .B(n16286), .A(n16287), .Z(n16284) );
  XOR U19196 ( .A(n16288), .B(n16285), .Z(n16286) );
  XNOR U19197 ( .A(n16289), .B(n16290), .Z(n16197) );
  ANDN U19198 ( .B(n16291), .A(n16292), .Z(n16289) );
  XOR U19199 ( .A(n16290), .B(n16293), .Z(n16291) );
  IV U19200 ( .A(n16196), .Z(n16281) );
  XOR U19201 ( .A(n16194), .B(n16294), .Z(n16196) );
  XOR U19202 ( .A(n16295), .B(n16296), .Z(n16294) );
  ANDN U19203 ( .B(n16297), .A(n16298), .Z(n16295) );
  XOR U19204 ( .A(n16299), .B(n16296), .Z(n16297) );
  IV U19205 ( .A(n16198), .Z(n16194) );
  XOR U19206 ( .A(n16300), .B(n16301), .Z(n16198) );
  ANDN U19207 ( .B(n16302), .A(n16303), .Z(n16300) );
  XOR U19208 ( .A(n16304), .B(n16301), .Z(n16302) );
  IV U19209 ( .A(n16208), .Z(n16212) );
  XOR U19210 ( .A(n16208), .B(n16111), .Z(n16210) );
  XOR U19211 ( .A(n16305), .B(n16306), .Z(n16111) );
  AND U19212 ( .A(n92), .B(n16307), .Z(n16305) );
  XOR U19213 ( .A(n16308), .B(n16306), .Z(n16307) );
  NANDN U19214 ( .A(n16113), .B(n16115), .Z(n16208) );
  XOR U19215 ( .A(n16309), .B(n16310), .Z(n16115) );
  AND U19216 ( .A(n92), .B(n16311), .Z(n16309) );
  XOR U19217 ( .A(n16310), .B(n16312), .Z(n16311) );
  XNOR U19218 ( .A(n16313), .B(n16314), .Z(n92) );
  AND U19219 ( .A(n16315), .B(n16316), .Z(n16313) );
  XOR U19220 ( .A(n16314), .B(n16126), .Z(n16316) );
  XNOR U19221 ( .A(n16317), .B(n16318), .Z(n16126) );
  ANDN U19222 ( .B(n16319), .A(n16320), .Z(n16317) );
  XOR U19223 ( .A(n16318), .B(n16321), .Z(n16319) );
  XNOR U19224 ( .A(n16314), .B(n16128), .Z(n16315) );
  XOR U19225 ( .A(n16322), .B(n16323), .Z(n16128) );
  AND U19226 ( .A(n96), .B(n16324), .Z(n16322) );
  XOR U19227 ( .A(n16325), .B(n16323), .Z(n16324) );
  XOR U19228 ( .A(n16326), .B(n16327), .Z(n16314) );
  AND U19229 ( .A(n16328), .B(n16329), .Z(n16326) );
  XOR U19230 ( .A(n16327), .B(n16153), .Z(n16329) );
  XOR U19231 ( .A(n16320), .B(n16321), .Z(n16153) );
  XNOR U19232 ( .A(n16330), .B(n16331), .Z(n16321) );
  ANDN U19233 ( .B(n16332), .A(n16333), .Z(n16330) );
  XOR U19234 ( .A(n16334), .B(n16335), .Z(n16332) );
  XOR U19235 ( .A(n16336), .B(n16337), .Z(n16320) );
  XNOR U19236 ( .A(n16338), .B(n16339), .Z(n16337) );
  ANDN U19237 ( .B(n16340), .A(n16341), .Z(n16338) );
  XNOR U19238 ( .A(n16342), .B(n16343), .Z(n16340) );
  IV U19239 ( .A(n16318), .Z(n16336) );
  XOR U19240 ( .A(n16344), .B(n16345), .Z(n16318) );
  ANDN U19241 ( .B(n16346), .A(n16347), .Z(n16344) );
  XOR U19242 ( .A(n16345), .B(n16348), .Z(n16346) );
  XNOR U19243 ( .A(n16327), .B(n16155), .Z(n16328) );
  XOR U19244 ( .A(n16349), .B(n16350), .Z(n16155) );
  AND U19245 ( .A(n96), .B(n16351), .Z(n16349) );
  XOR U19246 ( .A(n16352), .B(n16350), .Z(n16351) );
  XNOR U19247 ( .A(n16353), .B(n16354), .Z(n16327) );
  AND U19248 ( .A(n16355), .B(n16356), .Z(n16353) );
  XNOR U19249 ( .A(n16354), .B(n16205), .Z(n16356) );
  XOR U19250 ( .A(n16347), .B(n16348), .Z(n16205) );
  XOR U19251 ( .A(n16357), .B(n16335), .Z(n16348) );
  XNOR U19252 ( .A(n16358), .B(n16359), .Z(n16335) );
  ANDN U19253 ( .B(n16360), .A(n16361), .Z(n16358) );
  XOR U19254 ( .A(n16362), .B(n16363), .Z(n16360) );
  IV U19255 ( .A(n16333), .Z(n16357) );
  XOR U19256 ( .A(n16331), .B(n16364), .Z(n16333) );
  XNOR U19257 ( .A(n16365), .B(n16366), .Z(n16364) );
  ANDN U19258 ( .B(n16367), .A(n16368), .Z(n16365) );
  XNOR U19259 ( .A(n16369), .B(n16370), .Z(n16367) );
  IV U19260 ( .A(n16334), .Z(n16331) );
  XOR U19261 ( .A(n16371), .B(n16372), .Z(n16334) );
  ANDN U19262 ( .B(n16373), .A(n16374), .Z(n16371) );
  XOR U19263 ( .A(n16372), .B(n16375), .Z(n16373) );
  XOR U19264 ( .A(n16376), .B(n16377), .Z(n16347) );
  XNOR U19265 ( .A(n16342), .B(n16378), .Z(n16377) );
  IV U19266 ( .A(n16345), .Z(n16378) );
  XOR U19267 ( .A(n16379), .B(n16380), .Z(n16345) );
  ANDN U19268 ( .B(n16381), .A(n16382), .Z(n16379) );
  XOR U19269 ( .A(n16380), .B(n16383), .Z(n16381) );
  XNOR U19270 ( .A(n16384), .B(n16385), .Z(n16342) );
  ANDN U19271 ( .B(n16386), .A(n16387), .Z(n16384) );
  XOR U19272 ( .A(n16385), .B(n16388), .Z(n16386) );
  IV U19273 ( .A(n16341), .Z(n16376) );
  XOR U19274 ( .A(n16339), .B(n16389), .Z(n16341) );
  XNOR U19275 ( .A(n16390), .B(n16391), .Z(n16389) );
  ANDN U19276 ( .B(n16392), .A(n16393), .Z(n16390) );
  XNOR U19277 ( .A(n16394), .B(n16395), .Z(n16392) );
  IV U19278 ( .A(n16343), .Z(n16339) );
  XOR U19279 ( .A(n16396), .B(n16397), .Z(n16343) );
  ANDN U19280 ( .B(n16398), .A(n16399), .Z(n16396) );
  XOR U19281 ( .A(n16400), .B(n16397), .Z(n16398) );
  XOR U19282 ( .A(n16354), .B(n16207), .Z(n16355) );
  XOR U19283 ( .A(n16401), .B(n16402), .Z(n16207) );
  AND U19284 ( .A(n96), .B(n16403), .Z(n16401) );
  XOR U19285 ( .A(n16404), .B(n16402), .Z(n16403) );
  XNOR U19286 ( .A(n16405), .B(n16406), .Z(n16354) );
  NAND U19287 ( .A(n16407), .B(n16408), .Z(n16406) );
  XOR U19288 ( .A(n16409), .B(n16306), .Z(n16408) );
  XOR U19289 ( .A(n16382), .B(n16383), .Z(n16306) );
  XOR U19290 ( .A(n16410), .B(n16375), .Z(n16383) );
  XOR U19291 ( .A(n16411), .B(n16363), .Z(n16375) );
  XOR U19292 ( .A(n16412), .B(n16413), .Z(n16363) );
  ANDN U19293 ( .B(n16414), .A(n16415), .Z(n16412) );
  XOR U19294 ( .A(n16413), .B(n16416), .Z(n16414) );
  IV U19295 ( .A(n16361), .Z(n16411) );
  XOR U19296 ( .A(n16359), .B(n16417), .Z(n16361) );
  XOR U19297 ( .A(n16418), .B(n16419), .Z(n16417) );
  ANDN U19298 ( .B(n16420), .A(n16421), .Z(n16418) );
  XOR U19299 ( .A(n16422), .B(n16419), .Z(n16420) );
  IV U19300 ( .A(n16362), .Z(n16359) );
  XOR U19301 ( .A(n16423), .B(n16424), .Z(n16362) );
  ANDN U19302 ( .B(n16425), .A(n16426), .Z(n16423) );
  XOR U19303 ( .A(n16424), .B(n16427), .Z(n16425) );
  IV U19304 ( .A(n16374), .Z(n16410) );
  XOR U19305 ( .A(n16428), .B(n16429), .Z(n16374) );
  XNOR U19306 ( .A(n16369), .B(n16430), .Z(n16429) );
  IV U19307 ( .A(n16372), .Z(n16430) );
  XOR U19308 ( .A(n16431), .B(n16432), .Z(n16372) );
  ANDN U19309 ( .B(n16433), .A(n16434), .Z(n16431) );
  XOR U19310 ( .A(n16432), .B(n16435), .Z(n16433) );
  XNOR U19311 ( .A(n16436), .B(n16437), .Z(n16369) );
  ANDN U19312 ( .B(n16438), .A(n16439), .Z(n16436) );
  XOR U19313 ( .A(n16437), .B(n16440), .Z(n16438) );
  IV U19314 ( .A(n16368), .Z(n16428) );
  XOR U19315 ( .A(n16366), .B(n16441), .Z(n16368) );
  XOR U19316 ( .A(n16442), .B(n16443), .Z(n16441) );
  ANDN U19317 ( .B(n16444), .A(n16445), .Z(n16442) );
  XOR U19318 ( .A(n16446), .B(n16443), .Z(n16444) );
  IV U19319 ( .A(n16370), .Z(n16366) );
  XOR U19320 ( .A(n16447), .B(n16448), .Z(n16370) );
  ANDN U19321 ( .B(n16449), .A(n16450), .Z(n16447) );
  XOR U19322 ( .A(n16451), .B(n16448), .Z(n16449) );
  XOR U19323 ( .A(n16452), .B(n16453), .Z(n16382) );
  XOR U19324 ( .A(n16400), .B(n16454), .Z(n16453) );
  IV U19325 ( .A(n16380), .Z(n16454) );
  XOR U19326 ( .A(n16455), .B(n16456), .Z(n16380) );
  ANDN U19327 ( .B(n16457), .A(n16458), .Z(n16455) );
  XOR U19328 ( .A(n16456), .B(n16459), .Z(n16457) );
  XOR U19329 ( .A(n16460), .B(n16388), .Z(n16400) );
  XOR U19330 ( .A(n16461), .B(n16462), .Z(n16388) );
  ANDN U19331 ( .B(n16463), .A(n16464), .Z(n16461) );
  XOR U19332 ( .A(n16462), .B(n16465), .Z(n16463) );
  IV U19333 ( .A(n16387), .Z(n16460) );
  XOR U19334 ( .A(n16466), .B(n16467), .Z(n16387) );
  XOR U19335 ( .A(n16468), .B(n16469), .Z(n16467) );
  ANDN U19336 ( .B(n16470), .A(n16471), .Z(n16468) );
  XOR U19337 ( .A(n16472), .B(n16469), .Z(n16470) );
  IV U19338 ( .A(n16385), .Z(n16466) );
  XOR U19339 ( .A(n16473), .B(n16474), .Z(n16385) );
  ANDN U19340 ( .B(n16475), .A(n16476), .Z(n16473) );
  XOR U19341 ( .A(n16474), .B(n16477), .Z(n16475) );
  IV U19342 ( .A(n16399), .Z(n16452) );
  XOR U19343 ( .A(n16478), .B(n16479), .Z(n16399) );
  XNOR U19344 ( .A(n16394), .B(n16480), .Z(n16479) );
  IV U19345 ( .A(n16397), .Z(n16480) );
  XOR U19346 ( .A(n16481), .B(n16482), .Z(n16397) );
  ANDN U19347 ( .B(n16483), .A(n16484), .Z(n16481) );
  XOR U19348 ( .A(n16485), .B(n16482), .Z(n16483) );
  XNOR U19349 ( .A(n16486), .B(n16487), .Z(n16394) );
  ANDN U19350 ( .B(n16488), .A(n16489), .Z(n16486) );
  XOR U19351 ( .A(n16487), .B(n16490), .Z(n16488) );
  IV U19352 ( .A(n16393), .Z(n16478) );
  XOR U19353 ( .A(n16391), .B(n16491), .Z(n16393) );
  XOR U19354 ( .A(n16492), .B(n16493), .Z(n16491) );
  ANDN U19355 ( .B(n16494), .A(n16495), .Z(n16492) );
  XOR U19356 ( .A(n16496), .B(n16493), .Z(n16494) );
  IV U19357 ( .A(n16395), .Z(n16391) );
  XOR U19358 ( .A(n16497), .B(n16498), .Z(n16395) );
  ANDN U19359 ( .B(n16499), .A(n16500), .Z(n16497) );
  XOR U19360 ( .A(n16501), .B(n16498), .Z(n16499) );
  IV U19361 ( .A(n16405), .Z(n16409) );
  XOR U19362 ( .A(n16405), .B(n16308), .Z(n16407) );
  XOR U19363 ( .A(n16502), .B(n16503), .Z(n16308) );
  AND U19364 ( .A(n96), .B(n16504), .Z(n16502) );
  XOR U19365 ( .A(n16505), .B(n16503), .Z(n16504) );
  NANDN U19366 ( .A(n16310), .B(n16312), .Z(n16405) );
  XOR U19367 ( .A(n16506), .B(n16507), .Z(n16312) );
  AND U19368 ( .A(n96), .B(n16508), .Z(n16506) );
  XOR U19369 ( .A(n16507), .B(n16509), .Z(n16508) );
  XNOR U19370 ( .A(n16510), .B(n16511), .Z(n96) );
  AND U19371 ( .A(n16512), .B(n16513), .Z(n16510) );
  XOR U19372 ( .A(n16511), .B(n16323), .Z(n16513) );
  XNOR U19373 ( .A(n16514), .B(n16515), .Z(n16323) );
  ANDN U19374 ( .B(n16516), .A(n16517), .Z(n16514) );
  XOR U19375 ( .A(n16515), .B(n16518), .Z(n16516) );
  XNOR U19376 ( .A(n16511), .B(n16325), .Z(n16512) );
  XOR U19377 ( .A(n16519), .B(n16520), .Z(n16325) );
  AND U19378 ( .A(n100), .B(n16521), .Z(n16519) );
  XOR U19379 ( .A(n16522), .B(n16520), .Z(n16521) );
  XOR U19380 ( .A(n16523), .B(n16524), .Z(n16511) );
  AND U19381 ( .A(n16525), .B(n16526), .Z(n16523) );
  XOR U19382 ( .A(n16524), .B(n16350), .Z(n16526) );
  XOR U19383 ( .A(n16517), .B(n16518), .Z(n16350) );
  XNOR U19384 ( .A(n16527), .B(n16528), .Z(n16518) );
  ANDN U19385 ( .B(n16529), .A(n16530), .Z(n16527) );
  XOR U19386 ( .A(n16531), .B(n16532), .Z(n16529) );
  XOR U19387 ( .A(n16533), .B(n16534), .Z(n16517) );
  XNOR U19388 ( .A(n16535), .B(n16536), .Z(n16534) );
  ANDN U19389 ( .B(n16537), .A(n16538), .Z(n16535) );
  XNOR U19390 ( .A(n16539), .B(n16540), .Z(n16537) );
  IV U19391 ( .A(n16515), .Z(n16533) );
  XOR U19392 ( .A(n16541), .B(n16542), .Z(n16515) );
  ANDN U19393 ( .B(n16543), .A(n16544), .Z(n16541) );
  XOR U19394 ( .A(n16542), .B(n16545), .Z(n16543) );
  XNOR U19395 ( .A(n16524), .B(n16352), .Z(n16525) );
  XOR U19396 ( .A(n16546), .B(n16547), .Z(n16352) );
  AND U19397 ( .A(n100), .B(n16548), .Z(n16546) );
  XOR U19398 ( .A(n16549), .B(n16547), .Z(n16548) );
  XNOR U19399 ( .A(n16550), .B(n16551), .Z(n16524) );
  AND U19400 ( .A(n16552), .B(n16553), .Z(n16550) );
  XNOR U19401 ( .A(n16551), .B(n16402), .Z(n16553) );
  XOR U19402 ( .A(n16544), .B(n16545), .Z(n16402) );
  XOR U19403 ( .A(n16554), .B(n16532), .Z(n16545) );
  XNOR U19404 ( .A(n16555), .B(n16556), .Z(n16532) );
  ANDN U19405 ( .B(n16557), .A(n16558), .Z(n16555) );
  XOR U19406 ( .A(n16559), .B(n16560), .Z(n16557) );
  IV U19407 ( .A(n16530), .Z(n16554) );
  XOR U19408 ( .A(n16528), .B(n16561), .Z(n16530) );
  XNOR U19409 ( .A(n16562), .B(n16563), .Z(n16561) );
  ANDN U19410 ( .B(n16564), .A(n16565), .Z(n16562) );
  XNOR U19411 ( .A(n16566), .B(n16567), .Z(n16564) );
  IV U19412 ( .A(n16531), .Z(n16528) );
  XOR U19413 ( .A(n16568), .B(n16569), .Z(n16531) );
  ANDN U19414 ( .B(n16570), .A(n16571), .Z(n16568) );
  XOR U19415 ( .A(n16569), .B(n16572), .Z(n16570) );
  XOR U19416 ( .A(n16573), .B(n16574), .Z(n16544) );
  XNOR U19417 ( .A(n16539), .B(n16575), .Z(n16574) );
  IV U19418 ( .A(n16542), .Z(n16575) );
  XOR U19419 ( .A(n16576), .B(n16577), .Z(n16542) );
  ANDN U19420 ( .B(n16578), .A(n16579), .Z(n16576) );
  XOR U19421 ( .A(n16577), .B(n16580), .Z(n16578) );
  XNOR U19422 ( .A(n16581), .B(n16582), .Z(n16539) );
  ANDN U19423 ( .B(n16583), .A(n16584), .Z(n16581) );
  XOR U19424 ( .A(n16582), .B(n16585), .Z(n16583) );
  IV U19425 ( .A(n16538), .Z(n16573) );
  XOR U19426 ( .A(n16536), .B(n16586), .Z(n16538) );
  XNOR U19427 ( .A(n16587), .B(n16588), .Z(n16586) );
  ANDN U19428 ( .B(n16589), .A(n16590), .Z(n16587) );
  XNOR U19429 ( .A(n16591), .B(n16592), .Z(n16589) );
  IV U19430 ( .A(n16540), .Z(n16536) );
  XOR U19431 ( .A(n16593), .B(n16594), .Z(n16540) );
  ANDN U19432 ( .B(n16595), .A(n16596), .Z(n16593) );
  XOR U19433 ( .A(n16597), .B(n16594), .Z(n16595) );
  XOR U19434 ( .A(n16551), .B(n16404), .Z(n16552) );
  XOR U19435 ( .A(n16598), .B(n16599), .Z(n16404) );
  AND U19436 ( .A(n100), .B(n16600), .Z(n16598) );
  XOR U19437 ( .A(n16601), .B(n16599), .Z(n16600) );
  XNOR U19438 ( .A(n16602), .B(n16603), .Z(n16551) );
  NAND U19439 ( .A(n16604), .B(n16605), .Z(n16603) );
  XOR U19440 ( .A(n16606), .B(n16503), .Z(n16605) );
  XOR U19441 ( .A(n16579), .B(n16580), .Z(n16503) );
  XOR U19442 ( .A(n16607), .B(n16572), .Z(n16580) );
  XOR U19443 ( .A(n16608), .B(n16560), .Z(n16572) );
  XOR U19444 ( .A(n16609), .B(n16610), .Z(n16560) );
  ANDN U19445 ( .B(n16611), .A(n16612), .Z(n16609) );
  XOR U19446 ( .A(n16610), .B(n16613), .Z(n16611) );
  IV U19447 ( .A(n16558), .Z(n16608) );
  XOR U19448 ( .A(n16556), .B(n16614), .Z(n16558) );
  XOR U19449 ( .A(n16615), .B(n16616), .Z(n16614) );
  ANDN U19450 ( .B(n16617), .A(n16618), .Z(n16615) );
  XOR U19451 ( .A(n16619), .B(n16616), .Z(n16617) );
  IV U19452 ( .A(n16559), .Z(n16556) );
  XOR U19453 ( .A(n16620), .B(n16621), .Z(n16559) );
  ANDN U19454 ( .B(n16622), .A(n16623), .Z(n16620) );
  XOR U19455 ( .A(n16621), .B(n16624), .Z(n16622) );
  IV U19456 ( .A(n16571), .Z(n16607) );
  XOR U19457 ( .A(n16625), .B(n16626), .Z(n16571) );
  XNOR U19458 ( .A(n16566), .B(n16627), .Z(n16626) );
  IV U19459 ( .A(n16569), .Z(n16627) );
  XOR U19460 ( .A(n16628), .B(n16629), .Z(n16569) );
  ANDN U19461 ( .B(n16630), .A(n16631), .Z(n16628) );
  XOR U19462 ( .A(n16629), .B(n16632), .Z(n16630) );
  XNOR U19463 ( .A(n16633), .B(n16634), .Z(n16566) );
  ANDN U19464 ( .B(n16635), .A(n16636), .Z(n16633) );
  XOR U19465 ( .A(n16634), .B(n16637), .Z(n16635) );
  IV U19466 ( .A(n16565), .Z(n16625) );
  XOR U19467 ( .A(n16563), .B(n16638), .Z(n16565) );
  XOR U19468 ( .A(n16639), .B(n16640), .Z(n16638) );
  ANDN U19469 ( .B(n16641), .A(n16642), .Z(n16639) );
  XOR U19470 ( .A(n16643), .B(n16640), .Z(n16641) );
  IV U19471 ( .A(n16567), .Z(n16563) );
  XOR U19472 ( .A(n16644), .B(n16645), .Z(n16567) );
  ANDN U19473 ( .B(n16646), .A(n16647), .Z(n16644) );
  XOR U19474 ( .A(n16648), .B(n16645), .Z(n16646) );
  XOR U19475 ( .A(n16649), .B(n16650), .Z(n16579) );
  XOR U19476 ( .A(n16597), .B(n16651), .Z(n16650) );
  IV U19477 ( .A(n16577), .Z(n16651) );
  XOR U19478 ( .A(n16652), .B(n16653), .Z(n16577) );
  ANDN U19479 ( .B(n16654), .A(n16655), .Z(n16652) );
  XOR U19480 ( .A(n16653), .B(n16656), .Z(n16654) );
  XOR U19481 ( .A(n16657), .B(n16585), .Z(n16597) );
  XOR U19482 ( .A(n16658), .B(n16659), .Z(n16585) );
  ANDN U19483 ( .B(n16660), .A(n16661), .Z(n16658) );
  XOR U19484 ( .A(n16659), .B(n16662), .Z(n16660) );
  IV U19485 ( .A(n16584), .Z(n16657) );
  XOR U19486 ( .A(n16663), .B(n16664), .Z(n16584) );
  XOR U19487 ( .A(n16665), .B(n16666), .Z(n16664) );
  ANDN U19488 ( .B(n16667), .A(n16668), .Z(n16665) );
  XOR U19489 ( .A(n16669), .B(n16666), .Z(n16667) );
  IV U19490 ( .A(n16582), .Z(n16663) );
  XOR U19491 ( .A(n16670), .B(n16671), .Z(n16582) );
  ANDN U19492 ( .B(n16672), .A(n16673), .Z(n16670) );
  XOR U19493 ( .A(n16671), .B(n16674), .Z(n16672) );
  IV U19494 ( .A(n16596), .Z(n16649) );
  XOR U19495 ( .A(n16675), .B(n16676), .Z(n16596) );
  XNOR U19496 ( .A(n16591), .B(n16677), .Z(n16676) );
  IV U19497 ( .A(n16594), .Z(n16677) );
  XOR U19498 ( .A(n16678), .B(n16679), .Z(n16594) );
  ANDN U19499 ( .B(n16680), .A(n16681), .Z(n16678) );
  XOR U19500 ( .A(n16682), .B(n16679), .Z(n16680) );
  XNOR U19501 ( .A(n16683), .B(n16684), .Z(n16591) );
  ANDN U19502 ( .B(n16685), .A(n16686), .Z(n16683) );
  XOR U19503 ( .A(n16684), .B(n16687), .Z(n16685) );
  IV U19504 ( .A(n16590), .Z(n16675) );
  XOR U19505 ( .A(n16588), .B(n16688), .Z(n16590) );
  XOR U19506 ( .A(n16689), .B(n16690), .Z(n16688) );
  ANDN U19507 ( .B(n16691), .A(n16692), .Z(n16689) );
  XOR U19508 ( .A(n16693), .B(n16690), .Z(n16691) );
  IV U19509 ( .A(n16592), .Z(n16588) );
  XOR U19510 ( .A(n16694), .B(n16695), .Z(n16592) );
  ANDN U19511 ( .B(n16696), .A(n16697), .Z(n16694) );
  XOR U19512 ( .A(n16698), .B(n16695), .Z(n16696) );
  IV U19513 ( .A(n16602), .Z(n16606) );
  XOR U19514 ( .A(n16602), .B(n16505), .Z(n16604) );
  XOR U19515 ( .A(n16699), .B(n16700), .Z(n16505) );
  AND U19516 ( .A(n100), .B(n16701), .Z(n16699) );
  XOR U19517 ( .A(n16702), .B(n16700), .Z(n16701) );
  NANDN U19518 ( .A(n16507), .B(n16509), .Z(n16602) );
  XOR U19519 ( .A(n16703), .B(n16704), .Z(n16509) );
  AND U19520 ( .A(n100), .B(n16705), .Z(n16703) );
  XOR U19521 ( .A(n16704), .B(n16706), .Z(n16705) );
  XNOR U19522 ( .A(n16707), .B(n16708), .Z(n100) );
  AND U19523 ( .A(n16709), .B(n16710), .Z(n16707) );
  XOR U19524 ( .A(n16708), .B(n16520), .Z(n16710) );
  XNOR U19525 ( .A(n16711), .B(n16712), .Z(n16520) );
  ANDN U19526 ( .B(n16713), .A(n16714), .Z(n16711) );
  XOR U19527 ( .A(n16712), .B(n16715), .Z(n16713) );
  XNOR U19528 ( .A(n16708), .B(n16522), .Z(n16709) );
  XOR U19529 ( .A(n16716), .B(n16717), .Z(n16522) );
  AND U19530 ( .A(n104), .B(n16718), .Z(n16716) );
  XOR U19531 ( .A(n16719), .B(n16717), .Z(n16718) );
  XOR U19532 ( .A(n16720), .B(n16721), .Z(n16708) );
  AND U19533 ( .A(n16722), .B(n16723), .Z(n16720) );
  XOR U19534 ( .A(n16721), .B(n16547), .Z(n16723) );
  XOR U19535 ( .A(n16714), .B(n16715), .Z(n16547) );
  XNOR U19536 ( .A(n16724), .B(n16725), .Z(n16715) );
  ANDN U19537 ( .B(n16726), .A(n16727), .Z(n16724) );
  XOR U19538 ( .A(n16728), .B(n16729), .Z(n16726) );
  XOR U19539 ( .A(n16730), .B(n16731), .Z(n16714) );
  XNOR U19540 ( .A(n16732), .B(n16733), .Z(n16731) );
  ANDN U19541 ( .B(n16734), .A(n16735), .Z(n16732) );
  XNOR U19542 ( .A(n16736), .B(n16737), .Z(n16734) );
  IV U19543 ( .A(n16712), .Z(n16730) );
  XOR U19544 ( .A(n16738), .B(n16739), .Z(n16712) );
  ANDN U19545 ( .B(n16740), .A(n16741), .Z(n16738) );
  XOR U19546 ( .A(n16739), .B(n16742), .Z(n16740) );
  XNOR U19547 ( .A(n16721), .B(n16549), .Z(n16722) );
  XOR U19548 ( .A(n16743), .B(n16744), .Z(n16549) );
  AND U19549 ( .A(n104), .B(n16745), .Z(n16743) );
  XOR U19550 ( .A(n16746), .B(n16744), .Z(n16745) );
  XNOR U19551 ( .A(n16747), .B(n16748), .Z(n16721) );
  AND U19552 ( .A(n16749), .B(n16750), .Z(n16747) );
  XNOR U19553 ( .A(n16748), .B(n16599), .Z(n16750) );
  XOR U19554 ( .A(n16741), .B(n16742), .Z(n16599) );
  XOR U19555 ( .A(n16751), .B(n16729), .Z(n16742) );
  XNOR U19556 ( .A(n16752), .B(n16753), .Z(n16729) );
  ANDN U19557 ( .B(n16754), .A(n16755), .Z(n16752) );
  XOR U19558 ( .A(n16756), .B(n16757), .Z(n16754) );
  IV U19559 ( .A(n16727), .Z(n16751) );
  XOR U19560 ( .A(n16725), .B(n16758), .Z(n16727) );
  XNOR U19561 ( .A(n16759), .B(n16760), .Z(n16758) );
  ANDN U19562 ( .B(n16761), .A(n16762), .Z(n16759) );
  XNOR U19563 ( .A(n16763), .B(n16764), .Z(n16761) );
  IV U19564 ( .A(n16728), .Z(n16725) );
  XOR U19565 ( .A(n16765), .B(n16766), .Z(n16728) );
  ANDN U19566 ( .B(n16767), .A(n16768), .Z(n16765) );
  XOR U19567 ( .A(n16766), .B(n16769), .Z(n16767) );
  XOR U19568 ( .A(n16770), .B(n16771), .Z(n16741) );
  XNOR U19569 ( .A(n16736), .B(n16772), .Z(n16771) );
  IV U19570 ( .A(n16739), .Z(n16772) );
  XOR U19571 ( .A(n16773), .B(n16774), .Z(n16739) );
  ANDN U19572 ( .B(n16775), .A(n16776), .Z(n16773) );
  XOR U19573 ( .A(n16774), .B(n16777), .Z(n16775) );
  XNOR U19574 ( .A(n16778), .B(n16779), .Z(n16736) );
  ANDN U19575 ( .B(n16780), .A(n16781), .Z(n16778) );
  XOR U19576 ( .A(n16779), .B(n16782), .Z(n16780) );
  IV U19577 ( .A(n16735), .Z(n16770) );
  XOR U19578 ( .A(n16733), .B(n16783), .Z(n16735) );
  XNOR U19579 ( .A(n16784), .B(n16785), .Z(n16783) );
  ANDN U19580 ( .B(n16786), .A(n16787), .Z(n16784) );
  XNOR U19581 ( .A(n16788), .B(n16789), .Z(n16786) );
  IV U19582 ( .A(n16737), .Z(n16733) );
  XOR U19583 ( .A(n16790), .B(n16791), .Z(n16737) );
  ANDN U19584 ( .B(n16792), .A(n16793), .Z(n16790) );
  XOR U19585 ( .A(n16794), .B(n16791), .Z(n16792) );
  XOR U19586 ( .A(n16748), .B(n16601), .Z(n16749) );
  XOR U19587 ( .A(n16795), .B(n16796), .Z(n16601) );
  AND U19588 ( .A(n104), .B(n16797), .Z(n16795) );
  XOR U19589 ( .A(n16798), .B(n16796), .Z(n16797) );
  XNOR U19590 ( .A(n16799), .B(n16800), .Z(n16748) );
  NAND U19591 ( .A(n16801), .B(n16802), .Z(n16800) );
  XOR U19592 ( .A(n16803), .B(n16700), .Z(n16802) );
  XOR U19593 ( .A(n16776), .B(n16777), .Z(n16700) );
  XOR U19594 ( .A(n16804), .B(n16769), .Z(n16777) );
  XOR U19595 ( .A(n16805), .B(n16757), .Z(n16769) );
  XOR U19596 ( .A(n16806), .B(n16807), .Z(n16757) );
  ANDN U19597 ( .B(n16808), .A(n16809), .Z(n16806) );
  XOR U19598 ( .A(n16807), .B(n16810), .Z(n16808) );
  IV U19599 ( .A(n16755), .Z(n16805) );
  XOR U19600 ( .A(n16753), .B(n16811), .Z(n16755) );
  XOR U19601 ( .A(n16812), .B(n16813), .Z(n16811) );
  ANDN U19602 ( .B(n16814), .A(n16815), .Z(n16812) );
  XOR U19603 ( .A(n16816), .B(n16813), .Z(n16814) );
  IV U19604 ( .A(n16756), .Z(n16753) );
  XOR U19605 ( .A(n16817), .B(n16818), .Z(n16756) );
  ANDN U19606 ( .B(n16819), .A(n16820), .Z(n16817) );
  XOR U19607 ( .A(n16818), .B(n16821), .Z(n16819) );
  IV U19608 ( .A(n16768), .Z(n16804) );
  XOR U19609 ( .A(n16822), .B(n16823), .Z(n16768) );
  XNOR U19610 ( .A(n16763), .B(n16824), .Z(n16823) );
  IV U19611 ( .A(n16766), .Z(n16824) );
  XOR U19612 ( .A(n16825), .B(n16826), .Z(n16766) );
  ANDN U19613 ( .B(n16827), .A(n16828), .Z(n16825) );
  XOR U19614 ( .A(n16826), .B(n16829), .Z(n16827) );
  XNOR U19615 ( .A(n16830), .B(n16831), .Z(n16763) );
  ANDN U19616 ( .B(n16832), .A(n16833), .Z(n16830) );
  XOR U19617 ( .A(n16831), .B(n16834), .Z(n16832) );
  IV U19618 ( .A(n16762), .Z(n16822) );
  XOR U19619 ( .A(n16760), .B(n16835), .Z(n16762) );
  XOR U19620 ( .A(n16836), .B(n16837), .Z(n16835) );
  ANDN U19621 ( .B(n16838), .A(n16839), .Z(n16836) );
  XOR U19622 ( .A(n16840), .B(n16837), .Z(n16838) );
  IV U19623 ( .A(n16764), .Z(n16760) );
  XOR U19624 ( .A(n16841), .B(n16842), .Z(n16764) );
  ANDN U19625 ( .B(n16843), .A(n16844), .Z(n16841) );
  XOR U19626 ( .A(n16845), .B(n16842), .Z(n16843) );
  XOR U19627 ( .A(n16846), .B(n16847), .Z(n16776) );
  XOR U19628 ( .A(n16794), .B(n16848), .Z(n16847) );
  IV U19629 ( .A(n16774), .Z(n16848) );
  XOR U19630 ( .A(n16849), .B(n16850), .Z(n16774) );
  ANDN U19631 ( .B(n16851), .A(n16852), .Z(n16849) );
  XOR U19632 ( .A(n16850), .B(n16853), .Z(n16851) );
  XOR U19633 ( .A(n16854), .B(n16782), .Z(n16794) );
  XOR U19634 ( .A(n16855), .B(n16856), .Z(n16782) );
  ANDN U19635 ( .B(n16857), .A(n16858), .Z(n16855) );
  XOR U19636 ( .A(n16856), .B(n16859), .Z(n16857) );
  IV U19637 ( .A(n16781), .Z(n16854) );
  XOR U19638 ( .A(n16860), .B(n16861), .Z(n16781) );
  XOR U19639 ( .A(n16862), .B(n16863), .Z(n16861) );
  ANDN U19640 ( .B(n16864), .A(n16865), .Z(n16862) );
  XOR U19641 ( .A(n16866), .B(n16863), .Z(n16864) );
  IV U19642 ( .A(n16779), .Z(n16860) );
  XOR U19643 ( .A(n16867), .B(n16868), .Z(n16779) );
  ANDN U19644 ( .B(n16869), .A(n16870), .Z(n16867) );
  XOR U19645 ( .A(n16868), .B(n16871), .Z(n16869) );
  IV U19646 ( .A(n16793), .Z(n16846) );
  XOR U19647 ( .A(n16872), .B(n16873), .Z(n16793) );
  XNOR U19648 ( .A(n16788), .B(n16874), .Z(n16873) );
  IV U19649 ( .A(n16791), .Z(n16874) );
  XOR U19650 ( .A(n16875), .B(n16876), .Z(n16791) );
  ANDN U19651 ( .B(n16877), .A(n16878), .Z(n16875) );
  XOR U19652 ( .A(n16879), .B(n16876), .Z(n16877) );
  XNOR U19653 ( .A(n16880), .B(n16881), .Z(n16788) );
  ANDN U19654 ( .B(n16882), .A(n16883), .Z(n16880) );
  XOR U19655 ( .A(n16881), .B(n16884), .Z(n16882) );
  IV U19656 ( .A(n16787), .Z(n16872) );
  XOR U19657 ( .A(n16785), .B(n16885), .Z(n16787) );
  XOR U19658 ( .A(n16886), .B(n16887), .Z(n16885) );
  ANDN U19659 ( .B(n16888), .A(n16889), .Z(n16886) );
  XOR U19660 ( .A(n16890), .B(n16887), .Z(n16888) );
  IV U19661 ( .A(n16789), .Z(n16785) );
  XOR U19662 ( .A(n16891), .B(n16892), .Z(n16789) );
  ANDN U19663 ( .B(n16893), .A(n16894), .Z(n16891) );
  XOR U19664 ( .A(n16895), .B(n16892), .Z(n16893) );
  IV U19665 ( .A(n16799), .Z(n16803) );
  XOR U19666 ( .A(n16799), .B(n16702), .Z(n16801) );
  XOR U19667 ( .A(n16896), .B(n16897), .Z(n16702) );
  AND U19668 ( .A(n104), .B(n16898), .Z(n16896) );
  XOR U19669 ( .A(n16899), .B(n16897), .Z(n16898) );
  NANDN U19670 ( .A(n16704), .B(n16706), .Z(n16799) );
  XOR U19671 ( .A(n16900), .B(n16901), .Z(n16706) );
  AND U19672 ( .A(n104), .B(n16902), .Z(n16900) );
  XOR U19673 ( .A(n16901), .B(n16903), .Z(n16902) );
  XNOR U19674 ( .A(n16904), .B(n16905), .Z(n104) );
  AND U19675 ( .A(n16906), .B(n16907), .Z(n16904) );
  XOR U19676 ( .A(n16905), .B(n16717), .Z(n16907) );
  XNOR U19677 ( .A(n16908), .B(n16909), .Z(n16717) );
  ANDN U19678 ( .B(n16910), .A(n16911), .Z(n16908) );
  XOR U19679 ( .A(n16909), .B(n16912), .Z(n16910) );
  XNOR U19680 ( .A(n16905), .B(n16719), .Z(n16906) );
  XOR U19681 ( .A(n16913), .B(n16914), .Z(n16719) );
  AND U19682 ( .A(n108), .B(n16915), .Z(n16913) );
  XOR U19683 ( .A(n16916), .B(n16914), .Z(n16915) );
  XOR U19684 ( .A(n16917), .B(n16918), .Z(n16905) );
  AND U19685 ( .A(n16919), .B(n16920), .Z(n16917) );
  XOR U19686 ( .A(n16918), .B(n16744), .Z(n16920) );
  XOR U19687 ( .A(n16911), .B(n16912), .Z(n16744) );
  XNOR U19688 ( .A(n16921), .B(n16922), .Z(n16912) );
  ANDN U19689 ( .B(n16923), .A(n16924), .Z(n16921) );
  XOR U19690 ( .A(n16925), .B(n16926), .Z(n16923) );
  XOR U19691 ( .A(n16927), .B(n16928), .Z(n16911) );
  XNOR U19692 ( .A(n16929), .B(n16930), .Z(n16928) );
  ANDN U19693 ( .B(n16931), .A(n16932), .Z(n16929) );
  XNOR U19694 ( .A(n16933), .B(n16934), .Z(n16931) );
  IV U19695 ( .A(n16909), .Z(n16927) );
  XOR U19696 ( .A(n16935), .B(n16936), .Z(n16909) );
  ANDN U19697 ( .B(n16937), .A(n16938), .Z(n16935) );
  XOR U19698 ( .A(n16936), .B(n16939), .Z(n16937) );
  XNOR U19699 ( .A(n16918), .B(n16746), .Z(n16919) );
  XOR U19700 ( .A(n16940), .B(n16941), .Z(n16746) );
  AND U19701 ( .A(n108), .B(n16942), .Z(n16940) );
  XOR U19702 ( .A(n16943), .B(n16941), .Z(n16942) );
  XNOR U19703 ( .A(n16944), .B(n16945), .Z(n16918) );
  AND U19704 ( .A(n16946), .B(n16947), .Z(n16944) );
  XNOR U19705 ( .A(n16945), .B(n16796), .Z(n16947) );
  XOR U19706 ( .A(n16938), .B(n16939), .Z(n16796) );
  XOR U19707 ( .A(n16948), .B(n16926), .Z(n16939) );
  XNOR U19708 ( .A(n16949), .B(n16950), .Z(n16926) );
  ANDN U19709 ( .B(n16951), .A(n16952), .Z(n16949) );
  XOR U19710 ( .A(n16953), .B(n16954), .Z(n16951) );
  IV U19711 ( .A(n16924), .Z(n16948) );
  XOR U19712 ( .A(n16922), .B(n16955), .Z(n16924) );
  XNOR U19713 ( .A(n16956), .B(n16957), .Z(n16955) );
  ANDN U19714 ( .B(n16958), .A(n16959), .Z(n16956) );
  XNOR U19715 ( .A(n16960), .B(n16961), .Z(n16958) );
  IV U19716 ( .A(n16925), .Z(n16922) );
  XOR U19717 ( .A(n16962), .B(n16963), .Z(n16925) );
  ANDN U19718 ( .B(n16964), .A(n16965), .Z(n16962) );
  XOR U19719 ( .A(n16963), .B(n16966), .Z(n16964) );
  XOR U19720 ( .A(n16967), .B(n16968), .Z(n16938) );
  XNOR U19721 ( .A(n16933), .B(n16969), .Z(n16968) );
  IV U19722 ( .A(n16936), .Z(n16969) );
  XOR U19723 ( .A(n16970), .B(n16971), .Z(n16936) );
  ANDN U19724 ( .B(n16972), .A(n16973), .Z(n16970) );
  XOR U19725 ( .A(n16971), .B(n16974), .Z(n16972) );
  XNOR U19726 ( .A(n16975), .B(n16976), .Z(n16933) );
  ANDN U19727 ( .B(n16977), .A(n16978), .Z(n16975) );
  XOR U19728 ( .A(n16976), .B(n16979), .Z(n16977) );
  IV U19729 ( .A(n16932), .Z(n16967) );
  XOR U19730 ( .A(n16930), .B(n16980), .Z(n16932) );
  XNOR U19731 ( .A(n16981), .B(n16982), .Z(n16980) );
  ANDN U19732 ( .B(n16983), .A(n16984), .Z(n16981) );
  XNOR U19733 ( .A(n16985), .B(n16986), .Z(n16983) );
  IV U19734 ( .A(n16934), .Z(n16930) );
  XOR U19735 ( .A(n16987), .B(n16988), .Z(n16934) );
  ANDN U19736 ( .B(n16989), .A(n16990), .Z(n16987) );
  XOR U19737 ( .A(n16991), .B(n16988), .Z(n16989) );
  XOR U19738 ( .A(n16945), .B(n16798), .Z(n16946) );
  XOR U19739 ( .A(n16992), .B(n16993), .Z(n16798) );
  AND U19740 ( .A(n108), .B(n16994), .Z(n16992) );
  XOR U19741 ( .A(n16995), .B(n16993), .Z(n16994) );
  XNOR U19742 ( .A(n16996), .B(n16997), .Z(n16945) );
  NAND U19743 ( .A(n16998), .B(n16999), .Z(n16997) );
  XOR U19744 ( .A(n17000), .B(n16897), .Z(n16999) );
  XOR U19745 ( .A(n16973), .B(n16974), .Z(n16897) );
  XOR U19746 ( .A(n17001), .B(n16966), .Z(n16974) );
  XOR U19747 ( .A(n17002), .B(n16954), .Z(n16966) );
  XOR U19748 ( .A(n17003), .B(n17004), .Z(n16954) );
  ANDN U19749 ( .B(n17005), .A(n17006), .Z(n17003) );
  XOR U19750 ( .A(n17004), .B(n17007), .Z(n17005) );
  IV U19751 ( .A(n16952), .Z(n17002) );
  XOR U19752 ( .A(n16950), .B(n17008), .Z(n16952) );
  XOR U19753 ( .A(n17009), .B(n17010), .Z(n17008) );
  ANDN U19754 ( .B(n17011), .A(n17012), .Z(n17009) );
  XOR U19755 ( .A(n17013), .B(n17010), .Z(n17011) );
  IV U19756 ( .A(n16953), .Z(n16950) );
  XOR U19757 ( .A(n17014), .B(n17015), .Z(n16953) );
  ANDN U19758 ( .B(n17016), .A(n17017), .Z(n17014) );
  XOR U19759 ( .A(n17015), .B(n17018), .Z(n17016) );
  IV U19760 ( .A(n16965), .Z(n17001) );
  XOR U19761 ( .A(n17019), .B(n17020), .Z(n16965) );
  XNOR U19762 ( .A(n16960), .B(n17021), .Z(n17020) );
  IV U19763 ( .A(n16963), .Z(n17021) );
  XOR U19764 ( .A(n17022), .B(n17023), .Z(n16963) );
  ANDN U19765 ( .B(n17024), .A(n17025), .Z(n17022) );
  XOR U19766 ( .A(n17023), .B(n17026), .Z(n17024) );
  XNOR U19767 ( .A(n17027), .B(n17028), .Z(n16960) );
  ANDN U19768 ( .B(n17029), .A(n17030), .Z(n17027) );
  XOR U19769 ( .A(n17028), .B(n17031), .Z(n17029) );
  IV U19770 ( .A(n16959), .Z(n17019) );
  XOR U19771 ( .A(n16957), .B(n17032), .Z(n16959) );
  XOR U19772 ( .A(n17033), .B(n17034), .Z(n17032) );
  ANDN U19773 ( .B(n17035), .A(n17036), .Z(n17033) );
  XOR U19774 ( .A(n17037), .B(n17034), .Z(n17035) );
  IV U19775 ( .A(n16961), .Z(n16957) );
  XOR U19776 ( .A(n17038), .B(n17039), .Z(n16961) );
  ANDN U19777 ( .B(n17040), .A(n17041), .Z(n17038) );
  XOR U19778 ( .A(n17042), .B(n17039), .Z(n17040) );
  XOR U19779 ( .A(n17043), .B(n17044), .Z(n16973) );
  XOR U19780 ( .A(n16991), .B(n17045), .Z(n17044) );
  IV U19781 ( .A(n16971), .Z(n17045) );
  XOR U19782 ( .A(n17046), .B(n17047), .Z(n16971) );
  ANDN U19783 ( .B(n17048), .A(n17049), .Z(n17046) );
  XOR U19784 ( .A(n17047), .B(n17050), .Z(n17048) );
  XOR U19785 ( .A(n17051), .B(n16979), .Z(n16991) );
  XOR U19786 ( .A(n17052), .B(n17053), .Z(n16979) );
  ANDN U19787 ( .B(n17054), .A(n17055), .Z(n17052) );
  XOR U19788 ( .A(n17053), .B(n17056), .Z(n17054) );
  IV U19789 ( .A(n16978), .Z(n17051) );
  XOR U19790 ( .A(n17057), .B(n17058), .Z(n16978) );
  XOR U19791 ( .A(n17059), .B(n17060), .Z(n17058) );
  ANDN U19792 ( .B(n17061), .A(n17062), .Z(n17059) );
  XOR U19793 ( .A(n17063), .B(n17060), .Z(n17061) );
  IV U19794 ( .A(n16976), .Z(n17057) );
  XOR U19795 ( .A(n17064), .B(n17065), .Z(n16976) );
  ANDN U19796 ( .B(n17066), .A(n17067), .Z(n17064) );
  XOR U19797 ( .A(n17065), .B(n17068), .Z(n17066) );
  IV U19798 ( .A(n16990), .Z(n17043) );
  XOR U19799 ( .A(n17069), .B(n17070), .Z(n16990) );
  XNOR U19800 ( .A(n16985), .B(n17071), .Z(n17070) );
  IV U19801 ( .A(n16988), .Z(n17071) );
  XOR U19802 ( .A(n17072), .B(n17073), .Z(n16988) );
  ANDN U19803 ( .B(n17074), .A(n17075), .Z(n17072) );
  XOR U19804 ( .A(n17076), .B(n17073), .Z(n17074) );
  XNOR U19805 ( .A(n17077), .B(n17078), .Z(n16985) );
  ANDN U19806 ( .B(n17079), .A(n17080), .Z(n17077) );
  XOR U19807 ( .A(n17078), .B(n17081), .Z(n17079) );
  IV U19808 ( .A(n16984), .Z(n17069) );
  XOR U19809 ( .A(n16982), .B(n17082), .Z(n16984) );
  XOR U19810 ( .A(n17083), .B(n17084), .Z(n17082) );
  ANDN U19811 ( .B(n17085), .A(n17086), .Z(n17083) );
  XOR U19812 ( .A(n17087), .B(n17084), .Z(n17085) );
  IV U19813 ( .A(n16986), .Z(n16982) );
  XOR U19814 ( .A(n17088), .B(n17089), .Z(n16986) );
  ANDN U19815 ( .B(n17090), .A(n17091), .Z(n17088) );
  XOR U19816 ( .A(n17092), .B(n17089), .Z(n17090) );
  IV U19817 ( .A(n16996), .Z(n17000) );
  XOR U19818 ( .A(n16996), .B(n16899), .Z(n16998) );
  XOR U19819 ( .A(n17093), .B(n17094), .Z(n16899) );
  AND U19820 ( .A(n108), .B(n17095), .Z(n17093) );
  XOR U19821 ( .A(n17096), .B(n17094), .Z(n17095) );
  NANDN U19822 ( .A(n16901), .B(n16903), .Z(n16996) );
  XOR U19823 ( .A(n17097), .B(n17098), .Z(n16903) );
  AND U19824 ( .A(n108), .B(n17099), .Z(n17097) );
  XOR U19825 ( .A(n17098), .B(n17100), .Z(n17099) );
  XNOR U19826 ( .A(n17101), .B(n17102), .Z(n108) );
  AND U19827 ( .A(n17103), .B(n17104), .Z(n17101) );
  XOR U19828 ( .A(n17102), .B(n16914), .Z(n17104) );
  XNOR U19829 ( .A(n17105), .B(n17106), .Z(n16914) );
  ANDN U19830 ( .B(n17107), .A(n17108), .Z(n17105) );
  XOR U19831 ( .A(n17106), .B(n17109), .Z(n17107) );
  XNOR U19832 ( .A(n17102), .B(n16916), .Z(n17103) );
  XOR U19833 ( .A(n17110), .B(n17111), .Z(n16916) );
  AND U19834 ( .A(n112), .B(n17112), .Z(n17110) );
  XOR U19835 ( .A(n17113), .B(n17111), .Z(n17112) );
  XOR U19836 ( .A(n17114), .B(n17115), .Z(n17102) );
  AND U19837 ( .A(n17116), .B(n17117), .Z(n17114) );
  XOR U19838 ( .A(n17115), .B(n16941), .Z(n17117) );
  XOR U19839 ( .A(n17108), .B(n17109), .Z(n16941) );
  XNOR U19840 ( .A(n17118), .B(n17119), .Z(n17109) );
  ANDN U19841 ( .B(n17120), .A(n17121), .Z(n17118) );
  XOR U19842 ( .A(n17122), .B(n17123), .Z(n17120) );
  XOR U19843 ( .A(n17124), .B(n17125), .Z(n17108) );
  XNOR U19844 ( .A(n17126), .B(n17127), .Z(n17125) );
  ANDN U19845 ( .B(n17128), .A(n17129), .Z(n17126) );
  XNOR U19846 ( .A(n17130), .B(n17131), .Z(n17128) );
  IV U19847 ( .A(n17106), .Z(n17124) );
  XOR U19848 ( .A(n17132), .B(n17133), .Z(n17106) );
  ANDN U19849 ( .B(n17134), .A(n17135), .Z(n17132) );
  XOR U19850 ( .A(n17133), .B(n17136), .Z(n17134) );
  XNOR U19851 ( .A(n17115), .B(n16943), .Z(n17116) );
  XOR U19852 ( .A(n17137), .B(n17138), .Z(n16943) );
  AND U19853 ( .A(n112), .B(n17139), .Z(n17137) );
  XOR U19854 ( .A(n17140), .B(n17138), .Z(n17139) );
  XNOR U19855 ( .A(n17141), .B(n17142), .Z(n17115) );
  AND U19856 ( .A(n17143), .B(n17144), .Z(n17141) );
  XNOR U19857 ( .A(n17142), .B(n16993), .Z(n17144) );
  XOR U19858 ( .A(n17135), .B(n17136), .Z(n16993) );
  XOR U19859 ( .A(n17145), .B(n17123), .Z(n17136) );
  XNOR U19860 ( .A(n17146), .B(n17147), .Z(n17123) );
  ANDN U19861 ( .B(n17148), .A(n17149), .Z(n17146) );
  XOR U19862 ( .A(n17150), .B(n17151), .Z(n17148) );
  IV U19863 ( .A(n17121), .Z(n17145) );
  XOR U19864 ( .A(n17119), .B(n17152), .Z(n17121) );
  XNOR U19865 ( .A(n17153), .B(n17154), .Z(n17152) );
  ANDN U19866 ( .B(n17155), .A(n17156), .Z(n17153) );
  XNOR U19867 ( .A(n17157), .B(n17158), .Z(n17155) );
  IV U19868 ( .A(n17122), .Z(n17119) );
  XOR U19869 ( .A(n17159), .B(n17160), .Z(n17122) );
  ANDN U19870 ( .B(n17161), .A(n17162), .Z(n17159) );
  XOR U19871 ( .A(n17160), .B(n17163), .Z(n17161) );
  XOR U19872 ( .A(n17164), .B(n17165), .Z(n17135) );
  XNOR U19873 ( .A(n17130), .B(n17166), .Z(n17165) );
  IV U19874 ( .A(n17133), .Z(n17166) );
  XOR U19875 ( .A(n17167), .B(n17168), .Z(n17133) );
  ANDN U19876 ( .B(n17169), .A(n17170), .Z(n17167) );
  XOR U19877 ( .A(n17168), .B(n17171), .Z(n17169) );
  XNOR U19878 ( .A(n17172), .B(n17173), .Z(n17130) );
  ANDN U19879 ( .B(n17174), .A(n17175), .Z(n17172) );
  XOR U19880 ( .A(n17173), .B(n17176), .Z(n17174) );
  IV U19881 ( .A(n17129), .Z(n17164) );
  XOR U19882 ( .A(n17127), .B(n17177), .Z(n17129) );
  XNOR U19883 ( .A(n17178), .B(n17179), .Z(n17177) );
  ANDN U19884 ( .B(n17180), .A(n17181), .Z(n17178) );
  XNOR U19885 ( .A(n17182), .B(n17183), .Z(n17180) );
  IV U19886 ( .A(n17131), .Z(n17127) );
  XOR U19887 ( .A(n17184), .B(n17185), .Z(n17131) );
  ANDN U19888 ( .B(n17186), .A(n17187), .Z(n17184) );
  XOR U19889 ( .A(n17188), .B(n17185), .Z(n17186) );
  XOR U19890 ( .A(n17142), .B(n16995), .Z(n17143) );
  XOR U19891 ( .A(n17189), .B(n17190), .Z(n16995) );
  AND U19892 ( .A(n112), .B(n17191), .Z(n17189) );
  XOR U19893 ( .A(n17192), .B(n17190), .Z(n17191) );
  XNOR U19894 ( .A(n17193), .B(n17194), .Z(n17142) );
  NAND U19895 ( .A(n17195), .B(n17196), .Z(n17194) );
  XOR U19896 ( .A(n17197), .B(n17094), .Z(n17196) );
  XOR U19897 ( .A(n17170), .B(n17171), .Z(n17094) );
  XOR U19898 ( .A(n17198), .B(n17163), .Z(n17171) );
  XOR U19899 ( .A(n17199), .B(n17151), .Z(n17163) );
  XOR U19900 ( .A(n17200), .B(n17201), .Z(n17151) );
  ANDN U19901 ( .B(n17202), .A(n17203), .Z(n17200) );
  XOR U19902 ( .A(n17201), .B(n17204), .Z(n17202) );
  IV U19903 ( .A(n17149), .Z(n17199) );
  XOR U19904 ( .A(n17147), .B(n17205), .Z(n17149) );
  XOR U19905 ( .A(n17206), .B(n17207), .Z(n17205) );
  ANDN U19906 ( .B(n17208), .A(n17209), .Z(n17206) );
  XOR U19907 ( .A(n17210), .B(n17207), .Z(n17208) );
  IV U19908 ( .A(n17150), .Z(n17147) );
  XOR U19909 ( .A(n17211), .B(n17212), .Z(n17150) );
  ANDN U19910 ( .B(n17213), .A(n17214), .Z(n17211) );
  XOR U19911 ( .A(n17212), .B(n17215), .Z(n17213) );
  IV U19912 ( .A(n17162), .Z(n17198) );
  XOR U19913 ( .A(n17216), .B(n17217), .Z(n17162) );
  XNOR U19914 ( .A(n17157), .B(n17218), .Z(n17217) );
  IV U19915 ( .A(n17160), .Z(n17218) );
  XOR U19916 ( .A(n17219), .B(n17220), .Z(n17160) );
  ANDN U19917 ( .B(n17221), .A(n17222), .Z(n17219) );
  XOR U19918 ( .A(n17220), .B(n17223), .Z(n17221) );
  XNOR U19919 ( .A(n17224), .B(n17225), .Z(n17157) );
  ANDN U19920 ( .B(n17226), .A(n17227), .Z(n17224) );
  XOR U19921 ( .A(n17225), .B(n17228), .Z(n17226) );
  IV U19922 ( .A(n17156), .Z(n17216) );
  XOR U19923 ( .A(n17154), .B(n17229), .Z(n17156) );
  XOR U19924 ( .A(n17230), .B(n17231), .Z(n17229) );
  ANDN U19925 ( .B(n17232), .A(n17233), .Z(n17230) );
  XOR U19926 ( .A(n17234), .B(n17231), .Z(n17232) );
  IV U19927 ( .A(n17158), .Z(n17154) );
  XOR U19928 ( .A(n17235), .B(n17236), .Z(n17158) );
  ANDN U19929 ( .B(n17237), .A(n17238), .Z(n17235) );
  XOR U19930 ( .A(n17239), .B(n17236), .Z(n17237) );
  XOR U19931 ( .A(n17240), .B(n17241), .Z(n17170) );
  XOR U19932 ( .A(n17188), .B(n17242), .Z(n17241) );
  IV U19933 ( .A(n17168), .Z(n17242) );
  XOR U19934 ( .A(n17243), .B(n17244), .Z(n17168) );
  ANDN U19935 ( .B(n17245), .A(n17246), .Z(n17243) );
  XOR U19936 ( .A(n17244), .B(n17247), .Z(n17245) );
  XOR U19937 ( .A(n17248), .B(n17176), .Z(n17188) );
  XOR U19938 ( .A(n17249), .B(n17250), .Z(n17176) );
  ANDN U19939 ( .B(n17251), .A(n17252), .Z(n17249) );
  XOR U19940 ( .A(n17250), .B(n17253), .Z(n17251) );
  IV U19941 ( .A(n17175), .Z(n17248) );
  XOR U19942 ( .A(n17254), .B(n17255), .Z(n17175) );
  XOR U19943 ( .A(n17256), .B(n17257), .Z(n17255) );
  ANDN U19944 ( .B(n17258), .A(n17259), .Z(n17256) );
  XOR U19945 ( .A(n17260), .B(n17257), .Z(n17258) );
  IV U19946 ( .A(n17173), .Z(n17254) );
  XOR U19947 ( .A(n17261), .B(n17262), .Z(n17173) );
  ANDN U19948 ( .B(n17263), .A(n17264), .Z(n17261) );
  XOR U19949 ( .A(n17262), .B(n17265), .Z(n17263) );
  IV U19950 ( .A(n17187), .Z(n17240) );
  XOR U19951 ( .A(n17266), .B(n17267), .Z(n17187) );
  XNOR U19952 ( .A(n17182), .B(n17268), .Z(n17267) );
  IV U19953 ( .A(n17185), .Z(n17268) );
  XOR U19954 ( .A(n17269), .B(n17270), .Z(n17185) );
  ANDN U19955 ( .B(n17271), .A(n17272), .Z(n17269) );
  XOR U19956 ( .A(n17273), .B(n17270), .Z(n17271) );
  XNOR U19957 ( .A(n17274), .B(n17275), .Z(n17182) );
  ANDN U19958 ( .B(n17276), .A(n17277), .Z(n17274) );
  XOR U19959 ( .A(n17275), .B(n17278), .Z(n17276) );
  IV U19960 ( .A(n17181), .Z(n17266) );
  XOR U19961 ( .A(n17179), .B(n17279), .Z(n17181) );
  XOR U19962 ( .A(n17280), .B(n17281), .Z(n17279) );
  ANDN U19963 ( .B(n17282), .A(n17283), .Z(n17280) );
  XOR U19964 ( .A(n17284), .B(n17281), .Z(n17282) );
  IV U19965 ( .A(n17183), .Z(n17179) );
  XOR U19966 ( .A(n17285), .B(n17286), .Z(n17183) );
  ANDN U19967 ( .B(n17287), .A(n17288), .Z(n17285) );
  XOR U19968 ( .A(n17289), .B(n17286), .Z(n17287) );
  IV U19969 ( .A(n17193), .Z(n17197) );
  XOR U19970 ( .A(n17193), .B(n17096), .Z(n17195) );
  XOR U19971 ( .A(n17290), .B(n17291), .Z(n17096) );
  AND U19972 ( .A(n112), .B(n17292), .Z(n17290) );
  XOR U19973 ( .A(n17293), .B(n17291), .Z(n17292) );
  NANDN U19974 ( .A(n17098), .B(n17100), .Z(n17193) );
  XOR U19975 ( .A(n17294), .B(n17295), .Z(n17100) );
  AND U19976 ( .A(n112), .B(n17296), .Z(n17294) );
  XOR U19977 ( .A(n17295), .B(n17297), .Z(n17296) );
  XNOR U19978 ( .A(n17298), .B(n17299), .Z(n112) );
  AND U19979 ( .A(n17300), .B(n17301), .Z(n17298) );
  XOR U19980 ( .A(n17299), .B(n17111), .Z(n17301) );
  XNOR U19981 ( .A(n17302), .B(n17303), .Z(n17111) );
  ANDN U19982 ( .B(n17304), .A(n17305), .Z(n17302) );
  XOR U19983 ( .A(n17303), .B(n17306), .Z(n17304) );
  XNOR U19984 ( .A(n17299), .B(n17113), .Z(n17300) );
  XOR U19985 ( .A(n17307), .B(n17308), .Z(n17113) );
  AND U19986 ( .A(n116), .B(n17309), .Z(n17307) );
  XOR U19987 ( .A(n17310), .B(n17308), .Z(n17309) );
  XOR U19988 ( .A(n17311), .B(n17312), .Z(n17299) );
  AND U19989 ( .A(n17313), .B(n17314), .Z(n17311) );
  XOR U19990 ( .A(n17312), .B(n17138), .Z(n17314) );
  XOR U19991 ( .A(n17305), .B(n17306), .Z(n17138) );
  XNOR U19992 ( .A(n17315), .B(n17316), .Z(n17306) );
  ANDN U19993 ( .B(n17317), .A(n17318), .Z(n17315) );
  XOR U19994 ( .A(n17319), .B(n17320), .Z(n17317) );
  XOR U19995 ( .A(n17321), .B(n17322), .Z(n17305) );
  XNOR U19996 ( .A(n17323), .B(n17324), .Z(n17322) );
  ANDN U19997 ( .B(n17325), .A(n17326), .Z(n17323) );
  XNOR U19998 ( .A(n17327), .B(n17328), .Z(n17325) );
  IV U19999 ( .A(n17303), .Z(n17321) );
  XOR U20000 ( .A(n17329), .B(n17330), .Z(n17303) );
  ANDN U20001 ( .B(n17331), .A(n17332), .Z(n17329) );
  XOR U20002 ( .A(n17330), .B(n17333), .Z(n17331) );
  XNOR U20003 ( .A(n17312), .B(n17140), .Z(n17313) );
  XOR U20004 ( .A(n17334), .B(n17335), .Z(n17140) );
  AND U20005 ( .A(n116), .B(n17336), .Z(n17334) );
  XOR U20006 ( .A(n17337), .B(n17335), .Z(n17336) );
  XNOR U20007 ( .A(n17338), .B(n17339), .Z(n17312) );
  AND U20008 ( .A(n17340), .B(n17341), .Z(n17338) );
  XNOR U20009 ( .A(n17339), .B(n17190), .Z(n17341) );
  XOR U20010 ( .A(n17332), .B(n17333), .Z(n17190) );
  XOR U20011 ( .A(n17342), .B(n17320), .Z(n17333) );
  XNOR U20012 ( .A(n17343), .B(n17344), .Z(n17320) );
  ANDN U20013 ( .B(n17345), .A(n17346), .Z(n17343) );
  XOR U20014 ( .A(n17347), .B(n17348), .Z(n17345) );
  IV U20015 ( .A(n17318), .Z(n17342) );
  XOR U20016 ( .A(n17316), .B(n17349), .Z(n17318) );
  XNOR U20017 ( .A(n17350), .B(n17351), .Z(n17349) );
  ANDN U20018 ( .B(n17352), .A(n17353), .Z(n17350) );
  XNOR U20019 ( .A(n17354), .B(n17355), .Z(n17352) );
  IV U20020 ( .A(n17319), .Z(n17316) );
  XOR U20021 ( .A(n17356), .B(n17357), .Z(n17319) );
  ANDN U20022 ( .B(n17358), .A(n17359), .Z(n17356) );
  XOR U20023 ( .A(n17357), .B(n17360), .Z(n17358) );
  XOR U20024 ( .A(n17361), .B(n17362), .Z(n17332) );
  XNOR U20025 ( .A(n17327), .B(n17363), .Z(n17362) );
  IV U20026 ( .A(n17330), .Z(n17363) );
  XOR U20027 ( .A(n17364), .B(n17365), .Z(n17330) );
  ANDN U20028 ( .B(n17366), .A(n17367), .Z(n17364) );
  XOR U20029 ( .A(n17365), .B(n17368), .Z(n17366) );
  XNOR U20030 ( .A(n17369), .B(n17370), .Z(n17327) );
  ANDN U20031 ( .B(n17371), .A(n17372), .Z(n17369) );
  XOR U20032 ( .A(n17370), .B(n17373), .Z(n17371) );
  IV U20033 ( .A(n17326), .Z(n17361) );
  XOR U20034 ( .A(n17324), .B(n17374), .Z(n17326) );
  XNOR U20035 ( .A(n17375), .B(n17376), .Z(n17374) );
  ANDN U20036 ( .B(n17377), .A(n17378), .Z(n17375) );
  XNOR U20037 ( .A(n17379), .B(n17380), .Z(n17377) );
  IV U20038 ( .A(n17328), .Z(n17324) );
  XOR U20039 ( .A(n17381), .B(n17382), .Z(n17328) );
  ANDN U20040 ( .B(n17383), .A(n17384), .Z(n17381) );
  XOR U20041 ( .A(n17385), .B(n17382), .Z(n17383) );
  XOR U20042 ( .A(n17339), .B(n17192), .Z(n17340) );
  XOR U20043 ( .A(n17386), .B(n17387), .Z(n17192) );
  AND U20044 ( .A(n116), .B(n17388), .Z(n17386) );
  XOR U20045 ( .A(n17389), .B(n17387), .Z(n17388) );
  XNOR U20046 ( .A(n17390), .B(n17391), .Z(n17339) );
  NAND U20047 ( .A(n17392), .B(n17393), .Z(n17391) );
  XOR U20048 ( .A(n17394), .B(n17291), .Z(n17393) );
  XOR U20049 ( .A(n17367), .B(n17368), .Z(n17291) );
  XOR U20050 ( .A(n17395), .B(n17360), .Z(n17368) );
  XOR U20051 ( .A(n17396), .B(n17348), .Z(n17360) );
  XOR U20052 ( .A(n17397), .B(n17398), .Z(n17348) );
  ANDN U20053 ( .B(n17399), .A(n17400), .Z(n17397) );
  XOR U20054 ( .A(n17398), .B(n17401), .Z(n17399) );
  IV U20055 ( .A(n17346), .Z(n17396) );
  XOR U20056 ( .A(n17344), .B(n17402), .Z(n17346) );
  XOR U20057 ( .A(n17403), .B(n17404), .Z(n17402) );
  ANDN U20058 ( .B(n17405), .A(n17406), .Z(n17403) );
  XOR U20059 ( .A(n17407), .B(n17404), .Z(n17405) );
  IV U20060 ( .A(n17347), .Z(n17344) );
  XOR U20061 ( .A(n17408), .B(n17409), .Z(n17347) );
  ANDN U20062 ( .B(n17410), .A(n17411), .Z(n17408) );
  XOR U20063 ( .A(n17409), .B(n17412), .Z(n17410) );
  IV U20064 ( .A(n17359), .Z(n17395) );
  XOR U20065 ( .A(n17413), .B(n17414), .Z(n17359) );
  XNOR U20066 ( .A(n17354), .B(n17415), .Z(n17414) );
  IV U20067 ( .A(n17357), .Z(n17415) );
  XOR U20068 ( .A(n17416), .B(n17417), .Z(n17357) );
  ANDN U20069 ( .B(n17418), .A(n17419), .Z(n17416) );
  XOR U20070 ( .A(n17417), .B(n17420), .Z(n17418) );
  XNOR U20071 ( .A(n17421), .B(n17422), .Z(n17354) );
  ANDN U20072 ( .B(n17423), .A(n17424), .Z(n17421) );
  XOR U20073 ( .A(n17422), .B(n17425), .Z(n17423) );
  IV U20074 ( .A(n17353), .Z(n17413) );
  XOR U20075 ( .A(n17351), .B(n17426), .Z(n17353) );
  XOR U20076 ( .A(n17427), .B(n17428), .Z(n17426) );
  ANDN U20077 ( .B(n17429), .A(n17430), .Z(n17427) );
  XOR U20078 ( .A(n17431), .B(n17428), .Z(n17429) );
  IV U20079 ( .A(n17355), .Z(n17351) );
  XOR U20080 ( .A(n17432), .B(n17433), .Z(n17355) );
  ANDN U20081 ( .B(n17434), .A(n17435), .Z(n17432) );
  XOR U20082 ( .A(n17436), .B(n17433), .Z(n17434) );
  XOR U20083 ( .A(n17437), .B(n17438), .Z(n17367) );
  XOR U20084 ( .A(n17385), .B(n17439), .Z(n17438) );
  IV U20085 ( .A(n17365), .Z(n17439) );
  XOR U20086 ( .A(n17440), .B(n17441), .Z(n17365) );
  ANDN U20087 ( .B(n17442), .A(n17443), .Z(n17440) );
  XOR U20088 ( .A(n17441), .B(n17444), .Z(n17442) );
  XOR U20089 ( .A(n17445), .B(n17373), .Z(n17385) );
  XOR U20090 ( .A(n17446), .B(n17447), .Z(n17373) );
  ANDN U20091 ( .B(n17448), .A(n17449), .Z(n17446) );
  XOR U20092 ( .A(n17447), .B(n17450), .Z(n17448) );
  IV U20093 ( .A(n17372), .Z(n17445) );
  XOR U20094 ( .A(n17451), .B(n17452), .Z(n17372) );
  XOR U20095 ( .A(n17453), .B(n17454), .Z(n17452) );
  ANDN U20096 ( .B(n17455), .A(n17456), .Z(n17453) );
  XOR U20097 ( .A(n17457), .B(n17454), .Z(n17455) );
  IV U20098 ( .A(n17370), .Z(n17451) );
  XOR U20099 ( .A(n17458), .B(n17459), .Z(n17370) );
  ANDN U20100 ( .B(n17460), .A(n17461), .Z(n17458) );
  XOR U20101 ( .A(n17459), .B(n17462), .Z(n17460) );
  IV U20102 ( .A(n17384), .Z(n17437) );
  XOR U20103 ( .A(n17463), .B(n17464), .Z(n17384) );
  XNOR U20104 ( .A(n17379), .B(n17465), .Z(n17464) );
  IV U20105 ( .A(n17382), .Z(n17465) );
  XOR U20106 ( .A(n17466), .B(n17467), .Z(n17382) );
  ANDN U20107 ( .B(n17468), .A(n17469), .Z(n17466) );
  XOR U20108 ( .A(n17470), .B(n17467), .Z(n17468) );
  XNOR U20109 ( .A(n17471), .B(n17472), .Z(n17379) );
  ANDN U20110 ( .B(n17473), .A(n17474), .Z(n17471) );
  XOR U20111 ( .A(n17472), .B(n17475), .Z(n17473) );
  IV U20112 ( .A(n17378), .Z(n17463) );
  XOR U20113 ( .A(n17376), .B(n17476), .Z(n17378) );
  XOR U20114 ( .A(n17477), .B(n17478), .Z(n17476) );
  ANDN U20115 ( .B(n17479), .A(n17480), .Z(n17477) );
  XOR U20116 ( .A(n17481), .B(n17478), .Z(n17479) );
  IV U20117 ( .A(n17380), .Z(n17376) );
  XOR U20118 ( .A(n17482), .B(n17483), .Z(n17380) );
  ANDN U20119 ( .B(n17484), .A(n17485), .Z(n17482) );
  XOR U20120 ( .A(n17486), .B(n17483), .Z(n17484) );
  IV U20121 ( .A(n17390), .Z(n17394) );
  XOR U20122 ( .A(n17390), .B(n17293), .Z(n17392) );
  XOR U20123 ( .A(n17487), .B(n17488), .Z(n17293) );
  AND U20124 ( .A(n116), .B(n17489), .Z(n17487) );
  XOR U20125 ( .A(n17490), .B(n17488), .Z(n17489) );
  NANDN U20126 ( .A(n17295), .B(n17297), .Z(n17390) );
  XOR U20127 ( .A(n17491), .B(n17492), .Z(n17297) );
  AND U20128 ( .A(n116), .B(n17493), .Z(n17491) );
  XOR U20129 ( .A(n17492), .B(n17494), .Z(n17493) );
  XNOR U20130 ( .A(n17495), .B(n17496), .Z(n116) );
  AND U20131 ( .A(n17497), .B(n17498), .Z(n17495) );
  XOR U20132 ( .A(n17496), .B(n17308), .Z(n17498) );
  XNOR U20133 ( .A(n17499), .B(n17500), .Z(n17308) );
  ANDN U20134 ( .B(n17501), .A(n17502), .Z(n17499) );
  XOR U20135 ( .A(n17500), .B(n17503), .Z(n17501) );
  XNOR U20136 ( .A(n17496), .B(n17310), .Z(n17497) );
  XOR U20137 ( .A(n17504), .B(n17505), .Z(n17310) );
  AND U20138 ( .A(n120), .B(n17506), .Z(n17504) );
  XOR U20139 ( .A(n17507), .B(n17505), .Z(n17506) );
  XOR U20140 ( .A(n17508), .B(n17509), .Z(n17496) );
  AND U20141 ( .A(n17510), .B(n17511), .Z(n17508) );
  XOR U20142 ( .A(n17509), .B(n17335), .Z(n17511) );
  XOR U20143 ( .A(n17502), .B(n17503), .Z(n17335) );
  XNOR U20144 ( .A(n17512), .B(n17513), .Z(n17503) );
  ANDN U20145 ( .B(n17514), .A(n17515), .Z(n17512) );
  XOR U20146 ( .A(n17516), .B(n17517), .Z(n17514) );
  XOR U20147 ( .A(n17518), .B(n17519), .Z(n17502) );
  XNOR U20148 ( .A(n17520), .B(n17521), .Z(n17519) );
  ANDN U20149 ( .B(n17522), .A(n17523), .Z(n17520) );
  XNOR U20150 ( .A(n17524), .B(n17525), .Z(n17522) );
  IV U20151 ( .A(n17500), .Z(n17518) );
  XOR U20152 ( .A(n17526), .B(n17527), .Z(n17500) );
  ANDN U20153 ( .B(n17528), .A(n17529), .Z(n17526) );
  XOR U20154 ( .A(n17527), .B(n17530), .Z(n17528) );
  XNOR U20155 ( .A(n17509), .B(n17337), .Z(n17510) );
  XOR U20156 ( .A(n17531), .B(n17532), .Z(n17337) );
  AND U20157 ( .A(n120), .B(n17533), .Z(n17531) );
  XOR U20158 ( .A(n17534), .B(n17532), .Z(n17533) );
  XNOR U20159 ( .A(n17535), .B(n17536), .Z(n17509) );
  AND U20160 ( .A(n17537), .B(n17538), .Z(n17535) );
  XNOR U20161 ( .A(n17536), .B(n17387), .Z(n17538) );
  XOR U20162 ( .A(n17529), .B(n17530), .Z(n17387) );
  XOR U20163 ( .A(n17539), .B(n17517), .Z(n17530) );
  XNOR U20164 ( .A(n17540), .B(n17541), .Z(n17517) );
  ANDN U20165 ( .B(n17542), .A(n17543), .Z(n17540) );
  XOR U20166 ( .A(n17544), .B(n17545), .Z(n17542) );
  IV U20167 ( .A(n17515), .Z(n17539) );
  XOR U20168 ( .A(n17513), .B(n17546), .Z(n17515) );
  XNOR U20169 ( .A(n17547), .B(n17548), .Z(n17546) );
  ANDN U20170 ( .B(n17549), .A(n17550), .Z(n17547) );
  XNOR U20171 ( .A(n17551), .B(n17552), .Z(n17549) );
  IV U20172 ( .A(n17516), .Z(n17513) );
  XOR U20173 ( .A(n17553), .B(n17554), .Z(n17516) );
  ANDN U20174 ( .B(n17555), .A(n17556), .Z(n17553) );
  XOR U20175 ( .A(n17554), .B(n17557), .Z(n17555) );
  XOR U20176 ( .A(n17558), .B(n17559), .Z(n17529) );
  XNOR U20177 ( .A(n17524), .B(n17560), .Z(n17559) );
  IV U20178 ( .A(n17527), .Z(n17560) );
  XOR U20179 ( .A(n17561), .B(n17562), .Z(n17527) );
  ANDN U20180 ( .B(n17563), .A(n17564), .Z(n17561) );
  XOR U20181 ( .A(n17562), .B(n17565), .Z(n17563) );
  XNOR U20182 ( .A(n17566), .B(n17567), .Z(n17524) );
  ANDN U20183 ( .B(n17568), .A(n17569), .Z(n17566) );
  XOR U20184 ( .A(n17567), .B(n17570), .Z(n17568) );
  IV U20185 ( .A(n17523), .Z(n17558) );
  XOR U20186 ( .A(n17521), .B(n17571), .Z(n17523) );
  XNOR U20187 ( .A(n17572), .B(n17573), .Z(n17571) );
  ANDN U20188 ( .B(n17574), .A(n17575), .Z(n17572) );
  XNOR U20189 ( .A(n17576), .B(n17577), .Z(n17574) );
  IV U20190 ( .A(n17525), .Z(n17521) );
  XOR U20191 ( .A(n17578), .B(n17579), .Z(n17525) );
  ANDN U20192 ( .B(n17580), .A(n17581), .Z(n17578) );
  XOR U20193 ( .A(n17582), .B(n17579), .Z(n17580) );
  XOR U20194 ( .A(n17536), .B(n17389), .Z(n17537) );
  XOR U20195 ( .A(n17583), .B(n17584), .Z(n17389) );
  AND U20196 ( .A(n120), .B(n17585), .Z(n17583) );
  XOR U20197 ( .A(n17586), .B(n17584), .Z(n17585) );
  XNOR U20198 ( .A(n17587), .B(n17588), .Z(n17536) );
  NAND U20199 ( .A(n17589), .B(n17590), .Z(n17588) );
  XOR U20200 ( .A(n17591), .B(n17488), .Z(n17590) );
  XOR U20201 ( .A(n17564), .B(n17565), .Z(n17488) );
  XOR U20202 ( .A(n17592), .B(n17557), .Z(n17565) );
  XOR U20203 ( .A(n17593), .B(n17545), .Z(n17557) );
  XOR U20204 ( .A(n17594), .B(n17595), .Z(n17545) );
  ANDN U20205 ( .B(n17596), .A(n17597), .Z(n17594) );
  XOR U20206 ( .A(n17595), .B(n17598), .Z(n17596) );
  IV U20207 ( .A(n17543), .Z(n17593) );
  XOR U20208 ( .A(n17541), .B(n17599), .Z(n17543) );
  XOR U20209 ( .A(n17600), .B(n17601), .Z(n17599) );
  ANDN U20210 ( .B(n17602), .A(n17603), .Z(n17600) );
  XOR U20211 ( .A(n17604), .B(n17601), .Z(n17602) );
  IV U20212 ( .A(n17544), .Z(n17541) );
  XOR U20213 ( .A(n17605), .B(n17606), .Z(n17544) );
  ANDN U20214 ( .B(n17607), .A(n17608), .Z(n17605) );
  XOR U20215 ( .A(n17606), .B(n17609), .Z(n17607) );
  IV U20216 ( .A(n17556), .Z(n17592) );
  XOR U20217 ( .A(n17610), .B(n17611), .Z(n17556) );
  XNOR U20218 ( .A(n17551), .B(n17612), .Z(n17611) );
  IV U20219 ( .A(n17554), .Z(n17612) );
  XOR U20220 ( .A(n17613), .B(n17614), .Z(n17554) );
  ANDN U20221 ( .B(n17615), .A(n17616), .Z(n17613) );
  XOR U20222 ( .A(n17614), .B(n17617), .Z(n17615) );
  XNOR U20223 ( .A(n17618), .B(n17619), .Z(n17551) );
  ANDN U20224 ( .B(n17620), .A(n17621), .Z(n17618) );
  XOR U20225 ( .A(n17619), .B(n17622), .Z(n17620) );
  IV U20226 ( .A(n17550), .Z(n17610) );
  XOR U20227 ( .A(n17548), .B(n17623), .Z(n17550) );
  XOR U20228 ( .A(n17624), .B(n17625), .Z(n17623) );
  ANDN U20229 ( .B(n17626), .A(n17627), .Z(n17624) );
  XOR U20230 ( .A(n17628), .B(n17625), .Z(n17626) );
  IV U20231 ( .A(n17552), .Z(n17548) );
  XOR U20232 ( .A(n17629), .B(n17630), .Z(n17552) );
  ANDN U20233 ( .B(n17631), .A(n17632), .Z(n17629) );
  XOR U20234 ( .A(n17633), .B(n17630), .Z(n17631) );
  XOR U20235 ( .A(n17634), .B(n17635), .Z(n17564) );
  XOR U20236 ( .A(n17582), .B(n17636), .Z(n17635) );
  IV U20237 ( .A(n17562), .Z(n17636) );
  XOR U20238 ( .A(n17637), .B(n17638), .Z(n17562) );
  ANDN U20239 ( .B(n17639), .A(n17640), .Z(n17637) );
  XOR U20240 ( .A(n17638), .B(n17641), .Z(n17639) );
  XOR U20241 ( .A(n17642), .B(n17570), .Z(n17582) );
  XOR U20242 ( .A(n17643), .B(n17644), .Z(n17570) );
  ANDN U20243 ( .B(n17645), .A(n17646), .Z(n17643) );
  XOR U20244 ( .A(n17644), .B(n17647), .Z(n17645) );
  IV U20245 ( .A(n17569), .Z(n17642) );
  XOR U20246 ( .A(n17648), .B(n17649), .Z(n17569) );
  XOR U20247 ( .A(n17650), .B(n17651), .Z(n17649) );
  ANDN U20248 ( .B(n17652), .A(n17653), .Z(n17650) );
  XOR U20249 ( .A(n17654), .B(n17651), .Z(n17652) );
  IV U20250 ( .A(n17567), .Z(n17648) );
  XOR U20251 ( .A(n17655), .B(n17656), .Z(n17567) );
  ANDN U20252 ( .B(n17657), .A(n17658), .Z(n17655) );
  XOR U20253 ( .A(n17656), .B(n17659), .Z(n17657) );
  IV U20254 ( .A(n17581), .Z(n17634) );
  XOR U20255 ( .A(n17660), .B(n17661), .Z(n17581) );
  XNOR U20256 ( .A(n17576), .B(n17662), .Z(n17661) );
  IV U20257 ( .A(n17579), .Z(n17662) );
  XOR U20258 ( .A(n17663), .B(n17664), .Z(n17579) );
  ANDN U20259 ( .B(n17665), .A(n17666), .Z(n17663) );
  XOR U20260 ( .A(n17667), .B(n17664), .Z(n17665) );
  XNOR U20261 ( .A(n17668), .B(n17669), .Z(n17576) );
  ANDN U20262 ( .B(n17670), .A(n17671), .Z(n17668) );
  XOR U20263 ( .A(n17669), .B(n17672), .Z(n17670) );
  IV U20264 ( .A(n17575), .Z(n17660) );
  XOR U20265 ( .A(n17573), .B(n17673), .Z(n17575) );
  XOR U20266 ( .A(n17674), .B(n17675), .Z(n17673) );
  ANDN U20267 ( .B(n17676), .A(n17677), .Z(n17674) );
  XOR U20268 ( .A(n17678), .B(n17675), .Z(n17676) );
  IV U20269 ( .A(n17577), .Z(n17573) );
  XOR U20270 ( .A(n17679), .B(n17680), .Z(n17577) );
  ANDN U20271 ( .B(n17681), .A(n17682), .Z(n17679) );
  XOR U20272 ( .A(n17683), .B(n17680), .Z(n17681) );
  IV U20273 ( .A(n17587), .Z(n17591) );
  XOR U20274 ( .A(n17587), .B(n17490), .Z(n17589) );
  XOR U20275 ( .A(n17684), .B(n17685), .Z(n17490) );
  AND U20276 ( .A(n120), .B(n17686), .Z(n17684) );
  XOR U20277 ( .A(n17687), .B(n17685), .Z(n17686) );
  NANDN U20278 ( .A(n17492), .B(n17494), .Z(n17587) );
  XOR U20279 ( .A(n17688), .B(n17689), .Z(n17494) );
  AND U20280 ( .A(n120), .B(n17690), .Z(n17688) );
  XOR U20281 ( .A(n17689), .B(n17691), .Z(n17690) );
  XNOR U20282 ( .A(n17692), .B(n17693), .Z(n120) );
  AND U20283 ( .A(n17694), .B(n17695), .Z(n17692) );
  XOR U20284 ( .A(n17693), .B(n17505), .Z(n17695) );
  XNOR U20285 ( .A(n17696), .B(n17697), .Z(n17505) );
  ANDN U20286 ( .B(n17698), .A(n17699), .Z(n17696) );
  XOR U20287 ( .A(n17697), .B(n17700), .Z(n17698) );
  XNOR U20288 ( .A(n17693), .B(n17507), .Z(n17694) );
  XOR U20289 ( .A(n17701), .B(n17702), .Z(n17507) );
  AND U20290 ( .A(n124), .B(n17703), .Z(n17701) );
  XOR U20291 ( .A(n17704), .B(n17702), .Z(n17703) );
  XOR U20292 ( .A(n17705), .B(n17706), .Z(n17693) );
  AND U20293 ( .A(n17707), .B(n17708), .Z(n17705) );
  XOR U20294 ( .A(n17706), .B(n17532), .Z(n17708) );
  XOR U20295 ( .A(n17699), .B(n17700), .Z(n17532) );
  XNOR U20296 ( .A(n17709), .B(n17710), .Z(n17700) );
  ANDN U20297 ( .B(n17711), .A(n17712), .Z(n17709) );
  XOR U20298 ( .A(n17713), .B(n17714), .Z(n17711) );
  XOR U20299 ( .A(n17715), .B(n17716), .Z(n17699) );
  XNOR U20300 ( .A(n17717), .B(n17718), .Z(n17716) );
  ANDN U20301 ( .B(n17719), .A(n17720), .Z(n17717) );
  XNOR U20302 ( .A(n17721), .B(n17722), .Z(n17719) );
  IV U20303 ( .A(n17697), .Z(n17715) );
  XOR U20304 ( .A(n17723), .B(n17724), .Z(n17697) );
  ANDN U20305 ( .B(n17725), .A(n17726), .Z(n17723) );
  XOR U20306 ( .A(n17724), .B(n17727), .Z(n17725) );
  XNOR U20307 ( .A(n17706), .B(n17534), .Z(n17707) );
  XOR U20308 ( .A(n17728), .B(n17729), .Z(n17534) );
  AND U20309 ( .A(n124), .B(n17730), .Z(n17728) );
  XOR U20310 ( .A(n17731), .B(n17729), .Z(n17730) );
  XNOR U20311 ( .A(n17732), .B(n17733), .Z(n17706) );
  AND U20312 ( .A(n17734), .B(n17735), .Z(n17732) );
  XNOR U20313 ( .A(n17733), .B(n17584), .Z(n17735) );
  XOR U20314 ( .A(n17726), .B(n17727), .Z(n17584) );
  XOR U20315 ( .A(n17736), .B(n17714), .Z(n17727) );
  XNOR U20316 ( .A(n17737), .B(n17738), .Z(n17714) );
  ANDN U20317 ( .B(n17739), .A(n17740), .Z(n17737) );
  XOR U20318 ( .A(n17741), .B(n17742), .Z(n17739) );
  IV U20319 ( .A(n17712), .Z(n17736) );
  XOR U20320 ( .A(n17710), .B(n17743), .Z(n17712) );
  XNOR U20321 ( .A(n17744), .B(n17745), .Z(n17743) );
  ANDN U20322 ( .B(n17746), .A(n17747), .Z(n17744) );
  XNOR U20323 ( .A(n17748), .B(n17749), .Z(n17746) );
  IV U20324 ( .A(n17713), .Z(n17710) );
  XOR U20325 ( .A(n17750), .B(n17751), .Z(n17713) );
  ANDN U20326 ( .B(n17752), .A(n17753), .Z(n17750) );
  XOR U20327 ( .A(n17751), .B(n17754), .Z(n17752) );
  XOR U20328 ( .A(n17755), .B(n17756), .Z(n17726) );
  XNOR U20329 ( .A(n17721), .B(n17757), .Z(n17756) );
  IV U20330 ( .A(n17724), .Z(n17757) );
  XOR U20331 ( .A(n17758), .B(n17759), .Z(n17724) );
  ANDN U20332 ( .B(n17760), .A(n17761), .Z(n17758) );
  XOR U20333 ( .A(n17759), .B(n17762), .Z(n17760) );
  XNOR U20334 ( .A(n17763), .B(n17764), .Z(n17721) );
  ANDN U20335 ( .B(n17765), .A(n17766), .Z(n17763) );
  XOR U20336 ( .A(n17764), .B(n17767), .Z(n17765) );
  IV U20337 ( .A(n17720), .Z(n17755) );
  XOR U20338 ( .A(n17718), .B(n17768), .Z(n17720) );
  XNOR U20339 ( .A(n17769), .B(n17770), .Z(n17768) );
  ANDN U20340 ( .B(n17771), .A(n17772), .Z(n17769) );
  XNOR U20341 ( .A(n17773), .B(n17774), .Z(n17771) );
  IV U20342 ( .A(n17722), .Z(n17718) );
  XOR U20343 ( .A(n17775), .B(n17776), .Z(n17722) );
  ANDN U20344 ( .B(n17777), .A(n17778), .Z(n17775) );
  XOR U20345 ( .A(n17779), .B(n17776), .Z(n17777) );
  XOR U20346 ( .A(n17733), .B(n17586), .Z(n17734) );
  XOR U20347 ( .A(n17780), .B(n17781), .Z(n17586) );
  AND U20348 ( .A(n124), .B(n17782), .Z(n17780) );
  XOR U20349 ( .A(n17783), .B(n17781), .Z(n17782) );
  XNOR U20350 ( .A(n17784), .B(n17785), .Z(n17733) );
  NAND U20351 ( .A(n17786), .B(n17787), .Z(n17785) );
  XOR U20352 ( .A(n17788), .B(n17685), .Z(n17787) );
  XOR U20353 ( .A(n17761), .B(n17762), .Z(n17685) );
  XOR U20354 ( .A(n17789), .B(n17754), .Z(n17762) );
  XOR U20355 ( .A(n17790), .B(n17742), .Z(n17754) );
  XOR U20356 ( .A(n17791), .B(n17792), .Z(n17742) );
  ANDN U20357 ( .B(n17793), .A(n17794), .Z(n17791) );
  XOR U20358 ( .A(n17792), .B(n17795), .Z(n17793) );
  IV U20359 ( .A(n17740), .Z(n17790) );
  XOR U20360 ( .A(n17738), .B(n17796), .Z(n17740) );
  XOR U20361 ( .A(n17797), .B(n17798), .Z(n17796) );
  ANDN U20362 ( .B(n17799), .A(n17800), .Z(n17797) );
  XOR U20363 ( .A(n17801), .B(n17798), .Z(n17799) );
  IV U20364 ( .A(n17741), .Z(n17738) );
  XOR U20365 ( .A(n17802), .B(n17803), .Z(n17741) );
  ANDN U20366 ( .B(n17804), .A(n17805), .Z(n17802) );
  XOR U20367 ( .A(n17803), .B(n17806), .Z(n17804) );
  IV U20368 ( .A(n17753), .Z(n17789) );
  XOR U20369 ( .A(n17807), .B(n17808), .Z(n17753) );
  XNOR U20370 ( .A(n17748), .B(n17809), .Z(n17808) );
  IV U20371 ( .A(n17751), .Z(n17809) );
  XOR U20372 ( .A(n17810), .B(n17811), .Z(n17751) );
  ANDN U20373 ( .B(n17812), .A(n17813), .Z(n17810) );
  XOR U20374 ( .A(n17811), .B(n17814), .Z(n17812) );
  XNOR U20375 ( .A(n17815), .B(n17816), .Z(n17748) );
  ANDN U20376 ( .B(n17817), .A(n17818), .Z(n17815) );
  XOR U20377 ( .A(n17816), .B(n17819), .Z(n17817) );
  IV U20378 ( .A(n17747), .Z(n17807) );
  XOR U20379 ( .A(n17745), .B(n17820), .Z(n17747) );
  XOR U20380 ( .A(n17821), .B(n17822), .Z(n17820) );
  ANDN U20381 ( .B(n17823), .A(n17824), .Z(n17821) );
  XOR U20382 ( .A(n17825), .B(n17822), .Z(n17823) );
  IV U20383 ( .A(n17749), .Z(n17745) );
  XOR U20384 ( .A(n17826), .B(n17827), .Z(n17749) );
  ANDN U20385 ( .B(n17828), .A(n17829), .Z(n17826) );
  XOR U20386 ( .A(n17830), .B(n17827), .Z(n17828) );
  XOR U20387 ( .A(n17831), .B(n17832), .Z(n17761) );
  XOR U20388 ( .A(n17779), .B(n17833), .Z(n17832) );
  IV U20389 ( .A(n17759), .Z(n17833) );
  XOR U20390 ( .A(n17834), .B(n17835), .Z(n17759) );
  ANDN U20391 ( .B(n17836), .A(n17837), .Z(n17834) );
  XOR U20392 ( .A(n17835), .B(n17838), .Z(n17836) );
  XOR U20393 ( .A(n17839), .B(n17767), .Z(n17779) );
  XOR U20394 ( .A(n17840), .B(n17841), .Z(n17767) );
  ANDN U20395 ( .B(n17842), .A(n17843), .Z(n17840) );
  XOR U20396 ( .A(n17841), .B(n17844), .Z(n17842) );
  IV U20397 ( .A(n17766), .Z(n17839) );
  XOR U20398 ( .A(n17845), .B(n17846), .Z(n17766) );
  XOR U20399 ( .A(n17847), .B(n17848), .Z(n17846) );
  ANDN U20400 ( .B(n17849), .A(n17850), .Z(n17847) );
  XOR U20401 ( .A(n17851), .B(n17848), .Z(n17849) );
  IV U20402 ( .A(n17764), .Z(n17845) );
  XOR U20403 ( .A(n17852), .B(n17853), .Z(n17764) );
  ANDN U20404 ( .B(n17854), .A(n17855), .Z(n17852) );
  XOR U20405 ( .A(n17853), .B(n17856), .Z(n17854) );
  IV U20406 ( .A(n17778), .Z(n17831) );
  XOR U20407 ( .A(n17857), .B(n17858), .Z(n17778) );
  XNOR U20408 ( .A(n17773), .B(n17859), .Z(n17858) );
  IV U20409 ( .A(n17776), .Z(n17859) );
  XOR U20410 ( .A(n17860), .B(n17861), .Z(n17776) );
  ANDN U20411 ( .B(n17862), .A(n17863), .Z(n17860) );
  XOR U20412 ( .A(n17864), .B(n17861), .Z(n17862) );
  XNOR U20413 ( .A(n17865), .B(n17866), .Z(n17773) );
  ANDN U20414 ( .B(n17867), .A(n17868), .Z(n17865) );
  XOR U20415 ( .A(n17866), .B(n17869), .Z(n17867) );
  IV U20416 ( .A(n17772), .Z(n17857) );
  XOR U20417 ( .A(n17770), .B(n17870), .Z(n17772) );
  XOR U20418 ( .A(n17871), .B(n17872), .Z(n17870) );
  ANDN U20419 ( .B(n17873), .A(n17874), .Z(n17871) );
  XOR U20420 ( .A(n17875), .B(n17872), .Z(n17873) );
  IV U20421 ( .A(n17774), .Z(n17770) );
  XOR U20422 ( .A(n17876), .B(n17877), .Z(n17774) );
  ANDN U20423 ( .B(n17878), .A(n17879), .Z(n17876) );
  XOR U20424 ( .A(n17880), .B(n17877), .Z(n17878) );
  IV U20425 ( .A(n17784), .Z(n17788) );
  XOR U20426 ( .A(n17784), .B(n17687), .Z(n17786) );
  XOR U20427 ( .A(n17881), .B(n17882), .Z(n17687) );
  AND U20428 ( .A(n124), .B(n17883), .Z(n17881) );
  XOR U20429 ( .A(n17884), .B(n17882), .Z(n17883) );
  NANDN U20430 ( .A(n17689), .B(n17691), .Z(n17784) );
  XOR U20431 ( .A(n17885), .B(n17886), .Z(n17691) );
  AND U20432 ( .A(n124), .B(n17887), .Z(n17885) );
  XOR U20433 ( .A(n17886), .B(n17888), .Z(n17887) );
  XNOR U20434 ( .A(n17889), .B(n17890), .Z(n124) );
  AND U20435 ( .A(n17891), .B(n17892), .Z(n17889) );
  XOR U20436 ( .A(n17890), .B(n17702), .Z(n17892) );
  XNOR U20437 ( .A(n17893), .B(n17894), .Z(n17702) );
  ANDN U20438 ( .B(n17895), .A(n17896), .Z(n17893) );
  XOR U20439 ( .A(n17894), .B(n17897), .Z(n17895) );
  XNOR U20440 ( .A(n17890), .B(n17704), .Z(n17891) );
  XOR U20441 ( .A(n17898), .B(n17899), .Z(n17704) );
  AND U20442 ( .A(n128), .B(n17900), .Z(n17898) );
  XOR U20443 ( .A(n17901), .B(n17899), .Z(n17900) );
  XOR U20444 ( .A(n17902), .B(n17903), .Z(n17890) );
  AND U20445 ( .A(n17904), .B(n17905), .Z(n17902) );
  XOR U20446 ( .A(n17903), .B(n17729), .Z(n17905) );
  XOR U20447 ( .A(n17896), .B(n17897), .Z(n17729) );
  XNOR U20448 ( .A(n17906), .B(n17907), .Z(n17897) );
  ANDN U20449 ( .B(n17908), .A(n17909), .Z(n17906) );
  XOR U20450 ( .A(n17910), .B(n17911), .Z(n17908) );
  XOR U20451 ( .A(n17912), .B(n17913), .Z(n17896) );
  XNOR U20452 ( .A(n17914), .B(n17915), .Z(n17913) );
  ANDN U20453 ( .B(n17916), .A(n17917), .Z(n17914) );
  XNOR U20454 ( .A(n17918), .B(n17919), .Z(n17916) );
  IV U20455 ( .A(n17894), .Z(n17912) );
  XOR U20456 ( .A(n17920), .B(n17921), .Z(n17894) );
  ANDN U20457 ( .B(n17922), .A(n17923), .Z(n17920) );
  XOR U20458 ( .A(n17921), .B(n17924), .Z(n17922) );
  XNOR U20459 ( .A(n17903), .B(n17731), .Z(n17904) );
  XOR U20460 ( .A(n17925), .B(n17926), .Z(n17731) );
  AND U20461 ( .A(n128), .B(n17927), .Z(n17925) );
  XOR U20462 ( .A(n17928), .B(n17926), .Z(n17927) );
  XNOR U20463 ( .A(n17929), .B(n17930), .Z(n17903) );
  AND U20464 ( .A(n17931), .B(n17932), .Z(n17929) );
  XNOR U20465 ( .A(n17930), .B(n17781), .Z(n17932) );
  XOR U20466 ( .A(n17923), .B(n17924), .Z(n17781) );
  XOR U20467 ( .A(n17933), .B(n17911), .Z(n17924) );
  XNOR U20468 ( .A(n17934), .B(n17935), .Z(n17911) );
  ANDN U20469 ( .B(n17936), .A(n17937), .Z(n17934) );
  XOR U20470 ( .A(n17938), .B(n17939), .Z(n17936) );
  IV U20471 ( .A(n17909), .Z(n17933) );
  XOR U20472 ( .A(n17907), .B(n17940), .Z(n17909) );
  XNOR U20473 ( .A(n17941), .B(n17942), .Z(n17940) );
  ANDN U20474 ( .B(n17943), .A(n17944), .Z(n17941) );
  XNOR U20475 ( .A(n17945), .B(n17946), .Z(n17943) );
  IV U20476 ( .A(n17910), .Z(n17907) );
  XOR U20477 ( .A(n17947), .B(n17948), .Z(n17910) );
  ANDN U20478 ( .B(n17949), .A(n17950), .Z(n17947) );
  XOR U20479 ( .A(n17948), .B(n17951), .Z(n17949) );
  XOR U20480 ( .A(n17952), .B(n17953), .Z(n17923) );
  XNOR U20481 ( .A(n17918), .B(n17954), .Z(n17953) );
  IV U20482 ( .A(n17921), .Z(n17954) );
  XOR U20483 ( .A(n17955), .B(n17956), .Z(n17921) );
  ANDN U20484 ( .B(n17957), .A(n17958), .Z(n17955) );
  XOR U20485 ( .A(n17956), .B(n17959), .Z(n17957) );
  XNOR U20486 ( .A(n17960), .B(n17961), .Z(n17918) );
  ANDN U20487 ( .B(n17962), .A(n17963), .Z(n17960) );
  XOR U20488 ( .A(n17961), .B(n17964), .Z(n17962) );
  IV U20489 ( .A(n17917), .Z(n17952) );
  XOR U20490 ( .A(n17915), .B(n17965), .Z(n17917) );
  XNOR U20491 ( .A(n17966), .B(n17967), .Z(n17965) );
  ANDN U20492 ( .B(n17968), .A(n17969), .Z(n17966) );
  XNOR U20493 ( .A(n17970), .B(n17971), .Z(n17968) );
  IV U20494 ( .A(n17919), .Z(n17915) );
  XOR U20495 ( .A(n17972), .B(n17973), .Z(n17919) );
  ANDN U20496 ( .B(n17974), .A(n17975), .Z(n17972) );
  XOR U20497 ( .A(n17976), .B(n17973), .Z(n17974) );
  XOR U20498 ( .A(n17930), .B(n17783), .Z(n17931) );
  XOR U20499 ( .A(n17977), .B(n17978), .Z(n17783) );
  AND U20500 ( .A(n128), .B(n17979), .Z(n17977) );
  XOR U20501 ( .A(n17980), .B(n17978), .Z(n17979) );
  XNOR U20502 ( .A(n17981), .B(n17982), .Z(n17930) );
  NAND U20503 ( .A(n17983), .B(n17984), .Z(n17982) );
  XOR U20504 ( .A(n17985), .B(n17882), .Z(n17984) );
  XOR U20505 ( .A(n17958), .B(n17959), .Z(n17882) );
  XOR U20506 ( .A(n17986), .B(n17951), .Z(n17959) );
  XOR U20507 ( .A(n17987), .B(n17939), .Z(n17951) );
  XOR U20508 ( .A(n17988), .B(n17989), .Z(n17939) );
  ANDN U20509 ( .B(n17990), .A(n17991), .Z(n17988) );
  XOR U20510 ( .A(n17989), .B(n17992), .Z(n17990) );
  IV U20511 ( .A(n17937), .Z(n17987) );
  XOR U20512 ( .A(n17935), .B(n17993), .Z(n17937) );
  XOR U20513 ( .A(n17994), .B(n17995), .Z(n17993) );
  ANDN U20514 ( .B(n17996), .A(n17997), .Z(n17994) );
  XOR U20515 ( .A(n17998), .B(n17995), .Z(n17996) );
  IV U20516 ( .A(n17938), .Z(n17935) );
  XOR U20517 ( .A(n17999), .B(n18000), .Z(n17938) );
  ANDN U20518 ( .B(n18001), .A(n18002), .Z(n17999) );
  XOR U20519 ( .A(n18000), .B(n18003), .Z(n18001) );
  IV U20520 ( .A(n17950), .Z(n17986) );
  XOR U20521 ( .A(n18004), .B(n18005), .Z(n17950) );
  XNOR U20522 ( .A(n17945), .B(n18006), .Z(n18005) );
  IV U20523 ( .A(n17948), .Z(n18006) );
  XOR U20524 ( .A(n18007), .B(n18008), .Z(n17948) );
  ANDN U20525 ( .B(n18009), .A(n18010), .Z(n18007) );
  XOR U20526 ( .A(n18008), .B(n18011), .Z(n18009) );
  XNOR U20527 ( .A(n18012), .B(n18013), .Z(n17945) );
  ANDN U20528 ( .B(n18014), .A(n18015), .Z(n18012) );
  XOR U20529 ( .A(n18013), .B(n18016), .Z(n18014) );
  IV U20530 ( .A(n17944), .Z(n18004) );
  XOR U20531 ( .A(n17942), .B(n18017), .Z(n17944) );
  XOR U20532 ( .A(n18018), .B(n18019), .Z(n18017) );
  ANDN U20533 ( .B(n18020), .A(n18021), .Z(n18018) );
  XOR U20534 ( .A(n18022), .B(n18019), .Z(n18020) );
  IV U20535 ( .A(n17946), .Z(n17942) );
  XOR U20536 ( .A(n18023), .B(n18024), .Z(n17946) );
  ANDN U20537 ( .B(n18025), .A(n18026), .Z(n18023) );
  XOR U20538 ( .A(n18027), .B(n18024), .Z(n18025) );
  XOR U20539 ( .A(n18028), .B(n18029), .Z(n17958) );
  XOR U20540 ( .A(n17976), .B(n18030), .Z(n18029) );
  IV U20541 ( .A(n17956), .Z(n18030) );
  XOR U20542 ( .A(n18031), .B(n18032), .Z(n17956) );
  ANDN U20543 ( .B(n18033), .A(n18034), .Z(n18031) );
  XOR U20544 ( .A(n18032), .B(n18035), .Z(n18033) );
  XOR U20545 ( .A(n18036), .B(n17964), .Z(n17976) );
  XOR U20546 ( .A(n18037), .B(n18038), .Z(n17964) );
  ANDN U20547 ( .B(n18039), .A(n18040), .Z(n18037) );
  XOR U20548 ( .A(n18038), .B(n18041), .Z(n18039) );
  IV U20549 ( .A(n17963), .Z(n18036) );
  XOR U20550 ( .A(n18042), .B(n18043), .Z(n17963) );
  XOR U20551 ( .A(n18044), .B(n18045), .Z(n18043) );
  ANDN U20552 ( .B(n18046), .A(n18047), .Z(n18044) );
  XOR U20553 ( .A(n18048), .B(n18045), .Z(n18046) );
  IV U20554 ( .A(n17961), .Z(n18042) );
  XOR U20555 ( .A(n18049), .B(n18050), .Z(n17961) );
  ANDN U20556 ( .B(n18051), .A(n18052), .Z(n18049) );
  XOR U20557 ( .A(n18050), .B(n18053), .Z(n18051) );
  IV U20558 ( .A(n17975), .Z(n18028) );
  XOR U20559 ( .A(n18054), .B(n18055), .Z(n17975) );
  XNOR U20560 ( .A(n17970), .B(n18056), .Z(n18055) );
  IV U20561 ( .A(n17973), .Z(n18056) );
  XOR U20562 ( .A(n18057), .B(n18058), .Z(n17973) );
  ANDN U20563 ( .B(n18059), .A(n18060), .Z(n18057) );
  XOR U20564 ( .A(n18061), .B(n18058), .Z(n18059) );
  XNOR U20565 ( .A(n18062), .B(n18063), .Z(n17970) );
  ANDN U20566 ( .B(n18064), .A(n18065), .Z(n18062) );
  XOR U20567 ( .A(n18063), .B(n18066), .Z(n18064) );
  IV U20568 ( .A(n17969), .Z(n18054) );
  XOR U20569 ( .A(n17967), .B(n18067), .Z(n17969) );
  XOR U20570 ( .A(n18068), .B(n18069), .Z(n18067) );
  ANDN U20571 ( .B(n18070), .A(n18071), .Z(n18068) );
  XOR U20572 ( .A(n18072), .B(n18069), .Z(n18070) );
  IV U20573 ( .A(n17971), .Z(n17967) );
  XOR U20574 ( .A(n18073), .B(n18074), .Z(n17971) );
  ANDN U20575 ( .B(n18075), .A(n18076), .Z(n18073) );
  XOR U20576 ( .A(n18077), .B(n18074), .Z(n18075) );
  IV U20577 ( .A(n17981), .Z(n17985) );
  XOR U20578 ( .A(n17981), .B(n17884), .Z(n17983) );
  XOR U20579 ( .A(n18078), .B(n18079), .Z(n17884) );
  AND U20580 ( .A(n128), .B(n18080), .Z(n18078) );
  XOR U20581 ( .A(n18081), .B(n18079), .Z(n18080) );
  NANDN U20582 ( .A(n17886), .B(n17888), .Z(n17981) );
  XOR U20583 ( .A(n18082), .B(n18083), .Z(n17888) );
  AND U20584 ( .A(n128), .B(n18084), .Z(n18082) );
  XOR U20585 ( .A(n18083), .B(n18085), .Z(n18084) );
  XNOR U20586 ( .A(n18086), .B(n18087), .Z(n128) );
  AND U20587 ( .A(n18088), .B(n18089), .Z(n18086) );
  XOR U20588 ( .A(n18087), .B(n17899), .Z(n18089) );
  XNOR U20589 ( .A(n18090), .B(n18091), .Z(n17899) );
  ANDN U20590 ( .B(n18092), .A(n18093), .Z(n18090) );
  XOR U20591 ( .A(n18091), .B(n18094), .Z(n18092) );
  XNOR U20592 ( .A(n18087), .B(n17901), .Z(n18088) );
  XOR U20593 ( .A(n18095), .B(n18096), .Z(n17901) );
  AND U20594 ( .A(n132), .B(n18097), .Z(n18095) );
  XOR U20595 ( .A(n18098), .B(n18096), .Z(n18097) );
  XOR U20596 ( .A(n18099), .B(n18100), .Z(n18087) );
  AND U20597 ( .A(n18101), .B(n18102), .Z(n18099) );
  XOR U20598 ( .A(n18100), .B(n17926), .Z(n18102) );
  XOR U20599 ( .A(n18093), .B(n18094), .Z(n17926) );
  XNOR U20600 ( .A(n18103), .B(n18104), .Z(n18094) );
  ANDN U20601 ( .B(n18105), .A(n18106), .Z(n18103) );
  XOR U20602 ( .A(n18107), .B(n18108), .Z(n18105) );
  XOR U20603 ( .A(n18109), .B(n18110), .Z(n18093) );
  XNOR U20604 ( .A(n18111), .B(n18112), .Z(n18110) );
  ANDN U20605 ( .B(n18113), .A(n18114), .Z(n18111) );
  XNOR U20606 ( .A(n18115), .B(n18116), .Z(n18113) );
  IV U20607 ( .A(n18091), .Z(n18109) );
  XOR U20608 ( .A(n18117), .B(n18118), .Z(n18091) );
  ANDN U20609 ( .B(n18119), .A(n18120), .Z(n18117) );
  XOR U20610 ( .A(n18118), .B(n18121), .Z(n18119) );
  XNOR U20611 ( .A(n18100), .B(n17928), .Z(n18101) );
  XOR U20612 ( .A(n18122), .B(n18123), .Z(n17928) );
  AND U20613 ( .A(n132), .B(n18124), .Z(n18122) );
  XOR U20614 ( .A(n18125), .B(n18123), .Z(n18124) );
  XNOR U20615 ( .A(n18126), .B(n18127), .Z(n18100) );
  AND U20616 ( .A(n18128), .B(n18129), .Z(n18126) );
  XNOR U20617 ( .A(n18127), .B(n17978), .Z(n18129) );
  XOR U20618 ( .A(n18120), .B(n18121), .Z(n17978) );
  XOR U20619 ( .A(n18130), .B(n18108), .Z(n18121) );
  XNOR U20620 ( .A(n18131), .B(n18132), .Z(n18108) );
  ANDN U20621 ( .B(n18133), .A(n18134), .Z(n18131) );
  XOR U20622 ( .A(n18135), .B(n18136), .Z(n18133) );
  IV U20623 ( .A(n18106), .Z(n18130) );
  XOR U20624 ( .A(n18104), .B(n18137), .Z(n18106) );
  XNOR U20625 ( .A(n18138), .B(n18139), .Z(n18137) );
  ANDN U20626 ( .B(n18140), .A(n18141), .Z(n18138) );
  XNOR U20627 ( .A(n18142), .B(n18143), .Z(n18140) );
  IV U20628 ( .A(n18107), .Z(n18104) );
  XOR U20629 ( .A(n18144), .B(n18145), .Z(n18107) );
  ANDN U20630 ( .B(n18146), .A(n18147), .Z(n18144) );
  XOR U20631 ( .A(n18145), .B(n18148), .Z(n18146) );
  XOR U20632 ( .A(n18149), .B(n18150), .Z(n18120) );
  XNOR U20633 ( .A(n18115), .B(n18151), .Z(n18150) );
  IV U20634 ( .A(n18118), .Z(n18151) );
  XOR U20635 ( .A(n18152), .B(n18153), .Z(n18118) );
  ANDN U20636 ( .B(n18154), .A(n18155), .Z(n18152) );
  XOR U20637 ( .A(n18153), .B(n18156), .Z(n18154) );
  XNOR U20638 ( .A(n18157), .B(n18158), .Z(n18115) );
  ANDN U20639 ( .B(n18159), .A(n18160), .Z(n18157) );
  XOR U20640 ( .A(n18158), .B(n18161), .Z(n18159) );
  IV U20641 ( .A(n18114), .Z(n18149) );
  XOR U20642 ( .A(n18112), .B(n18162), .Z(n18114) );
  XNOR U20643 ( .A(n18163), .B(n18164), .Z(n18162) );
  ANDN U20644 ( .B(n18165), .A(n18166), .Z(n18163) );
  XNOR U20645 ( .A(n18167), .B(n18168), .Z(n18165) );
  IV U20646 ( .A(n18116), .Z(n18112) );
  XOR U20647 ( .A(n18169), .B(n18170), .Z(n18116) );
  ANDN U20648 ( .B(n18171), .A(n18172), .Z(n18169) );
  XOR U20649 ( .A(n18173), .B(n18170), .Z(n18171) );
  XOR U20650 ( .A(n18127), .B(n17980), .Z(n18128) );
  XOR U20651 ( .A(n18174), .B(n18175), .Z(n17980) );
  AND U20652 ( .A(n132), .B(n18176), .Z(n18174) );
  XOR U20653 ( .A(n18177), .B(n18175), .Z(n18176) );
  XNOR U20654 ( .A(n18178), .B(n18179), .Z(n18127) );
  NAND U20655 ( .A(n18180), .B(n18181), .Z(n18179) );
  XOR U20656 ( .A(n18182), .B(n18079), .Z(n18181) );
  XOR U20657 ( .A(n18155), .B(n18156), .Z(n18079) );
  XOR U20658 ( .A(n18183), .B(n18148), .Z(n18156) );
  XOR U20659 ( .A(n18184), .B(n18136), .Z(n18148) );
  XOR U20660 ( .A(n18185), .B(n18186), .Z(n18136) );
  ANDN U20661 ( .B(n18187), .A(n18188), .Z(n18185) );
  XOR U20662 ( .A(n18186), .B(n18189), .Z(n18187) );
  IV U20663 ( .A(n18134), .Z(n18184) );
  XOR U20664 ( .A(n18132), .B(n18190), .Z(n18134) );
  XOR U20665 ( .A(n18191), .B(n18192), .Z(n18190) );
  ANDN U20666 ( .B(n18193), .A(n18194), .Z(n18191) );
  XOR U20667 ( .A(n18195), .B(n18192), .Z(n18193) );
  IV U20668 ( .A(n18135), .Z(n18132) );
  XOR U20669 ( .A(n18196), .B(n18197), .Z(n18135) );
  ANDN U20670 ( .B(n18198), .A(n18199), .Z(n18196) );
  XOR U20671 ( .A(n18197), .B(n18200), .Z(n18198) );
  IV U20672 ( .A(n18147), .Z(n18183) );
  XOR U20673 ( .A(n18201), .B(n18202), .Z(n18147) );
  XNOR U20674 ( .A(n18142), .B(n18203), .Z(n18202) );
  IV U20675 ( .A(n18145), .Z(n18203) );
  XOR U20676 ( .A(n18204), .B(n18205), .Z(n18145) );
  ANDN U20677 ( .B(n18206), .A(n18207), .Z(n18204) );
  XOR U20678 ( .A(n18205), .B(n18208), .Z(n18206) );
  XNOR U20679 ( .A(n18209), .B(n18210), .Z(n18142) );
  ANDN U20680 ( .B(n18211), .A(n18212), .Z(n18209) );
  XOR U20681 ( .A(n18210), .B(n18213), .Z(n18211) );
  IV U20682 ( .A(n18141), .Z(n18201) );
  XOR U20683 ( .A(n18139), .B(n18214), .Z(n18141) );
  XOR U20684 ( .A(n18215), .B(n18216), .Z(n18214) );
  ANDN U20685 ( .B(n18217), .A(n18218), .Z(n18215) );
  XOR U20686 ( .A(n18219), .B(n18216), .Z(n18217) );
  IV U20687 ( .A(n18143), .Z(n18139) );
  XOR U20688 ( .A(n18220), .B(n18221), .Z(n18143) );
  ANDN U20689 ( .B(n18222), .A(n18223), .Z(n18220) );
  XOR U20690 ( .A(n18224), .B(n18221), .Z(n18222) );
  XOR U20691 ( .A(n18225), .B(n18226), .Z(n18155) );
  XOR U20692 ( .A(n18173), .B(n18227), .Z(n18226) );
  IV U20693 ( .A(n18153), .Z(n18227) );
  XOR U20694 ( .A(n18228), .B(n18229), .Z(n18153) );
  ANDN U20695 ( .B(n18230), .A(n18231), .Z(n18228) );
  XOR U20696 ( .A(n18229), .B(n18232), .Z(n18230) );
  XOR U20697 ( .A(n18233), .B(n18161), .Z(n18173) );
  XOR U20698 ( .A(n18234), .B(n18235), .Z(n18161) );
  ANDN U20699 ( .B(n18236), .A(n18237), .Z(n18234) );
  XOR U20700 ( .A(n18235), .B(n18238), .Z(n18236) );
  IV U20701 ( .A(n18160), .Z(n18233) );
  XOR U20702 ( .A(n18239), .B(n18240), .Z(n18160) );
  XOR U20703 ( .A(n18241), .B(n18242), .Z(n18240) );
  ANDN U20704 ( .B(n18243), .A(n18244), .Z(n18241) );
  XOR U20705 ( .A(n18245), .B(n18242), .Z(n18243) );
  IV U20706 ( .A(n18158), .Z(n18239) );
  XOR U20707 ( .A(n18246), .B(n18247), .Z(n18158) );
  ANDN U20708 ( .B(n18248), .A(n18249), .Z(n18246) );
  XOR U20709 ( .A(n18247), .B(n18250), .Z(n18248) );
  IV U20710 ( .A(n18172), .Z(n18225) );
  XOR U20711 ( .A(n18251), .B(n18252), .Z(n18172) );
  XNOR U20712 ( .A(n18167), .B(n18253), .Z(n18252) );
  IV U20713 ( .A(n18170), .Z(n18253) );
  XOR U20714 ( .A(n18254), .B(n18255), .Z(n18170) );
  ANDN U20715 ( .B(n18256), .A(n18257), .Z(n18254) );
  XOR U20716 ( .A(n18258), .B(n18255), .Z(n18256) );
  XNOR U20717 ( .A(n18259), .B(n18260), .Z(n18167) );
  ANDN U20718 ( .B(n18261), .A(n18262), .Z(n18259) );
  XOR U20719 ( .A(n18260), .B(n18263), .Z(n18261) );
  IV U20720 ( .A(n18166), .Z(n18251) );
  XOR U20721 ( .A(n18164), .B(n18264), .Z(n18166) );
  XOR U20722 ( .A(n18265), .B(n18266), .Z(n18264) );
  ANDN U20723 ( .B(n18267), .A(n18268), .Z(n18265) );
  XOR U20724 ( .A(n18269), .B(n18266), .Z(n18267) );
  IV U20725 ( .A(n18168), .Z(n18164) );
  XOR U20726 ( .A(n18270), .B(n18271), .Z(n18168) );
  ANDN U20727 ( .B(n18272), .A(n18273), .Z(n18270) );
  XOR U20728 ( .A(n18274), .B(n18271), .Z(n18272) );
  IV U20729 ( .A(n18178), .Z(n18182) );
  XOR U20730 ( .A(n18178), .B(n18081), .Z(n18180) );
  XOR U20731 ( .A(n18275), .B(n18276), .Z(n18081) );
  AND U20732 ( .A(n132), .B(n18277), .Z(n18275) );
  XOR U20733 ( .A(n18278), .B(n18276), .Z(n18277) );
  NANDN U20734 ( .A(n18083), .B(n18085), .Z(n18178) );
  XOR U20735 ( .A(n18279), .B(n18280), .Z(n18085) );
  AND U20736 ( .A(n132), .B(n18281), .Z(n18279) );
  XOR U20737 ( .A(n18280), .B(n18282), .Z(n18281) );
  XNOR U20738 ( .A(n18283), .B(n18284), .Z(n132) );
  AND U20739 ( .A(n18285), .B(n18286), .Z(n18283) );
  XOR U20740 ( .A(n18284), .B(n18096), .Z(n18286) );
  XNOR U20741 ( .A(n18287), .B(n18288), .Z(n18096) );
  ANDN U20742 ( .B(n18289), .A(n18290), .Z(n18287) );
  XOR U20743 ( .A(n18288), .B(n18291), .Z(n18289) );
  XNOR U20744 ( .A(n18284), .B(n18098), .Z(n18285) );
  XOR U20745 ( .A(n18292), .B(n18293), .Z(n18098) );
  AND U20746 ( .A(n136), .B(n18294), .Z(n18292) );
  XOR U20747 ( .A(n18295), .B(n18293), .Z(n18294) );
  XOR U20748 ( .A(n18296), .B(n18297), .Z(n18284) );
  AND U20749 ( .A(n18298), .B(n18299), .Z(n18296) );
  XOR U20750 ( .A(n18297), .B(n18123), .Z(n18299) );
  XOR U20751 ( .A(n18290), .B(n18291), .Z(n18123) );
  XNOR U20752 ( .A(n18300), .B(n18301), .Z(n18291) );
  ANDN U20753 ( .B(n18302), .A(n18303), .Z(n18300) );
  XOR U20754 ( .A(n18304), .B(n18305), .Z(n18302) );
  XOR U20755 ( .A(n18306), .B(n18307), .Z(n18290) );
  XNOR U20756 ( .A(n18308), .B(n18309), .Z(n18307) );
  ANDN U20757 ( .B(n18310), .A(n18311), .Z(n18308) );
  XNOR U20758 ( .A(n18312), .B(n18313), .Z(n18310) );
  IV U20759 ( .A(n18288), .Z(n18306) );
  XOR U20760 ( .A(n18314), .B(n18315), .Z(n18288) );
  ANDN U20761 ( .B(n18316), .A(n18317), .Z(n18314) );
  XOR U20762 ( .A(n18315), .B(n18318), .Z(n18316) );
  XNOR U20763 ( .A(n18297), .B(n18125), .Z(n18298) );
  XOR U20764 ( .A(n18319), .B(n18320), .Z(n18125) );
  AND U20765 ( .A(n136), .B(n18321), .Z(n18319) );
  XOR U20766 ( .A(n18322), .B(n18320), .Z(n18321) );
  XNOR U20767 ( .A(n18323), .B(n18324), .Z(n18297) );
  AND U20768 ( .A(n18325), .B(n18326), .Z(n18323) );
  XNOR U20769 ( .A(n18324), .B(n18175), .Z(n18326) );
  XOR U20770 ( .A(n18317), .B(n18318), .Z(n18175) );
  XOR U20771 ( .A(n18327), .B(n18305), .Z(n18318) );
  XNOR U20772 ( .A(n18328), .B(n18329), .Z(n18305) );
  ANDN U20773 ( .B(n18330), .A(n18331), .Z(n18328) );
  XOR U20774 ( .A(n18332), .B(n18333), .Z(n18330) );
  IV U20775 ( .A(n18303), .Z(n18327) );
  XOR U20776 ( .A(n18301), .B(n18334), .Z(n18303) );
  XNOR U20777 ( .A(n18335), .B(n18336), .Z(n18334) );
  ANDN U20778 ( .B(n18337), .A(n18338), .Z(n18335) );
  XNOR U20779 ( .A(n18339), .B(n18340), .Z(n18337) );
  IV U20780 ( .A(n18304), .Z(n18301) );
  XOR U20781 ( .A(n18341), .B(n18342), .Z(n18304) );
  ANDN U20782 ( .B(n18343), .A(n18344), .Z(n18341) );
  XOR U20783 ( .A(n18342), .B(n18345), .Z(n18343) );
  XOR U20784 ( .A(n18346), .B(n18347), .Z(n18317) );
  XNOR U20785 ( .A(n18312), .B(n18348), .Z(n18347) );
  IV U20786 ( .A(n18315), .Z(n18348) );
  XOR U20787 ( .A(n18349), .B(n18350), .Z(n18315) );
  ANDN U20788 ( .B(n18351), .A(n18352), .Z(n18349) );
  XOR U20789 ( .A(n18350), .B(n18353), .Z(n18351) );
  XNOR U20790 ( .A(n18354), .B(n18355), .Z(n18312) );
  ANDN U20791 ( .B(n18356), .A(n18357), .Z(n18354) );
  XOR U20792 ( .A(n18355), .B(n18358), .Z(n18356) );
  IV U20793 ( .A(n18311), .Z(n18346) );
  XOR U20794 ( .A(n18309), .B(n18359), .Z(n18311) );
  XNOR U20795 ( .A(n18360), .B(n18361), .Z(n18359) );
  ANDN U20796 ( .B(n18362), .A(n18363), .Z(n18360) );
  XNOR U20797 ( .A(n18364), .B(n18365), .Z(n18362) );
  IV U20798 ( .A(n18313), .Z(n18309) );
  XOR U20799 ( .A(n18366), .B(n18367), .Z(n18313) );
  ANDN U20800 ( .B(n18368), .A(n18369), .Z(n18366) );
  XOR U20801 ( .A(n18370), .B(n18367), .Z(n18368) );
  XOR U20802 ( .A(n18324), .B(n18177), .Z(n18325) );
  XOR U20803 ( .A(n18371), .B(n18372), .Z(n18177) );
  AND U20804 ( .A(n136), .B(n18373), .Z(n18371) );
  XOR U20805 ( .A(n18374), .B(n18372), .Z(n18373) );
  XNOR U20806 ( .A(n18375), .B(n18376), .Z(n18324) );
  NAND U20807 ( .A(n18377), .B(n18378), .Z(n18376) );
  XOR U20808 ( .A(n18379), .B(n18276), .Z(n18378) );
  XOR U20809 ( .A(n18352), .B(n18353), .Z(n18276) );
  XOR U20810 ( .A(n18380), .B(n18345), .Z(n18353) );
  XOR U20811 ( .A(n18381), .B(n18333), .Z(n18345) );
  XOR U20812 ( .A(n18382), .B(n18383), .Z(n18333) );
  ANDN U20813 ( .B(n18384), .A(n18385), .Z(n18382) );
  XOR U20814 ( .A(n18383), .B(n18386), .Z(n18384) );
  IV U20815 ( .A(n18331), .Z(n18381) );
  XOR U20816 ( .A(n18329), .B(n18387), .Z(n18331) );
  XOR U20817 ( .A(n18388), .B(n18389), .Z(n18387) );
  ANDN U20818 ( .B(n18390), .A(n18391), .Z(n18388) );
  XOR U20819 ( .A(n18392), .B(n18389), .Z(n18390) );
  IV U20820 ( .A(n18332), .Z(n18329) );
  XOR U20821 ( .A(n18393), .B(n18394), .Z(n18332) );
  ANDN U20822 ( .B(n18395), .A(n18396), .Z(n18393) );
  XOR U20823 ( .A(n18394), .B(n18397), .Z(n18395) );
  IV U20824 ( .A(n18344), .Z(n18380) );
  XOR U20825 ( .A(n18398), .B(n18399), .Z(n18344) );
  XNOR U20826 ( .A(n18339), .B(n18400), .Z(n18399) );
  IV U20827 ( .A(n18342), .Z(n18400) );
  XOR U20828 ( .A(n18401), .B(n18402), .Z(n18342) );
  ANDN U20829 ( .B(n18403), .A(n18404), .Z(n18401) );
  XOR U20830 ( .A(n18402), .B(n18405), .Z(n18403) );
  XNOR U20831 ( .A(n18406), .B(n18407), .Z(n18339) );
  ANDN U20832 ( .B(n18408), .A(n18409), .Z(n18406) );
  XOR U20833 ( .A(n18407), .B(n18410), .Z(n18408) );
  IV U20834 ( .A(n18338), .Z(n18398) );
  XOR U20835 ( .A(n18336), .B(n18411), .Z(n18338) );
  XOR U20836 ( .A(n18412), .B(n18413), .Z(n18411) );
  ANDN U20837 ( .B(n18414), .A(n18415), .Z(n18412) );
  XOR U20838 ( .A(n18416), .B(n18413), .Z(n18414) );
  IV U20839 ( .A(n18340), .Z(n18336) );
  XOR U20840 ( .A(n18417), .B(n18418), .Z(n18340) );
  ANDN U20841 ( .B(n18419), .A(n18420), .Z(n18417) );
  XOR U20842 ( .A(n18421), .B(n18418), .Z(n18419) );
  XOR U20843 ( .A(n18422), .B(n18423), .Z(n18352) );
  XOR U20844 ( .A(n18370), .B(n18424), .Z(n18423) );
  IV U20845 ( .A(n18350), .Z(n18424) );
  XOR U20846 ( .A(n18425), .B(n18426), .Z(n18350) );
  ANDN U20847 ( .B(n18427), .A(n18428), .Z(n18425) );
  XOR U20848 ( .A(n18426), .B(n18429), .Z(n18427) );
  XOR U20849 ( .A(n18430), .B(n18358), .Z(n18370) );
  XOR U20850 ( .A(n18431), .B(n18432), .Z(n18358) );
  ANDN U20851 ( .B(n18433), .A(n18434), .Z(n18431) );
  XOR U20852 ( .A(n18432), .B(n18435), .Z(n18433) );
  IV U20853 ( .A(n18357), .Z(n18430) );
  XOR U20854 ( .A(n18436), .B(n18437), .Z(n18357) );
  XOR U20855 ( .A(n18438), .B(n18439), .Z(n18437) );
  ANDN U20856 ( .B(n18440), .A(n18441), .Z(n18438) );
  XOR U20857 ( .A(n18442), .B(n18439), .Z(n18440) );
  IV U20858 ( .A(n18355), .Z(n18436) );
  XOR U20859 ( .A(n18443), .B(n18444), .Z(n18355) );
  ANDN U20860 ( .B(n18445), .A(n18446), .Z(n18443) );
  XOR U20861 ( .A(n18444), .B(n18447), .Z(n18445) );
  IV U20862 ( .A(n18369), .Z(n18422) );
  XOR U20863 ( .A(n18448), .B(n18449), .Z(n18369) );
  XNOR U20864 ( .A(n18364), .B(n18450), .Z(n18449) );
  IV U20865 ( .A(n18367), .Z(n18450) );
  XOR U20866 ( .A(n18451), .B(n18452), .Z(n18367) );
  ANDN U20867 ( .B(n18453), .A(n18454), .Z(n18451) );
  XOR U20868 ( .A(n18455), .B(n18452), .Z(n18453) );
  XNOR U20869 ( .A(n18456), .B(n18457), .Z(n18364) );
  ANDN U20870 ( .B(n18458), .A(n18459), .Z(n18456) );
  XOR U20871 ( .A(n18457), .B(n18460), .Z(n18458) );
  IV U20872 ( .A(n18363), .Z(n18448) );
  XOR U20873 ( .A(n18361), .B(n18461), .Z(n18363) );
  XOR U20874 ( .A(n18462), .B(n18463), .Z(n18461) );
  ANDN U20875 ( .B(n18464), .A(n18465), .Z(n18462) );
  XOR U20876 ( .A(n18466), .B(n18463), .Z(n18464) );
  IV U20877 ( .A(n18365), .Z(n18361) );
  XOR U20878 ( .A(n18467), .B(n18468), .Z(n18365) );
  ANDN U20879 ( .B(n18469), .A(n18470), .Z(n18467) );
  XOR U20880 ( .A(n18471), .B(n18468), .Z(n18469) );
  IV U20881 ( .A(n18375), .Z(n18379) );
  XOR U20882 ( .A(n18375), .B(n18278), .Z(n18377) );
  XOR U20883 ( .A(n18472), .B(n18473), .Z(n18278) );
  AND U20884 ( .A(n136), .B(n18474), .Z(n18472) );
  XOR U20885 ( .A(n18475), .B(n18473), .Z(n18474) );
  NANDN U20886 ( .A(n18280), .B(n18282), .Z(n18375) );
  XOR U20887 ( .A(n18476), .B(n18477), .Z(n18282) );
  AND U20888 ( .A(n136), .B(n18478), .Z(n18476) );
  XOR U20889 ( .A(n18477), .B(n18479), .Z(n18478) );
  XNOR U20890 ( .A(n18480), .B(n18481), .Z(n136) );
  AND U20891 ( .A(n18482), .B(n18483), .Z(n18480) );
  XOR U20892 ( .A(n18481), .B(n18293), .Z(n18483) );
  XNOR U20893 ( .A(n18484), .B(n18485), .Z(n18293) );
  ANDN U20894 ( .B(n18486), .A(n18487), .Z(n18484) );
  XOR U20895 ( .A(n18485), .B(n18488), .Z(n18486) );
  XNOR U20896 ( .A(n18481), .B(n18295), .Z(n18482) );
  XOR U20897 ( .A(n18489), .B(n18490), .Z(n18295) );
  AND U20898 ( .A(n140), .B(n18491), .Z(n18489) );
  XOR U20899 ( .A(n18492), .B(n18490), .Z(n18491) );
  XOR U20900 ( .A(n18493), .B(n18494), .Z(n18481) );
  AND U20901 ( .A(n18495), .B(n18496), .Z(n18493) );
  XOR U20902 ( .A(n18494), .B(n18320), .Z(n18496) );
  XOR U20903 ( .A(n18487), .B(n18488), .Z(n18320) );
  XNOR U20904 ( .A(n18497), .B(n18498), .Z(n18488) );
  ANDN U20905 ( .B(n18499), .A(n18500), .Z(n18497) );
  XOR U20906 ( .A(n18501), .B(n18502), .Z(n18499) );
  XOR U20907 ( .A(n18503), .B(n18504), .Z(n18487) );
  XNOR U20908 ( .A(n18505), .B(n18506), .Z(n18504) );
  ANDN U20909 ( .B(n18507), .A(n18508), .Z(n18505) );
  XNOR U20910 ( .A(n18509), .B(n18510), .Z(n18507) );
  IV U20911 ( .A(n18485), .Z(n18503) );
  XOR U20912 ( .A(n18511), .B(n18512), .Z(n18485) );
  ANDN U20913 ( .B(n18513), .A(n18514), .Z(n18511) );
  XOR U20914 ( .A(n18512), .B(n18515), .Z(n18513) );
  XNOR U20915 ( .A(n18494), .B(n18322), .Z(n18495) );
  XOR U20916 ( .A(n18516), .B(n18517), .Z(n18322) );
  AND U20917 ( .A(n140), .B(n18518), .Z(n18516) );
  XOR U20918 ( .A(n18519), .B(n18517), .Z(n18518) );
  XNOR U20919 ( .A(n18520), .B(n18521), .Z(n18494) );
  AND U20920 ( .A(n18522), .B(n18523), .Z(n18520) );
  XNOR U20921 ( .A(n18521), .B(n18372), .Z(n18523) );
  XOR U20922 ( .A(n18514), .B(n18515), .Z(n18372) );
  XOR U20923 ( .A(n18524), .B(n18502), .Z(n18515) );
  XNOR U20924 ( .A(n18525), .B(n18526), .Z(n18502) );
  ANDN U20925 ( .B(n18527), .A(n18528), .Z(n18525) );
  XOR U20926 ( .A(n18529), .B(n18530), .Z(n18527) );
  IV U20927 ( .A(n18500), .Z(n18524) );
  XOR U20928 ( .A(n18498), .B(n18531), .Z(n18500) );
  XNOR U20929 ( .A(n18532), .B(n18533), .Z(n18531) );
  ANDN U20930 ( .B(n18534), .A(n18535), .Z(n18532) );
  XNOR U20931 ( .A(n18536), .B(n18537), .Z(n18534) );
  IV U20932 ( .A(n18501), .Z(n18498) );
  XOR U20933 ( .A(n18538), .B(n18539), .Z(n18501) );
  ANDN U20934 ( .B(n18540), .A(n18541), .Z(n18538) );
  XOR U20935 ( .A(n18539), .B(n18542), .Z(n18540) );
  XOR U20936 ( .A(n18543), .B(n18544), .Z(n18514) );
  XNOR U20937 ( .A(n18509), .B(n18545), .Z(n18544) );
  IV U20938 ( .A(n18512), .Z(n18545) );
  XOR U20939 ( .A(n18546), .B(n18547), .Z(n18512) );
  ANDN U20940 ( .B(n18548), .A(n18549), .Z(n18546) );
  XOR U20941 ( .A(n18547), .B(n18550), .Z(n18548) );
  XNOR U20942 ( .A(n18551), .B(n18552), .Z(n18509) );
  ANDN U20943 ( .B(n18553), .A(n18554), .Z(n18551) );
  XOR U20944 ( .A(n18552), .B(n18555), .Z(n18553) );
  IV U20945 ( .A(n18508), .Z(n18543) );
  XOR U20946 ( .A(n18506), .B(n18556), .Z(n18508) );
  XNOR U20947 ( .A(n18557), .B(n18558), .Z(n18556) );
  ANDN U20948 ( .B(n18559), .A(n18560), .Z(n18557) );
  XNOR U20949 ( .A(n18561), .B(n18562), .Z(n18559) );
  IV U20950 ( .A(n18510), .Z(n18506) );
  XOR U20951 ( .A(n18563), .B(n18564), .Z(n18510) );
  ANDN U20952 ( .B(n18565), .A(n18566), .Z(n18563) );
  XOR U20953 ( .A(n18567), .B(n18564), .Z(n18565) );
  XOR U20954 ( .A(n18521), .B(n18374), .Z(n18522) );
  XOR U20955 ( .A(n18568), .B(n18569), .Z(n18374) );
  AND U20956 ( .A(n140), .B(n18570), .Z(n18568) );
  XOR U20957 ( .A(n18571), .B(n18569), .Z(n18570) );
  XNOR U20958 ( .A(n18572), .B(n18573), .Z(n18521) );
  NAND U20959 ( .A(n18574), .B(n18575), .Z(n18573) );
  XOR U20960 ( .A(n18576), .B(n18473), .Z(n18575) );
  XOR U20961 ( .A(n18549), .B(n18550), .Z(n18473) );
  XOR U20962 ( .A(n18577), .B(n18542), .Z(n18550) );
  XOR U20963 ( .A(n18578), .B(n18530), .Z(n18542) );
  XOR U20964 ( .A(n18579), .B(n18580), .Z(n18530) );
  ANDN U20965 ( .B(n18581), .A(n18582), .Z(n18579) );
  XOR U20966 ( .A(n18580), .B(n18583), .Z(n18581) );
  IV U20967 ( .A(n18528), .Z(n18578) );
  XOR U20968 ( .A(n18526), .B(n18584), .Z(n18528) );
  XOR U20969 ( .A(n18585), .B(n18586), .Z(n18584) );
  ANDN U20970 ( .B(n18587), .A(n18588), .Z(n18585) );
  XOR U20971 ( .A(n18589), .B(n18586), .Z(n18587) );
  IV U20972 ( .A(n18529), .Z(n18526) );
  XOR U20973 ( .A(n18590), .B(n18591), .Z(n18529) );
  ANDN U20974 ( .B(n18592), .A(n18593), .Z(n18590) );
  XOR U20975 ( .A(n18591), .B(n18594), .Z(n18592) );
  IV U20976 ( .A(n18541), .Z(n18577) );
  XOR U20977 ( .A(n18595), .B(n18596), .Z(n18541) );
  XNOR U20978 ( .A(n18536), .B(n18597), .Z(n18596) );
  IV U20979 ( .A(n18539), .Z(n18597) );
  XOR U20980 ( .A(n18598), .B(n18599), .Z(n18539) );
  ANDN U20981 ( .B(n18600), .A(n18601), .Z(n18598) );
  XOR U20982 ( .A(n18599), .B(n18602), .Z(n18600) );
  XNOR U20983 ( .A(n18603), .B(n18604), .Z(n18536) );
  ANDN U20984 ( .B(n18605), .A(n18606), .Z(n18603) );
  XOR U20985 ( .A(n18604), .B(n18607), .Z(n18605) );
  IV U20986 ( .A(n18535), .Z(n18595) );
  XOR U20987 ( .A(n18533), .B(n18608), .Z(n18535) );
  XOR U20988 ( .A(n18609), .B(n18610), .Z(n18608) );
  ANDN U20989 ( .B(n18611), .A(n18612), .Z(n18609) );
  XOR U20990 ( .A(n18613), .B(n18610), .Z(n18611) );
  IV U20991 ( .A(n18537), .Z(n18533) );
  XOR U20992 ( .A(n18614), .B(n18615), .Z(n18537) );
  ANDN U20993 ( .B(n18616), .A(n18617), .Z(n18614) );
  XOR U20994 ( .A(n18618), .B(n18615), .Z(n18616) );
  XOR U20995 ( .A(n18619), .B(n18620), .Z(n18549) );
  XOR U20996 ( .A(n18567), .B(n18621), .Z(n18620) );
  IV U20997 ( .A(n18547), .Z(n18621) );
  XOR U20998 ( .A(n18622), .B(n18623), .Z(n18547) );
  ANDN U20999 ( .B(n18624), .A(n18625), .Z(n18622) );
  XOR U21000 ( .A(n18623), .B(n18626), .Z(n18624) );
  XOR U21001 ( .A(n18627), .B(n18555), .Z(n18567) );
  XOR U21002 ( .A(n18628), .B(n18629), .Z(n18555) );
  ANDN U21003 ( .B(n18630), .A(n18631), .Z(n18628) );
  XOR U21004 ( .A(n18629), .B(n18632), .Z(n18630) );
  IV U21005 ( .A(n18554), .Z(n18627) );
  XOR U21006 ( .A(n18633), .B(n18634), .Z(n18554) );
  XOR U21007 ( .A(n18635), .B(n18636), .Z(n18634) );
  ANDN U21008 ( .B(n18637), .A(n18638), .Z(n18635) );
  XOR U21009 ( .A(n18639), .B(n18636), .Z(n18637) );
  IV U21010 ( .A(n18552), .Z(n18633) );
  XOR U21011 ( .A(n18640), .B(n18641), .Z(n18552) );
  ANDN U21012 ( .B(n18642), .A(n18643), .Z(n18640) );
  XOR U21013 ( .A(n18641), .B(n18644), .Z(n18642) );
  IV U21014 ( .A(n18566), .Z(n18619) );
  XOR U21015 ( .A(n18645), .B(n18646), .Z(n18566) );
  XNOR U21016 ( .A(n18561), .B(n18647), .Z(n18646) );
  IV U21017 ( .A(n18564), .Z(n18647) );
  XOR U21018 ( .A(n18648), .B(n18649), .Z(n18564) );
  ANDN U21019 ( .B(n18650), .A(n18651), .Z(n18648) );
  XOR U21020 ( .A(n18652), .B(n18649), .Z(n18650) );
  XNOR U21021 ( .A(n18653), .B(n18654), .Z(n18561) );
  ANDN U21022 ( .B(n18655), .A(n18656), .Z(n18653) );
  XOR U21023 ( .A(n18654), .B(n18657), .Z(n18655) );
  IV U21024 ( .A(n18560), .Z(n18645) );
  XOR U21025 ( .A(n18558), .B(n18658), .Z(n18560) );
  XOR U21026 ( .A(n18659), .B(n18660), .Z(n18658) );
  ANDN U21027 ( .B(n18661), .A(n18662), .Z(n18659) );
  XOR U21028 ( .A(n18663), .B(n18660), .Z(n18661) );
  IV U21029 ( .A(n18562), .Z(n18558) );
  XOR U21030 ( .A(n18664), .B(n18665), .Z(n18562) );
  ANDN U21031 ( .B(n18666), .A(n18667), .Z(n18664) );
  XOR U21032 ( .A(n18668), .B(n18665), .Z(n18666) );
  IV U21033 ( .A(n18572), .Z(n18576) );
  XOR U21034 ( .A(n18572), .B(n18475), .Z(n18574) );
  XOR U21035 ( .A(n18669), .B(n18670), .Z(n18475) );
  AND U21036 ( .A(n140), .B(n18671), .Z(n18669) );
  XOR U21037 ( .A(n18672), .B(n18670), .Z(n18671) );
  NANDN U21038 ( .A(n18477), .B(n18479), .Z(n18572) );
  XOR U21039 ( .A(n18673), .B(n18674), .Z(n18479) );
  AND U21040 ( .A(n140), .B(n18675), .Z(n18673) );
  XOR U21041 ( .A(n18674), .B(n18676), .Z(n18675) );
  XNOR U21042 ( .A(n18677), .B(n18678), .Z(n140) );
  AND U21043 ( .A(n18679), .B(n18680), .Z(n18677) );
  XOR U21044 ( .A(n18678), .B(n18490), .Z(n18680) );
  XNOR U21045 ( .A(n18681), .B(n18682), .Z(n18490) );
  ANDN U21046 ( .B(n18683), .A(n18684), .Z(n18681) );
  XOR U21047 ( .A(n18682), .B(n18685), .Z(n18683) );
  XNOR U21048 ( .A(n18678), .B(n18492), .Z(n18679) );
  XOR U21049 ( .A(n18686), .B(n18687), .Z(n18492) );
  AND U21050 ( .A(n144), .B(n18688), .Z(n18686) );
  XOR U21051 ( .A(n18689), .B(n18687), .Z(n18688) );
  XOR U21052 ( .A(n18690), .B(n18691), .Z(n18678) );
  AND U21053 ( .A(n18692), .B(n18693), .Z(n18690) );
  XOR U21054 ( .A(n18691), .B(n18517), .Z(n18693) );
  XOR U21055 ( .A(n18684), .B(n18685), .Z(n18517) );
  XNOR U21056 ( .A(n18694), .B(n18695), .Z(n18685) );
  ANDN U21057 ( .B(n18696), .A(n18697), .Z(n18694) );
  XOR U21058 ( .A(n18698), .B(n18699), .Z(n18696) );
  XOR U21059 ( .A(n18700), .B(n18701), .Z(n18684) );
  XNOR U21060 ( .A(n18702), .B(n18703), .Z(n18701) );
  ANDN U21061 ( .B(n18704), .A(n18705), .Z(n18702) );
  XNOR U21062 ( .A(n18706), .B(n18707), .Z(n18704) );
  IV U21063 ( .A(n18682), .Z(n18700) );
  XOR U21064 ( .A(n18708), .B(n18709), .Z(n18682) );
  ANDN U21065 ( .B(n18710), .A(n18711), .Z(n18708) );
  XOR U21066 ( .A(n18709), .B(n18712), .Z(n18710) );
  XNOR U21067 ( .A(n18691), .B(n18519), .Z(n18692) );
  XOR U21068 ( .A(n18713), .B(n18714), .Z(n18519) );
  AND U21069 ( .A(n144), .B(n18715), .Z(n18713) );
  XOR U21070 ( .A(n18716), .B(n18714), .Z(n18715) );
  XNOR U21071 ( .A(n18717), .B(n18718), .Z(n18691) );
  AND U21072 ( .A(n18719), .B(n18720), .Z(n18717) );
  XNOR U21073 ( .A(n18718), .B(n18569), .Z(n18720) );
  XOR U21074 ( .A(n18711), .B(n18712), .Z(n18569) );
  XOR U21075 ( .A(n18721), .B(n18699), .Z(n18712) );
  XNOR U21076 ( .A(n18722), .B(n18723), .Z(n18699) );
  ANDN U21077 ( .B(n18724), .A(n18725), .Z(n18722) );
  XOR U21078 ( .A(n18726), .B(n18727), .Z(n18724) );
  IV U21079 ( .A(n18697), .Z(n18721) );
  XOR U21080 ( .A(n18695), .B(n18728), .Z(n18697) );
  XNOR U21081 ( .A(n18729), .B(n18730), .Z(n18728) );
  ANDN U21082 ( .B(n18731), .A(n18732), .Z(n18729) );
  XNOR U21083 ( .A(n18733), .B(n18734), .Z(n18731) );
  IV U21084 ( .A(n18698), .Z(n18695) );
  XOR U21085 ( .A(n18735), .B(n18736), .Z(n18698) );
  ANDN U21086 ( .B(n18737), .A(n18738), .Z(n18735) );
  XOR U21087 ( .A(n18736), .B(n18739), .Z(n18737) );
  XOR U21088 ( .A(n18740), .B(n18741), .Z(n18711) );
  XNOR U21089 ( .A(n18706), .B(n18742), .Z(n18741) );
  IV U21090 ( .A(n18709), .Z(n18742) );
  XOR U21091 ( .A(n18743), .B(n18744), .Z(n18709) );
  ANDN U21092 ( .B(n18745), .A(n18746), .Z(n18743) );
  XOR U21093 ( .A(n18744), .B(n18747), .Z(n18745) );
  XNOR U21094 ( .A(n18748), .B(n18749), .Z(n18706) );
  ANDN U21095 ( .B(n18750), .A(n18751), .Z(n18748) );
  XOR U21096 ( .A(n18749), .B(n18752), .Z(n18750) );
  IV U21097 ( .A(n18705), .Z(n18740) );
  XOR U21098 ( .A(n18703), .B(n18753), .Z(n18705) );
  XNOR U21099 ( .A(n18754), .B(n18755), .Z(n18753) );
  ANDN U21100 ( .B(n18756), .A(n18757), .Z(n18754) );
  XNOR U21101 ( .A(n18758), .B(n18759), .Z(n18756) );
  IV U21102 ( .A(n18707), .Z(n18703) );
  XOR U21103 ( .A(n18760), .B(n18761), .Z(n18707) );
  ANDN U21104 ( .B(n18762), .A(n18763), .Z(n18760) );
  XOR U21105 ( .A(n18764), .B(n18761), .Z(n18762) );
  XOR U21106 ( .A(n18718), .B(n18571), .Z(n18719) );
  XOR U21107 ( .A(n18765), .B(n18766), .Z(n18571) );
  AND U21108 ( .A(n144), .B(n18767), .Z(n18765) );
  XOR U21109 ( .A(n18768), .B(n18766), .Z(n18767) );
  XNOR U21110 ( .A(n18769), .B(n18770), .Z(n18718) );
  NAND U21111 ( .A(n18771), .B(n18772), .Z(n18770) );
  XOR U21112 ( .A(n18773), .B(n18670), .Z(n18772) );
  XOR U21113 ( .A(n18746), .B(n18747), .Z(n18670) );
  XOR U21114 ( .A(n18774), .B(n18739), .Z(n18747) );
  XOR U21115 ( .A(n18775), .B(n18727), .Z(n18739) );
  XOR U21116 ( .A(n18776), .B(n18777), .Z(n18727) );
  ANDN U21117 ( .B(n18778), .A(n18779), .Z(n18776) );
  XOR U21118 ( .A(n18777), .B(n18780), .Z(n18778) );
  IV U21119 ( .A(n18725), .Z(n18775) );
  XOR U21120 ( .A(n18723), .B(n18781), .Z(n18725) );
  XOR U21121 ( .A(n18782), .B(n18783), .Z(n18781) );
  ANDN U21122 ( .B(n18784), .A(n18785), .Z(n18782) );
  XOR U21123 ( .A(n18786), .B(n18783), .Z(n18784) );
  IV U21124 ( .A(n18726), .Z(n18723) );
  XOR U21125 ( .A(n18787), .B(n18788), .Z(n18726) );
  ANDN U21126 ( .B(n18789), .A(n18790), .Z(n18787) );
  XOR U21127 ( .A(n18788), .B(n18791), .Z(n18789) );
  IV U21128 ( .A(n18738), .Z(n18774) );
  XOR U21129 ( .A(n18792), .B(n18793), .Z(n18738) );
  XNOR U21130 ( .A(n18733), .B(n18794), .Z(n18793) );
  IV U21131 ( .A(n18736), .Z(n18794) );
  XOR U21132 ( .A(n18795), .B(n18796), .Z(n18736) );
  ANDN U21133 ( .B(n18797), .A(n18798), .Z(n18795) );
  XOR U21134 ( .A(n18796), .B(n18799), .Z(n18797) );
  XNOR U21135 ( .A(n18800), .B(n18801), .Z(n18733) );
  ANDN U21136 ( .B(n18802), .A(n18803), .Z(n18800) );
  XOR U21137 ( .A(n18801), .B(n18804), .Z(n18802) );
  IV U21138 ( .A(n18732), .Z(n18792) );
  XOR U21139 ( .A(n18730), .B(n18805), .Z(n18732) );
  XOR U21140 ( .A(n18806), .B(n18807), .Z(n18805) );
  ANDN U21141 ( .B(n18808), .A(n18809), .Z(n18806) );
  XOR U21142 ( .A(n18810), .B(n18807), .Z(n18808) );
  IV U21143 ( .A(n18734), .Z(n18730) );
  XOR U21144 ( .A(n18811), .B(n18812), .Z(n18734) );
  ANDN U21145 ( .B(n18813), .A(n18814), .Z(n18811) );
  XOR U21146 ( .A(n18815), .B(n18812), .Z(n18813) );
  XOR U21147 ( .A(n18816), .B(n18817), .Z(n18746) );
  XOR U21148 ( .A(n18764), .B(n18818), .Z(n18817) );
  IV U21149 ( .A(n18744), .Z(n18818) );
  XOR U21150 ( .A(n18819), .B(n18820), .Z(n18744) );
  ANDN U21151 ( .B(n18821), .A(n18822), .Z(n18819) );
  XOR U21152 ( .A(n18820), .B(n18823), .Z(n18821) );
  XOR U21153 ( .A(n18824), .B(n18752), .Z(n18764) );
  XOR U21154 ( .A(n18825), .B(n18826), .Z(n18752) );
  ANDN U21155 ( .B(n18827), .A(n18828), .Z(n18825) );
  XOR U21156 ( .A(n18826), .B(n18829), .Z(n18827) );
  IV U21157 ( .A(n18751), .Z(n18824) );
  XOR U21158 ( .A(n18830), .B(n18831), .Z(n18751) );
  XOR U21159 ( .A(n18832), .B(n18833), .Z(n18831) );
  ANDN U21160 ( .B(n18834), .A(n18835), .Z(n18832) );
  XOR U21161 ( .A(n18836), .B(n18833), .Z(n18834) );
  IV U21162 ( .A(n18749), .Z(n18830) );
  XOR U21163 ( .A(n18837), .B(n18838), .Z(n18749) );
  ANDN U21164 ( .B(n18839), .A(n18840), .Z(n18837) );
  XOR U21165 ( .A(n18838), .B(n18841), .Z(n18839) );
  IV U21166 ( .A(n18763), .Z(n18816) );
  XOR U21167 ( .A(n18842), .B(n18843), .Z(n18763) );
  XNOR U21168 ( .A(n18758), .B(n18844), .Z(n18843) );
  IV U21169 ( .A(n18761), .Z(n18844) );
  XOR U21170 ( .A(n18845), .B(n18846), .Z(n18761) );
  ANDN U21171 ( .B(n18847), .A(n18848), .Z(n18845) );
  XOR U21172 ( .A(n18849), .B(n18846), .Z(n18847) );
  XNOR U21173 ( .A(n18850), .B(n18851), .Z(n18758) );
  ANDN U21174 ( .B(n18852), .A(n18853), .Z(n18850) );
  XOR U21175 ( .A(n18851), .B(n18854), .Z(n18852) );
  IV U21176 ( .A(n18757), .Z(n18842) );
  XOR U21177 ( .A(n18755), .B(n18855), .Z(n18757) );
  XOR U21178 ( .A(n18856), .B(n18857), .Z(n18855) );
  ANDN U21179 ( .B(n18858), .A(n18859), .Z(n18856) );
  XOR U21180 ( .A(n18860), .B(n18857), .Z(n18858) );
  IV U21181 ( .A(n18759), .Z(n18755) );
  XOR U21182 ( .A(n18861), .B(n18862), .Z(n18759) );
  ANDN U21183 ( .B(n18863), .A(n18864), .Z(n18861) );
  XOR U21184 ( .A(n18865), .B(n18862), .Z(n18863) );
  IV U21185 ( .A(n18769), .Z(n18773) );
  XOR U21186 ( .A(n18769), .B(n18672), .Z(n18771) );
  XOR U21187 ( .A(n18866), .B(n18867), .Z(n18672) );
  AND U21188 ( .A(n144), .B(n18868), .Z(n18866) );
  XOR U21189 ( .A(n18869), .B(n18867), .Z(n18868) );
  NANDN U21190 ( .A(n18674), .B(n18676), .Z(n18769) );
  XOR U21191 ( .A(n18870), .B(n18871), .Z(n18676) );
  AND U21192 ( .A(n144), .B(n18872), .Z(n18870) );
  XOR U21193 ( .A(n18871), .B(n18873), .Z(n18872) );
  XNOR U21194 ( .A(n18874), .B(n18875), .Z(n144) );
  AND U21195 ( .A(n18876), .B(n18877), .Z(n18874) );
  XOR U21196 ( .A(n18875), .B(n18687), .Z(n18877) );
  XNOR U21197 ( .A(n18878), .B(n18879), .Z(n18687) );
  ANDN U21198 ( .B(n18880), .A(n18881), .Z(n18878) );
  XOR U21199 ( .A(n18879), .B(n18882), .Z(n18880) );
  XNOR U21200 ( .A(n18875), .B(n18689), .Z(n18876) );
  XOR U21201 ( .A(n18883), .B(n18884), .Z(n18689) );
  AND U21202 ( .A(n148), .B(n18885), .Z(n18883) );
  XOR U21203 ( .A(n18886), .B(n18884), .Z(n18885) );
  XOR U21204 ( .A(n18887), .B(n18888), .Z(n18875) );
  AND U21205 ( .A(n18889), .B(n18890), .Z(n18887) );
  XOR U21206 ( .A(n18888), .B(n18714), .Z(n18890) );
  XOR U21207 ( .A(n18881), .B(n18882), .Z(n18714) );
  XNOR U21208 ( .A(n18891), .B(n18892), .Z(n18882) );
  ANDN U21209 ( .B(n18893), .A(n18894), .Z(n18891) );
  XOR U21210 ( .A(n18895), .B(n18896), .Z(n18893) );
  XOR U21211 ( .A(n18897), .B(n18898), .Z(n18881) );
  XNOR U21212 ( .A(n18899), .B(n18900), .Z(n18898) );
  ANDN U21213 ( .B(n18901), .A(n18902), .Z(n18899) );
  XNOR U21214 ( .A(n18903), .B(n18904), .Z(n18901) );
  IV U21215 ( .A(n18879), .Z(n18897) );
  XOR U21216 ( .A(n18905), .B(n18906), .Z(n18879) );
  ANDN U21217 ( .B(n18907), .A(n18908), .Z(n18905) );
  XOR U21218 ( .A(n18906), .B(n18909), .Z(n18907) );
  XNOR U21219 ( .A(n18888), .B(n18716), .Z(n18889) );
  XOR U21220 ( .A(n18910), .B(n18911), .Z(n18716) );
  AND U21221 ( .A(n148), .B(n18912), .Z(n18910) );
  XOR U21222 ( .A(n18913), .B(n18911), .Z(n18912) );
  XNOR U21223 ( .A(n18914), .B(n18915), .Z(n18888) );
  AND U21224 ( .A(n18916), .B(n18917), .Z(n18914) );
  XNOR U21225 ( .A(n18915), .B(n18766), .Z(n18917) );
  XOR U21226 ( .A(n18908), .B(n18909), .Z(n18766) );
  XOR U21227 ( .A(n18918), .B(n18896), .Z(n18909) );
  XNOR U21228 ( .A(n18919), .B(n18920), .Z(n18896) );
  ANDN U21229 ( .B(n18921), .A(n18922), .Z(n18919) );
  XOR U21230 ( .A(n18923), .B(n18924), .Z(n18921) );
  IV U21231 ( .A(n18894), .Z(n18918) );
  XOR U21232 ( .A(n18892), .B(n18925), .Z(n18894) );
  XNOR U21233 ( .A(n18926), .B(n18927), .Z(n18925) );
  ANDN U21234 ( .B(n18928), .A(n18929), .Z(n18926) );
  XNOR U21235 ( .A(n18930), .B(n18931), .Z(n18928) );
  IV U21236 ( .A(n18895), .Z(n18892) );
  XOR U21237 ( .A(n18932), .B(n18933), .Z(n18895) );
  ANDN U21238 ( .B(n18934), .A(n18935), .Z(n18932) );
  XOR U21239 ( .A(n18933), .B(n18936), .Z(n18934) );
  XOR U21240 ( .A(n18937), .B(n18938), .Z(n18908) );
  XNOR U21241 ( .A(n18903), .B(n18939), .Z(n18938) );
  IV U21242 ( .A(n18906), .Z(n18939) );
  XOR U21243 ( .A(n18940), .B(n18941), .Z(n18906) );
  ANDN U21244 ( .B(n18942), .A(n18943), .Z(n18940) );
  XOR U21245 ( .A(n18941), .B(n18944), .Z(n18942) );
  XNOR U21246 ( .A(n18945), .B(n18946), .Z(n18903) );
  ANDN U21247 ( .B(n18947), .A(n18948), .Z(n18945) );
  XOR U21248 ( .A(n18946), .B(n18949), .Z(n18947) );
  IV U21249 ( .A(n18902), .Z(n18937) );
  XOR U21250 ( .A(n18900), .B(n18950), .Z(n18902) );
  XNOR U21251 ( .A(n18951), .B(n18952), .Z(n18950) );
  ANDN U21252 ( .B(n18953), .A(n18954), .Z(n18951) );
  XNOR U21253 ( .A(n18955), .B(n18956), .Z(n18953) );
  IV U21254 ( .A(n18904), .Z(n18900) );
  XOR U21255 ( .A(n18957), .B(n18958), .Z(n18904) );
  ANDN U21256 ( .B(n18959), .A(n18960), .Z(n18957) );
  XOR U21257 ( .A(n18961), .B(n18958), .Z(n18959) );
  XOR U21258 ( .A(n18915), .B(n18768), .Z(n18916) );
  XOR U21259 ( .A(n18962), .B(n18963), .Z(n18768) );
  AND U21260 ( .A(n148), .B(n18964), .Z(n18962) );
  XOR U21261 ( .A(n18965), .B(n18963), .Z(n18964) );
  XNOR U21262 ( .A(n18966), .B(n18967), .Z(n18915) );
  NAND U21263 ( .A(n18968), .B(n18969), .Z(n18967) );
  XOR U21264 ( .A(n18970), .B(n18867), .Z(n18969) );
  XOR U21265 ( .A(n18943), .B(n18944), .Z(n18867) );
  XOR U21266 ( .A(n18971), .B(n18936), .Z(n18944) );
  XOR U21267 ( .A(n18972), .B(n18924), .Z(n18936) );
  XOR U21268 ( .A(n18973), .B(n18974), .Z(n18924) );
  ANDN U21269 ( .B(n18975), .A(n18976), .Z(n18973) );
  XOR U21270 ( .A(n18974), .B(n18977), .Z(n18975) );
  IV U21271 ( .A(n18922), .Z(n18972) );
  XOR U21272 ( .A(n18920), .B(n18978), .Z(n18922) );
  XOR U21273 ( .A(n18979), .B(n18980), .Z(n18978) );
  ANDN U21274 ( .B(n18981), .A(n18982), .Z(n18979) );
  XOR U21275 ( .A(n18983), .B(n18980), .Z(n18981) );
  IV U21276 ( .A(n18923), .Z(n18920) );
  XOR U21277 ( .A(n18984), .B(n18985), .Z(n18923) );
  ANDN U21278 ( .B(n18986), .A(n18987), .Z(n18984) );
  XOR U21279 ( .A(n18985), .B(n18988), .Z(n18986) );
  IV U21280 ( .A(n18935), .Z(n18971) );
  XOR U21281 ( .A(n18989), .B(n18990), .Z(n18935) );
  XNOR U21282 ( .A(n18930), .B(n18991), .Z(n18990) );
  IV U21283 ( .A(n18933), .Z(n18991) );
  XOR U21284 ( .A(n18992), .B(n18993), .Z(n18933) );
  ANDN U21285 ( .B(n18994), .A(n18995), .Z(n18992) );
  XOR U21286 ( .A(n18993), .B(n18996), .Z(n18994) );
  XNOR U21287 ( .A(n18997), .B(n18998), .Z(n18930) );
  ANDN U21288 ( .B(n18999), .A(n19000), .Z(n18997) );
  XOR U21289 ( .A(n18998), .B(n19001), .Z(n18999) );
  IV U21290 ( .A(n18929), .Z(n18989) );
  XOR U21291 ( .A(n18927), .B(n19002), .Z(n18929) );
  XOR U21292 ( .A(n19003), .B(n19004), .Z(n19002) );
  ANDN U21293 ( .B(n19005), .A(n19006), .Z(n19003) );
  XOR U21294 ( .A(n19007), .B(n19004), .Z(n19005) );
  IV U21295 ( .A(n18931), .Z(n18927) );
  XOR U21296 ( .A(n19008), .B(n19009), .Z(n18931) );
  ANDN U21297 ( .B(n19010), .A(n19011), .Z(n19008) );
  XOR U21298 ( .A(n19012), .B(n19009), .Z(n19010) );
  XOR U21299 ( .A(n19013), .B(n19014), .Z(n18943) );
  XOR U21300 ( .A(n18961), .B(n19015), .Z(n19014) );
  IV U21301 ( .A(n18941), .Z(n19015) );
  XOR U21302 ( .A(n19016), .B(n19017), .Z(n18941) );
  ANDN U21303 ( .B(n19018), .A(n19019), .Z(n19016) );
  XOR U21304 ( .A(n19017), .B(n19020), .Z(n19018) );
  XOR U21305 ( .A(n19021), .B(n18949), .Z(n18961) );
  XOR U21306 ( .A(n19022), .B(n19023), .Z(n18949) );
  ANDN U21307 ( .B(n19024), .A(n19025), .Z(n19022) );
  XOR U21308 ( .A(n19023), .B(n19026), .Z(n19024) );
  IV U21309 ( .A(n18948), .Z(n19021) );
  XOR U21310 ( .A(n19027), .B(n19028), .Z(n18948) );
  XOR U21311 ( .A(n19029), .B(n19030), .Z(n19028) );
  ANDN U21312 ( .B(n19031), .A(n19032), .Z(n19029) );
  XOR U21313 ( .A(n19033), .B(n19030), .Z(n19031) );
  IV U21314 ( .A(n18946), .Z(n19027) );
  XOR U21315 ( .A(n19034), .B(n19035), .Z(n18946) );
  ANDN U21316 ( .B(n19036), .A(n19037), .Z(n19034) );
  XOR U21317 ( .A(n19035), .B(n19038), .Z(n19036) );
  IV U21318 ( .A(n18960), .Z(n19013) );
  XOR U21319 ( .A(n19039), .B(n19040), .Z(n18960) );
  XNOR U21320 ( .A(n18955), .B(n19041), .Z(n19040) );
  IV U21321 ( .A(n18958), .Z(n19041) );
  XOR U21322 ( .A(n19042), .B(n19043), .Z(n18958) );
  ANDN U21323 ( .B(n19044), .A(n19045), .Z(n19042) );
  XOR U21324 ( .A(n19046), .B(n19043), .Z(n19044) );
  XNOR U21325 ( .A(n19047), .B(n19048), .Z(n18955) );
  ANDN U21326 ( .B(n19049), .A(n19050), .Z(n19047) );
  XOR U21327 ( .A(n19048), .B(n19051), .Z(n19049) );
  IV U21328 ( .A(n18954), .Z(n19039) );
  XOR U21329 ( .A(n18952), .B(n19052), .Z(n18954) );
  XOR U21330 ( .A(n19053), .B(n19054), .Z(n19052) );
  ANDN U21331 ( .B(n19055), .A(n19056), .Z(n19053) );
  XOR U21332 ( .A(n19057), .B(n19054), .Z(n19055) );
  IV U21333 ( .A(n18956), .Z(n18952) );
  XOR U21334 ( .A(n19058), .B(n19059), .Z(n18956) );
  ANDN U21335 ( .B(n19060), .A(n19061), .Z(n19058) );
  XOR U21336 ( .A(n19062), .B(n19059), .Z(n19060) );
  IV U21337 ( .A(n18966), .Z(n18970) );
  XOR U21338 ( .A(n18966), .B(n18869), .Z(n18968) );
  XOR U21339 ( .A(n19063), .B(n19064), .Z(n18869) );
  AND U21340 ( .A(n148), .B(n19065), .Z(n19063) );
  XOR U21341 ( .A(n19066), .B(n19064), .Z(n19065) );
  NANDN U21342 ( .A(n18871), .B(n18873), .Z(n18966) );
  XOR U21343 ( .A(n19067), .B(n19068), .Z(n18873) );
  AND U21344 ( .A(n148), .B(n19069), .Z(n19067) );
  XOR U21345 ( .A(n19068), .B(n19070), .Z(n19069) );
  XNOR U21346 ( .A(n19071), .B(n19072), .Z(n148) );
  AND U21347 ( .A(n19073), .B(n19074), .Z(n19071) );
  XOR U21348 ( .A(n19072), .B(n18884), .Z(n19074) );
  XNOR U21349 ( .A(n19075), .B(n19076), .Z(n18884) );
  ANDN U21350 ( .B(n19077), .A(n19078), .Z(n19075) );
  XOR U21351 ( .A(n19076), .B(n19079), .Z(n19077) );
  XNOR U21352 ( .A(n19072), .B(n18886), .Z(n19073) );
  XOR U21353 ( .A(n19080), .B(n19081), .Z(n18886) );
  AND U21354 ( .A(n152), .B(n19082), .Z(n19080) );
  XOR U21355 ( .A(n19083), .B(n19081), .Z(n19082) );
  XOR U21356 ( .A(n19084), .B(n19085), .Z(n19072) );
  AND U21357 ( .A(n19086), .B(n19087), .Z(n19084) );
  XOR U21358 ( .A(n19085), .B(n18911), .Z(n19087) );
  XOR U21359 ( .A(n19078), .B(n19079), .Z(n18911) );
  XNOR U21360 ( .A(n19088), .B(n19089), .Z(n19079) );
  ANDN U21361 ( .B(n19090), .A(n19091), .Z(n19088) );
  XOR U21362 ( .A(n19092), .B(n19093), .Z(n19090) );
  XOR U21363 ( .A(n19094), .B(n19095), .Z(n19078) );
  XNOR U21364 ( .A(n19096), .B(n19097), .Z(n19095) );
  ANDN U21365 ( .B(n19098), .A(n19099), .Z(n19096) );
  XNOR U21366 ( .A(n19100), .B(n19101), .Z(n19098) );
  IV U21367 ( .A(n19076), .Z(n19094) );
  XOR U21368 ( .A(n19102), .B(n19103), .Z(n19076) );
  ANDN U21369 ( .B(n19104), .A(n19105), .Z(n19102) );
  XOR U21370 ( .A(n19103), .B(n19106), .Z(n19104) );
  XNOR U21371 ( .A(n19085), .B(n18913), .Z(n19086) );
  XOR U21372 ( .A(n19107), .B(n19108), .Z(n18913) );
  AND U21373 ( .A(n152), .B(n19109), .Z(n19107) );
  XOR U21374 ( .A(n19110), .B(n19108), .Z(n19109) );
  XNOR U21375 ( .A(n19111), .B(n19112), .Z(n19085) );
  AND U21376 ( .A(n19113), .B(n19114), .Z(n19111) );
  XNOR U21377 ( .A(n19112), .B(n18963), .Z(n19114) );
  XOR U21378 ( .A(n19105), .B(n19106), .Z(n18963) );
  XOR U21379 ( .A(n19115), .B(n19093), .Z(n19106) );
  XNOR U21380 ( .A(n19116), .B(n19117), .Z(n19093) );
  ANDN U21381 ( .B(n19118), .A(n19119), .Z(n19116) );
  XOR U21382 ( .A(n19120), .B(n19121), .Z(n19118) );
  IV U21383 ( .A(n19091), .Z(n19115) );
  XOR U21384 ( .A(n19089), .B(n19122), .Z(n19091) );
  XNOR U21385 ( .A(n19123), .B(n19124), .Z(n19122) );
  ANDN U21386 ( .B(n19125), .A(n19126), .Z(n19123) );
  XNOR U21387 ( .A(n19127), .B(n19128), .Z(n19125) );
  IV U21388 ( .A(n19092), .Z(n19089) );
  XOR U21389 ( .A(n19129), .B(n19130), .Z(n19092) );
  ANDN U21390 ( .B(n19131), .A(n19132), .Z(n19129) );
  XOR U21391 ( .A(n19130), .B(n19133), .Z(n19131) );
  XOR U21392 ( .A(n19134), .B(n19135), .Z(n19105) );
  XNOR U21393 ( .A(n19100), .B(n19136), .Z(n19135) );
  IV U21394 ( .A(n19103), .Z(n19136) );
  XOR U21395 ( .A(n19137), .B(n19138), .Z(n19103) );
  ANDN U21396 ( .B(n19139), .A(n19140), .Z(n19137) );
  XOR U21397 ( .A(n19138), .B(n19141), .Z(n19139) );
  XNOR U21398 ( .A(n19142), .B(n19143), .Z(n19100) );
  ANDN U21399 ( .B(n19144), .A(n19145), .Z(n19142) );
  XOR U21400 ( .A(n19143), .B(n19146), .Z(n19144) );
  IV U21401 ( .A(n19099), .Z(n19134) );
  XOR U21402 ( .A(n19097), .B(n19147), .Z(n19099) );
  XNOR U21403 ( .A(n19148), .B(n19149), .Z(n19147) );
  ANDN U21404 ( .B(n19150), .A(n19151), .Z(n19148) );
  XNOR U21405 ( .A(n19152), .B(n19153), .Z(n19150) );
  IV U21406 ( .A(n19101), .Z(n19097) );
  XOR U21407 ( .A(n19154), .B(n19155), .Z(n19101) );
  ANDN U21408 ( .B(n19156), .A(n19157), .Z(n19154) );
  XOR U21409 ( .A(n19158), .B(n19155), .Z(n19156) );
  XOR U21410 ( .A(n19112), .B(n18965), .Z(n19113) );
  XOR U21411 ( .A(n19159), .B(n19160), .Z(n18965) );
  AND U21412 ( .A(n152), .B(n19161), .Z(n19159) );
  XOR U21413 ( .A(n19162), .B(n19160), .Z(n19161) );
  XNOR U21414 ( .A(n19163), .B(n19164), .Z(n19112) );
  NAND U21415 ( .A(n19165), .B(n19166), .Z(n19164) );
  XOR U21416 ( .A(n19167), .B(n19064), .Z(n19166) );
  XOR U21417 ( .A(n19140), .B(n19141), .Z(n19064) );
  XOR U21418 ( .A(n19168), .B(n19133), .Z(n19141) );
  XOR U21419 ( .A(n19169), .B(n19121), .Z(n19133) );
  XOR U21420 ( .A(n19170), .B(n19171), .Z(n19121) );
  ANDN U21421 ( .B(n19172), .A(n19173), .Z(n19170) );
  XOR U21422 ( .A(n19171), .B(n19174), .Z(n19172) );
  IV U21423 ( .A(n19119), .Z(n19169) );
  XOR U21424 ( .A(n19117), .B(n19175), .Z(n19119) );
  XOR U21425 ( .A(n19176), .B(n19177), .Z(n19175) );
  ANDN U21426 ( .B(n19178), .A(n19179), .Z(n19176) );
  XOR U21427 ( .A(n19180), .B(n19177), .Z(n19178) );
  IV U21428 ( .A(n19120), .Z(n19117) );
  XOR U21429 ( .A(n19181), .B(n19182), .Z(n19120) );
  ANDN U21430 ( .B(n19183), .A(n19184), .Z(n19181) );
  XOR U21431 ( .A(n19182), .B(n19185), .Z(n19183) );
  IV U21432 ( .A(n19132), .Z(n19168) );
  XOR U21433 ( .A(n19186), .B(n19187), .Z(n19132) );
  XNOR U21434 ( .A(n19127), .B(n19188), .Z(n19187) );
  IV U21435 ( .A(n19130), .Z(n19188) );
  XOR U21436 ( .A(n19189), .B(n19190), .Z(n19130) );
  ANDN U21437 ( .B(n19191), .A(n19192), .Z(n19189) );
  XOR U21438 ( .A(n19190), .B(n19193), .Z(n19191) );
  XNOR U21439 ( .A(n19194), .B(n19195), .Z(n19127) );
  ANDN U21440 ( .B(n19196), .A(n19197), .Z(n19194) );
  XOR U21441 ( .A(n19195), .B(n19198), .Z(n19196) );
  IV U21442 ( .A(n19126), .Z(n19186) );
  XOR U21443 ( .A(n19124), .B(n19199), .Z(n19126) );
  XOR U21444 ( .A(n19200), .B(n19201), .Z(n19199) );
  ANDN U21445 ( .B(n19202), .A(n19203), .Z(n19200) );
  XOR U21446 ( .A(n19204), .B(n19201), .Z(n19202) );
  IV U21447 ( .A(n19128), .Z(n19124) );
  XOR U21448 ( .A(n19205), .B(n19206), .Z(n19128) );
  ANDN U21449 ( .B(n19207), .A(n19208), .Z(n19205) );
  XOR U21450 ( .A(n19209), .B(n19206), .Z(n19207) );
  XOR U21451 ( .A(n19210), .B(n19211), .Z(n19140) );
  XOR U21452 ( .A(n19158), .B(n19212), .Z(n19211) );
  IV U21453 ( .A(n19138), .Z(n19212) );
  XOR U21454 ( .A(n19213), .B(n19214), .Z(n19138) );
  ANDN U21455 ( .B(n19215), .A(n19216), .Z(n19213) );
  XOR U21456 ( .A(n19214), .B(n19217), .Z(n19215) );
  XOR U21457 ( .A(n19218), .B(n19146), .Z(n19158) );
  XOR U21458 ( .A(n19219), .B(n19220), .Z(n19146) );
  ANDN U21459 ( .B(n19221), .A(n19222), .Z(n19219) );
  XOR U21460 ( .A(n19220), .B(n19223), .Z(n19221) );
  IV U21461 ( .A(n19145), .Z(n19218) );
  XOR U21462 ( .A(n19224), .B(n19225), .Z(n19145) );
  XOR U21463 ( .A(n19226), .B(n19227), .Z(n19225) );
  ANDN U21464 ( .B(n19228), .A(n19229), .Z(n19226) );
  XOR U21465 ( .A(n19230), .B(n19227), .Z(n19228) );
  IV U21466 ( .A(n19143), .Z(n19224) );
  XOR U21467 ( .A(n19231), .B(n19232), .Z(n19143) );
  ANDN U21468 ( .B(n19233), .A(n19234), .Z(n19231) );
  XOR U21469 ( .A(n19232), .B(n19235), .Z(n19233) );
  IV U21470 ( .A(n19157), .Z(n19210) );
  XOR U21471 ( .A(n19236), .B(n19237), .Z(n19157) );
  XNOR U21472 ( .A(n19152), .B(n19238), .Z(n19237) );
  IV U21473 ( .A(n19155), .Z(n19238) );
  XOR U21474 ( .A(n19239), .B(n19240), .Z(n19155) );
  ANDN U21475 ( .B(n19241), .A(n19242), .Z(n19239) );
  XOR U21476 ( .A(n19243), .B(n19240), .Z(n19241) );
  XNOR U21477 ( .A(n19244), .B(n19245), .Z(n19152) );
  ANDN U21478 ( .B(n19246), .A(n19247), .Z(n19244) );
  XOR U21479 ( .A(n19245), .B(n19248), .Z(n19246) );
  IV U21480 ( .A(n19151), .Z(n19236) );
  XOR U21481 ( .A(n19149), .B(n19249), .Z(n19151) );
  XOR U21482 ( .A(n19250), .B(n19251), .Z(n19249) );
  ANDN U21483 ( .B(n19252), .A(n19253), .Z(n19250) );
  XOR U21484 ( .A(n19254), .B(n19251), .Z(n19252) );
  IV U21485 ( .A(n19153), .Z(n19149) );
  XOR U21486 ( .A(n19255), .B(n19256), .Z(n19153) );
  ANDN U21487 ( .B(n19257), .A(n19258), .Z(n19255) );
  XOR U21488 ( .A(n19259), .B(n19256), .Z(n19257) );
  IV U21489 ( .A(n19163), .Z(n19167) );
  XOR U21490 ( .A(n19163), .B(n19066), .Z(n19165) );
  XOR U21491 ( .A(n19260), .B(n19261), .Z(n19066) );
  AND U21492 ( .A(n152), .B(n19262), .Z(n19260) );
  XOR U21493 ( .A(n19263), .B(n19261), .Z(n19262) );
  NANDN U21494 ( .A(n19068), .B(n19070), .Z(n19163) );
  XOR U21495 ( .A(n19264), .B(n19265), .Z(n19070) );
  AND U21496 ( .A(n152), .B(n19266), .Z(n19264) );
  XOR U21497 ( .A(n19265), .B(n19267), .Z(n19266) );
  XNOR U21498 ( .A(n19268), .B(n19269), .Z(n152) );
  AND U21499 ( .A(n19270), .B(n19271), .Z(n19268) );
  XOR U21500 ( .A(n19269), .B(n19081), .Z(n19271) );
  XNOR U21501 ( .A(n19272), .B(n19273), .Z(n19081) );
  ANDN U21502 ( .B(n19274), .A(n19275), .Z(n19272) );
  XOR U21503 ( .A(n19273), .B(n19276), .Z(n19274) );
  XNOR U21504 ( .A(n19269), .B(n19083), .Z(n19270) );
  XOR U21505 ( .A(n19277), .B(n19278), .Z(n19083) );
  AND U21506 ( .A(n156), .B(n19279), .Z(n19277) );
  XOR U21507 ( .A(n19280), .B(n19278), .Z(n19279) );
  XOR U21508 ( .A(n19281), .B(n19282), .Z(n19269) );
  AND U21509 ( .A(n19283), .B(n19284), .Z(n19281) );
  XOR U21510 ( .A(n19282), .B(n19108), .Z(n19284) );
  XOR U21511 ( .A(n19275), .B(n19276), .Z(n19108) );
  XNOR U21512 ( .A(n19285), .B(n19286), .Z(n19276) );
  ANDN U21513 ( .B(n19287), .A(n19288), .Z(n19285) );
  XOR U21514 ( .A(n19289), .B(n19290), .Z(n19287) );
  XOR U21515 ( .A(n19291), .B(n19292), .Z(n19275) );
  XNOR U21516 ( .A(n19293), .B(n19294), .Z(n19292) );
  ANDN U21517 ( .B(n19295), .A(n19296), .Z(n19293) );
  XNOR U21518 ( .A(n19297), .B(n19298), .Z(n19295) );
  IV U21519 ( .A(n19273), .Z(n19291) );
  XOR U21520 ( .A(n19299), .B(n19300), .Z(n19273) );
  ANDN U21521 ( .B(n19301), .A(n19302), .Z(n19299) );
  XOR U21522 ( .A(n19300), .B(n19303), .Z(n19301) );
  XNOR U21523 ( .A(n19282), .B(n19110), .Z(n19283) );
  XOR U21524 ( .A(n19304), .B(n19305), .Z(n19110) );
  AND U21525 ( .A(n156), .B(n19306), .Z(n19304) );
  XOR U21526 ( .A(n19307), .B(n19305), .Z(n19306) );
  XNOR U21527 ( .A(n19308), .B(n19309), .Z(n19282) );
  AND U21528 ( .A(n19310), .B(n19311), .Z(n19308) );
  XNOR U21529 ( .A(n19309), .B(n19160), .Z(n19311) );
  XOR U21530 ( .A(n19302), .B(n19303), .Z(n19160) );
  XOR U21531 ( .A(n19312), .B(n19290), .Z(n19303) );
  XNOR U21532 ( .A(n19313), .B(n19314), .Z(n19290) );
  ANDN U21533 ( .B(n19315), .A(n19316), .Z(n19313) );
  XOR U21534 ( .A(n19317), .B(n19318), .Z(n19315) );
  IV U21535 ( .A(n19288), .Z(n19312) );
  XOR U21536 ( .A(n19286), .B(n19319), .Z(n19288) );
  XNOR U21537 ( .A(n19320), .B(n19321), .Z(n19319) );
  ANDN U21538 ( .B(n19322), .A(n19323), .Z(n19320) );
  XNOR U21539 ( .A(n19324), .B(n19325), .Z(n19322) );
  IV U21540 ( .A(n19289), .Z(n19286) );
  XOR U21541 ( .A(n19326), .B(n19327), .Z(n19289) );
  ANDN U21542 ( .B(n19328), .A(n19329), .Z(n19326) );
  XOR U21543 ( .A(n19327), .B(n19330), .Z(n19328) );
  XOR U21544 ( .A(n19331), .B(n19332), .Z(n19302) );
  XNOR U21545 ( .A(n19297), .B(n19333), .Z(n19332) );
  IV U21546 ( .A(n19300), .Z(n19333) );
  XOR U21547 ( .A(n19334), .B(n19335), .Z(n19300) );
  ANDN U21548 ( .B(n19336), .A(n19337), .Z(n19334) );
  XOR U21549 ( .A(n19335), .B(n19338), .Z(n19336) );
  XNOR U21550 ( .A(n19339), .B(n19340), .Z(n19297) );
  ANDN U21551 ( .B(n19341), .A(n19342), .Z(n19339) );
  XOR U21552 ( .A(n19340), .B(n19343), .Z(n19341) );
  IV U21553 ( .A(n19296), .Z(n19331) );
  XOR U21554 ( .A(n19294), .B(n19344), .Z(n19296) );
  XNOR U21555 ( .A(n19345), .B(n19346), .Z(n19344) );
  ANDN U21556 ( .B(n19347), .A(n19348), .Z(n19345) );
  XNOR U21557 ( .A(n19349), .B(n19350), .Z(n19347) );
  IV U21558 ( .A(n19298), .Z(n19294) );
  XOR U21559 ( .A(n19351), .B(n19352), .Z(n19298) );
  ANDN U21560 ( .B(n19353), .A(n19354), .Z(n19351) );
  XOR U21561 ( .A(n19355), .B(n19352), .Z(n19353) );
  XOR U21562 ( .A(n19309), .B(n19162), .Z(n19310) );
  XOR U21563 ( .A(n19356), .B(n19357), .Z(n19162) );
  AND U21564 ( .A(n156), .B(n19358), .Z(n19356) );
  XOR U21565 ( .A(n19359), .B(n19357), .Z(n19358) );
  XNOR U21566 ( .A(n19360), .B(n19361), .Z(n19309) );
  NAND U21567 ( .A(n19362), .B(n19363), .Z(n19361) );
  XOR U21568 ( .A(n19364), .B(n19261), .Z(n19363) );
  XOR U21569 ( .A(n19337), .B(n19338), .Z(n19261) );
  XOR U21570 ( .A(n19365), .B(n19330), .Z(n19338) );
  XOR U21571 ( .A(n19366), .B(n19318), .Z(n19330) );
  XOR U21572 ( .A(n19367), .B(n19368), .Z(n19318) );
  ANDN U21573 ( .B(n19369), .A(n19370), .Z(n19367) );
  XOR U21574 ( .A(n19368), .B(n19371), .Z(n19369) );
  IV U21575 ( .A(n19316), .Z(n19366) );
  XOR U21576 ( .A(n19314), .B(n19372), .Z(n19316) );
  XOR U21577 ( .A(n19373), .B(n19374), .Z(n19372) );
  ANDN U21578 ( .B(n19375), .A(n19376), .Z(n19373) );
  XOR U21579 ( .A(n19377), .B(n19374), .Z(n19375) );
  IV U21580 ( .A(n19317), .Z(n19314) );
  XOR U21581 ( .A(n19378), .B(n19379), .Z(n19317) );
  ANDN U21582 ( .B(n19380), .A(n19381), .Z(n19378) );
  XOR U21583 ( .A(n19379), .B(n19382), .Z(n19380) );
  IV U21584 ( .A(n19329), .Z(n19365) );
  XOR U21585 ( .A(n19383), .B(n19384), .Z(n19329) );
  XNOR U21586 ( .A(n19324), .B(n19385), .Z(n19384) );
  IV U21587 ( .A(n19327), .Z(n19385) );
  XOR U21588 ( .A(n19386), .B(n19387), .Z(n19327) );
  ANDN U21589 ( .B(n19388), .A(n19389), .Z(n19386) );
  XOR U21590 ( .A(n19387), .B(n19390), .Z(n19388) );
  XNOR U21591 ( .A(n19391), .B(n19392), .Z(n19324) );
  ANDN U21592 ( .B(n19393), .A(n19394), .Z(n19391) );
  XOR U21593 ( .A(n19392), .B(n19395), .Z(n19393) );
  IV U21594 ( .A(n19323), .Z(n19383) );
  XOR U21595 ( .A(n19321), .B(n19396), .Z(n19323) );
  XOR U21596 ( .A(n19397), .B(n19398), .Z(n19396) );
  ANDN U21597 ( .B(n19399), .A(n19400), .Z(n19397) );
  XOR U21598 ( .A(n19401), .B(n19398), .Z(n19399) );
  IV U21599 ( .A(n19325), .Z(n19321) );
  XOR U21600 ( .A(n19402), .B(n19403), .Z(n19325) );
  ANDN U21601 ( .B(n19404), .A(n19405), .Z(n19402) );
  XOR U21602 ( .A(n19406), .B(n19403), .Z(n19404) );
  XOR U21603 ( .A(n19407), .B(n19408), .Z(n19337) );
  XOR U21604 ( .A(n19355), .B(n19409), .Z(n19408) );
  IV U21605 ( .A(n19335), .Z(n19409) );
  XOR U21606 ( .A(n19410), .B(n19411), .Z(n19335) );
  ANDN U21607 ( .B(n19412), .A(n19413), .Z(n19410) );
  XOR U21608 ( .A(n19411), .B(n19414), .Z(n19412) );
  XOR U21609 ( .A(n19415), .B(n19343), .Z(n19355) );
  XOR U21610 ( .A(n19416), .B(n19417), .Z(n19343) );
  ANDN U21611 ( .B(n19418), .A(n19419), .Z(n19416) );
  XOR U21612 ( .A(n19417), .B(n19420), .Z(n19418) );
  IV U21613 ( .A(n19342), .Z(n19415) );
  XOR U21614 ( .A(n19421), .B(n19422), .Z(n19342) );
  XOR U21615 ( .A(n19423), .B(n19424), .Z(n19422) );
  ANDN U21616 ( .B(n19425), .A(n19426), .Z(n19423) );
  XOR U21617 ( .A(n19427), .B(n19424), .Z(n19425) );
  IV U21618 ( .A(n19340), .Z(n19421) );
  XOR U21619 ( .A(n19428), .B(n19429), .Z(n19340) );
  ANDN U21620 ( .B(n19430), .A(n19431), .Z(n19428) );
  XOR U21621 ( .A(n19429), .B(n19432), .Z(n19430) );
  IV U21622 ( .A(n19354), .Z(n19407) );
  XOR U21623 ( .A(n19433), .B(n19434), .Z(n19354) );
  XNOR U21624 ( .A(n19349), .B(n19435), .Z(n19434) );
  IV U21625 ( .A(n19352), .Z(n19435) );
  XOR U21626 ( .A(n19436), .B(n19437), .Z(n19352) );
  ANDN U21627 ( .B(n19438), .A(n19439), .Z(n19436) );
  XOR U21628 ( .A(n19440), .B(n19437), .Z(n19438) );
  XNOR U21629 ( .A(n19441), .B(n19442), .Z(n19349) );
  ANDN U21630 ( .B(n19443), .A(n19444), .Z(n19441) );
  XOR U21631 ( .A(n19442), .B(n19445), .Z(n19443) );
  IV U21632 ( .A(n19348), .Z(n19433) );
  XOR U21633 ( .A(n19346), .B(n19446), .Z(n19348) );
  XOR U21634 ( .A(n19447), .B(n19448), .Z(n19446) );
  ANDN U21635 ( .B(n19449), .A(n19450), .Z(n19447) );
  XOR U21636 ( .A(n19451), .B(n19448), .Z(n19449) );
  IV U21637 ( .A(n19350), .Z(n19346) );
  XOR U21638 ( .A(n19452), .B(n19453), .Z(n19350) );
  ANDN U21639 ( .B(n19454), .A(n19455), .Z(n19452) );
  XOR U21640 ( .A(n19456), .B(n19453), .Z(n19454) );
  IV U21641 ( .A(n19360), .Z(n19364) );
  XOR U21642 ( .A(n19360), .B(n19263), .Z(n19362) );
  XOR U21643 ( .A(n19457), .B(n19458), .Z(n19263) );
  AND U21644 ( .A(n156), .B(n19459), .Z(n19457) );
  XOR U21645 ( .A(n19460), .B(n19458), .Z(n19459) );
  NANDN U21646 ( .A(n19265), .B(n19267), .Z(n19360) );
  XOR U21647 ( .A(n19461), .B(n19462), .Z(n19267) );
  AND U21648 ( .A(n156), .B(n19463), .Z(n19461) );
  XOR U21649 ( .A(n19462), .B(n19464), .Z(n19463) );
  XNOR U21650 ( .A(n19465), .B(n19466), .Z(n156) );
  AND U21651 ( .A(n19467), .B(n19468), .Z(n19465) );
  XOR U21652 ( .A(n19466), .B(n19278), .Z(n19468) );
  XNOR U21653 ( .A(n19469), .B(n19470), .Z(n19278) );
  ANDN U21654 ( .B(n19471), .A(n19472), .Z(n19469) );
  XOR U21655 ( .A(n19470), .B(n19473), .Z(n19471) );
  XNOR U21656 ( .A(n19466), .B(n19280), .Z(n19467) );
  XOR U21657 ( .A(n19474), .B(n19475), .Z(n19280) );
  AND U21658 ( .A(n160), .B(n19476), .Z(n19474) );
  XOR U21659 ( .A(n19477), .B(n19475), .Z(n19476) );
  XOR U21660 ( .A(n19478), .B(n19479), .Z(n19466) );
  AND U21661 ( .A(n19480), .B(n19481), .Z(n19478) );
  XOR U21662 ( .A(n19479), .B(n19305), .Z(n19481) );
  XOR U21663 ( .A(n19472), .B(n19473), .Z(n19305) );
  XNOR U21664 ( .A(n19482), .B(n19483), .Z(n19473) );
  ANDN U21665 ( .B(n19484), .A(n19485), .Z(n19482) );
  XOR U21666 ( .A(n19486), .B(n19487), .Z(n19484) );
  XOR U21667 ( .A(n19488), .B(n19489), .Z(n19472) );
  XNOR U21668 ( .A(n19490), .B(n19491), .Z(n19489) );
  ANDN U21669 ( .B(n19492), .A(n19493), .Z(n19490) );
  XNOR U21670 ( .A(n19494), .B(n19495), .Z(n19492) );
  IV U21671 ( .A(n19470), .Z(n19488) );
  XOR U21672 ( .A(n19496), .B(n19497), .Z(n19470) );
  ANDN U21673 ( .B(n19498), .A(n19499), .Z(n19496) );
  XOR U21674 ( .A(n19497), .B(n19500), .Z(n19498) );
  XNOR U21675 ( .A(n19479), .B(n19307), .Z(n19480) );
  XOR U21676 ( .A(n19501), .B(n19502), .Z(n19307) );
  AND U21677 ( .A(n160), .B(n19503), .Z(n19501) );
  XOR U21678 ( .A(n19504), .B(n19502), .Z(n19503) );
  XNOR U21679 ( .A(n19505), .B(n19506), .Z(n19479) );
  AND U21680 ( .A(n19507), .B(n19508), .Z(n19505) );
  XNOR U21681 ( .A(n19506), .B(n19357), .Z(n19508) );
  XOR U21682 ( .A(n19499), .B(n19500), .Z(n19357) );
  XOR U21683 ( .A(n19509), .B(n19487), .Z(n19500) );
  XNOR U21684 ( .A(n19510), .B(n19511), .Z(n19487) );
  ANDN U21685 ( .B(n19512), .A(n19513), .Z(n19510) );
  XOR U21686 ( .A(n19514), .B(n19515), .Z(n19512) );
  IV U21687 ( .A(n19485), .Z(n19509) );
  XOR U21688 ( .A(n19483), .B(n19516), .Z(n19485) );
  XNOR U21689 ( .A(n19517), .B(n19518), .Z(n19516) );
  ANDN U21690 ( .B(n19519), .A(n19520), .Z(n19517) );
  XNOR U21691 ( .A(n19521), .B(n19522), .Z(n19519) );
  IV U21692 ( .A(n19486), .Z(n19483) );
  XOR U21693 ( .A(n19523), .B(n19524), .Z(n19486) );
  ANDN U21694 ( .B(n19525), .A(n19526), .Z(n19523) );
  XOR U21695 ( .A(n19524), .B(n19527), .Z(n19525) );
  XOR U21696 ( .A(n19528), .B(n19529), .Z(n19499) );
  XNOR U21697 ( .A(n19494), .B(n19530), .Z(n19529) );
  IV U21698 ( .A(n19497), .Z(n19530) );
  XOR U21699 ( .A(n19531), .B(n19532), .Z(n19497) );
  ANDN U21700 ( .B(n19533), .A(n19534), .Z(n19531) );
  XOR U21701 ( .A(n19532), .B(n19535), .Z(n19533) );
  XNOR U21702 ( .A(n19536), .B(n19537), .Z(n19494) );
  ANDN U21703 ( .B(n19538), .A(n19539), .Z(n19536) );
  XOR U21704 ( .A(n19537), .B(n19540), .Z(n19538) );
  IV U21705 ( .A(n19493), .Z(n19528) );
  XOR U21706 ( .A(n19491), .B(n19541), .Z(n19493) );
  XNOR U21707 ( .A(n19542), .B(n19543), .Z(n19541) );
  ANDN U21708 ( .B(n19544), .A(n19545), .Z(n19542) );
  XNOR U21709 ( .A(n19546), .B(n19547), .Z(n19544) );
  IV U21710 ( .A(n19495), .Z(n19491) );
  XOR U21711 ( .A(n19548), .B(n19549), .Z(n19495) );
  ANDN U21712 ( .B(n19550), .A(n19551), .Z(n19548) );
  XOR U21713 ( .A(n19552), .B(n19549), .Z(n19550) );
  XOR U21714 ( .A(n19506), .B(n19359), .Z(n19507) );
  XOR U21715 ( .A(n19553), .B(n19554), .Z(n19359) );
  AND U21716 ( .A(n160), .B(n19555), .Z(n19553) );
  XOR U21717 ( .A(n19556), .B(n19554), .Z(n19555) );
  XNOR U21718 ( .A(n19557), .B(n19558), .Z(n19506) );
  NAND U21719 ( .A(n19559), .B(n19560), .Z(n19558) );
  XOR U21720 ( .A(n19561), .B(n19458), .Z(n19560) );
  XOR U21721 ( .A(n19534), .B(n19535), .Z(n19458) );
  XOR U21722 ( .A(n19562), .B(n19527), .Z(n19535) );
  XOR U21723 ( .A(n19563), .B(n19515), .Z(n19527) );
  XOR U21724 ( .A(n19564), .B(n19565), .Z(n19515) );
  ANDN U21725 ( .B(n19566), .A(n19567), .Z(n19564) );
  XOR U21726 ( .A(n19565), .B(n19568), .Z(n19566) );
  IV U21727 ( .A(n19513), .Z(n19563) );
  XOR U21728 ( .A(n19511), .B(n19569), .Z(n19513) );
  XOR U21729 ( .A(n19570), .B(n19571), .Z(n19569) );
  ANDN U21730 ( .B(n19572), .A(n19573), .Z(n19570) );
  XOR U21731 ( .A(n19574), .B(n19571), .Z(n19572) );
  IV U21732 ( .A(n19514), .Z(n19511) );
  XOR U21733 ( .A(n19575), .B(n19576), .Z(n19514) );
  ANDN U21734 ( .B(n19577), .A(n19578), .Z(n19575) );
  XOR U21735 ( .A(n19576), .B(n19579), .Z(n19577) );
  IV U21736 ( .A(n19526), .Z(n19562) );
  XOR U21737 ( .A(n19580), .B(n19581), .Z(n19526) );
  XNOR U21738 ( .A(n19521), .B(n19582), .Z(n19581) );
  IV U21739 ( .A(n19524), .Z(n19582) );
  XOR U21740 ( .A(n19583), .B(n19584), .Z(n19524) );
  ANDN U21741 ( .B(n19585), .A(n19586), .Z(n19583) );
  XOR U21742 ( .A(n19584), .B(n19587), .Z(n19585) );
  XNOR U21743 ( .A(n19588), .B(n19589), .Z(n19521) );
  ANDN U21744 ( .B(n19590), .A(n19591), .Z(n19588) );
  XOR U21745 ( .A(n19589), .B(n19592), .Z(n19590) );
  IV U21746 ( .A(n19520), .Z(n19580) );
  XOR U21747 ( .A(n19518), .B(n19593), .Z(n19520) );
  XOR U21748 ( .A(n19594), .B(n19595), .Z(n19593) );
  ANDN U21749 ( .B(n19596), .A(n19597), .Z(n19594) );
  XOR U21750 ( .A(n19598), .B(n19595), .Z(n19596) );
  IV U21751 ( .A(n19522), .Z(n19518) );
  XOR U21752 ( .A(n19599), .B(n19600), .Z(n19522) );
  ANDN U21753 ( .B(n19601), .A(n19602), .Z(n19599) );
  XOR U21754 ( .A(n19603), .B(n19600), .Z(n19601) );
  XOR U21755 ( .A(n19604), .B(n19605), .Z(n19534) );
  XOR U21756 ( .A(n19552), .B(n19606), .Z(n19605) );
  IV U21757 ( .A(n19532), .Z(n19606) );
  XOR U21758 ( .A(n19607), .B(n19608), .Z(n19532) );
  ANDN U21759 ( .B(n19609), .A(n19610), .Z(n19607) );
  XOR U21760 ( .A(n19608), .B(n19611), .Z(n19609) );
  XOR U21761 ( .A(n19612), .B(n19540), .Z(n19552) );
  XOR U21762 ( .A(n19613), .B(n19614), .Z(n19540) );
  ANDN U21763 ( .B(n19615), .A(n19616), .Z(n19613) );
  XOR U21764 ( .A(n19614), .B(n19617), .Z(n19615) );
  IV U21765 ( .A(n19539), .Z(n19612) );
  XOR U21766 ( .A(n19618), .B(n19619), .Z(n19539) );
  XOR U21767 ( .A(n19620), .B(n19621), .Z(n19619) );
  ANDN U21768 ( .B(n19622), .A(n19623), .Z(n19620) );
  XOR U21769 ( .A(n19624), .B(n19621), .Z(n19622) );
  IV U21770 ( .A(n19537), .Z(n19618) );
  XOR U21771 ( .A(n19625), .B(n19626), .Z(n19537) );
  ANDN U21772 ( .B(n19627), .A(n19628), .Z(n19625) );
  XOR U21773 ( .A(n19626), .B(n19629), .Z(n19627) );
  IV U21774 ( .A(n19551), .Z(n19604) );
  XOR U21775 ( .A(n19630), .B(n19631), .Z(n19551) );
  XNOR U21776 ( .A(n19546), .B(n19632), .Z(n19631) );
  IV U21777 ( .A(n19549), .Z(n19632) );
  XOR U21778 ( .A(n19633), .B(n19634), .Z(n19549) );
  ANDN U21779 ( .B(n19635), .A(n19636), .Z(n19633) );
  XOR U21780 ( .A(n19637), .B(n19634), .Z(n19635) );
  XNOR U21781 ( .A(n19638), .B(n19639), .Z(n19546) );
  ANDN U21782 ( .B(n19640), .A(n19641), .Z(n19638) );
  XOR U21783 ( .A(n19639), .B(n19642), .Z(n19640) );
  IV U21784 ( .A(n19545), .Z(n19630) );
  XOR U21785 ( .A(n19543), .B(n19643), .Z(n19545) );
  XOR U21786 ( .A(n19644), .B(n19645), .Z(n19643) );
  ANDN U21787 ( .B(n19646), .A(n19647), .Z(n19644) );
  XOR U21788 ( .A(n19648), .B(n19645), .Z(n19646) );
  IV U21789 ( .A(n19547), .Z(n19543) );
  XOR U21790 ( .A(n19649), .B(n19650), .Z(n19547) );
  ANDN U21791 ( .B(n19651), .A(n19652), .Z(n19649) );
  XOR U21792 ( .A(n19653), .B(n19650), .Z(n19651) );
  IV U21793 ( .A(n19557), .Z(n19561) );
  XOR U21794 ( .A(n19557), .B(n19460), .Z(n19559) );
  XOR U21795 ( .A(n19654), .B(n19655), .Z(n19460) );
  AND U21796 ( .A(n160), .B(n19656), .Z(n19654) );
  XOR U21797 ( .A(n19657), .B(n19655), .Z(n19656) );
  NANDN U21798 ( .A(n19462), .B(n19464), .Z(n19557) );
  XOR U21799 ( .A(n19658), .B(n19659), .Z(n19464) );
  AND U21800 ( .A(n160), .B(n19660), .Z(n19658) );
  XOR U21801 ( .A(n19659), .B(n19661), .Z(n19660) );
  XNOR U21802 ( .A(n19662), .B(n19663), .Z(n160) );
  AND U21803 ( .A(n19664), .B(n19665), .Z(n19662) );
  XOR U21804 ( .A(n19663), .B(n19475), .Z(n19665) );
  XNOR U21805 ( .A(n19666), .B(n19667), .Z(n19475) );
  ANDN U21806 ( .B(n19668), .A(n19669), .Z(n19666) );
  XOR U21807 ( .A(n19667), .B(n19670), .Z(n19668) );
  XNOR U21808 ( .A(n19663), .B(n19477), .Z(n19664) );
  XOR U21809 ( .A(n19671), .B(n19672), .Z(n19477) );
  AND U21810 ( .A(n164), .B(n19673), .Z(n19671) );
  XOR U21811 ( .A(n19674), .B(n19672), .Z(n19673) );
  XOR U21812 ( .A(n19675), .B(n19676), .Z(n19663) );
  AND U21813 ( .A(n19677), .B(n19678), .Z(n19675) );
  XOR U21814 ( .A(n19676), .B(n19502), .Z(n19678) );
  XOR U21815 ( .A(n19669), .B(n19670), .Z(n19502) );
  XNOR U21816 ( .A(n19679), .B(n19680), .Z(n19670) );
  ANDN U21817 ( .B(n19681), .A(n19682), .Z(n19679) );
  XOR U21818 ( .A(n19683), .B(n19684), .Z(n19681) );
  XOR U21819 ( .A(n19685), .B(n19686), .Z(n19669) );
  XNOR U21820 ( .A(n19687), .B(n19688), .Z(n19686) );
  ANDN U21821 ( .B(n19689), .A(n19690), .Z(n19687) );
  XNOR U21822 ( .A(n19691), .B(n19692), .Z(n19689) );
  IV U21823 ( .A(n19667), .Z(n19685) );
  XOR U21824 ( .A(n19693), .B(n19694), .Z(n19667) );
  ANDN U21825 ( .B(n19695), .A(n19696), .Z(n19693) );
  XOR U21826 ( .A(n19694), .B(n19697), .Z(n19695) );
  XNOR U21827 ( .A(n19676), .B(n19504), .Z(n19677) );
  XOR U21828 ( .A(n19698), .B(n19699), .Z(n19504) );
  AND U21829 ( .A(n164), .B(n19700), .Z(n19698) );
  XOR U21830 ( .A(n19701), .B(n19699), .Z(n19700) );
  XNOR U21831 ( .A(n19702), .B(n19703), .Z(n19676) );
  AND U21832 ( .A(n19704), .B(n19705), .Z(n19702) );
  XNOR U21833 ( .A(n19703), .B(n19554), .Z(n19705) );
  XOR U21834 ( .A(n19696), .B(n19697), .Z(n19554) );
  XOR U21835 ( .A(n19706), .B(n19684), .Z(n19697) );
  XNOR U21836 ( .A(n19707), .B(n19708), .Z(n19684) );
  ANDN U21837 ( .B(n19709), .A(n19710), .Z(n19707) );
  XOR U21838 ( .A(n19711), .B(n19712), .Z(n19709) );
  IV U21839 ( .A(n19682), .Z(n19706) );
  XOR U21840 ( .A(n19680), .B(n19713), .Z(n19682) );
  XNOR U21841 ( .A(n19714), .B(n19715), .Z(n19713) );
  ANDN U21842 ( .B(n19716), .A(n19717), .Z(n19714) );
  XNOR U21843 ( .A(n19718), .B(n19719), .Z(n19716) );
  IV U21844 ( .A(n19683), .Z(n19680) );
  XOR U21845 ( .A(n19720), .B(n19721), .Z(n19683) );
  ANDN U21846 ( .B(n19722), .A(n19723), .Z(n19720) );
  XOR U21847 ( .A(n19721), .B(n19724), .Z(n19722) );
  XOR U21848 ( .A(n19725), .B(n19726), .Z(n19696) );
  XNOR U21849 ( .A(n19691), .B(n19727), .Z(n19726) );
  IV U21850 ( .A(n19694), .Z(n19727) );
  XOR U21851 ( .A(n19728), .B(n19729), .Z(n19694) );
  ANDN U21852 ( .B(n19730), .A(n19731), .Z(n19728) );
  XOR U21853 ( .A(n19729), .B(n19732), .Z(n19730) );
  XNOR U21854 ( .A(n19733), .B(n19734), .Z(n19691) );
  ANDN U21855 ( .B(n19735), .A(n19736), .Z(n19733) );
  XOR U21856 ( .A(n19734), .B(n19737), .Z(n19735) );
  IV U21857 ( .A(n19690), .Z(n19725) );
  XOR U21858 ( .A(n19688), .B(n19738), .Z(n19690) );
  XNOR U21859 ( .A(n19739), .B(n19740), .Z(n19738) );
  ANDN U21860 ( .B(n19741), .A(n19742), .Z(n19739) );
  XNOR U21861 ( .A(n19743), .B(n19744), .Z(n19741) );
  IV U21862 ( .A(n19692), .Z(n19688) );
  XOR U21863 ( .A(n19745), .B(n19746), .Z(n19692) );
  ANDN U21864 ( .B(n19747), .A(n19748), .Z(n19745) );
  XOR U21865 ( .A(n19749), .B(n19746), .Z(n19747) );
  XOR U21866 ( .A(n19703), .B(n19556), .Z(n19704) );
  XOR U21867 ( .A(n19750), .B(n19751), .Z(n19556) );
  AND U21868 ( .A(n164), .B(n19752), .Z(n19750) );
  XOR U21869 ( .A(n19753), .B(n19751), .Z(n19752) );
  XNOR U21870 ( .A(n19754), .B(n19755), .Z(n19703) );
  NAND U21871 ( .A(n19756), .B(n19757), .Z(n19755) );
  XOR U21872 ( .A(n19758), .B(n19655), .Z(n19757) );
  XOR U21873 ( .A(n19731), .B(n19732), .Z(n19655) );
  XOR U21874 ( .A(n19759), .B(n19724), .Z(n19732) );
  XOR U21875 ( .A(n19760), .B(n19712), .Z(n19724) );
  XOR U21876 ( .A(n19761), .B(n19762), .Z(n19712) );
  ANDN U21877 ( .B(n19763), .A(n19764), .Z(n19761) );
  XOR U21878 ( .A(n19762), .B(n19765), .Z(n19763) );
  IV U21879 ( .A(n19710), .Z(n19760) );
  XOR U21880 ( .A(n19708), .B(n19766), .Z(n19710) );
  XOR U21881 ( .A(n19767), .B(n19768), .Z(n19766) );
  ANDN U21882 ( .B(n19769), .A(n19770), .Z(n19767) );
  XOR U21883 ( .A(n19771), .B(n19768), .Z(n19769) );
  IV U21884 ( .A(n19711), .Z(n19708) );
  XOR U21885 ( .A(n19772), .B(n19773), .Z(n19711) );
  ANDN U21886 ( .B(n19774), .A(n19775), .Z(n19772) );
  XOR U21887 ( .A(n19773), .B(n19776), .Z(n19774) );
  IV U21888 ( .A(n19723), .Z(n19759) );
  XOR U21889 ( .A(n19777), .B(n19778), .Z(n19723) );
  XNOR U21890 ( .A(n19718), .B(n19779), .Z(n19778) );
  IV U21891 ( .A(n19721), .Z(n19779) );
  XOR U21892 ( .A(n19780), .B(n19781), .Z(n19721) );
  ANDN U21893 ( .B(n19782), .A(n19783), .Z(n19780) );
  XOR U21894 ( .A(n19781), .B(n19784), .Z(n19782) );
  XNOR U21895 ( .A(n19785), .B(n19786), .Z(n19718) );
  ANDN U21896 ( .B(n19787), .A(n19788), .Z(n19785) );
  XOR U21897 ( .A(n19786), .B(n19789), .Z(n19787) );
  IV U21898 ( .A(n19717), .Z(n19777) );
  XOR U21899 ( .A(n19715), .B(n19790), .Z(n19717) );
  XOR U21900 ( .A(n19791), .B(n19792), .Z(n19790) );
  ANDN U21901 ( .B(n19793), .A(n19794), .Z(n19791) );
  XOR U21902 ( .A(n19795), .B(n19792), .Z(n19793) );
  IV U21903 ( .A(n19719), .Z(n19715) );
  XOR U21904 ( .A(n19796), .B(n19797), .Z(n19719) );
  ANDN U21905 ( .B(n19798), .A(n19799), .Z(n19796) );
  XOR U21906 ( .A(n19800), .B(n19797), .Z(n19798) );
  XOR U21907 ( .A(n19801), .B(n19802), .Z(n19731) );
  XOR U21908 ( .A(n19749), .B(n19803), .Z(n19802) );
  IV U21909 ( .A(n19729), .Z(n19803) );
  XOR U21910 ( .A(n19804), .B(n19805), .Z(n19729) );
  ANDN U21911 ( .B(n19806), .A(n19807), .Z(n19804) );
  XOR U21912 ( .A(n19805), .B(n19808), .Z(n19806) );
  XOR U21913 ( .A(n19809), .B(n19737), .Z(n19749) );
  XOR U21914 ( .A(n19810), .B(n19811), .Z(n19737) );
  ANDN U21915 ( .B(n19812), .A(n19813), .Z(n19810) );
  XOR U21916 ( .A(n19811), .B(n19814), .Z(n19812) );
  IV U21917 ( .A(n19736), .Z(n19809) );
  XOR U21918 ( .A(n19815), .B(n19816), .Z(n19736) );
  XOR U21919 ( .A(n19817), .B(n19818), .Z(n19816) );
  ANDN U21920 ( .B(n19819), .A(n19820), .Z(n19817) );
  XOR U21921 ( .A(n19821), .B(n19818), .Z(n19819) );
  IV U21922 ( .A(n19734), .Z(n19815) );
  XOR U21923 ( .A(n19822), .B(n19823), .Z(n19734) );
  ANDN U21924 ( .B(n19824), .A(n19825), .Z(n19822) );
  XOR U21925 ( .A(n19823), .B(n19826), .Z(n19824) );
  IV U21926 ( .A(n19748), .Z(n19801) );
  XOR U21927 ( .A(n19827), .B(n19828), .Z(n19748) );
  XNOR U21928 ( .A(n19743), .B(n19829), .Z(n19828) );
  IV U21929 ( .A(n19746), .Z(n19829) );
  XOR U21930 ( .A(n19830), .B(n19831), .Z(n19746) );
  ANDN U21931 ( .B(n19832), .A(n19833), .Z(n19830) );
  XOR U21932 ( .A(n19834), .B(n19831), .Z(n19832) );
  XNOR U21933 ( .A(n19835), .B(n19836), .Z(n19743) );
  ANDN U21934 ( .B(n19837), .A(n19838), .Z(n19835) );
  XOR U21935 ( .A(n19836), .B(n19839), .Z(n19837) );
  IV U21936 ( .A(n19742), .Z(n19827) );
  XOR U21937 ( .A(n19740), .B(n19840), .Z(n19742) );
  XOR U21938 ( .A(n19841), .B(n19842), .Z(n19840) );
  ANDN U21939 ( .B(n19843), .A(n19844), .Z(n19841) );
  XOR U21940 ( .A(n19845), .B(n19842), .Z(n19843) );
  IV U21941 ( .A(n19744), .Z(n19740) );
  XOR U21942 ( .A(n19846), .B(n19847), .Z(n19744) );
  ANDN U21943 ( .B(n19848), .A(n19849), .Z(n19846) );
  XOR U21944 ( .A(n19850), .B(n19847), .Z(n19848) );
  IV U21945 ( .A(n19754), .Z(n19758) );
  XOR U21946 ( .A(n19754), .B(n19657), .Z(n19756) );
  XOR U21947 ( .A(n19851), .B(n19852), .Z(n19657) );
  AND U21948 ( .A(n164), .B(n19853), .Z(n19851) );
  XOR U21949 ( .A(n19854), .B(n19852), .Z(n19853) );
  NANDN U21950 ( .A(n19659), .B(n19661), .Z(n19754) );
  XOR U21951 ( .A(n19855), .B(n19856), .Z(n19661) );
  AND U21952 ( .A(n164), .B(n19857), .Z(n19855) );
  XOR U21953 ( .A(n19856), .B(n19858), .Z(n19857) );
  XNOR U21954 ( .A(n19859), .B(n19860), .Z(n164) );
  AND U21955 ( .A(n19861), .B(n19862), .Z(n19859) );
  XOR U21956 ( .A(n19860), .B(n19672), .Z(n19862) );
  XNOR U21957 ( .A(n19863), .B(n19864), .Z(n19672) );
  ANDN U21958 ( .B(n19865), .A(n19866), .Z(n19863) );
  XOR U21959 ( .A(n19864), .B(n19867), .Z(n19865) );
  XNOR U21960 ( .A(n19860), .B(n19674), .Z(n19861) );
  XOR U21961 ( .A(n19868), .B(n19869), .Z(n19674) );
  AND U21962 ( .A(n168), .B(n19870), .Z(n19868) );
  XOR U21963 ( .A(n19871), .B(n19869), .Z(n19870) );
  XOR U21964 ( .A(n19872), .B(n19873), .Z(n19860) );
  AND U21965 ( .A(n19874), .B(n19875), .Z(n19872) );
  XOR U21966 ( .A(n19873), .B(n19699), .Z(n19875) );
  XOR U21967 ( .A(n19866), .B(n19867), .Z(n19699) );
  XNOR U21968 ( .A(n19876), .B(n19877), .Z(n19867) );
  ANDN U21969 ( .B(n19878), .A(n19879), .Z(n19876) );
  XOR U21970 ( .A(n19880), .B(n19881), .Z(n19878) );
  XOR U21971 ( .A(n19882), .B(n19883), .Z(n19866) );
  XNOR U21972 ( .A(n19884), .B(n19885), .Z(n19883) );
  ANDN U21973 ( .B(n19886), .A(n19887), .Z(n19884) );
  XNOR U21974 ( .A(n19888), .B(n19889), .Z(n19886) );
  IV U21975 ( .A(n19864), .Z(n19882) );
  XOR U21976 ( .A(n19890), .B(n19891), .Z(n19864) );
  ANDN U21977 ( .B(n19892), .A(n19893), .Z(n19890) );
  XOR U21978 ( .A(n19891), .B(n19894), .Z(n19892) );
  XNOR U21979 ( .A(n19873), .B(n19701), .Z(n19874) );
  XOR U21980 ( .A(n19895), .B(n19896), .Z(n19701) );
  AND U21981 ( .A(n168), .B(n19897), .Z(n19895) );
  XOR U21982 ( .A(n19898), .B(n19896), .Z(n19897) );
  XNOR U21983 ( .A(n19899), .B(n19900), .Z(n19873) );
  AND U21984 ( .A(n19901), .B(n19902), .Z(n19899) );
  XNOR U21985 ( .A(n19900), .B(n19751), .Z(n19902) );
  XOR U21986 ( .A(n19893), .B(n19894), .Z(n19751) );
  XOR U21987 ( .A(n19903), .B(n19881), .Z(n19894) );
  XNOR U21988 ( .A(n19904), .B(n19905), .Z(n19881) );
  ANDN U21989 ( .B(n19906), .A(n19907), .Z(n19904) );
  XOR U21990 ( .A(n19908), .B(n19909), .Z(n19906) );
  IV U21991 ( .A(n19879), .Z(n19903) );
  XOR U21992 ( .A(n19877), .B(n19910), .Z(n19879) );
  XNOR U21993 ( .A(n19911), .B(n19912), .Z(n19910) );
  ANDN U21994 ( .B(n19913), .A(n19914), .Z(n19911) );
  XNOR U21995 ( .A(n19915), .B(n19916), .Z(n19913) );
  IV U21996 ( .A(n19880), .Z(n19877) );
  XOR U21997 ( .A(n19917), .B(n19918), .Z(n19880) );
  ANDN U21998 ( .B(n19919), .A(n19920), .Z(n19917) );
  XOR U21999 ( .A(n19918), .B(n19921), .Z(n19919) );
  XOR U22000 ( .A(n19922), .B(n19923), .Z(n19893) );
  XNOR U22001 ( .A(n19888), .B(n19924), .Z(n19923) );
  IV U22002 ( .A(n19891), .Z(n19924) );
  XOR U22003 ( .A(n19925), .B(n19926), .Z(n19891) );
  ANDN U22004 ( .B(n19927), .A(n19928), .Z(n19925) );
  XOR U22005 ( .A(n19926), .B(n19929), .Z(n19927) );
  XNOR U22006 ( .A(n19930), .B(n19931), .Z(n19888) );
  ANDN U22007 ( .B(n19932), .A(n19933), .Z(n19930) );
  XOR U22008 ( .A(n19931), .B(n19934), .Z(n19932) );
  IV U22009 ( .A(n19887), .Z(n19922) );
  XOR U22010 ( .A(n19885), .B(n19935), .Z(n19887) );
  XNOR U22011 ( .A(n19936), .B(n19937), .Z(n19935) );
  ANDN U22012 ( .B(n19938), .A(n19939), .Z(n19936) );
  XNOR U22013 ( .A(n19940), .B(n19941), .Z(n19938) );
  IV U22014 ( .A(n19889), .Z(n19885) );
  XOR U22015 ( .A(n19942), .B(n19943), .Z(n19889) );
  ANDN U22016 ( .B(n19944), .A(n19945), .Z(n19942) );
  XOR U22017 ( .A(n19946), .B(n19943), .Z(n19944) );
  XOR U22018 ( .A(n19900), .B(n19753), .Z(n19901) );
  XOR U22019 ( .A(n19947), .B(n19948), .Z(n19753) );
  AND U22020 ( .A(n168), .B(n19949), .Z(n19947) );
  XOR U22021 ( .A(n19950), .B(n19948), .Z(n19949) );
  XNOR U22022 ( .A(n19951), .B(n19952), .Z(n19900) );
  NAND U22023 ( .A(n19953), .B(n19954), .Z(n19952) );
  XOR U22024 ( .A(n19955), .B(n19852), .Z(n19954) );
  XOR U22025 ( .A(n19928), .B(n19929), .Z(n19852) );
  XOR U22026 ( .A(n19956), .B(n19921), .Z(n19929) );
  XOR U22027 ( .A(n19957), .B(n19909), .Z(n19921) );
  XOR U22028 ( .A(n19958), .B(n19959), .Z(n19909) );
  ANDN U22029 ( .B(n19960), .A(n19961), .Z(n19958) );
  XOR U22030 ( .A(n19959), .B(n19962), .Z(n19960) );
  IV U22031 ( .A(n19907), .Z(n19957) );
  XOR U22032 ( .A(n19905), .B(n19963), .Z(n19907) );
  XOR U22033 ( .A(n19964), .B(n19965), .Z(n19963) );
  ANDN U22034 ( .B(n19966), .A(n19967), .Z(n19964) );
  XOR U22035 ( .A(n19968), .B(n19965), .Z(n19966) );
  IV U22036 ( .A(n19908), .Z(n19905) );
  XOR U22037 ( .A(n19969), .B(n19970), .Z(n19908) );
  ANDN U22038 ( .B(n19971), .A(n19972), .Z(n19969) );
  XOR U22039 ( .A(n19970), .B(n19973), .Z(n19971) );
  IV U22040 ( .A(n19920), .Z(n19956) );
  XOR U22041 ( .A(n19974), .B(n19975), .Z(n19920) );
  XNOR U22042 ( .A(n19915), .B(n19976), .Z(n19975) );
  IV U22043 ( .A(n19918), .Z(n19976) );
  XOR U22044 ( .A(n19977), .B(n19978), .Z(n19918) );
  ANDN U22045 ( .B(n19979), .A(n19980), .Z(n19977) );
  XOR U22046 ( .A(n19978), .B(n19981), .Z(n19979) );
  XNOR U22047 ( .A(n19982), .B(n19983), .Z(n19915) );
  ANDN U22048 ( .B(n19984), .A(n19985), .Z(n19982) );
  XOR U22049 ( .A(n19983), .B(n19986), .Z(n19984) );
  IV U22050 ( .A(n19914), .Z(n19974) );
  XOR U22051 ( .A(n19912), .B(n19987), .Z(n19914) );
  XOR U22052 ( .A(n19988), .B(n19989), .Z(n19987) );
  ANDN U22053 ( .B(n19990), .A(n19991), .Z(n19988) );
  XOR U22054 ( .A(n19992), .B(n19989), .Z(n19990) );
  IV U22055 ( .A(n19916), .Z(n19912) );
  XOR U22056 ( .A(n19993), .B(n19994), .Z(n19916) );
  ANDN U22057 ( .B(n19995), .A(n19996), .Z(n19993) );
  XOR U22058 ( .A(n19997), .B(n19994), .Z(n19995) );
  XOR U22059 ( .A(n19998), .B(n19999), .Z(n19928) );
  XOR U22060 ( .A(n19946), .B(n20000), .Z(n19999) );
  IV U22061 ( .A(n19926), .Z(n20000) );
  XOR U22062 ( .A(n20001), .B(n20002), .Z(n19926) );
  ANDN U22063 ( .B(n20003), .A(n20004), .Z(n20001) );
  XOR U22064 ( .A(n20002), .B(n20005), .Z(n20003) );
  XOR U22065 ( .A(n20006), .B(n19934), .Z(n19946) );
  XOR U22066 ( .A(n20007), .B(n20008), .Z(n19934) );
  ANDN U22067 ( .B(n20009), .A(n20010), .Z(n20007) );
  XOR U22068 ( .A(n20008), .B(n20011), .Z(n20009) );
  IV U22069 ( .A(n19933), .Z(n20006) );
  XOR U22070 ( .A(n20012), .B(n20013), .Z(n19933) );
  XOR U22071 ( .A(n20014), .B(n20015), .Z(n20013) );
  ANDN U22072 ( .B(n20016), .A(n20017), .Z(n20014) );
  XOR U22073 ( .A(n20018), .B(n20015), .Z(n20016) );
  IV U22074 ( .A(n19931), .Z(n20012) );
  XOR U22075 ( .A(n20019), .B(n20020), .Z(n19931) );
  ANDN U22076 ( .B(n20021), .A(n20022), .Z(n20019) );
  XOR U22077 ( .A(n20020), .B(n20023), .Z(n20021) );
  IV U22078 ( .A(n19945), .Z(n19998) );
  XOR U22079 ( .A(n20024), .B(n20025), .Z(n19945) );
  XNOR U22080 ( .A(n19940), .B(n20026), .Z(n20025) );
  IV U22081 ( .A(n19943), .Z(n20026) );
  XOR U22082 ( .A(n20027), .B(n20028), .Z(n19943) );
  ANDN U22083 ( .B(n20029), .A(n20030), .Z(n20027) );
  XOR U22084 ( .A(n20031), .B(n20028), .Z(n20029) );
  XNOR U22085 ( .A(n20032), .B(n20033), .Z(n19940) );
  ANDN U22086 ( .B(n20034), .A(n20035), .Z(n20032) );
  XOR U22087 ( .A(n20033), .B(n20036), .Z(n20034) );
  IV U22088 ( .A(n19939), .Z(n20024) );
  XOR U22089 ( .A(n19937), .B(n20037), .Z(n19939) );
  XOR U22090 ( .A(n20038), .B(n20039), .Z(n20037) );
  ANDN U22091 ( .B(n20040), .A(n20041), .Z(n20038) );
  XOR U22092 ( .A(n20042), .B(n20039), .Z(n20040) );
  IV U22093 ( .A(n19941), .Z(n19937) );
  XOR U22094 ( .A(n20043), .B(n20044), .Z(n19941) );
  ANDN U22095 ( .B(n20045), .A(n20046), .Z(n20043) );
  XOR U22096 ( .A(n20047), .B(n20044), .Z(n20045) );
  IV U22097 ( .A(n19951), .Z(n19955) );
  XOR U22098 ( .A(n19951), .B(n19854), .Z(n19953) );
  XOR U22099 ( .A(n20048), .B(n20049), .Z(n19854) );
  AND U22100 ( .A(n168), .B(n20050), .Z(n20048) );
  XOR U22101 ( .A(n20051), .B(n20049), .Z(n20050) );
  NANDN U22102 ( .A(n19856), .B(n19858), .Z(n19951) );
  XOR U22103 ( .A(n20052), .B(n20053), .Z(n19858) );
  AND U22104 ( .A(n168), .B(n20054), .Z(n20052) );
  XOR U22105 ( .A(n20053), .B(n20055), .Z(n20054) );
  XNOR U22106 ( .A(n20056), .B(n20057), .Z(n168) );
  AND U22107 ( .A(n20058), .B(n20059), .Z(n20056) );
  XOR U22108 ( .A(n20057), .B(n19869), .Z(n20059) );
  XNOR U22109 ( .A(n20060), .B(n20061), .Z(n19869) );
  ANDN U22110 ( .B(n20062), .A(n20063), .Z(n20060) );
  XOR U22111 ( .A(n20061), .B(n20064), .Z(n20062) );
  XNOR U22112 ( .A(n20057), .B(n19871), .Z(n20058) );
  XOR U22113 ( .A(n20065), .B(n20066), .Z(n19871) );
  AND U22114 ( .A(n172), .B(n20067), .Z(n20065) );
  XOR U22115 ( .A(n20068), .B(n20066), .Z(n20067) );
  XOR U22116 ( .A(n20069), .B(n20070), .Z(n20057) );
  AND U22117 ( .A(n20071), .B(n20072), .Z(n20069) );
  XOR U22118 ( .A(n20070), .B(n19896), .Z(n20072) );
  XOR U22119 ( .A(n20063), .B(n20064), .Z(n19896) );
  XNOR U22120 ( .A(n20073), .B(n20074), .Z(n20064) );
  ANDN U22121 ( .B(n20075), .A(n20076), .Z(n20073) );
  XOR U22122 ( .A(n20077), .B(n20078), .Z(n20075) );
  XOR U22123 ( .A(n20079), .B(n20080), .Z(n20063) );
  XNOR U22124 ( .A(n20081), .B(n20082), .Z(n20080) );
  ANDN U22125 ( .B(n20083), .A(n20084), .Z(n20081) );
  XNOR U22126 ( .A(n20085), .B(n20086), .Z(n20083) );
  IV U22127 ( .A(n20061), .Z(n20079) );
  XOR U22128 ( .A(n20087), .B(n20088), .Z(n20061) );
  ANDN U22129 ( .B(n20089), .A(n20090), .Z(n20087) );
  XOR U22130 ( .A(n20088), .B(n20091), .Z(n20089) );
  XNOR U22131 ( .A(n20070), .B(n19898), .Z(n20071) );
  XOR U22132 ( .A(n20092), .B(n20093), .Z(n19898) );
  AND U22133 ( .A(n172), .B(n20094), .Z(n20092) );
  XOR U22134 ( .A(n20095), .B(n20093), .Z(n20094) );
  XNOR U22135 ( .A(n20096), .B(n20097), .Z(n20070) );
  AND U22136 ( .A(n20098), .B(n20099), .Z(n20096) );
  XNOR U22137 ( .A(n20097), .B(n19948), .Z(n20099) );
  XOR U22138 ( .A(n20090), .B(n20091), .Z(n19948) );
  XOR U22139 ( .A(n20100), .B(n20078), .Z(n20091) );
  XNOR U22140 ( .A(n20101), .B(n20102), .Z(n20078) );
  ANDN U22141 ( .B(n20103), .A(n20104), .Z(n20101) );
  XOR U22142 ( .A(n20105), .B(n20106), .Z(n20103) );
  IV U22143 ( .A(n20076), .Z(n20100) );
  XOR U22144 ( .A(n20074), .B(n20107), .Z(n20076) );
  XNOR U22145 ( .A(n20108), .B(n20109), .Z(n20107) );
  ANDN U22146 ( .B(n20110), .A(n20111), .Z(n20108) );
  XNOR U22147 ( .A(n20112), .B(n20113), .Z(n20110) );
  IV U22148 ( .A(n20077), .Z(n20074) );
  XOR U22149 ( .A(n20114), .B(n20115), .Z(n20077) );
  ANDN U22150 ( .B(n20116), .A(n20117), .Z(n20114) );
  XOR U22151 ( .A(n20115), .B(n20118), .Z(n20116) );
  XOR U22152 ( .A(n20119), .B(n20120), .Z(n20090) );
  XNOR U22153 ( .A(n20085), .B(n20121), .Z(n20120) );
  IV U22154 ( .A(n20088), .Z(n20121) );
  XOR U22155 ( .A(n20122), .B(n20123), .Z(n20088) );
  ANDN U22156 ( .B(n20124), .A(n20125), .Z(n20122) );
  XOR U22157 ( .A(n20123), .B(n20126), .Z(n20124) );
  XNOR U22158 ( .A(n20127), .B(n20128), .Z(n20085) );
  ANDN U22159 ( .B(n20129), .A(n20130), .Z(n20127) );
  XOR U22160 ( .A(n20128), .B(n20131), .Z(n20129) );
  IV U22161 ( .A(n20084), .Z(n20119) );
  XOR U22162 ( .A(n20082), .B(n20132), .Z(n20084) );
  XNOR U22163 ( .A(n20133), .B(n20134), .Z(n20132) );
  ANDN U22164 ( .B(n20135), .A(n20136), .Z(n20133) );
  XNOR U22165 ( .A(n20137), .B(n20138), .Z(n20135) );
  IV U22166 ( .A(n20086), .Z(n20082) );
  XOR U22167 ( .A(n20139), .B(n20140), .Z(n20086) );
  ANDN U22168 ( .B(n20141), .A(n20142), .Z(n20139) );
  XOR U22169 ( .A(n20143), .B(n20140), .Z(n20141) );
  XOR U22170 ( .A(n20097), .B(n19950), .Z(n20098) );
  XOR U22171 ( .A(n20144), .B(n20145), .Z(n19950) );
  AND U22172 ( .A(n172), .B(n20146), .Z(n20144) );
  XOR U22173 ( .A(n20147), .B(n20145), .Z(n20146) );
  XNOR U22174 ( .A(n20148), .B(n20149), .Z(n20097) );
  NAND U22175 ( .A(n20150), .B(n20151), .Z(n20149) );
  XOR U22176 ( .A(n20152), .B(n20049), .Z(n20151) );
  XOR U22177 ( .A(n20125), .B(n20126), .Z(n20049) );
  XOR U22178 ( .A(n20153), .B(n20118), .Z(n20126) );
  XOR U22179 ( .A(n20154), .B(n20106), .Z(n20118) );
  XOR U22180 ( .A(n20155), .B(n20156), .Z(n20106) );
  ANDN U22181 ( .B(n20157), .A(n20158), .Z(n20155) );
  XOR U22182 ( .A(n20156), .B(n20159), .Z(n20157) );
  IV U22183 ( .A(n20104), .Z(n20154) );
  XOR U22184 ( .A(n20102), .B(n20160), .Z(n20104) );
  XOR U22185 ( .A(n20161), .B(n20162), .Z(n20160) );
  ANDN U22186 ( .B(n20163), .A(n20164), .Z(n20161) );
  XOR U22187 ( .A(n20165), .B(n20162), .Z(n20163) );
  IV U22188 ( .A(n20105), .Z(n20102) );
  XOR U22189 ( .A(n20166), .B(n20167), .Z(n20105) );
  ANDN U22190 ( .B(n20168), .A(n20169), .Z(n20166) );
  XOR U22191 ( .A(n20167), .B(n20170), .Z(n20168) );
  IV U22192 ( .A(n20117), .Z(n20153) );
  XOR U22193 ( .A(n20171), .B(n20172), .Z(n20117) );
  XNOR U22194 ( .A(n20112), .B(n20173), .Z(n20172) );
  IV U22195 ( .A(n20115), .Z(n20173) );
  XOR U22196 ( .A(n20174), .B(n20175), .Z(n20115) );
  ANDN U22197 ( .B(n20176), .A(n20177), .Z(n20174) );
  XOR U22198 ( .A(n20175), .B(n20178), .Z(n20176) );
  XNOR U22199 ( .A(n20179), .B(n20180), .Z(n20112) );
  ANDN U22200 ( .B(n20181), .A(n20182), .Z(n20179) );
  XOR U22201 ( .A(n20180), .B(n20183), .Z(n20181) );
  IV U22202 ( .A(n20111), .Z(n20171) );
  XOR U22203 ( .A(n20109), .B(n20184), .Z(n20111) );
  XOR U22204 ( .A(n20185), .B(n20186), .Z(n20184) );
  ANDN U22205 ( .B(n20187), .A(n20188), .Z(n20185) );
  XOR U22206 ( .A(n20189), .B(n20186), .Z(n20187) );
  IV U22207 ( .A(n20113), .Z(n20109) );
  XOR U22208 ( .A(n20190), .B(n20191), .Z(n20113) );
  ANDN U22209 ( .B(n20192), .A(n20193), .Z(n20190) );
  XOR U22210 ( .A(n20194), .B(n20191), .Z(n20192) );
  XOR U22211 ( .A(n20195), .B(n20196), .Z(n20125) );
  XOR U22212 ( .A(n20143), .B(n20197), .Z(n20196) );
  IV U22213 ( .A(n20123), .Z(n20197) );
  XOR U22214 ( .A(n20198), .B(n20199), .Z(n20123) );
  ANDN U22215 ( .B(n20200), .A(n20201), .Z(n20198) );
  XOR U22216 ( .A(n20199), .B(n20202), .Z(n20200) );
  XOR U22217 ( .A(n20203), .B(n20131), .Z(n20143) );
  XOR U22218 ( .A(n20204), .B(n20205), .Z(n20131) );
  ANDN U22219 ( .B(n20206), .A(n20207), .Z(n20204) );
  XOR U22220 ( .A(n20205), .B(n20208), .Z(n20206) );
  IV U22221 ( .A(n20130), .Z(n20203) );
  XOR U22222 ( .A(n20209), .B(n20210), .Z(n20130) );
  XOR U22223 ( .A(n20211), .B(n20212), .Z(n20210) );
  ANDN U22224 ( .B(n20213), .A(n20214), .Z(n20211) );
  XOR U22225 ( .A(n20215), .B(n20212), .Z(n20213) );
  IV U22226 ( .A(n20128), .Z(n20209) );
  XOR U22227 ( .A(n20216), .B(n20217), .Z(n20128) );
  ANDN U22228 ( .B(n20218), .A(n20219), .Z(n20216) );
  XOR U22229 ( .A(n20217), .B(n20220), .Z(n20218) );
  IV U22230 ( .A(n20142), .Z(n20195) );
  XOR U22231 ( .A(n20221), .B(n20222), .Z(n20142) );
  XNOR U22232 ( .A(n20137), .B(n20223), .Z(n20222) );
  IV U22233 ( .A(n20140), .Z(n20223) );
  XOR U22234 ( .A(n20224), .B(n20225), .Z(n20140) );
  ANDN U22235 ( .B(n20226), .A(n20227), .Z(n20224) );
  XOR U22236 ( .A(n20228), .B(n20225), .Z(n20226) );
  XNOR U22237 ( .A(n20229), .B(n20230), .Z(n20137) );
  ANDN U22238 ( .B(n20231), .A(n20232), .Z(n20229) );
  XOR U22239 ( .A(n20230), .B(n20233), .Z(n20231) );
  IV U22240 ( .A(n20136), .Z(n20221) );
  XOR U22241 ( .A(n20134), .B(n20234), .Z(n20136) );
  XOR U22242 ( .A(n20235), .B(n20236), .Z(n20234) );
  ANDN U22243 ( .B(n20237), .A(n20238), .Z(n20235) );
  XOR U22244 ( .A(n20239), .B(n20236), .Z(n20237) );
  IV U22245 ( .A(n20138), .Z(n20134) );
  XOR U22246 ( .A(n20240), .B(n20241), .Z(n20138) );
  ANDN U22247 ( .B(n20242), .A(n20243), .Z(n20240) );
  XOR U22248 ( .A(n20244), .B(n20241), .Z(n20242) );
  IV U22249 ( .A(n20148), .Z(n20152) );
  XOR U22250 ( .A(n20148), .B(n20051), .Z(n20150) );
  XOR U22251 ( .A(n20245), .B(n20246), .Z(n20051) );
  AND U22252 ( .A(n172), .B(n20247), .Z(n20245) );
  XOR U22253 ( .A(n20248), .B(n20246), .Z(n20247) );
  NANDN U22254 ( .A(n20053), .B(n20055), .Z(n20148) );
  XOR U22255 ( .A(n20249), .B(n20250), .Z(n20055) );
  AND U22256 ( .A(n172), .B(n20251), .Z(n20249) );
  XOR U22257 ( .A(n20250), .B(n20252), .Z(n20251) );
  XNOR U22258 ( .A(n20253), .B(n20254), .Z(n172) );
  AND U22259 ( .A(n20255), .B(n20256), .Z(n20253) );
  XOR U22260 ( .A(n20254), .B(n20066), .Z(n20256) );
  XNOR U22261 ( .A(n20257), .B(n20258), .Z(n20066) );
  ANDN U22262 ( .B(n20259), .A(n20260), .Z(n20257) );
  XOR U22263 ( .A(n20258), .B(n20261), .Z(n20259) );
  XNOR U22264 ( .A(n20254), .B(n20068), .Z(n20255) );
  XOR U22265 ( .A(n20262), .B(n20263), .Z(n20068) );
  AND U22266 ( .A(n176), .B(n20264), .Z(n20262) );
  XOR U22267 ( .A(n20265), .B(n20263), .Z(n20264) );
  XOR U22268 ( .A(n20266), .B(n20267), .Z(n20254) );
  AND U22269 ( .A(n20268), .B(n20269), .Z(n20266) );
  XOR U22270 ( .A(n20267), .B(n20093), .Z(n20269) );
  XOR U22271 ( .A(n20260), .B(n20261), .Z(n20093) );
  XNOR U22272 ( .A(n20270), .B(n20271), .Z(n20261) );
  ANDN U22273 ( .B(n20272), .A(n20273), .Z(n20270) );
  XOR U22274 ( .A(n20274), .B(n20275), .Z(n20272) );
  XOR U22275 ( .A(n20276), .B(n20277), .Z(n20260) );
  XNOR U22276 ( .A(n20278), .B(n20279), .Z(n20277) );
  ANDN U22277 ( .B(n20280), .A(n20281), .Z(n20278) );
  XNOR U22278 ( .A(n20282), .B(n20283), .Z(n20280) );
  IV U22279 ( .A(n20258), .Z(n20276) );
  XOR U22280 ( .A(n20284), .B(n20285), .Z(n20258) );
  ANDN U22281 ( .B(n20286), .A(n20287), .Z(n20284) );
  XOR U22282 ( .A(n20285), .B(n20288), .Z(n20286) );
  XNOR U22283 ( .A(n20267), .B(n20095), .Z(n20268) );
  XOR U22284 ( .A(n20289), .B(n20290), .Z(n20095) );
  AND U22285 ( .A(n176), .B(n20291), .Z(n20289) );
  XOR U22286 ( .A(n20292), .B(n20290), .Z(n20291) );
  XNOR U22287 ( .A(n20293), .B(n20294), .Z(n20267) );
  AND U22288 ( .A(n20295), .B(n20296), .Z(n20293) );
  XNOR U22289 ( .A(n20294), .B(n20145), .Z(n20296) );
  XOR U22290 ( .A(n20287), .B(n20288), .Z(n20145) );
  XOR U22291 ( .A(n20297), .B(n20275), .Z(n20288) );
  XNOR U22292 ( .A(n20298), .B(n20299), .Z(n20275) );
  ANDN U22293 ( .B(n20300), .A(n20301), .Z(n20298) );
  XOR U22294 ( .A(n20302), .B(n20303), .Z(n20300) );
  IV U22295 ( .A(n20273), .Z(n20297) );
  XOR U22296 ( .A(n20271), .B(n20304), .Z(n20273) );
  XNOR U22297 ( .A(n20305), .B(n20306), .Z(n20304) );
  ANDN U22298 ( .B(n20307), .A(n20308), .Z(n20305) );
  XNOR U22299 ( .A(n20309), .B(n20310), .Z(n20307) );
  IV U22300 ( .A(n20274), .Z(n20271) );
  XOR U22301 ( .A(n20311), .B(n20312), .Z(n20274) );
  ANDN U22302 ( .B(n20313), .A(n20314), .Z(n20311) );
  XOR U22303 ( .A(n20312), .B(n20315), .Z(n20313) );
  XOR U22304 ( .A(n20316), .B(n20317), .Z(n20287) );
  XNOR U22305 ( .A(n20282), .B(n20318), .Z(n20317) );
  IV U22306 ( .A(n20285), .Z(n20318) );
  XOR U22307 ( .A(n20319), .B(n20320), .Z(n20285) );
  ANDN U22308 ( .B(n20321), .A(n20322), .Z(n20319) );
  XOR U22309 ( .A(n20320), .B(n20323), .Z(n20321) );
  XNOR U22310 ( .A(n20324), .B(n20325), .Z(n20282) );
  ANDN U22311 ( .B(n20326), .A(n20327), .Z(n20324) );
  XOR U22312 ( .A(n20325), .B(n20328), .Z(n20326) );
  IV U22313 ( .A(n20281), .Z(n20316) );
  XOR U22314 ( .A(n20279), .B(n20329), .Z(n20281) );
  XNOR U22315 ( .A(n20330), .B(n20331), .Z(n20329) );
  ANDN U22316 ( .B(n20332), .A(n20333), .Z(n20330) );
  XNOR U22317 ( .A(n20334), .B(n20335), .Z(n20332) );
  IV U22318 ( .A(n20283), .Z(n20279) );
  XOR U22319 ( .A(n20336), .B(n20337), .Z(n20283) );
  ANDN U22320 ( .B(n20338), .A(n20339), .Z(n20336) );
  XOR U22321 ( .A(n20340), .B(n20337), .Z(n20338) );
  XOR U22322 ( .A(n20294), .B(n20147), .Z(n20295) );
  XOR U22323 ( .A(n20341), .B(n20342), .Z(n20147) );
  AND U22324 ( .A(n176), .B(n20343), .Z(n20341) );
  XOR U22325 ( .A(n20344), .B(n20342), .Z(n20343) );
  XNOR U22326 ( .A(n20345), .B(n20346), .Z(n20294) );
  NAND U22327 ( .A(n20347), .B(n20348), .Z(n20346) );
  XOR U22328 ( .A(n20349), .B(n20246), .Z(n20348) );
  XOR U22329 ( .A(n20322), .B(n20323), .Z(n20246) );
  XOR U22330 ( .A(n20350), .B(n20315), .Z(n20323) );
  XOR U22331 ( .A(n20351), .B(n20303), .Z(n20315) );
  XOR U22332 ( .A(n20352), .B(n20353), .Z(n20303) );
  ANDN U22333 ( .B(n20354), .A(n20355), .Z(n20352) );
  XOR U22334 ( .A(n20353), .B(n20356), .Z(n20354) );
  IV U22335 ( .A(n20301), .Z(n20351) );
  XOR U22336 ( .A(n20299), .B(n20357), .Z(n20301) );
  XOR U22337 ( .A(n20358), .B(n20359), .Z(n20357) );
  ANDN U22338 ( .B(n20360), .A(n20361), .Z(n20358) );
  XOR U22339 ( .A(n20362), .B(n20359), .Z(n20360) );
  IV U22340 ( .A(n20302), .Z(n20299) );
  XOR U22341 ( .A(n20363), .B(n20364), .Z(n20302) );
  ANDN U22342 ( .B(n20365), .A(n20366), .Z(n20363) );
  XOR U22343 ( .A(n20364), .B(n20367), .Z(n20365) );
  IV U22344 ( .A(n20314), .Z(n20350) );
  XOR U22345 ( .A(n20368), .B(n20369), .Z(n20314) );
  XNOR U22346 ( .A(n20309), .B(n20370), .Z(n20369) );
  IV U22347 ( .A(n20312), .Z(n20370) );
  XOR U22348 ( .A(n20371), .B(n20372), .Z(n20312) );
  ANDN U22349 ( .B(n20373), .A(n20374), .Z(n20371) );
  XOR U22350 ( .A(n20372), .B(n20375), .Z(n20373) );
  XNOR U22351 ( .A(n20376), .B(n20377), .Z(n20309) );
  ANDN U22352 ( .B(n20378), .A(n20379), .Z(n20376) );
  XOR U22353 ( .A(n20377), .B(n20380), .Z(n20378) );
  IV U22354 ( .A(n20308), .Z(n20368) );
  XOR U22355 ( .A(n20306), .B(n20381), .Z(n20308) );
  XOR U22356 ( .A(n20382), .B(n20383), .Z(n20381) );
  ANDN U22357 ( .B(n20384), .A(n20385), .Z(n20382) );
  XOR U22358 ( .A(n20386), .B(n20383), .Z(n20384) );
  IV U22359 ( .A(n20310), .Z(n20306) );
  XOR U22360 ( .A(n20387), .B(n20388), .Z(n20310) );
  ANDN U22361 ( .B(n20389), .A(n20390), .Z(n20387) );
  XOR U22362 ( .A(n20391), .B(n20388), .Z(n20389) );
  XOR U22363 ( .A(n20392), .B(n20393), .Z(n20322) );
  XOR U22364 ( .A(n20340), .B(n20394), .Z(n20393) );
  IV U22365 ( .A(n20320), .Z(n20394) );
  XOR U22366 ( .A(n20395), .B(n20396), .Z(n20320) );
  ANDN U22367 ( .B(n20397), .A(n20398), .Z(n20395) );
  XOR U22368 ( .A(n20396), .B(n20399), .Z(n20397) );
  XOR U22369 ( .A(n20400), .B(n20328), .Z(n20340) );
  XOR U22370 ( .A(n20401), .B(n20402), .Z(n20328) );
  ANDN U22371 ( .B(n20403), .A(n20404), .Z(n20401) );
  XOR U22372 ( .A(n20402), .B(n20405), .Z(n20403) );
  IV U22373 ( .A(n20327), .Z(n20400) );
  XOR U22374 ( .A(n20406), .B(n20407), .Z(n20327) );
  XOR U22375 ( .A(n20408), .B(n20409), .Z(n20407) );
  ANDN U22376 ( .B(n20410), .A(n20411), .Z(n20408) );
  XOR U22377 ( .A(n20412), .B(n20409), .Z(n20410) );
  IV U22378 ( .A(n20325), .Z(n20406) );
  XOR U22379 ( .A(n20413), .B(n20414), .Z(n20325) );
  ANDN U22380 ( .B(n20415), .A(n20416), .Z(n20413) );
  XOR U22381 ( .A(n20414), .B(n20417), .Z(n20415) );
  IV U22382 ( .A(n20339), .Z(n20392) );
  XOR U22383 ( .A(n20418), .B(n20419), .Z(n20339) );
  XNOR U22384 ( .A(n20334), .B(n20420), .Z(n20419) );
  IV U22385 ( .A(n20337), .Z(n20420) );
  XOR U22386 ( .A(n20421), .B(n20422), .Z(n20337) );
  ANDN U22387 ( .B(n20423), .A(n20424), .Z(n20421) );
  XOR U22388 ( .A(n20425), .B(n20422), .Z(n20423) );
  XNOR U22389 ( .A(n20426), .B(n20427), .Z(n20334) );
  ANDN U22390 ( .B(n20428), .A(n20429), .Z(n20426) );
  XOR U22391 ( .A(n20427), .B(n20430), .Z(n20428) );
  IV U22392 ( .A(n20333), .Z(n20418) );
  XOR U22393 ( .A(n20331), .B(n20431), .Z(n20333) );
  XOR U22394 ( .A(n20432), .B(n20433), .Z(n20431) );
  ANDN U22395 ( .B(n20434), .A(n20435), .Z(n20432) );
  XOR U22396 ( .A(n20436), .B(n20433), .Z(n20434) );
  IV U22397 ( .A(n20335), .Z(n20331) );
  XOR U22398 ( .A(n20437), .B(n20438), .Z(n20335) );
  ANDN U22399 ( .B(n20439), .A(n20440), .Z(n20437) );
  XOR U22400 ( .A(n20441), .B(n20438), .Z(n20439) );
  IV U22401 ( .A(n20345), .Z(n20349) );
  XOR U22402 ( .A(n20345), .B(n20248), .Z(n20347) );
  XOR U22403 ( .A(n20442), .B(n20443), .Z(n20248) );
  AND U22404 ( .A(n176), .B(n20444), .Z(n20442) );
  XOR U22405 ( .A(n20445), .B(n20443), .Z(n20444) );
  NANDN U22406 ( .A(n20250), .B(n20252), .Z(n20345) );
  XOR U22407 ( .A(n20446), .B(n20447), .Z(n20252) );
  AND U22408 ( .A(n176), .B(n20448), .Z(n20446) );
  XOR U22409 ( .A(n20447), .B(n20449), .Z(n20448) );
  XNOR U22410 ( .A(n20450), .B(n20451), .Z(n176) );
  AND U22411 ( .A(n20452), .B(n20453), .Z(n20450) );
  XOR U22412 ( .A(n20451), .B(n20263), .Z(n20453) );
  XNOR U22413 ( .A(n20454), .B(n20455), .Z(n20263) );
  ANDN U22414 ( .B(n20456), .A(n20457), .Z(n20454) );
  XOR U22415 ( .A(n20455), .B(n20458), .Z(n20456) );
  XNOR U22416 ( .A(n20451), .B(n20265), .Z(n20452) );
  XOR U22417 ( .A(n20459), .B(n20460), .Z(n20265) );
  AND U22418 ( .A(n180), .B(n20461), .Z(n20459) );
  XOR U22419 ( .A(n20462), .B(n20460), .Z(n20461) );
  XOR U22420 ( .A(n20463), .B(n20464), .Z(n20451) );
  AND U22421 ( .A(n20465), .B(n20466), .Z(n20463) );
  XOR U22422 ( .A(n20464), .B(n20290), .Z(n20466) );
  XOR U22423 ( .A(n20457), .B(n20458), .Z(n20290) );
  XNOR U22424 ( .A(n20467), .B(n20468), .Z(n20458) );
  ANDN U22425 ( .B(n20469), .A(n20470), .Z(n20467) );
  XOR U22426 ( .A(n20471), .B(n20472), .Z(n20469) );
  XOR U22427 ( .A(n20473), .B(n20474), .Z(n20457) );
  XNOR U22428 ( .A(n20475), .B(n20476), .Z(n20474) );
  ANDN U22429 ( .B(n20477), .A(n20478), .Z(n20475) );
  XNOR U22430 ( .A(n20479), .B(n20480), .Z(n20477) );
  IV U22431 ( .A(n20455), .Z(n20473) );
  XOR U22432 ( .A(n20481), .B(n20482), .Z(n20455) );
  ANDN U22433 ( .B(n20483), .A(n20484), .Z(n20481) );
  XOR U22434 ( .A(n20482), .B(n20485), .Z(n20483) );
  XNOR U22435 ( .A(n20464), .B(n20292), .Z(n20465) );
  XOR U22436 ( .A(n20486), .B(n20487), .Z(n20292) );
  AND U22437 ( .A(n180), .B(n20488), .Z(n20486) );
  XOR U22438 ( .A(n20489), .B(n20487), .Z(n20488) );
  XNOR U22439 ( .A(n20490), .B(n20491), .Z(n20464) );
  AND U22440 ( .A(n20492), .B(n20493), .Z(n20490) );
  XNOR U22441 ( .A(n20491), .B(n20342), .Z(n20493) );
  XOR U22442 ( .A(n20484), .B(n20485), .Z(n20342) );
  XOR U22443 ( .A(n20494), .B(n20472), .Z(n20485) );
  XNOR U22444 ( .A(n20495), .B(n20496), .Z(n20472) );
  ANDN U22445 ( .B(n20497), .A(n20498), .Z(n20495) );
  XOR U22446 ( .A(n20499), .B(n20500), .Z(n20497) );
  IV U22447 ( .A(n20470), .Z(n20494) );
  XOR U22448 ( .A(n20468), .B(n20501), .Z(n20470) );
  XNOR U22449 ( .A(n20502), .B(n20503), .Z(n20501) );
  ANDN U22450 ( .B(n20504), .A(n20505), .Z(n20502) );
  XNOR U22451 ( .A(n20506), .B(n20507), .Z(n20504) );
  IV U22452 ( .A(n20471), .Z(n20468) );
  XOR U22453 ( .A(n20508), .B(n20509), .Z(n20471) );
  ANDN U22454 ( .B(n20510), .A(n20511), .Z(n20508) );
  XOR U22455 ( .A(n20509), .B(n20512), .Z(n20510) );
  XOR U22456 ( .A(n20513), .B(n20514), .Z(n20484) );
  XNOR U22457 ( .A(n20479), .B(n20515), .Z(n20514) );
  IV U22458 ( .A(n20482), .Z(n20515) );
  XOR U22459 ( .A(n20516), .B(n20517), .Z(n20482) );
  ANDN U22460 ( .B(n20518), .A(n20519), .Z(n20516) );
  XOR U22461 ( .A(n20517), .B(n20520), .Z(n20518) );
  XNOR U22462 ( .A(n20521), .B(n20522), .Z(n20479) );
  ANDN U22463 ( .B(n20523), .A(n20524), .Z(n20521) );
  XOR U22464 ( .A(n20522), .B(n20525), .Z(n20523) );
  IV U22465 ( .A(n20478), .Z(n20513) );
  XOR U22466 ( .A(n20476), .B(n20526), .Z(n20478) );
  XNOR U22467 ( .A(n20527), .B(n20528), .Z(n20526) );
  ANDN U22468 ( .B(n20529), .A(n20530), .Z(n20527) );
  XNOR U22469 ( .A(n20531), .B(n20532), .Z(n20529) );
  IV U22470 ( .A(n20480), .Z(n20476) );
  XOR U22471 ( .A(n20533), .B(n20534), .Z(n20480) );
  ANDN U22472 ( .B(n20535), .A(n20536), .Z(n20533) );
  XOR U22473 ( .A(n20537), .B(n20534), .Z(n20535) );
  XOR U22474 ( .A(n20491), .B(n20344), .Z(n20492) );
  XOR U22475 ( .A(n20538), .B(n20539), .Z(n20344) );
  AND U22476 ( .A(n180), .B(n20540), .Z(n20538) );
  XOR U22477 ( .A(n20541), .B(n20539), .Z(n20540) );
  XNOR U22478 ( .A(n20542), .B(n20543), .Z(n20491) );
  NAND U22479 ( .A(n20544), .B(n20545), .Z(n20543) );
  XOR U22480 ( .A(n20546), .B(n20443), .Z(n20545) );
  XOR U22481 ( .A(n20519), .B(n20520), .Z(n20443) );
  XOR U22482 ( .A(n20547), .B(n20512), .Z(n20520) );
  XOR U22483 ( .A(n20548), .B(n20500), .Z(n20512) );
  XOR U22484 ( .A(n20549), .B(n20550), .Z(n20500) );
  ANDN U22485 ( .B(n20551), .A(n20552), .Z(n20549) );
  XOR U22486 ( .A(n20550), .B(n20553), .Z(n20551) );
  IV U22487 ( .A(n20498), .Z(n20548) );
  XOR U22488 ( .A(n20496), .B(n20554), .Z(n20498) );
  XOR U22489 ( .A(n20555), .B(n20556), .Z(n20554) );
  ANDN U22490 ( .B(n20557), .A(n20558), .Z(n20555) );
  XOR U22491 ( .A(n20559), .B(n20556), .Z(n20557) );
  IV U22492 ( .A(n20499), .Z(n20496) );
  XOR U22493 ( .A(n20560), .B(n20561), .Z(n20499) );
  ANDN U22494 ( .B(n20562), .A(n20563), .Z(n20560) );
  XOR U22495 ( .A(n20561), .B(n20564), .Z(n20562) );
  IV U22496 ( .A(n20511), .Z(n20547) );
  XOR U22497 ( .A(n20565), .B(n20566), .Z(n20511) );
  XNOR U22498 ( .A(n20506), .B(n20567), .Z(n20566) );
  IV U22499 ( .A(n20509), .Z(n20567) );
  XOR U22500 ( .A(n20568), .B(n20569), .Z(n20509) );
  ANDN U22501 ( .B(n20570), .A(n20571), .Z(n20568) );
  XOR U22502 ( .A(n20569), .B(n20572), .Z(n20570) );
  XNOR U22503 ( .A(n20573), .B(n20574), .Z(n20506) );
  ANDN U22504 ( .B(n20575), .A(n20576), .Z(n20573) );
  XOR U22505 ( .A(n20574), .B(n20577), .Z(n20575) );
  IV U22506 ( .A(n20505), .Z(n20565) );
  XOR U22507 ( .A(n20503), .B(n20578), .Z(n20505) );
  XOR U22508 ( .A(n20579), .B(n20580), .Z(n20578) );
  ANDN U22509 ( .B(n20581), .A(n20582), .Z(n20579) );
  XOR U22510 ( .A(n20583), .B(n20580), .Z(n20581) );
  IV U22511 ( .A(n20507), .Z(n20503) );
  XOR U22512 ( .A(n20584), .B(n20585), .Z(n20507) );
  ANDN U22513 ( .B(n20586), .A(n20587), .Z(n20584) );
  XOR U22514 ( .A(n20588), .B(n20585), .Z(n20586) );
  XOR U22515 ( .A(n20589), .B(n20590), .Z(n20519) );
  XOR U22516 ( .A(n20537), .B(n20591), .Z(n20590) );
  IV U22517 ( .A(n20517), .Z(n20591) );
  XOR U22518 ( .A(n20592), .B(n20593), .Z(n20517) );
  ANDN U22519 ( .B(n20594), .A(n20595), .Z(n20592) );
  XOR U22520 ( .A(n20593), .B(n20596), .Z(n20594) );
  XOR U22521 ( .A(n20597), .B(n20525), .Z(n20537) );
  XOR U22522 ( .A(n20598), .B(n20599), .Z(n20525) );
  ANDN U22523 ( .B(n20600), .A(n20601), .Z(n20598) );
  XOR U22524 ( .A(n20599), .B(n20602), .Z(n20600) );
  IV U22525 ( .A(n20524), .Z(n20597) );
  XOR U22526 ( .A(n20603), .B(n20604), .Z(n20524) );
  XOR U22527 ( .A(n20605), .B(n20606), .Z(n20604) );
  ANDN U22528 ( .B(n20607), .A(n20608), .Z(n20605) );
  XOR U22529 ( .A(n20609), .B(n20606), .Z(n20607) );
  IV U22530 ( .A(n20522), .Z(n20603) );
  XOR U22531 ( .A(n20610), .B(n20611), .Z(n20522) );
  ANDN U22532 ( .B(n20612), .A(n20613), .Z(n20610) );
  XOR U22533 ( .A(n20611), .B(n20614), .Z(n20612) );
  IV U22534 ( .A(n20536), .Z(n20589) );
  XOR U22535 ( .A(n20615), .B(n20616), .Z(n20536) );
  XNOR U22536 ( .A(n20531), .B(n20617), .Z(n20616) );
  IV U22537 ( .A(n20534), .Z(n20617) );
  XOR U22538 ( .A(n20618), .B(n20619), .Z(n20534) );
  ANDN U22539 ( .B(n20620), .A(n20621), .Z(n20618) );
  XOR U22540 ( .A(n20622), .B(n20619), .Z(n20620) );
  XNOR U22541 ( .A(n20623), .B(n20624), .Z(n20531) );
  ANDN U22542 ( .B(n20625), .A(n20626), .Z(n20623) );
  XOR U22543 ( .A(n20624), .B(n20627), .Z(n20625) );
  IV U22544 ( .A(n20530), .Z(n20615) );
  XOR U22545 ( .A(n20528), .B(n20628), .Z(n20530) );
  XOR U22546 ( .A(n20629), .B(n20630), .Z(n20628) );
  ANDN U22547 ( .B(n20631), .A(n20632), .Z(n20629) );
  XOR U22548 ( .A(n20633), .B(n20630), .Z(n20631) );
  IV U22549 ( .A(n20532), .Z(n20528) );
  XOR U22550 ( .A(n20634), .B(n20635), .Z(n20532) );
  ANDN U22551 ( .B(n20636), .A(n20637), .Z(n20634) );
  XOR U22552 ( .A(n20638), .B(n20635), .Z(n20636) );
  IV U22553 ( .A(n20542), .Z(n20546) );
  XOR U22554 ( .A(n20542), .B(n20445), .Z(n20544) );
  XOR U22555 ( .A(n20639), .B(n20640), .Z(n20445) );
  AND U22556 ( .A(n180), .B(n20641), .Z(n20639) );
  XOR U22557 ( .A(n20642), .B(n20640), .Z(n20641) );
  NANDN U22558 ( .A(n20447), .B(n20449), .Z(n20542) );
  XOR U22559 ( .A(n20643), .B(n20644), .Z(n20449) );
  AND U22560 ( .A(n180), .B(n20645), .Z(n20643) );
  XOR U22561 ( .A(n20644), .B(n20646), .Z(n20645) );
  XNOR U22562 ( .A(n20647), .B(n20648), .Z(n180) );
  AND U22563 ( .A(n20649), .B(n20650), .Z(n20647) );
  XOR U22564 ( .A(n20648), .B(n20460), .Z(n20650) );
  XNOR U22565 ( .A(n20651), .B(n20652), .Z(n20460) );
  ANDN U22566 ( .B(n20653), .A(n20654), .Z(n20651) );
  XOR U22567 ( .A(n20652), .B(n20655), .Z(n20653) );
  XNOR U22568 ( .A(n20648), .B(n20462), .Z(n20649) );
  XOR U22569 ( .A(n20656), .B(n20657), .Z(n20462) );
  AND U22570 ( .A(n184), .B(n20658), .Z(n20656) );
  XOR U22571 ( .A(n20659), .B(n20657), .Z(n20658) );
  XOR U22572 ( .A(n20660), .B(n20661), .Z(n20648) );
  AND U22573 ( .A(n20662), .B(n20663), .Z(n20660) );
  XOR U22574 ( .A(n20661), .B(n20487), .Z(n20663) );
  XOR U22575 ( .A(n20654), .B(n20655), .Z(n20487) );
  XNOR U22576 ( .A(n20664), .B(n20665), .Z(n20655) );
  ANDN U22577 ( .B(n20666), .A(n20667), .Z(n20664) );
  XOR U22578 ( .A(n20668), .B(n20669), .Z(n20666) );
  XOR U22579 ( .A(n20670), .B(n20671), .Z(n20654) );
  XNOR U22580 ( .A(n20672), .B(n20673), .Z(n20671) );
  ANDN U22581 ( .B(n20674), .A(n20675), .Z(n20672) );
  XNOR U22582 ( .A(n20676), .B(n20677), .Z(n20674) );
  IV U22583 ( .A(n20652), .Z(n20670) );
  XOR U22584 ( .A(n20678), .B(n20679), .Z(n20652) );
  ANDN U22585 ( .B(n20680), .A(n20681), .Z(n20678) );
  XOR U22586 ( .A(n20679), .B(n20682), .Z(n20680) );
  XNOR U22587 ( .A(n20661), .B(n20489), .Z(n20662) );
  XOR U22588 ( .A(n20683), .B(n20684), .Z(n20489) );
  AND U22589 ( .A(n184), .B(n20685), .Z(n20683) );
  XOR U22590 ( .A(n20686), .B(n20684), .Z(n20685) );
  XNOR U22591 ( .A(n20687), .B(n20688), .Z(n20661) );
  AND U22592 ( .A(n20689), .B(n20690), .Z(n20687) );
  XNOR U22593 ( .A(n20688), .B(n20539), .Z(n20690) );
  XOR U22594 ( .A(n20681), .B(n20682), .Z(n20539) );
  XOR U22595 ( .A(n20691), .B(n20669), .Z(n20682) );
  XNOR U22596 ( .A(n20692), .B(n20693), .Z(n20669) );
  ANDN U22597 ( .B(n20694), .A(n20695), .Z(n20692) );
  XOR U22598 ( .A(n20696), .B(n20697), .Z(n20694) );
  IV U22599 ( .A(n20667), .Z(n20691) );
  XOR U22600 ( .A(n20665), .B(n20698), .Z(n20667) );
  XNOR U22601 ( .A(n20699), .B(n20700), .Z(n20698) );
  ANDN U22602 ( .B(n20701), .A(n20702), .Z(n20699) );
  XNOR U22603 ( .A(n20703), .B(n20704), .Z(n20701) );
  IV U22604 ( .A(n20668), .Z(n20665) );
  XOR U22605 ( .A(n20705), .B(n20706), .Z(n20668) );
  ANDN U22606 ( .B(n20707), .A(n20708), .Z(n20705) );
  XOR U22607 ( .A(n20706), .B(n20709), .Z(n20707) );
  XOR U22608 ( .A(n20710), .B(n20711), .Z(n20681) );
  XNOR U22609 ( .A(n20676), .B(n20712), .Z(n20711) );
  IV U22610 ( .A(n20679), .Z(n20712) );
  XOR U22611 ( .A(n20713), .B(n20714), .Z(n20679) );
  ANDN U22612 ( .B(n20715), .A(n20716), .Z(n20713) );
  XOR U22613 ( .A(n20714), .B(n20717), .Z(n20715) );
  XNOR U22614 ( .A(n20718), .B(n20719), .Z(n20676) );
  ANDN U22615 ( .B(n20720), .A(n20721), .Z(n20718) );
  XOR U22616 ( .A(n20719), .B(n20722), .Z(n20720) );
  IV U22617 ( .A(n20675), .Z(n20710) );
  XOR U22618 ( .A(n20673), .B(n20723), .Z(n20675) );
  XNOR U22619 ( .A(n20724), .B(n20725), .Z(n20723) );
  ANDN U22620 ( .B(n20726), .A(n20727), .Z(n20724) );
  XNOR U22621 ( .A(n20728), .B(n20729), .Z(n20726) );
  IV U22622 ( .A(n20677), .Z(n20673) );
  XOR U22623 ( .A(n20730), .B(n20731), .Z(n20677) );
  ANDN U22624 ( .B(n20732), .A(n20733), .Z(n20730) );
  XOR U22625 ( .A(n20734), .B(n20731), .Z(n20732) );
  XOR U22626 ( .A(n20688), .B(n20541), .Z(n20689) );
  XOR U22627 ( .A(n20735), .B(n20736), .Z(n20541) );
  AND U22628 ( .A(n184), .B(n20737), .Z(n20735) );
  XOR U22629 ( .A(n20738), .B(n20736), .Z(n20737) );
  XNOR U22630 ( .A(n20739), .B(n20740), .Z(n20688) );
  NAND U22631 ( .A(n20741), .B(n20742), .Z(n20740) );
  XOR U22632 ( .A(n20743), .B(n20640), .Z(n20742) );
  XOR U22633 ( .A(n20716), .B(n20717), .Z(n20640) );
  XOR U22634 ( .A(n20744), .B(n20709), .Z(n20717) );
  XOR U22635 ( .A(n20745), .B(n20697), .Z(n20709) );
  XOR U22636 ( .A(n20746), .B(n20747), .Z(n20697) );
  ANDN U22637 ( .B(n20748), .A(n20749), .Z(n20746) );
  XOR U22638 ( .A(n20747), .B(n20750), .Z(n20748) );
  IV U22639 ( .A(n20695), .Z(n20745) );
  XOR U22640 ( .A(n20693), .B(n20751), .Z(n20695) );
  XOR U22641 ( .A(n20752), .B(n20753), .Z(n20751) );
  ANDN U22642 ( .B(n20754), .A(n20755), .Z(n20752) );
  XOR U22643 ( .A(n20756), .B(n20753), .Z(n20754) );
  IV U22644 ( .A(n20696), .Z(n20693) );
  XOR U22645 ( .A(n20757), .B(n20758), .Z(n20696) );
  ANDN U22646 ( .B(n20759), .A(n20760), .Z(n20757) );
  XOR U22647 ( .A(n20758), .B(n20761), .Z(n20759) );
  IV U22648 ( .A(n20708), .Z(n20744) );
  XOR U22649 ( .A(n20762), .B(n20763), .Z(n20708) );
  XNOR U22650 ( .A(n20703), .B(n20764), .Z(n20763) );
  IV U22651 ( .A(n20706), .Z(n20764) );
  XOR U22652 ( .A(n20765), .B(n20766), .Z(n20706) );
  ANDN U22653 ( .B(n20767), .A(n20768), .Z(n20765) );
  XOR U22654 ( .A(n20766), .B(n20769), .Z(n20767) );
  XNOR U22655 ( .A(n20770), .B(n20771), .Z(n20703) );
  ANDN U22656 ( .B(n20772), .A(n20773), .Z(n20770) );
  XOR U22657 ( .A(n20771), .B(n20774), .Z(n20772) );
  IV U22658 ( .A(n20702), .Z(n20762) );
  XOR U22659 ( .A(n20700), .B(n20775), .Z(n20702) );
  XOR U22660 ( .A(n20776), .B(n20777), .Z(n20775) );
  ANDN U22661 ( .B(n20778), .A(n20779), .Z(n20776) );
  XOR U22662 ( .A(n20780), .B(n20777), .Z(n20778) );
  IV U22663 ( .A(n20704), .Z(n20700) );
  XOR U22664 ( .A(n20781), .B(n20782), .Z(n20704) );
  ANDN U22665 ( .B(n20783), .A(n20784), .Z(n20781) );
  XOR U22666 ( .A(n20785), .B(n20782), .Z(n20783) );
  XOR U22667 ( .A(n20786), .B(n20787), .Z(n20716) );
  XOR U22668 ( .A(n20734), .B(n20788), .Z(n20787) );
  IV U22669 ( .A(n20714), .Z(n20788) );
  XOR U22670 ( .A(n20789), .B(n20790), .Z(n20714) );
  ANDN U22671 ( .B(n20791), .A(n20792), .Z(n20789) );
  XOR U22672 ( .A(n20790), .B(n20793), .Z(n20791) );
  XOR U22673 ( .A(n20794), .B(n20722), .Z(n20734) );
  XOR U22674 ( .A(n20795), .B(n20796), .Z(n20722) );
  ANDN U22675 ( .B(n20797), .A(n20798), .Z(n20795) );
  XOR U22676 ( .A(n20796), .B(n20799), .Z(n20797) );
  IV U22677 ( .A(n20721), .Z(n20794) );
  XOR U22678 ( .A(n20800), .B(n20801), .Z(n20721) );
  XOR U22679 ( .A(n20802), .B(n20803), .Z(n20801) );
  ANDN U22680 ( .B(n20804), .A(n20805), .Z(n20802) );
  XOR U22681 ( .A(n20806), .B(n20803), .Z(n20804) );
  IV U22682 ( .A(n20719), .Z(n20800) );
  XOR U22683 ( .A(n20807), .B(n20808), .Z(n20719) );
  ANDN U22684 ( .B(n20809), .A(n20810), .Z(n20807) );
  XOR U22685 ( .A(n20808), .B(n20811), .Z(n20809) );
  IV U22686 ( .A(n20733), .Z(n20786) );
  XOR U22687 ( .A(n20812), .B(n20813), .Z(n20733) );
  XNOR U22688 ( .A(n20728), .B(n20814), .Z(n20813) );
  IV U22689 ( .A(n20731), .Z(n20814) );
  XOR U22690 ( .A(n20815), .B(n20816), .Z(n20731) );
  ANDN U22691 ( .B(n20817), .A(n20818), .Z(n20815) );
  XOR U22692 ( .A(n20819), .B(n20816), .Z(n20817) );
  XNOR U22693 ( .A(n20820), .B(n20821), .Z(n20728) );
  ANDN U22694 ( .B(n20822), .A(n20823), .Z(n20820) );
  XOR U22695 ( .A(n20821), .B(n20824), .Z(n20822) );
  IV U22696 ( .A(n20727), .Z(n20812) );
  XOR U22697 ( .A(n20725), .B(n20825), .Z(n20727) );
  XOR U22698 ( .A(n20826), .B(n20827), .Z(n20825) );
  ANDN U22699 ( .B(n20828), .A(n20829), .Z(n20826) );
  XOR U22700 ( .A(n20830), .B(n20827), .Z(n20828) );
  IV U22701 ( .A(n20729), .Z(n20725) );
  XOR U22702 ( .A(n20831), .B(n20832), .Z(n20729) );
  ANDN U22703 ( .B(n20833), .A(n20834), .Z(n20831) );
  XOR U22704 ( .A(n20835), .B(n20832), .Z(n20833) );
  IV U22705 ( .A(n20739), .Z(n20743) );
  XOR U22706 ( .A(n20739), .B(n20642), .Z(n20741) );
  XOR U22707 ( .A(n20836), .B(n20837), .Z(n20642) );
  AND U22708 ( .A(n184), .B(n20838), .Z(n20836) );
  XOR U22709 ( .A(n20839), .B(n20837), .Z(n20838) );
  NANDN U22710 ( .A(n20644), .B(n20646), .Z(n20739) );
  XOR U22711 ( .A(n20840), .B(n20841), .Z(n20646) );
  AND U22712 ( .A(n184), .B(n20842), .Z(n20840) );
  XOR U22713 ( .A(n20841), .B(n20843), .Z(n20842) );
  XNOR U22714 ( .A(n20844), .B(n20845), .Z(n184) );
  AND U22715 ( .A(n20846), .B(n20847), .Z(n20844) );
  XOR U22716 ( .A(n20845), .B(n20657), .Z(n20847) );
  XNOR U22717 ( .A(n20848), .B(n20849), .Z(n20657) );
  ANDN U22718 ( .B(n20850), .A(n20851), .Z(n20848) );
  XOR U22719 ( .A(n20849), .B(n20852), .Z(n20850) );
  XNOR U22720 ( .A(n20845), .B(n20659), .Z(n20846) );
  XOR U22721 ( .A(n20853), .B(n20854), .Z(n20659) );
  AND U22722 ( .A(n188), .B(n20855), .Z(n20853) );
  XOR U22723 ( .A(n20856), .B(n20854), .Z(n20855) );
  XOR U22724 ( .A(n20857), .B(n20858), .Z(n20845) );
  AND U22725 ( .A(n20859), .B(n20860), .Z(n20857) );
  XOR U22726 ( .A(n20858), .B(n20684), .Z(n20860) );
  XOR U22727 ( .A(n20851), .B(n20852), .Z(n20684) );
  XNOR U22728 ( .A(n20861), .B(n20862), .Z(n20852) );
  ANDN U22729 ( .B(n20863), .A(n20864), .Z(n20861) );
  XOR U22730 ( .A(n20865), .B(n20866), .Z(n20863) );
  XOR U22731 ( .A(n20867), .B(n20868), .Z(n20851) );
  XNOR U22732 ( .A(n20869), .B(n20870), .Z(n20868) );
  ANDN U22733 ( .B(n20871), .A(n20872), .Z(n20869) );
  XNOR U22734 ( .A(n20873), .B(n20874), .Z(n20871) );
  IV U22735 ( .A(n20849), .Z(n20867) );
  XOR U22736 ( .A(n20875), .B(n20876), .Z(n20849) );
  ANDN U22737 ( .B(n20877), .A(n20878), .Z(n20875) );
  XOR U22738 ( .A(n20876), .B(n20879), .Z(n20877) );
  XNOR U22739 ( .A(n20858), .B(n20686), .Z(n20859) );
  XOR U22740 ( .A(n20880), .B(n20881), .Z(n20686) );
  AND U22741 ( .A(n188), .B(n20882), .Z(n20880) );
  XOR U22742 ( .A(n20883), .B(n20881), .Z(n20882) );
  XNOR U22743 ( .A(n20884), .B(n20885), .Z(n20858) );
  AND U22744 ( .A(n20886), .B(n20887), .Z(n20884) );
  XNOR U22745 ( .A(n20885), .B(n20736), .Z(n20887) );
  XOR U22746 ( .A(n20878), .B(n20879), .Z(n20736) );
  XOR U22747 ( .A(n20888), .B(n20866), .Z(n20879) );
  XNOR U22748 ( .A(n20889), .B(n20890), .Z(n20866) );
  ANDN U22749 ( .B(n20891), .A(n20892), .Z(n20889) );
  XOR U22750 ( .A(n20893), .B(n20894), .Z(n20891) );
  IV U22751 ( .A(n20864), .Z(n20888) );
  XOR U22752 ( .A(n20862), .B(n20895), .Z(n20864) );
  XNOR U22753 ( .A(n20896), .B(n20897), .Z(n20895) );
  ANDN U22754 ( .B(n20898), .A(n20899), .Z(n20896) );
  XNOR U22755 ( .A(n20900), .B(n20901), .Z(n20898) );
  IV U22756 ( .A(n20865), .Z(n20862) );
  XOR U22757 ( .A(n20902), .B(n20903), .Z(n20865) );
  ANDN U22758 ( .B(n20904), .A(n20905), .Z(n20902) );
  XOR U22759 ( .A(n20903), .B(n20906), .Z(n20904) );
  XOR U22760 ( .A(n20907), .B(n20908), .Z(n20878) );
  XNOR U22761 ( .A(n20873), .B(n20909), .Z(n20908) );
  IV U22762 ( .A(n20876), .Z(n20909) );
  XOR U22763 ( .A(n20910), .B(n20911), .Z(n20876) );
  ANDN U22764 ( .B(n20912), .A(n20913), .Z(n20910) );
  XOR U22765 ( .A(n20911), .B(n20914), .Z(n20912) );
  XNOR U22766 ( .A(n20915), .B(n20916), .Z(n20873) );
  ANDN U22767 ( .B(n20917), .A(n20918), .Z(n20915) );
  XOR U22768 ( .A(n20916), .B(n20919), .Z(n20917) );
  IV U22769 ( .A(n20872), .Z(n20907) );
  XOR U22770 ( .A(n20870), .B(n20920), .Z(n20872) );
  XNOR U22771 ( .A(n20921), .B(n20922), .Z(n20920) );
  ANDN U22772 ( .B(n20923), .A(n20924), .Z(n20921) );
  XNOR U22773 ( .A(n20925), .B(n20926), .Z(n20923) );
  IV U22774 ( .A(n20874), .Z(n20870) );
  XOR U22775 ( .A(n20927), .B(n20928), .Z(n20874) );
  ANDN U22776 ( .B(n20929), .A(n20930), .Z(n20927) );
  XOR U22777 ( .A(n20931), .B(n20928), .Z(n20929) );
  XOR U22778 ( .A(n20885), .B(n20738), .Z(n20886) );
  XOR U22779 ( .A(n20932), .B(n20933), .Z(n20738) );
  AND U22780 ( .A(n188), .B(n20934), .Z(n20932) );
  XOR U22781 ( .A(n20935), .B(n20933), .Z(n20934) );
  XNOR U22782 ( .A(n20936), .B(n20937), .Z(n20885) );
  NAND U22783 ( .A(n20938), .B(n20939), .Z(n20937) );
  XOR U22784 ( .A(n20940), .B(n20837), .Z(n20939) );
  XOR U22785 ( .A(n20913), .B(n20914), .Z(n20837) );
  XOR U22786 ( .A(n20941), .B(n20906), .Z(n20914) );
  XOR U22787 ( .A(n20942), .B(n20894), .Z(n20906) );
  XOR U22788 ( .A(n20943), .B(n20944), .Z(n20894) );
  ANDN U22789 ( .B(n20945), .A(n20946), .Z(n20943) );
  XOR U22790 ( .A(n20944), .B(n20947), .Z(n20945) );
  IV U22791 ( .A(n20892), .Z(n20942) );
  XOR U22792 ( .A(n20890), .B(n20948), .Z(n20892) );
  XOR U22793 ( .A(n20949), .B(n20950), .Z(n20948) );
  ANDN U22794 ( .B(n20951), .A(n20952), .Z(n20949) );
  XOR U22795 ( .A(n20953), .B(n20950), .Z(n20951) );
  IV U22796 ( .A(n20893), .Z(n20890) );
  XOR U22797 ( .A(n20954), .B(n20955), .Z(n20893) );
  ANDN U22798 ( .B(n20956), .A(n20957), .Z(n20954) );
  XOR U22799 ( .A(n20955), .B(n20958), .Z(n20956) );
  IV U22800 ( .A(n20905), .Z(n20941) );
  XOR U22801 ( .A(n20959), .B(n20960), .Z(n20905) );
  XNOR U22802 ( .A(n20900), .B(n20961), .Z(n20960) );
  IV U22803 ( .A(n20903), .Z(n20961) );
  XOR U22804 ( .A(n20962), .B(n20963), .Z(n20903) );
  ANDN U22805 ( .B(n20964), .A(n20965), .Z(n20962) );
  XOR U22806 ( .A(n20963), .B(n20966), .Z(n20964) );
  XNOR U22807 ( .A(n20967), .B(n20968), .Z(n20900) );
  ANDN U22808 ( .B(n20969), .A(n20970), .Z(n20967) );
  XOR U22809 ( .A(n20968), .B(n20971), .Z(n20969) );
  IV U22810 ( .A(n20899), .Z(n20959) );
  XOR U22811 ( .A(n20897), .B(n20972), .Z(n20899) );
  XOR U22812 ( .A(n20973), .B(n20974), .Z(n20972) );
  ANDN U22813 ( .B(n20975), .A(n20976), .Z(n20973) );
  XOR U22814 ( .A(n20977), .B(n20974), .Z(n20975) );
  IV U22815 ( .A(n20901), .Z(n20897) );
  XOR U22816 ( .A(n20978), .B(n20979), .Z(n20901) );
  ANDN U22817 ( .B(n20980), .A(n20981), .Z(n20978) );
  XOR U22818 ( .A(n20982), .B(n20979), .Z(n20980) );
  XOR U22819 ( .A(n20983), .B(n20984), .Z(n20913) );
  XOR U22820 ( .A(n20931), .B(n20985), .Z(n20984) );
  IV U22821 ( .A(n20911), .Z(n20985) );
  XOR U22822 ( .A(n20986), .B(n20987), .Z(n20911) );
  ANDN U22823 ( .B(n20988), .A(n20989), .Z(n20986) );
  XOR U22824 ( .A(n20987), .B(n20990), .Z(n20988) );
  XOR U22825 ( .A(n20991), .B(n20919), .Z(n20931) );
  XOR U22826 ( .A(n20992), .B(n20993), .Z(n20919) );
  ANDN U22827 ( .B(n20994), .A(n20995), .Z(n20992) );
  XOR U22828 ( .A(n20993), .B(n20996), .Z(n20994) );
  IV U22829 ( .A(n20918), .Z(n20991) );
  XOR U22830 ( .A(n20997), .B(n20998), .Z(n20918) );
  XOR U22831 ( .A(n20999), .B(n21000), .Z(n20998) );
  ANDN U22832 ( .B(n21001), .A(n21002), .Z(n20999) );
  XOR U22833 ( .A(n21003), .B(n21000), .Z(n21001) );
  IV U22834 ( .A(n20916), .Z(n20997) );
  XOR U22835 ( .A(n21004), .B(n21005), .Z(n20916) );
  ANDN U22836 ( .B(n21006), .A(n21007), .Z(n21004) );
  XOR U22837 ( .A(n21005), .B(n21008), .Z(n21006) );
  IV U22838 ( .A(n20930), .Z(n20983) );
  XOR U22839 ( .A(n21009), .B(n21010), .Z(n20930) );
  XNOR U22840 ( .A(n20925), .B(n21011), .Z(n21010) );
  IV U22841 ( .A(n20928), .Z(n21011) );
  XOR U22842 ( .A(n21012), .B(n21013), .Z(n20928) );
  ANDN U22843 ( .B(n21014), .A(n21015), .Z(n21012) );
  XOR U22844 ( .A(n21016), .B(n21013), .Z(n21014) );
  XNOR U22845 ( .A(n21017), .B(n21018), .Z(n20925) );
  ANDN U22846 ( .B(n21019), .A(n21020), .Z(n21017) );
  XOR U22847 ( .A(n21018), .B(n21021), .Z(n21019) );
  IV U22848 ( .A(n20924), .Z(n21009) );
  XOR U22849 ( .A(n20922), .B(n21022), .Z(n20924) );
  XOR U22850 ( .A(n21023), .B(n21024), .Z(n21022) );
  ANDN U22851 ( .B(n21025), .A(n21026), .Z(n21023) );
  XOR U22852 ( .A(n21027), .B(n21024), .Z(n21025) );
  IV U22853 ( .A(n20926), .Z(n20922) );
  XOR U22854 ( .A(n21028), .B(n21029), .Z(n20926) );
  ANDN U22855 ( .B(n21030), .A(n21031), .Z(n21028) );
  XOR U22856 ( .A(n21032), .B(n21029), .Z(n21030) );
  IV U22857 ( .A(n20936), .Z(n20940) );
  XOR U22858 ( .A(n20936), .B(n20839), .Z(n20938) );
  XOR U22859 ( .A(n21033), .B(n21034), .Z(n20839) );
  AND U22860 ( .A(n188), .B(n21035), .Z(n21033) );
  XOR U22861 ( .A(n21036), .B(n21034), .Z(n21035) );
  NANDN U22862 ( .A(n20841), .B(n20843), .Z(n20936) );
  XOR U22863 ( .A(n21037), .B(n21038), .Z(n20843) );
  AND U22864 ( .A(n188), .B(n21039), .Z(n21037) );
  XOR U22865 ( .A(n21038), .B(n21040), .Z(n21039) );
  XNOR U22866 ( .A(n21041), .B(n21042), .Z(n188) );
  AND U22867 ( .A(n21043), .B(n21044), .Z(n21041) );
  XOR U22868 ( .A(n21042), .B(n20854), .Z(n21044) );
  XNOR U22869 ( .A(n21045), .B(n21046), .Z(n20854) );
  ANDN U22870 ( .B(n21047), .A(n21048), .Z(n21045) );
  XOR U22871 ( .A(n21046), .B(n21049), .Z(n21047) );
  XNOR U22872 ( .A(n21042), .B(n20856), .Z(n21043) );
  XOR U22873 ( .A(n21050), .B(n21051), .Z(n20856) );
  AND U22874 ( .A(n192), .B(n21052), .Z(n21050) );
  XOR U22875 ( .A(n21053), .B(n21051), .Z(n21052) );
  XOR U22876 ( .A(n21054), .B(n21055), .Z(n21042) );
  AND U22877 ( .A(n21056), .B(n21057), .Z(n21054) );
  XOR U22878 ( .A(n21055), .B(n20881), .Z(n21057) );
  XOR U22879 ( .A(n21048), .B(n21049), .Z(n20881) );
  XNOR U22880 ( .A(n21058), .B(n21059), .Z(n21049) );
  ANDN U22881 ( .B(n21060), .A(n21061), .Z(n21058) );
  XOR U22882 ( .A(n21062), .B(n21063), .Z(n21060) );
  XOR U22883 ( .A(n21064), .B(n21065), .Z(n21048) );
  XNOR U22884 ( .A(n21066), .B(n21067), .Z(n21065) );
  ANDN U22885 ( .B(n21068), .A(n21069), .Z(n21066) );
  XNOR U22886 ( .A(n21070), .B(n21071), .Z(n21068) );
  IV U22887 ( .A(n21046), .Z(n21064) );
  XOR U22888 ( .A(n21072), .B(n21073), .Z(n21046) );
  ANDN U22889 ( .B(n21074), .A(n21075), .Z(n21072) );
  XOR U22890 ( .A(n21073), .B(n21076), .Z(n21074) );
  XNOR U22891 ( .A(n21055), .B(n20883), .Z(n21056) );
  XOR U22892 ( .A(n21077), .B(n21078), .Z(n20883) );
  AND U22893 ( .A(n192), .B(n21079), .Z(n21077) );
  XOR U22894 ( .A(n21080), .B(n21078), .Z(n21079) );
  XNOR U22895 ( .A(n21081), .B(n21082), .Z(n21055) );
  AND U22896 ( .A(n21083), .B(n21084), .Z(n21081) );
  XNOR U22897 ( .A(n21082), .B(n20933), .Z(n21084) );
  XOR U22898 ( .A(n21075), .B(n21076), .Z(n20933) );
  XOR U22899 ( .A(n21085), .B(n21063), .Z(n21076) );
  XNOR U22900 ( .A(n21086), .B(n21087), .Z(n21063) );
  ANDN U22901 ( .B(n21088), .A(n21089), .Z(n21086) );
  XOR U22902 ( .A(n21090), .B(n21091), .Z(n21088) );
  IV U22903 ( .A(n21061), .Z(n21085) );
  XOR U22904 ( .A(n21059), .B(n21092), .Z(n21061) );
  XNOR U22905 ( .A(n21093), .B(n21094), .Z(n21092) );
  ANDN U22906 ( .B(n21095), .A(n21096), .Z(n21093) );
  XNOR U22907 ( .A(n21097), .B(n21098), .Z(n21095) );
  IV U22908 ( .A(n21062), .Z(n21059) );
  XOR U22909 ( .A(n21099), .B(n21100), .Z(n21062) );
  ANDN U22910 ( .B(n21101), .A(n21102), .Z(n21099) );
  XOR U22911 ( .A(n21100), .B(n21103), .Z(n21101) );
  XOR U22912 ( .A(n21104), .B(n21105), .Z(n21075) );
  XNOR U22913 ( .A(n21070), .B(n21106), .Z(n21105) );
  IV U22914 ( .A(n21073), .Z(n21106) );
  XOR U22915 ( .A(n21107), .B(n21108), .Z(n21073) );
  ANDN U22916 ( .B(n21109), .A(n21110), .Z(n21107) );
  XOR U22917 ( .A(n21108), .B(n21111), .Z(n21109) );
  XNOR U22918 ( .A(n21112), .B(n21113), .Z(n21070) );
  ANDN U22919 ( .B(n21114), .A(n21115), .Z(n21112) );
  XOR U22920 ( .A(n21113), .B(n21116), .Z(n21114) );
  IV U22921 ( .A(n21069), .Z(n21104) );
  XOR U22922 ( .A(n21067), .B(n21117), .Z(n21069) );
  XNOR U22923 ( .A(n21118), .B(n21119), .Z(n21117) );
  ANDN U22924 ( .B(n21120), .A(n21121), .Z(n21118) );
  XNOR U22925 ( .A(n21122), .B(n21123), .Z(n21120) );
  IV U22926 ( .A(n21071), .Z(n21067) );
  XOR U22927 ( .A(n21124), .B(n21125), .Z(n21071) );
  ANDN U22928 ( .B(n21126), .A(n21127), .Z(n21124) );
  XOR U22929 ( .A(n21128), .B(n21125), .Z(n21126) );
  XOR U22930 ( .A(n21082), .B(n20935), .Z(n21083) );
  XOR U22931 ( .A(n21129), .B(n21130), .Z(n20935) );
  AND U22932 ( .A(n192), .B(n21131), .Z(n21129) );
  XOR U22933 ( .A(n21132), .B(n21130), .Z(n21131) );
  XNOR U22934 ( .A(n21133), .B(n21134), .Z(n21082) );
  NAND U22935 ( .A(n21135), .B(n21136), .Z(n21134) );
  XOR U22936 ( .A(n21137), .B(n21034), .Z(n21136) );
  XOR U22937 ( .A(n21110), .B(n21111), .Z(n21034) );
  XOR U22938 ( .A(n21138), .B(n21103), .Z(n21111) );
  XOR U22939 ( .A(n21139), .B(n21091), .Z(n21103) );
  XOR U22940 ( .A(n21140), .B(n21141), .Z(n21091) );
  ANDN U22941 ( .B(n21142), .A(n21143), .Z(n21140) );
  XOR U22942 ( .A(n21141), .B(n21144), .Z(n21142) );
  IV U22943 ( .A(n21089), .Z(n21139) );
  XOR U22944 ( .A(n21087), .B(n21145), .Z(n21089) );
  XOR U22945 ( .A(n21146), .B(n21147), .Z(n21145) );
  ANDN U22946 ( .B(n21148), .A(n21149), .Z(n21146) );
  XOR U22947 ( .A(n21150), .B(n21147), .Z(n21148) );
  IV U22948 ( .A(n21090), .Z(n21087) );
  XOR U22949 ( .A(n21151), .B(n21152), .Z(n21090) );
  ANDN U22950 ( .B(n21153), .A(n21154), .Z(n21151) );
  XOR U22951 ( .A(n21152), .B(n21155), .Z(n21153) );
  IV U22952 ( .A(n21102), .Z(n21138) );
  XOR U22953 ( .A(n21156), .B(n21157), .Z(n21102) );
  XNOR U22954 ( .A(n21097), .B(n21158), .Z(n21157) );
  IV U22955 ( .A(n21100), .Z(n21158) );
  XOR U22956 ( .A(n21159), .B(n21160), .Z(n21100) );
  ANDN U22957 ( .B(n21161), .A(n21162), .Z(n21159) );
  XOR U22958 ( .A(n21160), .B(n21163), .Z(n21161) );
  XNOR U22959 ( .A(n21164), .B(n21165), .Z(n21097) );
  ANDN U22960 ( .B(n21166), .A(n21167), .Z(n21164) );
  XOR U22961 ( .A(n21165), .B(n21168), .Z(n21166) );
  IV U22962 ( .A(n21096), .Z(n21156) );
  XOR U22963 ( .A(n21094), .B(n21169), .Z(n21096) );
  XOR U22964 ( .A(n21170), .B(n21171), .Z(n21169) );
  ANDN U22965 ( .B(n21172), .A(n21173), .Z(n21170) );
  XOR U22966 ( .A(n21174), .B(n21171), .Z(n21172) );
  IV U22967 ( .A(n21098), .Z(n21094) );
  XOR U22968 ( .A(n21175), .B(n21176), .Z(n21098) );
  ANDN U22969 ( .B(n21177), .A(n21178), .Z(n21175) );
  XOR U22970 ( .A(n21179), .B(n21176), .Z(n21177) );
  XOR U22971 ( .A(n21180), .B(n21181), .Z(n21110) );
  XOR U22972 ( .A(n21128), .B(n21182), .Z(n21181) );
  IV U22973 ( .A(n21108), .Z(n21182) );
  XOR U22974 ( .A(n21183), .B(n21184), .Z(n21108) );
  ANDN U22975 ( .B(n21185), .A(n21186), .Z(n21183) );
  XOR U22976 ( .A(n21184), .B(n21187), .Z(n21185) );
  XOR U22977 ( .A(n21188), .B(n21116), .Z(n21128) );
  XOR U22978 ( .A(n21189), .B(n21190), .Z(n21116) );
  ANDN U22979 ( .B(n21191), .A(n21192), .Z(n21189) );
  XOR U22980 ( .A(n21190), .B(n21193), .Z(n21191) );
  IV U22981 ( .A(n21115), .Z(n21188) );
  XOR U22982 ( .A(n21194), .B(n21195), .Z(n21115) );
  XOR U22983 ( .A(n21196), .B(n21197), .Z(n21195) );
  ANDN U22984 ( .B(n21198), .A(n21199), .Z(n21196) );
  XOR U22985 ( .A(n21200), .B(n21197), .Z(n21198) );
  IV U22986 ( .A(n21113), .Z(n21194) );
  XOR U22987 ( .A(n21201), .B(n21202), .Z(n21113) );
  ANDN U22988 ( .B(n21203), .A(n21204), .Z(n21201) );
  XOR U22989 ( .A(n21202), .B(n21205), .Z(n21203) );
  IV U22990 ( .A(n21127), .Z(n21180) );
  XOR U22991 ( .A(n21206), .B(n21207), .Z(n21127) );
  XNOR U22992 ( .A(n21122), .B(n21208), .Z(n21207) );
  IV U22993 ( .A(n21125), .Z(n21208) );
  XOR U22994 ( .A(n21209), .B(n21210), .Z(n21125) );
  ANDN U22995 ( .B(n21211), .A(n21212), .Z(n21209) );
  XOR U22996 ( .A(n21213), .B(n21210), .Z(n21211) );
  XNOR U22997 ( .A(n21214), .B(n21215), .Z(n21122) );
  ANDN U22998 ( .B(n21216), .A(n21217), .Z(n21214) );
  XOR U22999 ( .A(n21215), .B(n21218), .Z(n21216) );
  IV U23000 ( .A(n21121), .Z(n21206) );
  XOR U23001 ( .A(n21119), .B(n21219), .Z(n21121) );
  XOR U23002 ( .A(n21220), .B(n21221), .Z(n21219) );
  ANDN U23003 ( .B(n21222), .A(n21223), .Z(n21220) );
  XOR U23004 ( .A(n21224), .B(n21221), .Z(n21222) );
  IV U23005 ( .A(n21123), .Z(n21119) );
  XOR U23006 ( .A(n21225), .B(n21226), .Z(n21123) );
  ANDN U23007 ( .B(n21227), .A(n21228), .Z(n21225) );
  XOR U23008 ( .A(n21229), .B(n21226), .Z(n21227) );
  IV U23009 ( .A(n21133), .Z(n21137) );
  XOR U23010 ( .A(n21133), .B(n21036), .Z(n21135) );
  XOR U23011 ( .A(n21230), .B(n21231), .Z(n21036) );
  AND U23012 ( .A(n192), .B(n21232), .Z(n21230) );
  XOR U23013 ( .A(n21233), .B(n21231), .Z(n21232) );
  NANDN U23014 ( .A(n21038), .B(n21040), .Z(n21133) );
  XOR U23015 ( .A(n21234), .B(n21235), .Z(n21040) );
  AND U23016 ( .A(n192), .B(n21236), .Z(n21234) );
  XOR U23017 ( .A(n21235), .B(n21237), .Z(n21236) );
  XNOR U23018 ( .A(n21238), .B(n21239), .Z(n192) );
  AND U23019 ( .A(n21240), .B(n21241), .Z(n21238) );
  XOR U23020 ( .A(n21239), .B(n21051), .Z(n21241) );
  XNOR U23021 ( .A(n21242), .B(n21243), .Z(n21051) );
  ANDN U23022 ( .B(n21244), .A(n21245), .Z(n21242) );
  XOR U23023 ( .A(n21243), .B(n21246), .Z(n21244) );
  XNOR U23024 ( .A(n21239), .B(n21053), .Z(n21240) );
  XOR U23025 ( .A(n21247), .B(n21248), .Z(n21053) );
  AND U23026 ( .A(n196), .B(n21249), .Z(n21247) );
  XOR U23027 ( .A(n21250), .B(n21248), .Z(n21249) );
  XOR U23028 ( .A(n21251), .B(n21252), .Z(n21239) );
  AND U23029 ( .A(n21253), .B(n21254), .Z(n21251) );
  XOR U23030 ( .A(n21252), .B(n21078), .Z(n21254) );
  XOR U23031 ( .A(n21245), .B(n21246), .Z(n21078) );
  XNOR U23032 ( .A(n21255), .B(n21256), .Z(n21246) );
  ANDN U23033 ( .B(n21257), .A(n21258), .Z(n21255) );
  XOR U23034 ( .A(n21259), .B(n21260), .Z(n21257) );
  XOR U23035 ( .A(n21261), .B(n21262), .Z(n21245) );
  XNOR U23036 ( .A(n21263), .B(n21264), .Z(n21262) );
  ANDN U23037 ( .B(n21265), .A(n21266), .Z(n21263) );
  XNOR U23038 ( .A(n21267), .B(n21268), .Z(n21265) );
  IV U23039 ( .A(n21243), .Z(n21261) );
  XOR U23040 ( .A(n21269), .B(n21270), .Z(n21243) );
  ANDN U23041 ( .B(n21271), .A(n21272), .Z(n21269) );
  XOR U23042 ( .A(n21270), .B(n21273), .Z(n21271) );
  XNOR U23043 ( .A(n21252), .B(n21080), .Z(n21253) );
  XOR U23044 ( .A(n21274), .B(n21275), .Z(n21080) );
  AND U23045 ( .A(n196), .B(n21276), .Z(n21274) );
  XOR U23046 ( .A(n21277), .B(n21275), .Z(n21276) );
  XNOR U23047 ( .A(n21278), .B(n21279), .Z(n21252) );
  AND U23048 ( .A(n21280), .B(n21281), .Z(n21278) );
  XNOR U23049 ( .A(n21279), .B(n21130), .Z(n21281) );
  XOR U23050 ( .A(n21272), .B(n21273), .Z(n21130) );
  XOR U23051 ( .A(n21282), .B(n21260), .Z(n21273) );
  XNOR U23052 ( .A(n21283), .B(n21284), .Z(n21260) );
  ANDN U23053 ( .B(n21285), .A(n21286), .Z(n21283) );
  XOR U23054 ( .A(n21287), .B(n21288), .Z(n21285) );
  IV U23055 ( .A(n21258), .Z(n21282) );
  XOR U23056 ( .A(n21256), .B(n21289), .Z(n21258) );
  XNOR U23057 ( .A(n21290), .B(n21291), .Z(n21289) );
  ANDN U23058 ( .B(n21292), .A(n21293), .Z(n21290) );
  XNOR U23059 ( .A(n21294), .B(n21295), .Z(n21292) );
  IV U23060 ( .A(n21259), .Z(n21256) );
  XOR U23061 ( .A(n21296), .B(n21297), .Z(n21259) );
  ANDN U23062 ( .B(n21298), .A(n21299), .Z(n21296) );
  XOR U23063 ( .A(n21297), .B(n21300), .Z(n21298) );
  XOR U23064 ( .A(n21301), .B(n21302), .Z(n21272) );
  XNOR U23065 ( .A(n21267), .B(n21303), .Z(n21302) );
  IV U23066 ( .A(n21270), .Z(n21303) );
  XOR U23067 ( .A(n21304), .B(n21305), .Z(n21270) );
  ANDN U23068 ( .B(n21306), .A(n21307), .Z(n21304) );
  XOR U23069 ( .A(n21305), .B(n21308), .Z(n21306) );
  XNOR U23070 ( .A(n21309), .B(n21310), .Z(n21267) );
  ANDN U23071 ( .B(n21311), .A(n21312), .Z(n21309) );
  XOR U23072 ( .A(n21310), .B(n21313), .Z(n21311) );
  IV U23073 ( .A(n21266), .Z(n21301) );
  XOR U23074 ( .A(n21264), .B(n21314), .Z(n21266) );
  XNOR U23075 ( .A(n21315), .B(n21316), .Z(n21314) );
  ANDN U23076 ( .B(n21317), .A(n21318), .Z(n21315) );
  XNOR U23077 ( .A(n21319), .B(n21320), .Z(n21317) );
  IV U23078 ( .A(n21268), .Z(n21264) );
  XOR U23079 ( .A(n21321), .B(n21322), .Z(n21268) );
  ANDN U23080 ( .B(n21323), .A(n21324), .Z(n21321) );
  XOR U23081 ( .A(n21325), .B(n21322), .Z(n21323) );
  XOR U23082 ( .A(n21279), .B(n21132), .Z(n21280) );
  XOR U23083 ( .A(n21326), .B(n21327), .Z(n21132) );
  AND U23084 ( .A(n196), .B(n21328), .Z(n21326) );
  XOR U23085 ( .A(n21329), .B(n21327), .Z(n21328) );
  XNOR U23086 ( .A(n21330), .B(n21331), .Z(n21279) );
  NAND U23087 ( .A(n21332), .B(n21333), .Z(n21331) );
  XOR U23088 ( .A(n21334), .B(n21231), .Z(n21333) );
  XOR U23089 ( .A(n21307), .B(n21308), .Z(n21231) );
  XOR U23090 ( .A(n21335), .B(n21300), .Z(n21308) );
  XOR U23091 ( .A(n21336), .B(n21288), .Z(n21300) );
  XOR U23092 ( .A(n21337), .B(n21338), .Z(n21288) );
  ANDN U23093 ( .B(n21339), .A(n21340), .Z(n21337) );
  XOR U23094 ( .A(n21338), .B(n21341), .Z(n21339) );
  IV U23095 ( .A(n21286), .Z(n21336) );
  XOR U23096 ( .A(n21284), .B(n21342), .Z(n21286) );
  XOR U23097 ( .A(n21343), .B(n21344), .Z(n21342) );
  ANDN U23098 ( .B(n21345), .A(n21346), .Z(n21343) );
  XOR U23099 ( .A(n21347), .B(n21344), .Z(n21345) );
  IV U23100 ( .A(n21287), .Z(n21284) );
  XOR U23101 ( .A(n21348), .B(n21349), .Z(n21287) );
  ANDN U23102 ( .B(n21350), .A(n21351), .Z(n21348) );
  XOR U23103 ( .A(n21349), .B(n21352), .Z(n21350) );
  IV U23104 ( .A(n21299), .Z(n21335) );
  XOR U23105 ( .A(n21353), .B(n21354), .Z(n21299) );
  XNOR U23106 ( .A(n21294), .B(n21355), .Z(n21354) );
  IV U23107 ( .A(n21297), .Z(n21355) );
  XOR U23108 ( .A(n21356), .B(n21357), .Z(n21297) );
  ANDN U23109 ( .B(n21358), .A(n21359), .Z(n21356) );
  XOR U23110 ( .A(n21357), .B(n21360), .Z(n21358) );
  XNOR U23111 ( .A(n21361), .B(n21362), .Z(n21294) );
  ANDN U23112 ( .B(n21363), .A(n21364), .Z(n21361) );
  XOR U23113 ( .A(n21362), .B(n21365), .Z(n21363) );
  IV U23114 ( .A(n21293), .Z(n21353) );
  XOR U23115 ( .A(n21291), .B(n21366), .Z(n21293) );
  XOR U23116 ( .A(n21367), .B(n21368), .Z(n21366) );
  ANDN U23117 ( .B(n21369), .A(n21370), .Z(n21367) );
  XOR U23118 ( .A(n21371), .B(n21368), .Z(n21369) );
  IV U23119 ( .A(n21295), .Z(n21291) );
  XOR U23120 ( .A(n21372), .B(n21373), .Z(n21295) );
  ANDN U23121 ( .B(n21374), .A(n21375), .Z(n21372) );
  XOR U23122 ( .A(n21376), .B(n21373), .Z(n21374) );
  XOR U23123 ( .A(n21377), .B(n21378), .Z(n21307) );
  XOR U23124 ( .A(n21325), .B(n21379), .Z(n21378) );
  IV U23125 ( .A(n21305), .Z(n21379) );
  XOR U23126 ( .A(n21380), .B(n21381), .Z(n21305) );
  ANDN U23127 ( .B(n21382), .A(n21383), .Z(n21380) );
  XOR U23128 ( .A(n21381), .B(n21384), .Z(n21382) );
  XOR U23129 ( .A(n21385), .B(n21313), .Z(n21325) );
  XOR U23130 ( .A(n21386), .B(n21387), .Z(n21313) );
  ANDN U23131 ( .B(n21388), .A(n21389), .Z(n21386) );
  XOR U23132 ( .A(n21387), .B(n21390), .Z(n21388) );
  IV U23133 ( .A(n21312), .Z(n21385) );
  XOR U23134 ( .A(n21391), .B(n21392), .Z(n21312) );
  XOR U23135 ( .A(n21393), .B(n21394), .Z(n21392) );
  ANDN U23136 ( .B(n21395), .A(n21396), .Z(n21393) );
  XOR U23137 ( .A(n21397), .B(n21394), .Z(n21395) );
  IV U23138 ( .A(n21310), .Z(n21391) );
  XOR U23139 ( .A(n21398), .B(n21399), .Z(n21310) );
  ANDN U23140 ( .B(n21400), .A(n21401), .Z(n21398) );
  XOR U23141 ( .A(n21399), .B(n21402), .Z(n21400) );
  IV U23142 ( .A(n21324), .Z(n21377) );
  XOR U23143 ( .A(n21403), .B(n21404), .Z(n21324) );
  XNOR U23144 ( .A(n21319), .B(n21405), .Z(n21404) );
  IV U23145 ( .A(n21322), .Z(n21405) );
  XOR U23146 ( .A(n21406), .B(n21407), .Z(n21322) );
  ANDN U23147 ( .B(n21408), .A(n21409), .Z(n21406) );
  XOR U23148 ( .A(n21410), .B(n21407), .Z(n21408) );
  XNOR U23149 ( .A(n21411), .B(n21412), .Z(n21319) );
  ANDN U23150 ( .B(n21413), .A(n21414), .Z(n21411) );
  XOR U23151 ( .A(n21412), .B(n21415), .Z(n21413) );
  IV U23152 ( .A(n21318), .Z(n21403) );
  XOR U23153 ( .A(n21316), .B(n21416), .Z(n21318) );
  XOR U23154 ( .A(n21417), .B(n21418), .Z(n21416) );
  ANDN U23155 ( .B(n21419), .A(n21420), .Z(n21417) );
  XOR U23156 ( .A(n21421), .B(n21418), .Z(n21419) );
  IV U23157 ( .A(n21320), .Z(n21316) );
  XOR U23158 ( .A(n21422), .B(n21423), .Z(n21320) );
  ANDN U23159 ( .B(n21424), .A(n21425), .Z(n21422) );
  XOR U23160 ( .A(n21426), .B(n21423), .Z(n21424) );
  IV U23161 ( .A(n21330), .Z(n21334) );
  XOR U23162 ( .A(n21330), .B(n21233), .Z(n21332) );
  XOR U23163 ( .A(n21427), .B(n21428), .Z(n21233) );
  AND U23164 ( .A(n196), .B(n21429), .Z(n21427) );
  XOR U23165 ( .A(n21430), .B(n21428), .Z(n21429) );
  NANDN U23166 ( .A(n21235), .B(n21237), .Z(n21330) );
  XOR U23167 ( .A(n21431), .B(n21432), .Z(n21237) );
  AND U23168 ( .A(n196), .B(n21433), .Z(n21431) );
  XOR U23169 ( .A(n21432), .B(n21434), .Z(n21433) );
  XNOR U23170 ( .A(n21435), .B(n21436), .Z(n196) );
  AND U23171 ( .A(n21437), .B(n21438), .Z(n21435) );
  XOR U23172 ( .A(n21436), .B(n21248), .Z(n21438) );
  XNOR U23173 ( .A(n21439), .B(n21440), .Z(n21248) );
  ANDN U23174 ( .B(n21441), .A(n21442), .Z(n21439) );
  XOR U23175 ( .A(n21440), .B(n21443), .Z(n21441) );
  XNOR U23176 ( .A(n21436), .B(n21250), .Z(n21437) );
  XOR U23177 ( .A(n21444), .B(n21445), .Z(n21250) );
  AND U23178 ( .A(n200), .B(n21446), .Z(n21444) );
  XOR U23179 ( .A(n21447), .B(n21445), .Z(n21446) );
  XOR U23180 ( .A(n21448), .B(n21449), .Z(n21436) );
  AND U23181 ( .A(n21450), .B(n21451), .Z(n21448) );
  XOR U23182 ( .A(n21449), .B(n21275), .Z(n21451) );
  XOR U23183 ( .A(n21442), .B(n21443), .Z(n21275) );
  XNOR U23184 ( .A(n21452), .B(n21453), .Z(n21443) );
  ANDN U23185 ( .B(n21454), .A(n21455), .Z(n21452) );
  XOR U23186 ( .A(n21456), .B(n21457), .Z(n21454) );
  XOR U23187 ( .A(n21458), .B(n21459), .Z(n21442) );
  XNOR U23188 ( .A(n21460), .B(n21461), .Z(n21459) );
  ANDN U23189 ( .B(n21462), .A(n21463), .Z(n21460) );
  XNOR U23190 ( .A(n21464), .B(n21465), .Z(n21462) );
  IV U23191 ( .A(n21440), .Z(n21458) );
  XOR U23192 ( .A(n21466), .B(n21467), .Z(n21440) );
  ANDN U23193 ( .B(n21468), .A(n21469), .Z(n21466) );
  XOR U23194 ( .A(n21467), .B(n21470), .Z(n21468) );
  XNOR U23195 ( .A(n21449), .B(n21277), .Z(n21450) );
  XOR U23196 ( .A(n21471), .B(n21472), .Z(n21277) );
  AND U23197 ( .A(n200), .B(n21473), .Z(n21471) );
  XOR U23198 ( .A(n21474), .B(n21472), .Z(n21473) );
  XNOR U23199 ( .A(n21475), .B(n21476), .Z(n21449) );
  AND U23200 ( .A(n21477), .B(n21478), .Z(n21475) );
  XNOR U23201 ( .A(n21476), .B(n21327), .Z(n21478) );
  XOR U23202 ( .A(n21469), .B(n21470), .Z(n21327) );
  XOR U23203 ( .A(n21479), .B(n21457), .Z(n21470) );
  XNOR U23204 ( .A(n21480), .B(n21481), .Z(n21457) );
  ANDN U23205 ( .B(n21482), .A(n21483), .Z(n21480) );
  XOR U23206 ( .A(n21484), .B(n21485), .Z(n21482) );
  IV U23207 ( .A(n21455), .Z(n21479) );
  XOR U23208 ( .A(n21453), .B(n21486), .Z(n21455) );
  XNOR U23209 ( .A(n21487), .B(n21488), .Z(n21486) );
  ANDN U23210 ( .B(n21489), .A(n21490), .Z(n21487) );
  XNOR U23211 ( .A(n21491), .B(n21492), .Z(n21489) );
  IV U23212 ( .A(n21456), .Z(n21453) );
  XOR U23213 ( .A(n21493), .B(n21494), .Z(n21456) );
  ANDN U23214 ( .B(n21495), .A(n21496), .Z(n21493) );
  XOR U23215 ( .A(n21494), .B(n21497), .Z(n21495) );
  XOR U23216 ( .A(n21498), .B(n21499), .Z(n21469) );
  XNOR U23217 ( .A(n21464), .B(n21500), .Z(n21499) );
  IV U23218 ( .A(n21467), .Z(n21500) );
  XOR U23219 ( .A(n21501), .B(n21502), .Z(n21467) );
  ANDN U23220 ( .B(n21503), .A(n21504), .Z(n21501) );
  XOR U23221 ( .A(n21502), .B(n21505), .Z(n21503) );
  XNOR U23222 ( .A(n21506), .B(n21507), .Z(n21464) );
  ANDN U23223 ( .B(n21508), .A(n21509), .Z(n21506) );
  XOR U23224 ( .A(n21507), .B(n21510), .Z(n21508) );
  IV U23225 ( .A(n21463), .Z(n21498) );
  XOR U23226 ( .A(n21461), .B(n21511), .Z(n21463) );
  XNOR U23227 ( .A(n21512), .B(n21513), .Z(n21511) );
  ANDN U23228 ( .B(n21514), .A(n21515), .Z(n21512) );
  XNOR U23229 ( .A(n21516), .B(n21517), .Z(n21514) );
  IV U23230 ( .A(n21465), .Z(n21461) );
  XOR U23231 ( .A(n21518), .B(n21519), .Z(n21465) );
  ANDN U23232 ( .B(n21520), .A(n21521), .Z(n21518) );
  XOR U23233 ( .A(n21522), .B(n21519), .Z(n21520) );
  XOR U23234 ( .A(n21476), .B(n21329), .Z(n21477) );
  XOR U23235 ( .A(n21523), .B(n21524), .Z(n21329) );
  AND U23236 ( .A(n200), .B(n21525), .Z(n21523) );
  XOR U23237 ( .A(n21526), .B(n21524), .Z(n21525) );
  XNOR U23238 ( .A(n21527), .B(n21528), .Z(n21476) );
  NAND U23239 ( .A(n21529), .B(n21530), .Z(n21528) );
  XOR U23240 ( .A(n21531), .B(n21428), .Z(n21530) );
  XOR U23241 ( .A(n21504), .B(n21505), .Z(n21428) );
  XOR U23242 ( .A(n21532), .B(n21497), .Z(n21505) );
  XOR U23243 ( .A(n21533), .B(n21485), .Z(n21497) );
  XOR U23244 ( .A(n21534), .B(n21535), .Z(n21485) );
  ANDN U23245 ( .B(n21536), .A(n21537), .Z(n21534) );
  XOR U23246 ( .A(n21535), .B(n21538), .Z(n21536) );
  IV U23247 ( .A(n21483), .Z(n21533) );
  XOR U23248 ( .A(n21481), .B(n21539), .Z(n21483) );
  XOR U23249 ( .A(n21540), .B(n21541), .Z(n21539) );
  ANDN U23250 ( .B(n21542), .A(n21543), .Z(n21540) );
  XOR U23251 ( .A(n21544), .B(n21541), .Z(n21542) );
  IV U23252 ( .A(n21484), .Z(n21481) );
  XOR U23253 ( .A(n21545), .B(n21546), .Z(n21484) );
  ANDN U23254 ( .B(n21547), .A(n21548), .Z(n21545) );
  XOR U23255 ( .A(n21546), .B(n21549), .Z(n21547) );
  IV U23256 ( .A(n21496), .Z(n21532) );
  XOR U23257 ( .A(n21550), .B(n21551), .Z(n21496) );
  XNOR U23258 ( .A(n21491), .B(n21552), .Z(n21551) );
  IV U23259 ( .A(n21494), .Z(n21552) );
  XOR U23260 ( .A(n21553), .B(n21554), .Z(n21494) );
  ANDN U23261 ( .B(n21555), .A(n21556), .Z(n21553) );
  XOR U23262 ( .A(n21554), .B(n21557), .Z(n21555) );
  XNOR U23263 ( .A(n21558), .B(n21559), .Z(n21491) );
  ANDN U23264 ( .B(n21560), .A(n21561), .Z(n21558) );
  XOR U23265 ( .A(n21559), .B(n21562), .Z(n21560) );
  IV U23266 ( .A(n21490), .Z(n21550) );
  XOR U23267 ( .A(n21488), .B(n21563), .Z(n21490) );
  XOR U23268 ( .A(n21564), .B(n21565), .Z(n21563) );
  ANDN U23269 ( .B(n21566), .A(n21567), .Z(n21564) );
  XOR U23270 ( .A(n21568), .B(n21565), .Z(n21566) );
  IV U23271 ( .A(n21492), .Z(n21488) );
  XOR U23272 ( .A(n21569), .B(n21570), .Z(n21492) );
  ANDN U23273 ( .B(n21571), .A(n21572), .Z(n21569) );
  XOR U23274 ( .A(n21573), .B(n21570), .Z(n21571) );
  XOR U23275 ( .A(n21574), .B(n21575), .Z(n21504) );
  XOR U23276 ( .A(n21522), .B(n21576), .Z(n21575) );
  IV U23277 ( .A(n21502), .Z(n21576) );
  XOR U23278 ( .A(n21577), .B(n21578), .Z(n21502) );
  ANDN U23279 ( .B(n21579), .A(n21580), .Z(n21577) );
  XOR U23280 ( .A(n21578), .B(n21581), .Z(n21579) );
  XOR U23281 ( .A(n21582), .B(n21510), .Z(n21522) );
  XOR U23282 ( .A(n21583), .B(n21584), .Z(n21510) );
  ANDN U23283 ( .B(n21585), .A(n21586), .Z(n21583) );
  XOR U23284 ( .A(n21584), .B(n21587), .Z(n21585) );
  IV U23285 ( .A(n21509), .Z(n21582) );
  XOR U23286 ( .A(n21588), .B(n21589), .Z(n21509) );
  XOR U23287 ( .A(n21590), .B(n21591), .Z(n21589) );
  ANDN U23288 ( .B(n21592), .A(n21593), .Z(n21590) );
  XOR U23289 ( .A(n21594), .B(n21591), .Z(n21592) );
  IV U23290 ( .A(n21507), .Z(n21588) );
  XOR U23291 ( .A(n21595), .B(n21596), .Z(n21507) );
  ANDN U23292 ( .B(n21597), .A(n21598), .Z(n21595) );
  XOR U23293 ( .A(n21596), .B(n21599), .Z(n21597) );
  IV U23294 ( .A(n21521), .Z(n21574) );
  XOR U23295 ( .A(n21600), .B(n21601), .Z(n21521) );
  XNOR U23296 ( .A(n21516), .B(n21602), .Z(n21601) );
  IV U23297 ( .A(n21519), .Z(n21602) );
  XOR U23298 ( .A(n21603), .B(n21604), .Z(n21519) );
  ANDN U23299 ( .B(n21605), .A(n21606), .Z(n21603) );
  XOR U23300 ( .A(n21607), .B(n21604), .Z(n21605) );
  XNOR U23301 ( .A(n21608), .B(n21609), .Z(n21516) );
  ANDN U23302 ( .B(n21610), .A(n21611), .Z(n21608) );
  XOR U23303 ( .A(n21609), .B(n21612), .Z(n21610) );
  IV U23304 ( .A(n21515), .Z(n21600) );
  XOR U23305 ( .A(n21513), .B(n21613), .Z(n21515) );
  XOR U23306 ( .A(n21614), .B(n21615), .Z(n21613) );
  ANDN U23307 ( .B(n21616), .A(n21617), .Z(n21614) );
  XOR U23308 ( .A(n21618), .B(n21615), .Z(n21616) );
  IV U23309 ( .A(n21517), .Z(n21513) );
  XOR U23310 ( .A(n21619), .B(n21620), .Z(n21517) );
  ANDN U23311 ( .B(n21621), .A(n21622), .Z(n21619) );
  XOR U23312 ( .A(n21623), .B(n21620), .Z(n21621) );
  IV U23313 ( .A(n21527), .Z(n21531) );
  XOR U23314 ( .A(n21527), .B(n21430), .Z(n21529) );
  XOR U23315 ( .A(n21624), .B(n21625), .Z(n21430) );
  AND U23316 ( .A(n200), .B(n21626), .Z(n21624) );
  XOR U23317 ( .A(n21627), .B(n21625), .Z(n21626) );
  NANDN U23318 ( .A(n21432), .B(n21434), .Z(n21527) );
  XOR U23319 ( .A(n21628), .B(n21629), .Z(n21434) );
  AND U23320 ( .A(n200), .B(n21630), .Z(n21628) );
  XOR U23321 ( .A(n21629), .B(n21631), .Z(n21630) );
  XNOR U23322 ( .A(n21632), .B(n21633), .Z(n200) );
  AND U23323 ( .A(n21634), .B(n21635), .Z(n21632) );
  XOR U23324 ( .A(n21633), .B(n21445), .Z(n21635) );
  XNOR U23325 ( .A(n21636), .B(n21637), .Z(n21445) );
  ANDN U23326 ( .B(n21638), .A(n21639), .Z(n21636) );
  XOR U23327 ( .A(n21637), .B(n21640), .Z(n21638) );
  XNOR U23328 ( .A(n21633), .B(n21447), .Z(n21634) );
  XOR U23329 ( .A(n21641), .B(n21642), .Z(n21447) );
  AND U23330 ( .A(n204), .B(n21643), .Z(n21641) );
  XOR U23331 ( .A(n21644), .B(n21642), .Z(n21643) );
  XOR U23332 ( .A(n21645), .B(n21646), .Z(n21633) );
  AND U23333 ( .A(n21647), .B(n21648), .Z(n21645) );
  XOR U23334 ( .A(n21646), .B(n21472), .Z(n21648) );
  XOR U23335 ( .A(n21639), .B(n21640), .Z(n21472) );
  XNOR U23336 ( .A(n21649), .B(n21650), .Z(n21640) );
  ANDN U23337 ( .B(n21651), .A(n21652), .Z(n21649) );
  XOR U23338 ( .A(n21653), .B(n21654), .Z(n21651) );
  XOR U23339 ( .A(n21655), .B(n21656), .Z(n21639) );
  XNOR U23340 ( .A(n21657), .B(n21658), .Z(n21656) );
  ANDN U23341 ( .B(n21659), .A(n21660), .Z(n21657) );
  XNOR U23342 ( .A(n21661), .B(n21662), .Z(n21659) );
  IV U23343 ( .A(n21637), .Z(n21655) );
  XOR U23344 ( .A(n21663), .B(n21664), .Z(n21637) );
  ANDN U23345 ( .B(n21665), .A(n21666), .Z(n21663) );
  XOR U23346 ( .A(n21664), .B(n21667), .Z(n21665) );
  XNOR U23347 ( .A(n21646), .B(n21474), .Z(n21647) );
  XOR U23348 ( .A(n21668), .B(n21669), .Z(n21474) );
  AND U23349 ( .A(n204), .B(n21670), .Z(n21668) );
  XOR U23350 ( .A(n21671), .B(n21669), .Z(n21670) );
  XNOR U23351 ( .A(n21672), .B(n21673), .Z(n21646) );
  AND U23352 ( .A(n21674), .B(n21675), .Z(n21672) );
  XNOR U23353 ( .A(n21673), .B(n21524), .Z(n21675) );
  XOR U23354 ( .A(n21666), .B(n21667), .Z(n21524) );
  XOR U23355 ( .A(n21676), .B(n21654), .Z(n21667) );
  XNOR U23356 ( .A(n21677), .B(n21678), .Z(n21654) );
  ANDN U23357 ( .B(n21679), .A(n21680), .Z(n21677) );
  XOR U23358 ( .A(n21681), .B(n21682), .Z(n21679) );
  IV U23359 ( .A(n21652), .Z(n21676) );
  XOR U23360 ( .A(n21650), .B(n21683), .Z(n21652) );
  XNOR U23361 ( .A(n21684), .B(n21685), .Z(n21683) );
  ANDN U23362 ( .B(n21686), .A(n21687), .Z(n21684) );
  XNOR U23363 ( .A(n21688), .B(n21689), .Z(n21686) );
  IV U23364 ( .A(n21653), .Z(n21650) );
  XOR U23365 ( .A(n21690), .B(n21691), .Z(n21653) );
  ANDN U23366 ( .B(n21692), .A(n21693), .Z(n21690) );
  XOR U23367 ( .A(n21691), .B(n21694), .Z(n21692) );
  XOR U23368 ( .A(n21695), .B(n21696), .Z(n21666) );
  XNOR U23369 ( .A(n21661), .B(n21697), .Z(n21696) );
  IV U23370 ( .A(n21664), .Z(n21697) );
  XOR U23371 ( .A(n21698), .B(n21699), .Z(n21664) );
  ANDN U23372 ( .B(n21700), .A(n21701), .Z(n21698) );
  XOR U23373 ( .A(n21699), .B(n21702), .Z(n21700) );
  XNOR U23374 ( .A(n21703), .B(n21704), .Z(n21661) );
  ANDN U23375 ( .B(n21705), .A(n21706), .Z(n21703) );
  XOR U23376 ( .A(n21704), .B(n21707), .Z(n21705) );
  IV U23377 ( .A(n21660), .Z(n21695) );
  XOR U23378 ( .A(n21658), .B(n21708), .Z(n21660) );
  XNOR U23379 ( .A(n21709), .B(n21710), .Z(n21708) );
  ANDN U23380 ( .B(n21711), .A(n21712), .Z(n21709) );
  XNOR U23381 ( .A(n21713), .B(n21714), .Z(n21711) );
  IV U23382 ( .A(n21662), .Z(n21658) );
  XOR U23383 ( .A(n21715), .B(n21716), .Z(n21662) );
  ANDN U23384 ( .B(n21717), .A(n21718), .Z(n21715) );
  XOR U23385 ( .A(n21719), .B(n21716), .Z(n21717) );
  XOR U23386 ( .A(n21673), .B(n21526), .Z(n21674) );
  XOR U23387 ( .A(n21720), .B(n21721), .Z(n21526) );
  AND U23388 ( .A(n204), .B(n21722), .Z(n21720) );
  XOR U23389 ( .A(n21723), .B(n21721), .Z(n21722) );
  XNOR U23390 ( .A(n21724), .B(n21725), .Z(n21673) );
  NAND U23391 ( .A(n21726), .B(n21727), .Z(n21725) );
  XOR U23392 ( .A(n21728), .B(n21625), .Z(n21727) );
  XOR U23393 ( .A(n21701), .B(n21702), .Z(n21625) );
  XOR U23394 ( .A(n21729), .B(n21694), .Z(n21702) );
  XOR U23395 ( .A(n21730), .B(n21682), .Z(n21694) );
  XOR U23396 ( .A(n21731), .B(n21732), .Z(n21682) );
  ANDN U23397 ( .B(n21733), .A(n21734), .Z(n21731) );
  XOR U23398 ( .A(n21732), .B(n21735), .Z(n21733) );
  IV U23399 ( .A(n21680), .Z(n21730) );
  XOR U23400 ( .A(n21678), .B(n21736), .Z(n21680) );
  XOR U23401 ( .A(n21737), .B(n21738), .Z(n21736) );
  ANDN U23402 ( .B(n21739), .A(n21740), .Z(n21737) );
  XOR U23403 ( .A(n21741), .B(n21738), .Z(n21739) );
  IV U23404 ( .A(n21681), .Z(n21678) );
  XOR U23405 ( .A(n21742), .B(n21743), .Z(n21681) );
  ANDN U23406 ( .B(n21744), .A(n21745), .Z(n21742) );
  XOR U23407 ( .A(n21743), .B(n21746), .Z(n21744) );
  IV U23408 ( .A(n21693), .Z(n21729) );
  XOR U23409 ( .A(n21747), .B(n21748), .Z(n21693) );
  XNOR U23410 ( .A(n21688), .B(n21749), .Z(n21748) );
  IV U23411 ( .A(n21691), .Z(n21749) );
  XOR U23412 ( .A(n21750), .B(n21751), .Z(n21691) );
  ANDN U23413 ( .B(n21752), .A(n21753), .Z(n21750) );
  XOR U23414 ( .A(n21751), .B(n21754), .Z(n21752) );
  XNOR U23415 ( .A(n21755), .B(n21756), .Z(n21688) );
  ANDN U23416 ( .B(n21757), .A(n21758), .Z(n21755) );
  XOR U23417 ( .A(n21756), .B(n21759), .Z(n21757) );
  IV U23418 ( .A(n21687), .Z(n21747) );
  XOR U23419 ( .A(n21685), .B(n21760), .Z(n21687) );
  XOR U23420 ( .A(n21761), .B(n21762), .Z(n21760) );
  ANDN U23421 ( .B(n21763), .A(n21764), .Z(n21761) );
  XOR U23422 ( .A(n21765), .B(n21762), .Z(n21763) );
  IV U23423 ( .A(n21689), .Z(n21685) );
  XOR U23424 ( .A(n21766), .B(n21767), .Z(n21689) );
  ANDN U23425 ( .B(n21768), .A(n21769), .Z(n21766) );
  XOR U23426 ( .A(n21770), .B(n21767), .Z(n21768) );
  XOR U23427 ( .A(n21771), .B(n21772), .Z(n21701) );
  XOR U23428 ( .A(n21719), .B(n21773), .Z(n21772) );
  IV U23429 ( .A(n21699), .Z(n21773) );
  XOR U23430 ( .A(n21774), .B(n21775), .Z(n21699) );
  ANDN U23431 ( .B(n21776), .A(n21777), .Z(n21774) );
  XOR U23432 ( .A(n21775), .B(n21778), .Z(n21776) );
  XOR U23433 ( .A(n21779), .B(n21707), .Z(n21719) );
  XOR U23434 ( .A(n21780), .B(n21781), .Z(n21707) );
  ANDN U23435 ( .B(n21782), .A(n21783), .Z(n21780) );
  XOR U23436 ( .A(n21781), .B(n21784), .Z(n21782) );
  IV U23437 ( .A(n21706), .Z(n21779) );
  XOR U23438 ( .A(n21785), .B(n21786), .Z(n21706) );
  XOR U23439 ( .A(n21787), .B(n21788), .Z(n21786) );
  ANDN U23440 ( .B(n21789), .A(n21790), .Z(n21787) );
  XOR U23441 ( .A(n21791), .B(n21788), .Z(n21789) );
  IV U23442 ( .A(n21704), .Z(n21785) );
  XOR U23443 ( .A(n21792), .B(n21793), .Z(n21704) );
  ANDN U23444 ( .B(n21794), .A(n21795), .Z(n21792) );
  XOR U23445 ( .A(n21793), .B(n21796), .Z(n21794) );
  IV U23446 ( .A(n21718), .Z(n21771) );
  XOR U23447 ( .A(n21797), .B(n21798), .Z(n21718) );
  XNOR U23448 ( .A(n21713), .B(n21799), .Z(n21798) );
  IV U23449 ( .A(n21716), .Z(n21799) );
  XOR U23450 ( .A(n21800), .B(n21801), .Z(n21716) );
  ANDN U23451 ( .B(n21802), .A(n21803), .Z(n21800) );
  XOR U23452 ( .A(n21804), .B(n21801), .Z(n21802) );
  XNOR U23453 ( .A(n21805), .B(n21806), .Z(n21713) );
  ANDN U23454 ( .B(n21807), .A(n21808), .Z(n21805) );
  XOR U23455 ( .A(n21806), .B(n21809), .Z(n21807) );
  IV U23456 ( .A(n21712), .Z(n21797) );
  XOR U23457 ( .A(n21710), .B(n21810), .Z(n21712) );
  XOR U23458 ( .A(n21811), .B(n21812), .Z(n21810) );
  ANDN U23459 ( .B(n21813), .A(n21814), .Z(n21811) );
  XOR U23460 ( .A(n21815), .B(n21812), .Z(n21813) );
  IV U23461 ( .A(n21714), .Z(n21710) );
  XOR U23462 ( .A(n21816), .B(n21817), .Z(n21714) );
  ANDN U23463 ( .B(n21818), .A(n21819), .Z(n21816) );
  XOR U23464 ( .A(n21820), .B(n21817), .Z(n21818) );
  IV U23465 ( .A(n21724), .Z(n21728) );
  XOR U23466 ( .A(n21724), .B(n21627), .Z(n21726) );
  XOR U23467 ( .A(n21821), .B(n21822), .Z(n21627) );
  AND U23468 ( .A(n204), .B(n21823), .Z(n21821) );
  XOR U23469 ( .A(n21824), .B(n21822), .Z(n21823) );
  NANDN U23470 ( .A(n21629), .B(n21631), .Z(n21724) );
  XOR U23471 ( .A(n21825), .B(n21826), .Z(n21631) );
  AND U23472 ( .A(n204), .B(n21827), .Z(n21825) );
  XOR U23473 ( .A(n21826), .B(n21828), .Z(n21827) );
  XNOR U23474 ( .A(n21829), .B(n21830), .Z(n204) );
  AND U23475 ( .A(n21831), .B(n21832), .Z(n21829) );
  XOR U23476 ( .A(n21830), .B(n21642), .Z(n21832) );
  XNOR U23477 ( .A(n21833), .B(n21834), .Z(n21642) );
  ANDN U23478 ( .B(n21835), .A(n21836), .Z(n21833) );
  XOR U23479 ( .A(n21834), .B(n21837), .Z(n21835) );
  XNOR U23480 ( .A(n21830), .B(n21644), .Z(n21831) );
  XOR U23481 ( .A(n21838), .B(n21839), .Z(n21644) );
  AND U23482 ( .A(n208), .B(n21840), .Z(n21838) );
  XOR U23483 ( .A(n21841), .B(n21839), .Z(n21840) );
  XOR U23484 ( .A(n21842), .B(n21843), .Z(n21830) );
  AND U23485 ( .A(n21844), .B(n21845), .Z(n21842) );
  XOR U23486 ( .A(n21843), .B(n21669), .Z(n21845) );
  XOR U23487 ( .A(n21836), .B(n21837), .Z(n21669) );
  XNOR U23488 ( .A(n21846), .B(n21847), .Z(n21837) );
  ANDN U23489 ( .B(n21848), .A(n21849), .Z(n21846) );
  XOR U23490 ( .A(n21850), .B(n21851), .Z(n21848) );
  XOR U23491 ( .A(n21852), .B(n21853), .Z(n21836) );
  XNOR U23492 ( .A(n21854), .B(n21855), .Z(n21853) );
  ANDN U23493 ( .B(n21856), .A(n21857), .Z(n21854) );
  XNOR U23494 ( .A(n21858), .B(n21859), .Z(n21856) );
  IV U23495 ( .A(n21834), .Z(n21852) );
  XOR U23496 ( .A(n21860), .B(n21861), .Z(n21834) );
  ANDN U23497 ( .B(n21862), .A(n21863), .Z(n21860) );
  XOR U23498 ( .A(n21861), .B(n21864), .Z(n21862) );
  XNOR U23499 ( .A(n21843), .B(n21671), .Z(n21844) );
  XOR U23500 ( .A(n21865), .B(n21866), .Z(n21671) );
  AND U23501 ( .A(n208), .B(n21867), .Z(n21865) );
  XOR U23502 ( .A(n21868), .B(n21866), .Z(n21867) );
  XNOR U23503 ( .A(n21869), .B(n21870), .Z(n21843) );
  AND U23504 ( .A(n21871), .B(n21872), .Z(n21869) );
  XNOR U23505 ( .A(n21870), .B(n21721), .Z(n21872) );
  XOR U23506 ( .A(n21863), .B(n21864), .Z(n21721) );
  XOR U23507 ( .A(n21873), .B(n21851), .Z(n21864) );
  XNOR U23508 ( .A(n21874), .B(n21875), .Z(n21851) );
  ANDN U23509 ( .B(n21876), .A(n21877), .Z(n21874) );
  XOR U23510 ( .A(n21878), .B(n21879), .Z(n21876) );
  IV U23511 ( .A(n21849), .Z(n21873) );
  XOR U23512 ( .A(n21847), .B(n21880), .Z(n21849) );
  XNOR U23513 ( .A(n21881), .B(n21882), .Z(n21880) );
  ANDN U23514 ( .B(n21883), .A(n21884), .Z(n21881) );
  XNOR U23515 ( .A(n21885), .B(n21886), .Z(n21883) );
  IV U23516 ( .A(n21850), .Z(n21847) );
  XOR U23517 ( .A(n21887), .B(n21888), .Z(n21850) );
  ANDN U23518 ( .B(n21889), .A(n21890), .Z(n21887) );
  XOR U23519 ( .A(n21888), .B(n21891), .Z(n21889) );
  XOR U23520 ( .A(n21892), .B(n21893), .Z(n21863) );
  XNOR U23521 ( .A(n21858), .B(n21894), .Z(n21893) );
  IV U23522 ( .A(n21861), .Z(n21894) );
  XOR U23523 ( .A(n21895), .B(n21896), .Z(n21861) );
  ANDN U23524 ( .B(n21897), .A(n21898), .Z(n21895) );
  XOR U23525 ( .A(n21896), .B(n21899), .Z(n21897) );
  XNOR U23526 ( .A(n21900), .B(n21901), .Z(n21858) );
  ANDN U23527 ( .B(n21902), .A(n21903), .Z(n21900) );
  XOR U23528 ( .A(n21901), .B(n21904), .Z(n21902) );
  IV U23529 ( .A(n21857), .Z(n21892) );
  XOR U23530 ( .A(n21855), .B(n21905), .Z(n21857) );
  XNOR U23531 ( .A(n21906), .B(n21907), .Z(n21905) );
  ANDN U23532 ( .B(n21908), .A(n21909), .Z(n21906) );
  XNOR U23533 ( .A(n21910), .B(n21911), .Z(n21908) );
  IV U23534 ( .A(n21859), .Z(n21855) );
  XOR U23535 ( .A(n21912), .B(n21913), .Z(n21859) );
  ANDN U23536 ( .B(n21914), .A(n21915), .Z(n21912) );
  XOR U23537 ( .A(n21916), .B(n21913), .Z(n21914) );
  XOR U23538 ( .A(n21870), .B(n21723), .Z(n21871) );
  XOR U23539 ( .A(n21917), .B(n21918), .Z(n21723) );
  AND U23540 ( .A(n208), .B(n21919), .Z(n21917) );
  XOR U23541 ( .A(n21920), .B(n21918), .Z(n21919) );
  XNOR U23542 ( .A(n21921), .B(n21922), .Z(n21870) );
  NAND U23543 ( .A(n21923), .B(n21924), .Z(n21922) );
  XOR U23544 ( .A(n21925), .B(n21822), .Z(n21924) );
  XOR U23545 ( .A(n21898), .B(n21899), .Z(n21822) );
  XOR U23546 ( .A(n21926), .B(n21891), .Z(n21899) );
  XOR U23547 ( .A(n21927), .B(n21879), .Z(n21891) );
  XOR U23548 ( .A(n21928), .B(n21929), .Z(n21879) );
  ANDN U23549 ( .B(n21930), .A(n21931), .Z(n21928) );
  XOR U23550 ( .A(n21929), .B(n21932), .Z(n21930) );
  IV U23551 ( .A(n21877), .Z(n21927) );
  XOR U23552 ( .A(n21875), .B(n21933), .Z(n21877) );
  XOR U23553 ( .A(n21934), .B(n21935), .Z(n21933) );
  ANDN U23554 ( .B(n21936), .A(n21937), .Z(n21934) );
  XOR U23555 ( .A(n21938), .B(n21935), .Z(n21936) );
  IV U23556 ( .A(n21878), .Z(n21875) );
  XOR U23557 ( .A(n21939), .B(n21940), .Z(n21878) );
  ANDN U23558 ( .B(n21941), .A(n21942), .Z(n21939) );
  XOR U23559 ( .A(n21940), .B(n21943), .Z(n21941) );
  IV U23560 ( .A(n21890), .Z(n21926) );
  XOR U23561 ( .A(n21944), .B(n21945), .Z(n21890) );
  XNOR U23562 ( .A(n21885), .B(n21946), .Z(n21945) );
  IV U23563 ( .A(n21888), .Z(n21946) );
  XOR U23564 ( .A(n21947), .B(n21948), .Z(n21888) );
  ANDN U23565 ( .B(n21949), .A(n21950), .Z(n21947) );
  XOR U23566 ( .A(n21948), .B(n21951), .Z(n21949) );
  XNOR U23567 ( .A(n21952), .B(n21953), .Z(n21885) );
  ANDN U23568 ( .B(n21954), .A(n21955), .Z(n21952) );
  XOR U23569 ( .A(n21953), .B(n21956), .Z(n21954) );
  IV U23570 ( .A(n21884), .Z(n21944) );
  XOR U23571 ( .A(n21882), .B(n21957), .Z(n21884) );
  XOR U23572 ( .A(n21958), .B(n21959), .Z(n21957) );
  ANDN U23573 ( .B(n21960), .A(n21961), .Z(n21958) );
  XOR U23574 ( .A(n21962), .B(n21959), .Z(n21960) );
  IV U23575 ( .A(n21886), .Z(n21882) );
  XOR U23576 ( .A(n21963), .B(n21964), .Z(n21886) );
  ANDN U23577 ( .B(n21965), .A(n21966), .Z(n21963) );
  XOR U23578 ( .A(n21967), .B(n21964), .Z(n21965) );
  XOR U23579 ( .A(n21968), .B(n21969), .Z(n21898) );
  XOR U23580 ( .A(n21916), .B(n21970), .Z(n21969) );
  IV U23581 ( .A(n21896), .Z(n21970) );
  XOR U23582 ( .A(n21971), .B(n21972), .Z(n21896) );
  ANDN U23583 ( .B(n21973), .A(n21974), .Z(n21971) );
  XOR U23584 ( .A(n21972), .B(n21975), .Z(n21973) );
  XOR U23585 ( .A(n21976), .B(n21904), .Z(n21916) );
  XOR U23586 ( .A(n21977), .B(n21978), .Z(n21904) );
  ANDN U23587 ( .B(n21979), .A(n21980), .Z(n21977) );
  XOR U23588 ( .A(n21978), .B(n21981), .Z(n21979) );
  IV U23589 ( .A(n21903), .Z(n21976) );
  XOR U23590 ( .A(n21982), .B(n21983), .Z(n21903) );
  XOR U23591 ( .A(n21984), .B(n21985), .Z(n21983) );
  ANDN U23592 ( .B(n21986), .A(n21987), .Z(n21984) );
  XOR U23593 ( .A(n21988), .B(n21985), .Z(n21986) );
  IV U23594 ( .A(n21901), .Z(n21982) );
  XOR U23595 ( .A(n21989), .B(n21990), .Z(n21901) );
  ANDN U23596 ( .B(n21991), .A(n21992), .Z(n21989) );
  XOR U23597 ( .A(n21990), .B(n21993), .Z(n21991) );
  IV U23598 ( .A(n21915), .Z(n21968) );
  XOR U23599 ( .A(n21994), .B(n21995), .Z(n21915) );
  XNOR U23600 ( .A(n21910), .B(n21996), .Z(n21995) );
  IV U23601 ( .A(n21913), .Z(n21996) );
  XOR U23602 ( .A(n21997), .B(n21998), .Z(n21913) );
  ANDN U23603 ( .B(n21999), .A(n22000), .Z(n21997) );
  XOR U23604 ( .A(n22001), .B(n21998), .Z(n21999) );
  XNOR U23605 ( .A(n22002), .B(n22003), .Z(n21910) );
  ANDN U23606 ( .B(n22004), .A(n22005), .Z(n22002) );
  XOR U23607 ( .A(n22003), .B(n22006), .Z(n22004) );
  IV U23608 ( .A(n21909), .Z(n21994) );
  XOR U23609 ( .A(n21907), .B(n22007), .Z(n21909) );
  XOR U23610 ( .A(n22008), .B(n22009), .Z(n22007) );
  ANDN U23611 ( .B(n22010), .A(n22011), .Z(n22008) );
  XOR U23612 ( .A(n22012), .B(n22009), .Z(n22010) );
  IV U23613 ( .A(n21911), .Z(n21907) );
  XOR U23614 ( .A(n22013), .B(n22014), .Z(n21911) );
  ANDN U23615 ( .B(n22015), .A(n22016), .Z(n22013) );
  XOR U23616 ( .A(n22017), .B(n22014), .Z(n22015) );
  IV U23617 ( .A(n21921), .Z(n21925) );
  XOR U23618 ( .A(n21921), .B(n21824), .Z(n21923) );
  XOR U23619 ( .A(n22018), .B(n22019), .Z(n21824) );
  AND U23620 ( .A(n208), .B(n22020), .Z(n22018) );
  XOR U23621 ( .A(n22021), .B(n22019), .Z(n22020) );
  NANDN U23622 ( .A(n21826), .B(n21828), .Z(n21921) );
  XOR U23623 ( .A(n22022), .B(n22023), .Z(n21828) );
  AND U23624 ( .A(n208), .B(n22024), .Z(n22022) );
  XOR U23625 ( .A(n22023), .B(n22025), .Z(n22024) );
  XNOR U23626 ( .A(n22026), .B(n22027), .Z(n208) );
  AND U23627 ( .A(n22028), .B(n22029), .Z(n22026) );
  XOR U23628 ( .A(n22027), .B(n21839), .Z(n22029) );
  XNOR U23629 ( .A(n22030), .B(n22031), .Z(n21839) );
  ANDN U23630 ( .B(n22032), .A(n22033), .Z(n22030) );
  XOR U23631 ( .A(n22031), .B(n22034), .Z(n22032) );
  XNOR U23632 ( .A(n22027), .B(n21841), .Z(n22028) );
  XOR U23633 ( .A(n22035), .B(n22036), .Z(n21841) );
  AND U23634 ( .A(n212), .B(n22037), .Z(n22035) );
  XOR U23635 ( .A(n22038), .B(n22036), .Z(n22037) );
  XOR U23636 ( .A(n22039), .B(n22040), .Z(n22027) );
  AND U23637 ( .A(n22041), .B(n22042), .Z(n22039) );
  XOR U23638 ( .A(n22040), .B(n21866), .Z(n22042) );
  XOR U23639 ( .A(n22033), .B(n22034), .Z(n21866) );
  XNOR U23640 ( .A(n22043), .B(n22044), .Z(n22034) );
  ANDN U23641 ( .B(n22045), .A(n22046), .Z(n22043) );
  XOR U23642 ( .A(n22047), .B(n22048), .Z(n22045) );
  XOR U23643 ( .A(n22049), .B(n22050), .Z(n22033) );
  XNOR U23644 ( .A(n22051), .B(n22052), .Z(n22050) );
  ANDN U23645 ( .B(n22053), .A(n22054), .Z(n22051) );
  XNOR U23646 ( .A(n22055), .B(n22056), .Z(n22053) );
  IV U23647 ( .A(n22031), .Z(n22049) );
  XOR U23648 ( .A(n22057), .B(n22058), .Z(n22031) );
  ANDN U23649 ( .B(n22059), .A(n22060), .Z(n22057) );
  XOR U23650 ( .A(n22058), .B(n22061), .Z(n22059) );
  XNOR U23651 ( .A(n22040), .B(n21868), .Z(n22041) );
  XOR U23652 ( .A(n22062), .B(n22063), .Z(n21868) );
  AND U23653 ( .A(n212), .B(n22064), .Z(n22062) );
  XOR U23654 ( .A(n22065), .B(n22063), .Z(n22064) );
  XNOR U23655 ( .A(n22066), .B(n22067), .Z(n22040) );
  AND U23656 ( .A(n22068), .B(n22069), .Z(n22066) );
  XNOR U23657 ( .A(n22067), .B(n21918), .Z(n22069) );
  XOR U23658 ( .A(n22060), .B(n22061), .Z(n21918) );
  XOR U23659 ( .A(n22070), .B(n22048), .Z(n22061) );
  XNOR U23660 ( .A(n22071), .B(n22072), .Z(n22048) );
  ANDN U23661 ( .B(n22073), .A(n22074), .Z(n22071) );
  XOR U23662 ( .A(n22075), .B(n22076), .Z(n22073) );
  IV U23663 ( .A(n22046), .Z(n22070) );
  XOR U23664 ( .A(n22044), .B(n22077), .Z(n22046) );
  XNOR U23665 ( .A(n22078), .B(n22079), .Z(n22077) );
  ANDN U23666 ( .B(n22080), .A(n22081), .Z(n22078) );
  XNOR U23667 ( .A(n22082), .B(n22083), .Z(n22080) );
  IV U23668 ( .A(n22047), .Z(n22044) );
  XOR U23669 ( .A(n22084), .B(n22085), .Z(n22047) );
  ANDN U23670 ( .B(n22086), .A(n22087), .Z(n22084) );
  XOR U23671 ( .A(n22085), .B(n22088), .Z(n22086) );
  XOR U23672 ( .A(n22089), .B(n22090), .Z(n22060) );
  XNOR U23673 ( .A(n22055), .B(n22091), .Z(n22090) );
  IV U23674 ( .A(n22058), .Z(n22091) );
  XOR U23675 ( .A(n22092), .B(n22093), .Z(n22058) );
  ANDN U23676 ( .B(n22094), .A(n22095), .Z(n22092) );
  XOR U23677 ( .A(n22093), .B(n22096), .Z(n22094) );
  XNOR U23678 ( .A(n22097), .B(n22098), .Z(n22055) );
  ANDN U23679 ( .B(n22099), .A(n22100), .Z(n22097) );
  XOR U23680 ( .A(n22098), .B(n22101), .Z(n22099) );
  IV U23681 ( .A(n22054), .Z(n22089) );
  XOR U23682 ( .A(n22052), .B(n22102), .Z(n22054) );
  XNOR U23683 ( .A(n22103), .B(n22104), .Z(n22102) );
  ANDN U23684 ( .B(n22105), .A(n22106), .Z(n22103) );
  XNOR U23685 ( .A(n22107), .B(n22108), .Z(n22105) );
  IV U23686 ( .A(n22056), .Z(n22052) );
  XOR U23687 ( .A(n22109), .B(n22110), .Z(n22056) );
  ANDN U23688 ( .B(n22111), .A(n22112), .Z(n22109) );
  XOR U23689 ( .A(n22113), .B(n22110), .Z(n22111) );
  XOR U23690 ( .A(n22067), .B(n21920), .Z(n22068) );
  XOR U23691 ( .A(n22114), .B(n22115), .Z(n21920) );
  AND U23692 ( .A(n212), .B(n22116), .Z(n22114) );
  XOR U23693 ( .A(n22117), .B(n22115), .Z(n22116) );
  XNOR U23694 ( .A(n22118), .B(n22119), .Z(n22067) );
  NAND U23695 ( .A(n22120), .B(n22121), .Z(n22119) );
  XOR U23696 ( .A(n22122), .B(n22019), .Z(n22121) );
  XOR U23697 ( .A(n22095), .B(n22096), .Z(n22019) );
  XOR U23698 ( .A(n22123), .B(n22088), .Z(n22096) );
  XOR U23699 ( .A(n22124), .B(n22076), .Z(n22088) );
  XOR U23700 ( .A(n22125), .B(n22126), .Z(n22076) );
  ANDN U23701 ( .B(n22127), .A(n22128), .Z(n22125) );
  XOR U23702 ( .A(n22126), .B(n22129), .Z(n22127) );
  IV U23703 ( .A(n22074), .Z(n22124) );
  XOR U23704 ( .A(n22072), .B(n22130), .Z(n22074) );
  XOR U23705 ( .A(n22131), .B(n22132), .Z(n22130) );
  ANDN U23706 ( .B(n22133), .A(n22134), .Z(n22131) );
  XOR U23707 ( .A(n22135), .B(n22132), .Z(n22133) );
  IV U23708 ( .A(n22075), .Z(n22072) );
  XOR U23709 ( .A(n22136), .B(n22137), .Z(n22075) );
  ANDN U23710 ( .B(n22138), .A(n22139), .Z(n22136) );
  XOR U23711 ( .A(n22137), .B(n22140), .Z(n22138) );
  IV U23712 ( .A(n22087), .Z(n22123) );
  XOR U23713 ( .A(n22141), .B(n22142), .Z(n22087) );
  XNOR U23714 ( .A(n22082), .B(n22143), .Z(n22142) );
  IV U23715 ( .A(n22085), .Z(n22143) );
  XOR U23716 ( .A(n22144), .B(n22145), .Z(n22085) );
  ANDN U23717 ( .B(n22146), .A(n22147), .Z(n22144) );
  XOR U23718 ( .A(n22145), .B(n22148), .Z(n22146) );
  XNOR U23719 ( .A(n22149), .B(n22150), .Z(n22082) );
  ANDN U23720 ( .B(n22151), .A(n22152), .Z(n22149) );
  XOR U23721 ( .A(n22150), .B(n22153), .Z(n22151) );
  IV U23722 ( .A(n22081), .Z(n22141) );
  XOR U23723 ( .A(n22079), .B(n22154), .Z(n22081) );
  XOR U23724 ( .A(n22155), .B(n22156), .Z(n22154) );
  ANDN U23725 ( .B(n22157), .A(n22158), .Z(n22155) );
  XOR U23726 ( .A(n22159), .B(n22156), .Z(n22157) );
  IV U23727 ( .A(n22083), .Z(n22079) );
  XOR U23728 ( .A(n22160), .B(n22161), .Z(n22083) );
  ANDN U23729 ( .B(n22162), .A(n22163), .Z(n22160) );
  XOR U23730 ( .A(n22164), .B(n22161), .Z(n22162) );
  XOR U23731 ( .A(n22165), .B(n22166), .Z(n22095) );
  XOR U23732 ( .A(n22113), .B(n22167), .Z(n22166) );
  IV U23733 ( .A(n22093), .Z(n22167) );
  XOR U23734 ( .A(n22168), .B(n22169), .Z(n22093) );
  ANDN U23735 ( .B(n22170), .A(n22171), .Z(n22168) );
  XOR U23736 ( .A(n22169), .B(n22172), .Z(n22170) );
  XOR U23737 ( .A(n22173), .B(n22101), .Z(n22113) );
  XOR U23738 ( .A(n22174), .B(n22175), .Z(n22101) );
  ANDN U23739 ( .B(n22176), .A(n22177), .Z(n22174) );
  XOR U23740 ( .A(n22175), .B(n22178), .Z(n22176) );
  IV U23741 ( .A(n22100), .Z(n22173) );
  XOR U23742 ( .A(n22179), .B(n22180), .Z(n22100) );
  XOR U23743 ( .A(n22181), .B(n22182), .Z(n22180) );
  ANDN U23744 ( .B(n22183), .A(n22184), .Z(n22181) );
  XOR U23745 ( .A(n22185), .B(n22182), .Z(n22183) );
  IV U23746 ( .A(n22098), .Z(n22179) );
  XOR U23747 ( .A(n22186), .B(n22187), .Z(n22098) );
  ANDN U23748 ( .B(n22188), .A(n22189), .Z(n22186) );
  XOR U23749 ( .A(n22187), .B(n22190), .Z(n22188) );
  IV U23750 ( .A(n22112), .Z(n22165) );
  XOR U23751 ( .A(n22191), .B(n22192), .Z(n22112) );
  XNOR U23752 ( .A(n22107), .B(n22193), .Z(n22192) );
  IV U23753 ( .A(n22110), .Z(n22193) );
  XOR U23754 ( .A(n22194), .B(n22195), .Z(n22110) );
  ANDN U23755 ( .B(n22196), .A(n22197), .Z(n22194) );
  XOR U23756 ( .A(n22198), .B(n22195), .Z(n22196) );
  XNOR U23757 ( .A(n22199), .B(n22200), .Z(n22107) );
  ANDN U23758 ( .B(n22201), .A(n22202), .Z(n22199) );
  XOR U23759 ( .A(n22200), .B(n22203), .Z(n22201) );
  IV U23760 ( .A(n22106), .Z(n22191) );
  XOR U23761 ( .A(n22104), .B(n22204), .Z(n22106) );
  XOR U23762 ( .A(n22205), .B(n22206), .Z(n22204) );
  ANDN U23763 ( .B(n22207), .A(n22208), .Z(n22205) );
  XOR U23764 ( .A(n22209), .B(n22206), .Z(n22207) );
  IV U23765 ( .A(n22108), .Z(n22104) );
  XOR U23766 ( .A(n22210), .B(n22211), .Z(n22108) );
  ANDN U23767 ( .B(n22212), .A(n22213), .Z(n22210) );
  XOR U23768 ( .A(n22214), .B(n22211), .Z(n22212) );
  IV U23769 ( .A(n22118), .Z(n22122) );
  XOR U23770 ( .A(n22118), .B(n22021), .Z(n22120) );
  XOR U23771 ( .A(n22215), .B(n22216), .Z(n22021) );
  AND U23772 ( .A(n212), .B(n22217), .Z(n22215) );
  XOR U23773 ( .A(n22218), .B(n22216), .Z(n22217) );
  NANDN U23774 ( .A(n22023), .B(n22025), .Z(n22118) );
  XOR U23775 ( .A(n22219), .B(n22220), .Z(n22025) );
  AND U23776 ( .A(n212), .B(n22221), .Z(n22219) );
  XOR U23777 ( .A(n22220), .B(n22222), .Z(n22221) );
  XNOR U23778 ( .A(n22223), .B(n22224), .Z(n212) );
  AND U23779 ( .A(n22225), .B(n22226), .Z(n22223) );
  XOR U23780 ( .A(n22224), .B(n22036), .Z(n22226) );
  XNOR U23781 ( .A(n22227), .B(n22228), .Z(n22036) );
  ANDN U23782 ( .B(n22229), .A(n22230), .Z(n22227) );
  XOR U23783 ( .A(n22228), .B(n22231), .Z(n22229) );
  XNOR U23784 ( .A(n22224), .B(n22038), .Z(n22225) );
  XOR U23785 ( .A(n22232), .B(n22233), .Z(n22038) );
  AND U23786 ( .A(n216), .B(n22234), .Z(n22232) );
  XOR U23787 ( .A(n22235), .B(n22233), .Z(n22234) );
  XOR U23788 ( .A(n22236), .B(n22237), .Z(n22224) );
  AND U23789 ( .A(n22238), .B(n22239), .Z(n22236) );
  XOR U23790 ( .A(n22237), .B(n22063), .Z(n22239) );
  XOR U23791 ( .A(n22230), .B(n22231), .Z(n22063) );
  XNOR U23792 ( .A(n22240), .B(n22241), .Z(n22231) );
  ANDN U23793 ( .B(n22242), .A(n22243), .Z(n22240) );
  XOR U23794 ( .A(n22244), .B(n22245), .Z(n22242) );
  XOR U23795 ( .A(n22246), .B(n22247), .Z(n22230) );
  XNOR U23796 ( .A(n22248), .B(n22249), .Z(n22247) );
  ANDN U23797 ( .B(n22250), .A(n22251), .Z(n22248) );
  XNOR U23798 ( .A(n22252), .B(n22253), .Z(n22250) );
  IV U23799 ( .A(n22228), .Z(n22246) );
  XOR U23800 ( .A(n22254), .B(n22255), .Z(n22228) );
  ANDN U23801 ( .B(n22256), .A(n22257), .Z(n22254) );
  XOR U23802 ( .A(n22255), .B(n22258), .Z(n22256) );
  XNOR U23803 ( .A(n22237), .B(n22065), .Z(n22238) );
  XOR U23804 ( .A(n22259), .B(n22260), .Z(n22065) );
  AND U23805 ( .A(n216), .B(n22261), .Z(n22259) );
  XOR U23806 ( .A(n22262), .B(n22260), .Z(n22261) );
  XNOR U23807 ( .A(n22263), .B(n22264), .Z(n22237) );
  AND U23808 ( .A(n22265), .B(n22266), .Z(n22263) );
  XNOR U23809 ( .A(n22264), .B(n22115), .Z(n22266) );
  XOR U23810 ( .A(n22257), .B(n22258), .Z(n22115) );
  XOR U23811 ( .A(n22267), .B(n22245), .Z(n22258) );
  XNOR U23812 ( .A(n22268), .B(n22269), .Z(n22245) );
  ANDN U23813 ( .B(n22270), .A(n22271), .Z(n22268) );
  XOR U23814 ( .A(n22272), .B(n22273), .Z(n22270) );
  IV U23815 ( .A(n22243), .Z(n22267) );
  XOR U23816 ( .A(n22241), .B(n22274), .Z(n22243) );
  XNOR U23817 ( .A(n22275), .B(n22276), .Z(n22274) );
  ANDN U23818 ( .B(n22277), .A(n22278), .Z(n22275) );
  XNOR U23819 ( .A(n22279), .B(n22280), .Z(n22277) );
  IV U23820 ( .A(n22244), .Z(n22241) );
  XOR U23821 ( .A(n22281), .B(n22282), .Z(n22244) );
  ANDN U23822 ( .B(n22283), .A(n22284), .Z(n22281) );
  XOR U23823 ( .A(n22282), .B(n22285), .Z(n22283) );
  XOR U23824 ( .A(n22286), .B(n22287), .Z(n22257) );
  XNOR U23825 ( .A(n22252), .B(n22288), .Z(n22287) );
  IV U23826 ( .A(n22255), .Z(n22288) );
  XOR U23827 ( .A(n22289), .B(n22290), .Z(n22255) );
  ANDN U23828 ( .B(n22291), .A(n22292), .Z(n22289) );
  XOR U23829 ( .A(n22290), .B(n22293), .Z(n22291) );
  XNOR U23830 ( .A(n22294), .B(n22295), .Z(n22252) );
  ANDN U23831 ( .B(n22296), .A(n22297), .Z(n22294) );
  XOR U23832 ( .A(n22295), .B(n22298), .Z(n22296) );
  IV U23833 ( .A(n22251), .Z(n22286) );
  XOR U23834 ( .A(n22249), .B(n22299), .Z(n22251) );
  XNOR U23835 ( .A(n22300), .B(n22301), .Z(n22299) );
  ANDN U23836 ( .B(n22302), .A(n22303), .Z(n22300) );
  XNOR U23837 ( .A(n22304), .B(n22305), .Z(n22302) );
  IV U23838 ( .A(n22253), .Z(n22249) );
  XOR U23839 ( .A(n22306), .B(n22307), .Z(n22253) );
  ANDN U23840 ( .B(n22308), .A(n22309), .Z(n22306) );
  XOR U23841 ( .A(n22310), .B(n22307), .Z(n22308) );
  XOR U23842 ( .A(n22264), .B(n22117), .Z(n22265) );
  XOR U23843 ( .A(n22311), .B(n22312), .Z(n22117) );
  AND U23844 ( .A(n216), .B(n22313), .Z(n22311) );
  XOR U23845 ( .A(n22314), .B(n22312), .Z(n22313) );
  XNOR U23846 ( .A(n22315), .B(n22316), .Z(n22264) );
  NAND U23847 ( .A(n22317), .B(n22318), .Z(n22316) );
  XOR U23848 ( .A(n22319), .B(n22216), .Z(n22318) );
  XOR U23849 ( .A(n22292), .B(n22293), .Z(n22216) );
  XOR U23850 ( .A(n22320), .B(n22285), .Z(n22293) );
  XOR U23851 ( .A(n22321), .B(n22273), .Z(n22285) );
  XOR U23852 ( .A(n22322), .B(n22323), .Z(n22273) );
  ANDN U23853 ( .B(n22324), .A(n22325), .Z(n22322) );
  XOR U23854 ( .A(n22323), .B(n22326), .Z(n22324) );
  IV U23855 ( .A(n22271), .Z(n22321) );
  XOR U23856 ( .A(n22269), .B(n22327), .Z(n22271) );
  XOR U23857 ( .A(n22328), .B(n22329), .Z(n22327) );
  ANDN U23858 ( .B(n22330), .A(n22331), .Z(n22328) );
  XOR U23859 ( .A(n22332), .B(n22329), .Z(n22330) );
  IV U23860 ( .A(n22272), .Z(n22269) );
  XOR U23861 ( .A(n22333), .B(n22334), .Z(n22272) );
  ANDN U23862 ( .B(n22335), .A(n22336), .Z(n22333) );
  XOR U23863 ( .A(n22334), .B(n22337), .Z(n22335) );
  IV U23864 ( .A(n22284), .Z(n22320) );
  XOR U23865 ( .A(n22338), .B(n22339), .Z(n22284) );
  XNOR U23866 ( .A(n22279), .B(n22340), .Z(n22339) );
  IV U23867 ( .A(n22282), .Z(n22340) );
  XOR U23868 ( .A(n22341), .B(n22342), .Z(n22282) );
  ANDN U23869 ( .B(n22343), .A(n22344), .Z(n22341) );
  XOR U23870 ( .A(n22342), .B(n22345), .Z(n22343) );
  XNOR U23871 ( .A(n22346), .B(n22347), .Z(n22279) );
  ANDN U23872 ( .B(n22348), .A(n22349), .Z(n22346) );
  XOR U23873 ( .A(n22347), .B(n22350), .Z(n22348) );
  IV U23874 ( .A(n22278), .Z(n22338) );
  XOR U23875 ( .A(n22276), .B(n22351), .Z(n22278) );
  XOR U23876 ( .A(n22352), .B(n22353), .Z(n22351) );
  ANDN U23877 ( .B(n22354), .A(n22355), .Z(n22352) );
  XOR U23878 ( .A(n22356), .B(n22353), .Z(n22354) );
  IV U23879 ( .A(n22280), .Z(n22276) );
  XOR U23880 ( .A(n22357), .B(n22358), .Z(n22280) );
  ANDN U23881 ( .B(n22359), .A(n22360), .Z(n22357) );
  XOR U23882 ( .A(n22361), .B(n22358), .Z(n22359) );
  XOR U23883 ( .A(n22362), .B(n22363), .Z(n22292) );
  XOR U23884 ( .A(n22310), .B(n22364), .Z(n22363) );
  IV U23885 ( .A(n22290), .Z(n22364) );
  XOR U23886 ( .A(n22365), .B(n22366), .Z(n22290) );
  ANDN U23887 ( .B(n22367), .A(n22368), .Z(n22365) );
  XOR U23888 ( .A(n22366), .B(n22369), .Z(n22367) );
  XOR U23889 ( .A(n22370), .B(n22298), .Z(n22310) );
  XOR U23890 ( .A(n22371), .B(n22372), .Z(n22298) );
  ANDN U23891 ( .B(n22373), .A(n22374), .Z(n22371) );
  XOR U23892 ( .A(n22372), .B(n22375), .Z(n22373) );
  IV U23893 ( .A(n22297), .Z(n22370) );
  XOR U23894 ( .A(n22376), .B(n22377), .Z(n22297) );
  XOR U23895 ( .A(n22378), .B(n22379), .Z(n22377) );
  ANDN U23896 ( .B(n22380), .A(n22381), .Z(n22378) );
  XOR U23897 ( .A(n22382), .B(n22379), .Z(n22380) );
  IV U23898 ( .A(n22295), .Z(n22376) );
  XOR U23899 ( .A(n22383), .B(n22384), .Z(n22295) );
  ANDN U23900 ( .B(n22385), .A(n22386), .Z(n22383) );
  XOR U23901 ( .A(n22384), .B(n22387), .Z(n22385) );
  IV U23902 ( .A(n22309), .Z(n22362) );
  XOR U23903 ( .A(n22388), .B(n22389), .Z(n22309) );
  XNOR U23904 ( .A(n22304), .B(n22390), .Z(n22389) );
  IV U23905 ( .A(n22307), .Z(n22390) );
  XOR U23906 ( .A(n22391), .B(n22392), .Z(n22307) );
  ANDN U23907 ( .B(n22393), .A(n22394), .Z(n22391) );
  XOR U23908 ( .A(n22395), .B(n22392), .Z(n22393) );
  XNOR U23909 ( .A(n22396), .B(n22397), .Z(n22304) );
  ANDN U23910 ( .B(n22398), .A(n22399), .Z(n22396) );
  XOR U23911 ( .A(n22397), .B(n22400), .Z(n22398) );
  IV U23912 ( .A(n22303), .Z(n22388) );
  XOR U23913 ( .A(n22301), .B(n22401), .Z(n22303) );
  XOR U23914 ( .A(n22402), .B(n22403), .Z(n22401) );
  ANDN U23915 ( .B(n22404), .A(n22405), .Z(n22402) );
  XOR U23916 ( .A(n22406), .B(n22403), .Z(n22404) );
  IV U23917 ( .A(n22305), .Z(n22301) );
  XOR U23918 ( .A(n22407), .B(n22408), .Z(n22305) );
  ANDN U23919 ( .B(n22409), .A(n22410), .Z(n22407) );
  XOR U23920 ( .A(n22411), .B(n22408), .Z(n22409) );
  IV U23921 ( .A(n22315), .Z(n22319) );
  XOR U23922 ( .A(n22315), .B(n22218), .Z(n22317) );
  XOR U23923 ( .A(n22412), .B(n22413), .Z(n22218) );
  AND U23924 ( .A(n216), .B(n22414), .Z(n22412) );
  XOR U23925 ( .A(n22415), .B(n22413), .Z(n22414) );
  NANDN U23926 ( .A(n22220), .B(n22222), .Z(n22315) );
  XOR U23927 ( .A(n22416), .B(n22417), .Z(n22222) );
  AND U23928 ( .A(n216), .B(n22418), .Z(n22416) );
  XOR U23929 ( .A(n22417), .B(n22419), .Z(n22418) );
  XNOR U23930 ( .A(n22420), .B(n22421), .Z(n216) );
  AND U23931 ( .A(n22422), .B(n22423), .Z(n22420) );
  XOR U23932 ( .A(n22421), .B(n22233), .Z(n22423) );
  XNOR U23933 ( .A(n22424), .B(n22425), .Z(n22233) );
  ANDN U23934 ( .B(n22426), .A(n22427), .Z(n22424) );
  XOR U23935 ( .A(n22425), .B(n22428), .Z(n22426) );
  XNOR U23936 ( .A(n22421), .B(n22235), .Z(n22422) );
  XOR U23937 ( .A(n22429), .B(n22430), .Z(n22235) );
  AND U23938 ( .A(n220), .B(n22431), .Z(n22429) );
  XOR U23939 ( .A(n22432), .B(n22430), .Z(n22431) );
  XOR U23940 ( .A(n22433), .B(n22434), .Z(n22421) );
  AND U23941 ( .A(n22435), .B(n22436), .Z(n22433) );
  XOR U23942 ( .A(n22434), .B(n22260), .Z(n22436) );
  XOR U23943 ( .A(n22427), .B(n22428), .Z(n22260) );
  XNOR U23944 ( .A(n22437), .B(n22438), .Z(n22428) );
  ANDN U23945 ( .B(n22439), .A(n22440), .Z(n22437) );
  XOR U23946 ( .A(n22441), .B(n22442), .Z(n22439) );
  XOR U23947 ( .A(n22443), .B(n22444), .Z(n22427) );
  XNOR U23948 ( .A(n22445), .B(n22446), .Z(n22444) );
  ANDN U23949 ( .B(n22447), .A(n22448), .Z(n22445) );
  XNOR U23950 ( .A(n22449), .B(n22450), .Z(n22447) );
  IV U23951 ( .A(n22425), .Z(n22443) );
  XOR U23952 ( .A(n22451), .B(n22452), .Z(n22425) );
  ANDN U23953 ( .B(n22453), .A(n22454), .Z(n22451) );
  XOR U23954 ( .A(n22452), .B(n22455), .Z(n22453) );
  XNOR U23955 ( .A(n22434), .B(n22262), .Z(n22435) );
  XOR U23956 ( .A(n22456), .B(n22457), .Z(n22262) );
  AND U23957 ( .A(n220), .B(n22458), .Z(n22456) );
  XOR U23958 ( .A(n22459), .B(n22457), .Z(n22458) );
  XNOR U23959 ( .A(n22460), .B(n22461), .Z(n22434) );
  AND U23960 ( .A(n22462), .B(n22463), .Z(n22460) );
  XNOR U23961 ( .A(n22461), .B(n22312), .Z(n22463) );
  XOR U23962 ( .A(n22454), .B(n22455), .Z(n22312) );
  XOR U23963 ( .A(n22464), .B(n22442), .Z(n22455) );
  XNOR U23964 ( .A(n22465), .B(n22466), .Z(n22442) );
  ANDN U23965 ( .B(n22467), .A(n22468), .Z(n22465) );
  XOR U23966 ( .A(n22469), .B(n22470), .Z(n22467) );
  IV U23967 ( .A(n22440), .Z(n22464) );
  XOR U23968 ( .A(n22438), .B(n22471), .Z(n22440) );
  XNOR U23969 ( .A(n22472), .B(n22473), .Z(n22471) );
  ANDN U23970 ( .B(n22474), .A(n22475), .Z(n22472) );
  XNOR U23971 ( .A(n22476), .B(n22477), .Z(n22474) );
  IV U23972 ( .A(n22441), .Z(n22438) );
  XOR U23973 ( .A(n22478), .B(n22479), .Z(n22441) );
  ANDN U23974 ( .B(n22480), .A(n22481), .Z(n22478) );
  XOR U23975 ( .A(n22479), .B(n22482), .Z(n22480) );
  XOR U23976 ( .A(n22483), .B(n22484), .Z(n22454) );
  XNOR U23977 ( .A(n22449), .B(n22485), .Z(n22484) );
  IV U23978 ( .A(n22452), .Z(n22485) );
  XOR U23979 ( .A(n22486), .B(n22487), .Z(n22452) );
  ANDN U23980 ( .B(n22488), .A(n22489), .Z(n22486) );
  XOR U23981 ( .A(n22487), .B(n22490), .Z(n22488) );
  XNOR U23982 ( .A(n22491), .B(n22492), .Z(n22449) );
  ANDN U23983 ( .B(n22493), .A(n22494), .Z(n22491) );
  XOR U23984 ( .A(n22492), .B(n22495), .Z(n22493) );
  IV U23985 ( .A(n22448), .Z(n22483) );
  XOR U23986 ( .A(n22446), .B(n22496), .Z(n22448) );
  XNOR U23987 ( .A(n22497), .B(n22498), .Z(n22496) );
  ANDN U23988 ( .B(n22499), .A(n22500), .Z(n22497) );
  XNOR U23989 ( .A(n22501), .B(n22502), .Z(n22499) );
  IV U23990 ( .A(n22450), .Z(n22446) );
  XOR U23991 ( .A(n22503), .B(n22504), .Z(n22450) );
  ANDN U23992 ( .B(n22505), .A(n22506), .Z(n22503) );
  XOR U23993 ( .A(n22507), .B(n22504), .Z(n22505) );
  XOR U23994 ( .A(n22461), .B(n22314), .Z(n22462) );
  XOR U23995 ( .A(n22508), .B(n22509), .Z(n22314) );
  AND U23996 ( .A(n220), .B(n22510), .Z(n22508) );
  XOR U23997 ( .A(n22511), .B(n22509), .Z(n22510) );
  XNOR U23998 ( .A(n22512), .B(n22513), .Z(n22461) );
  NAND U23999 ( .A(n22514), .B(n22515), .Z(n22513) );
  XOR U24000 ( .A(n22516), .B(n22413), .Z(n22515) );
  XOR U24001 ( .A(n22489), .B(n22490), .Z(n22413) );
  XOR U24002 ( .A(n22517), .B(n22482), .Z(n22490) );
  XOR U24003 ( .A(n22518), .B(n22470), .Z(n22482) );
  XOR U24004 ( .A(n22519), .B(n22520), .Z(n22470) );
  ANDN U24005 ( .B(n22521), .A(n22522), .Z(n22519) );
  XOR U24006 ( .A(n22520), .B(n22523), .Z(n22521) );
  IV U24007 ( .A(n22468), .Z(n22518) );
  XOR U24008 ( .A(n22466), .B(n22524), .Z(n22468) );
  XOR U24009 ( .A(n22525), .B(n22526), .Z(n22524) );
  ANDN U24010 ( .B(n22527), .A(n22528), .Z(n22525) );
  XOR U24011 ( .A(n22529), .B(n22526), .Z(n22527) );
  IV U24012 ( .A(n22469), .Z(n22466) );
  XOR U24013 ( .A(n22530), .B(n22531), .Z(n22469) );
  ANDN U24014 ( .B(n22532), .A(n22533), .Z(n22530) );
  XOR U24015 ( .A(n22531), .B(n22534), .Z(n22532) );
  IV U24016 ( .A(n22481), .Z(n22517) );
  XOR U24017 ( .A(n22535), .B(n22536), .Z(n22481) );
  XNOR U24018 ( .A(n22476), .B(n22537), .Z(n22536) );
  IV U24019 ( .A(n22479), .Z(n22537) );
  XOR U24020 ( .A(n22538), .B(n22539), .Z(n22479) );
  ANDN U24021 ( .B(n22540), .A(n22541), .Z(n22538) );
  XOR U24022 ( .A(n22539), .B(n22542), .Z(n22540) );
  XNOR U24023 ( .A(n22543), .B(n22544), .Z(n22476) );
  ANDN U24024 ( .B(n22545), .A(n22546), .Z(n22543) );
  XOR U24025 ( .A(n22544), .B(n22547), .Z(n22545) );
  IV U24026 ( .A(n22475), .Z(n22535) );
  XOR U24027 ( .A(n22473), .B(n22548), .Z(n22475) );
  XOR U24028 ( .A(n22549), .B(n22550), .Z(n22548) );
  ANDN U24029 ( .B(n22551), .A(n22552), .Z(n22549) );
  XOR U24030 ( .A(n22553), .B(n22550), .Z(n22551) );
  IV U24031 ( .A(n22477), .Z(n22473) );
  XOR U24032 ( .A(n22554), .B(n22555), .Z(n22477) );
  ANDN U24033 ( .B(n22556), .A(n22557), .Z(n22554) );
  XOR U24034 ( .A(n22558), .B(n22555), .Z(n22556) );
  XOR U24035 ( .A(n22559), .B(n22560), .Z(n22489) );
  XOR U24036 ( .A(n22507), .B(n22561), .Z(n22560) );
  IV U24037 ( .A(n22487), .Z(n22561) );
  XOR U24038 ( .A(n22562), .B(n22563), .Z(n22487) );
  ANDN U24039 ( .B(n22564), .A(n22565), .Z(n22562) );
  XOR U24040 ( .A(n22563), .B(n22566), .Z(n22564) );
  XOR U24041 ( .A(n22567), .B(n22495), .Z(n22507) );
  XOR U24042 ( .A(n22568), .B(n22569), .Z(n22495) );
  ANDN U24043 ( .B(n22570), .A(n22571), .Z(n22568) );
  XOR U24044 ( .A(n22569), .B(n22572), .Z(n22570) );
  IV U24045 ( .A(n22494), .Z(n22567) );
  XOR U24046 ( .A(n22573), .B(n22574), .Z(n22494) );
  XOR U24047 ( .A(n22575), .B(n22576), .Z(n22574) );
  ANDN U24048 ( .B(n22577), .A(n22578), .Z(n22575) );
  XOR U24049 ( .A(n22579), .B(n22576), .Z(n22577) );
  IV U24050 ( .A(n22492), .Z(n22573) );
  XOR U24051 ( .A(n22580), .B(n22581), .Z(n22492) );
  ANDN U24052 ( .B(n22582), .A(n22583), .Z(n22580) );
  XOR U24053 ( .A(n22581), .B(n22584), .Z(n22582) );
  IV U24054 ( .A(n22506), .Z(n22559) );
  XOR U24055 ( .A(n22585), .B(n22586), .Z(n22506) );
  XNOR U24056 ( .A(n22501), .B(n22587), .Z(n22586) );
  IV U24057 ( .A(n22504), .Z(n22587) );
  XOR U24058 ( .A(n22588), .B(n22589), .Z(n22504) );
  ANDN U24059 ( .B(n22590), .A(n22591), .Z(n22588) );
  XOR U24060 ( .A(n22592), .B(n22589), .Z(n22590) );
  XNOR U24061 ( .A(n22593), .B(n22594), .Z(n22501) );
  ANDN U24062 ( .B(n22595), .A(n22596), .Z(n22593) );
  XOR U24063 ( .A(n22594), .B(n22597), .Z(n22595) );
  IV U24064 ( .A(n22500), .Z(n22585) );
  XOR U24065 ( .A(n22498), .B(n22598), .Z(n22500) );
  XOR U24066 ( .A(n22599), .B(n22600), .Z(n22598) );
  ANDN U24067 ( .B(n22601), .A(n22602), .Z(n22599) );
  XOR U24068 ( .A(n22603), .B(n22600), .Z(n22601) );
  IV U24069 ( .A(n22502), .Z(n22498) );
  XOR U24070 ( .A(n22604), .B(n22605), .Z(n22502) );
  ANDN U24071 ( .B(n22606), .A(n22607), .Z(n22604) );
  XOR U24072 ( .A(n22608), .B(n22605), .Z(n22606) );
  IV U24073 ( .A(n22512), .Z(n22516) );
  XOR U24074 ( .A(n22512), .B(n22415), .Z(n22514) );
  XOR U24075 ( .A(n22609), .B(n22610), .Z(n22415) );
  AND U24076 ( .A(n220), .B(n22611), .Z(n22609) );
  XOR U24077 ( .A(n22612), .B(n22610), .Z(n22611) );
  NANDN U24078 ( .A(n22417), .B(n22419), .Z(n22512) );
  XOR U24079 ( .A(n22613), .B(n22614), .Z(n22419) );
  AND U24080 ( .A(n220), .B(n22615), .Z(n22613) );
  XOR U24081 ( .A(n22614), .B(n22616), .Z(n22615) );
  XNOR U24082 ( .A(n22617), .B(n22618), .Z(n220) );
  AND U24083 ( .A(n22619), .B(n22620), .Z(n22617) );
  XOR U24084 ( .A(n22618), .B(n22430), .Z(n22620) );
  XNOR U24085 ( .A(n22621), .B(n22622), .Z(n22430) );
  ANDN U24086 ( .B(n22623), .A(n22624), .Z(n22621) );
  XOR U24087 ( .A(n22622), .B(n22625), .Z(n22623) );
  XNOR U24088 ( .A(n22618), .B(n22432), .Z(n22619) );
  XOR U24089 ( .A(n22626), .B(n22627), .Z(n22432) );
  AND U24090 ( .A(n224), .B(n22628), .Z(n22626) );
  XOR U24091 ( .A(n22629), .B(n22627), .Z(n22628) );
  XOR U24092 ( .A(n22630), .B(n22631), .Z(n22618) );
  AND U24093 ( .A(n22632), .B(n22633), .Z(n22630) );
  XOR U24094 ( .A(n22631), .B(n22457), .Z(n22633) );
  XOR U24095 ( .A(n22624), .B(n22625), .Z(n22457) );
  XNOR U24096 ( .A(n22634), .B(n22635), .Z(n22625) );
  ANDN U24097 ( .B(n22636), .A(n22637), .Z(n22634) );
  XOR U24098 ( .A(n22638), .B(n22639), .Z(n22636) );
  XOR U24099 ( .A(n22640), .B(n22641), .Z(n22624) );
  XNOR U24100 ( .A(n22642), .B(n22643), .Z(n22641) );
  ANDN U24101 ( .B(n22644), .A(n22645), .Z(n22642) );
  XNOR U24102 ( .A(n22646), .B(n22647), .Z(n22644) );
  IV U24103 ( .A(n22622), .Z(n22640) );
  XOR U24104 ( .A(n22648), .B(n22649), .Z(n22622) );
  ANDN U24105 ( .B(n22650), .A(n22651), .Z(n22648) );
  XOR U24106 ( .A(n22649), .B(n22652), .Z(n22650) );
  XNOR U24107 ( .A(n22631), .B(n22459), .Z(n22632) );
  XOR U24108 ( .A(n22653), .B(n22654), .Z(n22459) );
  AND U24109 ( .A(n224), .B(n22655), .Z(n22653) );
  XOR U24110 ( .A(n22656), .B(n22654), .Z(n22655) );
  XNOR U24111 ( .A(n22657), .B(n22658), .Z(n22631) );
  AND U24112 ( .A(n22659), .B(n22660), .Z(n22657) );
  XNOR U24113 ( .A(n22658), .B(n22509), .Z(n22660) );
  XOR U24114 ( .A(n22651), .B(n22652), .Z(n22509) );
  XOR U24115 ( .A(n22661), .B(n22639), .Z(n22652) );
  XNOR U24116 ( .A(n22662), .B(n22663), .Z(n22639) );
  ANDN U24117 ( .B(n22664), .A(n22665), .Z(n22662) );
  XOR U24118 ( .A(n22666), .B(n22667), .Z(n22664) );
  IV U24119 ( .A(n22637), .Z(n22661) );
  XOR U24120 ( .A(n22635), .B(n22668), .Z(n22637) );
  XNOR U24121 ( .A(n22669), .B(n22670), .Z(n22668) );
  ANDN U24122 ( .B(n22671), .A(n22672), .Z(n22669) );
  XNOR U24123 ( .A(n22673), .B(n22674), .Z(n22671) );
  IV U24124 ( .A(n22638), .Z(n22635) );
  XOR U24125 ( .A(n22675), .B(n22676), .Z(n22638) );
  ANDN U24126 ( .B(n22677), .A(n22678), .Z(n22675) );
  XOR U24127 ( .A(n22676), .B(n22679), .Z(n22677) );
  XOR U24128 ( .A(n22680), .B(n22681), .Z(n22651) );
  XNOR U24129 ( .A(n22646), .B(n22682), .Z(n22681) );
  IV U24130 ( .A(n22649), .Z(n22682) );
  XOR U24131 ( .A(n22683), .B(n22684), .Z(n22649) );
  ANDN U24132 ( .B(n22685), .A(n22686), .Z(n22683) );
  XOR U24133 ( .A(n22684), .B(n22687), .Z(n22685) );
  XNOR U24134 ( .A(n22688), .B(n22689), .Z(n22646) );
  ANDN U24135 ( .B(n22690), .A(n22691), .Z(n22688) );
  XOR U24136 ( .A(n22689), .B(n22692), .Z(n22690) );
  IV U24137 ( .A(n22645), .Z(n22680) );
  XOR U24138 ( .A(n22643), .B(n22693), .Z(n22645) );
  XNOR U24139 ( .A(n22694), .B(n22695), .Z(n22693) );
  ANDN U24140 ( .B(n22696), .A(n22697), .Z(n22694) );
  XNOR U24141 ( .A(n22698), .B(n22699), .Z(n22696) );
  IV U24142 ( .A(n22647), .Z(n22643) );
  XOR U24143 ( .A(n22700), .B(n22701), .Z(n22647) );
  ANDN U24144 ( .B(n22702), .A(n22703), .Z(n22700) );
  XOR U24145 ( .A(n22704), .B(n22701), .Z(n22702) );
  XOR U24146 ( .A(n22658), .B(n22511), .Z(n22659) );
  XOR U24147 ( .A(n22705), .B(n22706), .Z(n22511) );
  AND U24148 ( .A(n224), .B(n22707), .Z(n22705) );
  XOR U24149 ( .A(n22708), .B(n22706), .Z(n22707) );
  XNOR U24150 ( .A(n22709), .B(n22710), .Z(n22658) );
  NAND U24151 ( .A(n22711), .B(n22712), .Z(n22710) );
  XOR U24152 ( .A(n22713), .B(n22610), .Z(n22712) );
  XOR U24153 ( .A(n22686), .B(n22687), .Z(n22610) );
  XOR U24154 ( .A(n22714), .B(n22679), .Z(n22687) );
  XOR U24155 ( .A(n22715), .B(n22667), .Z(n22679) );
  XOR U24156 ( .A(n22716), .B(n22717), .Z(n22667) );
  ANDN U24157 ( .B(n22718), .A(n22719), .Z(n22716) );
  XOR U24158 ( .A(n22717), .B(n22720), .Z(n22718) );
  IV U24159 ( .A(n22665), .Z(n22715) );
  XOR U24160 ( .A(n22663), .B(n22721), .Z(n22665) );
  XOR U24161 ( .A(n22722), .B(n22723), .Z(n22721) );
  ANDN U24162 ( .B(n22724), .A(n22725), .Z(n22722) );
  XOR U24163 ( .A(n22726), .B(n22723), .Z(n22724) );
  IV U24164 ( .A(n22666), .Z(n22663) );
  XOR U24165 ( .A(n22727), .B(n22728), .Z(n22666) );
  ANDN U24166 ( .B(n22729), .A(n22730), .Z(n22727) );
  XOR U24167 ( .A(n22728), .B(n22731), .Z(n22729) );
  IV U24168 ( .A(n22678), .Z(n22714) );
  XOR U24169 ( .A(n22732), .B(n22733), .Z(n22678) );
  XNOR U24170 ( .A(n22673), .B(n22734), .Z(n22733) );
  IV U24171 ( .A(n22676), .Z(n22734) );
  XOR U24172 ( .A(n22735), .B(n22736), .Z(n22676) );
  ANDN U24173 ( .B(n22737), .A(n22738), .Z(n22735) );
  XOR U24174 ( .A(n22736), .B(n22739), .Z(n22737) );
  XNOR U24175 ( .A(n22740), .B(n22741), .Z(n22673) );
  ANDN U24176 ( .B(n22742), .A(n22743), .Z(n22740) );
  XOR U24177 ( .A(n22741), .B(n22744), .Z(n22742) );
  IV U24178 ( .A(n22672), .Z(n22732) );
  XOR U24179 ( .A(n22670), .B(n22745), .Z(n22672) );
  XOR U24180 ( .A(n22746), .B(n22747), .Z(n22745) );
  ANDN U24181 ( .B(n22748), .A(n22749), .Z(n22746) );
  XOR U24182 ( .A(n22750), .B(n22747), .Z(n22748) );
  IV U24183 ( .A(n22674), .Z(n22670) );
  XOR U24184 ( .A(n22751), .B(n22752), .Z(n22674) );
  ANDN U24185 ( .B(n22753), .A(n22754), .Z(n22751) );
  XOR U24186 ( .A(n22755), .B(n22752), .Z(n22753) );
  XOR U24187 ( .A(n22756), .B(n22757), .Z(n22686) );
  XOR U24188 ( .A(n22704), .B(n22758), .Z(n22757) );
  IV U24189 ( .A(n22684), .Z(n22758) );
  XOR U24190 ( .A(n22759), .B(n22760), .Z(n22684) );
  ANDN U24191 ( .B(n22761), .A(n22762), .Z(n22759) );
  XOR U24192 ( .A(n22760), .B(n22763), .Z(n22761) );
  XOR U24193 ( .A(n22764), .B(n22692), .Z(n22704) );
  XOR U24194 ( .A(n22765), .B(n22766), .Z(n22692) );
  ANDN U24195 ( .B(n22767), .A(n22768), .Z(n22765) );
  XOR U24196 ( .A(n22766), .B(n22769), .Z(n22767) );
  IV U24197 ( .A(n22691), .Z(n22764) );
  XOR U24198 ( .A(n22770), .B(n22771), .Z(n22691) );
  XOR U24199 ( .A(n22772), .B(n22773), .Z(n22771) );
  ANDN U24200 ( .B(n22774), .A(n22775), .Z(n22772) );
  XOR U24201 ( .A(n22776), .B(n22773), .Z(n22774) );
  IV U24202 ( .A(n22689), .Z(n22770) );
  XOR U24203 ( .A(n22777), .B(n22778), .Z(n22689) );
  ANDN U24204 ( .B(n22779), .A(n22780), .Z(n22777) );
  XOR U24205 ( .A(n22778), .B(n22781), .Z(n22779) );
  IV U24206 ( .A(n22703), .Z(n22756) );
  XOR U24207 ( .A(n22782), .B(n22783), .Z(n22703) );
  XNOR U24208 ( .A(n22698), .B(n22784), .Z(n22783) );
  IV U24209 ( .A(n22701), .Z(n22784) );
  XOR U24210 ( .A(n22785), .B(n22786), .Z(n22701) );
  ANDN U24211 ( .B(n22787), .A(n22788), .Z(n22785) );
  XOR U24212 ( .A(n22789), .B(n22786), .Z(n22787) );
  XNOR U24213 ( .A(n22790), .B(n22791), .Z(n22698) );
  ANDN U24214 ( .B(n22792), .A(n22793), .Z(n22790) );
  XOR U24215 ( .A(n22791), .B(n22794), .Z(n22792) );
  IV U24216 ( .A(n22697), .Z(n22782) );
  XOR U24217 ( .A(n22695), .B(n22795), .Z(n22697) );
  XOR U24218 ( .A(n22796), .B(n22797), .Z(n22795) );
  ANDN U24219 ( .B(n22798), .A(n22799), .Z(n22796) );
  XOR U24220 ( .A(n22800), .B(n22797), .Z(n22798) );
  IV U24221 ( .A(n22699), .Z(n22695) );
  XOR U24222 ( .A(n22801), .B(n22802), .Z(n22699) );
  ANDN U24223 ( .B(n22803), .A(n22804), .Z(n22801) );
  XOR U24224 ( .A(n22805), .B(n22802), .Z(n22803) );
  IV U24225 ( .A(n22709), .Z(n22713) );
  XOR U24226 ( .A(n22709), .B(n22612), .Z(n22711) );
  XOR U24227 ( .A(n22806), .B(n22807), .Z(n22612) );
  AND U24228 ( .A(n224), .B(n22808), .Z(n22806) );
  XOR U24229 ( .A(n22809), .B(n22807), .Z(n22808) );
  NANDN U24230 ( .A(n22614), .B(n22616), .Z(n22709) );
  XOR U24231 ( .A(n22810), .B(n22811), .Z(n22616) );
  AND U24232 ( .A(n224), .B(n22812), .Z(n22810) );
  XOR U24233 ( .A(n22811), .B(n22813), .Z(n22812) );
  XNOR U24234 ( .A(n22814), .B(n22815), .Z(n224) );
  AND U24235 ( .A(n22816), .B(n22817), .Z(n22814) );
  XOR U24236 ( .A(n22815), .B(n22627), .Z(n22817) );
  XNOR U24237 ( .A(n22818), .B(n22819), .Z(n22627) );
  ANDN U24238 ( .B(n22820), .A(n22821), .Z(n22818) );
  XOR U24239 ( .A(n22819), .B(n22822), .Z(n22820) );
  XNOR U24240 ( .A(n22815), .B(n22629), .Z(n22816) );
  XOR U24241 ( .A(n22823), .B(n22824), .Z(n22629) );
  AND U24242 ( .A(n228), .B(n22825), .Z(n22823) );
  XOR U24243 ( .A(n22826), .B(n22824), .Z(n22825) );
  XOR U24244 ( .A(n22827), .B(n22828), .Z(n22815) );
  AND U24245 ( .A(n22829), .B(n22830), .Z(n22827) );
  XOR U24246 ( .A(n22828), .B(n22654), .Z(n22830) );
  XOR U24247 ( .A(n22821), .B(n22822), .Z(n22654) );
  XNOR U24248 ( .A(n22831), .B(n22832), .Z(n22822) );
  ANDN U24249 ( .B(n22833), .A(n22834), .Z(n22831) );
  XOR U24250 ( .A(n22835), .B(n22836), .Z(n22833) );
  XOR U24251 ( .A(n22837), .B(n22838), .Z(n22821) );
  XNOR U24252 ( .A(n22839), .B(n22840), .Z(n22838) );
  ANDN U24253 ( .B(n22841), .A(n22842), .Z(n22839) );
  XNOR U24254 ( .A(n22843), .B(n22844), .Z(n22841) );
  IV U24255 ( .A(n22819), .Z(n22837) );
  XOR U24256 ( .A(n22845), .B(n22846), .Z(n22819) );
  ANDN U24257 ( .B(n22847), .A(n22848), .Z(n22845) );
  XOR U24258 ( .A(n22846), .B(n22849), .Z(n22847) );
  XNOR U24259 ( .A(n22828), .B(n22656), .Z(n22829) );
  XOR U24260 ( .A(n22850), .B(n22851), .Z(n22656) );
  AND U24261 ( .A(n228), .B(n22852), .Z(n22850) );
  XOR U24262 ( .A(n22853), .B(n22851), .Z(n22852) );
  XNOR U24263 ( .A(n22854), .B(n22855), .Z(n22828) );
  AND U24264 ( .A(n22856), .B(n22857), .Z(n22854) );
  XNOR U24265 ( .A(n22855), .B(n22706), .Z(n22857) );
  XOR U24266 ( .A(n22848), .B(n22849), .Z(n22706) );
  XOR U24267 ( .A(n22858), .B(n22836), .Z(n22849) );
  XNOR U24268 ( .A(n22859), .B(n22860), .Z(n22836) );
  ANDN U24269 ( .B(n22861), .A(n22862), .Z(n22859) );
  XOR U24270 ( .A(n22863), .B(n22864), .Z(n22861) );
  IV U24271 ( .A(n22834), .Z(n22858) );
  XOR U24272 ( .A(n22832), .B(n22865), .Z(n22834) );
  XNOR U24273 ( .A(n22866), .B(n22867), .Z(n22865) );
  ANDN U24274 ( .B(n22868), .A(n22869), .Z(n22866) );
  XNOR U24275 ( .A(n22870), .B(n22871), .Z(n22868) );
  IV U24276 ( .A(n22835), .Z(n22832) );
  XOR U24277 ( .A(n22872), .B(n22873), .Z(n22835) );
  ANDN U24278 ( .B(n22874), .A(n22875), .Z(n22872) );
  XOR U24279 ( .A(n22873), .B(n22876), .Z(n22874) );
  XOR U24280 ( .A(n22877), .B(n22878), .Z(n22848) );
  XNOR U24281 ( .A(n22843), .B(n22879), .Z(n22878) );
  IV U24282 ( .A(n22846), .Z(n22879) );
  XOR U24283 ( .A(n22880), .B(n22881), .Z(n22846) );
  ANDN U24284 ( .B(n22882), .A(n22883), .Z(n22880) );
  XOR U24285 ( .A(n22881), .B(n22884), .Z(n22882) );
  XNOR U24286 ( .A(n22885), .B(n22886), .Z(n22843) );
  ANDN U24287 ( .B(n22887), .A(n22888), .Z(n22885) );
  XOR U24288 ( .A(n22886), .B(n22889), .Z(n22887) );
  IV U24289 ( .A(n22842), .Z(n22877) );
  XOR U24290 ( .A(n22840), .B(n22890), .Z(n22842) );
  XNOR U24291 ( .A(n22891), .B(n22892), .Z(n22890) );
  ANDN U24292 ( .B(n22893), .A(n22894), .Z(n22891) );
  XNOR U24293 ( .A(n22895), .B(n22896), .Z(n22893) );
  IV U24294 ( .A(n22844), .Z(n22840) );
  XOR U24295 ( .A(n22897), .B(n22898), .Z(n22844) );
  ANDN U24296 ( .B(n22899), .A(n22900), .Z(n22897) );
  XOR U24297 ( .A(n22901), .B(n22898), .Z(n22899) );
  XOR U24298 ( .A(n22855), .B(n22708), .Z(n22856) );
  XOR U24299 ( .A(n22902), .B(n22903), .Z(n22708) );
  AND U24300 ( .A(n228), .B(n22904), .Z(n22902) );
  XOR U24301 ( .A(n22905), .B(n22903), .Z(n22904) );
  XNOR U24302 ( .A(n22906), .B(n22907), .Z(n22855) );
  NAND U24303 ( .A(n22908), .B(n22909), .Z(n22907) );
  XOR U24304 ( .A(n22910), .B(n22807), .Z(n22909) );
  XOR U24305 ( .A(n22883), .B(n22884), .Z(n22807) );
  XOR U24306 ( .A(n22911), .B(n22876), .Z(n22884) );
  XOR U24307 ( .A(n22912), .B(n22864), .Z(n22876) );
  XOR U24308 ( .A(n22913), .B(n22914), .Z(n22864) );
  ANDN U24309 ( .B(n22915), .A(n22916), .Z(n22913) );
  XOR U24310 ( .A(n22914), .B(n22917), .Z(n22915) );
  IV U24311 ( .A(n22862), .Z(n22912) );
  XOR U24312 ( .A(n22860), .B(n22918), .Z(n22862) );
  XOR U24313 ( .A(n22919), .B(n22920), .Z(n22918) );
  ANDN U24314 ( .B(n22921), .A(n22922), .Z(n22919) );
  XOR U24315 ( .A(n22923), .B(n22920), .Z(n22921) );
  IV U24316 ( .A(n22863), .Z(n22860) );
  XOR U24317 ( .A(n22924), .B(n22925), .Z(n22863) );
  ANDN U24318 ( .B(n22926), .A(n22927), .Z(n22924) );
  XOR U24319 ( .A(n22925), .B(n22928), .Z(n22926) );
  IV U24320 ( .A(n22875), .Z(n22911) );
  XOR U24321 ( .A(n22929), .B(n22930), .Z(n22875) );
  XNOR U24322 ( .A(n22870), .B(n22931), .Z(n22930) );
  IV U24323 ( .A(n22873), .Z(n22931) );
  XOR U24324 ( .A(n22932), .B(n22933), .Z(n22873) );
  ANDN U24325 ( .B(n22934), .A(n22935), .Z(n22932) );
  XOR U24326 ( .A(n22933), .B(n22936), .Z(n22934) );
  XNOR U24327 ( .A(n22937), .B(n22938), .Z(n22870) );
  ANDN U24328 ( .B(n22939), .A(n22940), .Z(n22937) );
  XOR U24329 ( .A(n22938), .B(n22941), .Z(n22939) );
  IV U24330 ( .A(n22869), .Z(n22929) );
  XOR U24331 ( .A(n22867), .B(n22942), .Z(n22869) );
  XOR U24332 ( .A(n22943), .B(n22944), .Z(n22942) );
  ANDN U24333 ( .B(n22945), .A(n22946), .Z(n22943) );
  XOR U24334 ( .A(n22947), .B(n22944), .Z(n22945) );
  IV U24335 ( .A(n22871), .Z(n22867) );
  XOR U24336 ( .A(n22948), .B(n22949), .Z(n22871) );
  ANDN U24337 ( .B(n22950), .A(n22951), .Z(n22948) );
  XOR U24338 ( .A(n22952), .B(n22949), .Z(n22950) );
  XOR U24339 ( .A(n22953), .B(n22954), .Z(n22883) );
  XOR U24340 ( .A(n22901), .B(n22955), .Z(n22954) );
  IV U24341 ( .A(n22881), .Z(n22955) );
  XOR U24342 ( .A(n22956), .B(n22957), .Z(n22881) );
  ANDN U24343 ( .B(n22958), .A(n22959), .Z(n22956) );
  XOR U24344 ( .A(n22957), .B(n22960), .Z(n22958) );
  XOR U24345 ( .A(n22961), .B(n22889), .Z(n22901) );
  XOR U24346 ( .A(n22962), .B(n22963), .Z(n22889) );
  ANDN U24347 ( .B(n22964), .A(n22965), .Z(n22962) );
  XOR U24348 ( .A(n22963), .B(n22966), .Z(n22964) );
  IV U24349 ( .A(n22888), .Z(n22961) );
  XOR U24350 ( .A(n22967), .B(n22968), .Z(n22888) );
  XOR U24351 ( .A(n22969), .B(n22970), .Z(n22968) );
  ANDN U24352 ( .B(n22971), .A(n22972), .Z(n22969) );
  XOR U24353 ( .A(n22973), .B(n22970), .Z(n22971) );
  IV U24354 ( .A(n22886), .Z(n22967) );
  XOR U24355 ( .A(n22974), .B(n22975), .Z(n22886) );
  ANDN U24356 ( .B(n22976), .A(n22977), .Z(n22974) );
  XOR U24357 ( .A(n22975), .B(n22978), .Z(n22976) );
  IV U24358 ( .A(n22900), .Z(n22953) );
  XOR U24359 ( .A(n22979), .B(n22980), .Z(n22900) );
  XNOR U24360 ( .A(n22895), .B(n22981), .Z(n22980) );
  IV U24361 ( .A(n22898), .Z(n22981) );
  XOR U24362 ( .A(n22982), .B(n22983), .Z(n22898) );
  ANDN U24363 ( .B(n22984), .A(n22985), .Z(n22982) );
  XOR U24364 ( .A(n22986), .B(n22983), .Z(n22984) );
  XNOR U24365 ( .A(n22987), .B(n22988), .Z(n22895) );
  ANDN U24366 ( .B(n22989), .A(n22990), .Z(n22987) );
  XOR U24367 ( .A(n22988), .B(n22991), .Z(n22989) );
  IV U24368 ( .A(n22894), .Z(n22979) );
  XOR U24369 ( .A(n22892), .B(n22992), .Z(n22894) );
  XOR U24370 ( .A(n22993), .B(n22994), .Z(n22992) );
  ANDN U24371 ( .B(n22995), .A(n22996), .Z(n22993) );
  XOR U24372 ( .A(n22997), .B(n22994), .Z(n22995) );
  IV U24373 ( .A(n22896), .Z(n22892) );
  XOR U24374 ( .A(n22998), .B(n22999), .Z(n22896) );
  ANDN U24375 ( .B(n23000), .A(n23001), .Z(n22998) );
  XOR U24376 ( .A(n23002), .B(n22999), .Z(n23000) );
  IV U24377 ( .A(n22906), .Z(n22910) );
  XOR U24378 ( .A(n22906), .B(n22809), .Z(n22908) );
  XOR U24379 ( .A(n23003), .B(n23004), .Z(n22809) );
  AND U24380 ( .A(n228), .B(n23005), .Z(n23003) );
  XOR U24381 ( .A(n23006), .B(n23004), .Z(n23005) );
  NANDN U24382 ( .A(n22811), .B(n22813), .Z(n22906) );
  XOR U24383 ( .A(n23007), .B(n23008), .Z(n22813) );
  AND U24384 ( .A(n228), .B(n23009), .Z(n23007) );
  XOR U24385 ( .A(n23008), .B(n23010), .Z(n23009) );
  XNOR U24386 ( .A(n23011), .B(n23012), .Z(n228) );
  AND U24387 ( .A(n23013), .B(n23014), .Z(n23011) );
  XOR U24388 ( .A(n23012), .B(n22824), .Z(n23014) );
  XNOR U24389 ( .A(n23015), .B(n23016), .Z(n22824) );
  ANDN U24390 ( .B(n23017), .A(n23018), .Z(n23015) );
  XOR U24391 ( .A(n23016), .B(n23019), .Z(n23017) );
  XNOR U24392 ( .A(n23012), .B(n22826), .Z(n23013) );
  XOR U24393 ( .A(n23020), .B(n23021), .Z(n22826) );
  AND U24394 ( .A(n232), .B(n23022), .Z(n23020) );
  XOR U24395 ( .A(n23023), .B(n23021), .Z(n23022) );
  XOR U24396 ( .A(n23024), .B(n23025), .Z(n23012) );
  AND U24397 ( .A(n23026), .B(n23027), .Z(n23024) );
  XOR U24398 ( .A(n23025), .B(n22851), .Z(n23027) );
  XOR U24399 ( .A(n23018), .B(n23019), .Z(n22851) );
  XNOR U24400 ( .A(n23028), .B(n23029), .Z(n23019) );
  ANDN U24401 ( .B(n23030), .A(n23031), .Z(n23028) );
  XOR U24402 ( .A(n23032), .B(n23033), .Z(n23030) );
  XOR U24403 ( .A(n23034), .B(n23035), .Z(n23018) );
  XNOR U24404 ( .A(n23036), .B(n23037), .Z(n23035) );
  ANDN U24405 ( .B(n23038), .A(n23039), .Z(n23036) );
  XNOR U24406 ( .A(n23040), .B(n23041), .Z(n23038) );
  IV U24407 ( .A(n23016), .Z(n23034) );
  XOR U24408 ( .A(n23042), .B(n23043), .Z(n23016) );
  ANDN U24409 ( .B(n23044), .A(n23045), .Z(n23042) );
  XOR U24410 ( .A(n23043), .B(n23046), .Z(n23044) );
  XNOR U24411 ( .A(n23025), .B(n22853), .Z(n23026) );
  XOR U24412 ( .A(n23047), .B(n23048), .Z(n22853) );
  AND U24413 ( .A(n232), .B(n23049), .Z(n23047) );
  XOR U24414 ( .A(n23050), .B(n23048), .Z(n23049) );
  XNOR U24415 ( .A(n23051), .B(n23052), .Z(n23025) );
  AND U24416 ( .A(n23053), .B(n23054), .Z(n23051) );
  XNOR U24417 ( .A(n23052), .B(n22903), .Z(n23054) );
  XOR U24418 ( .A(n23045), .B(n23046), .Z(n22903) );
  XOR U24419 ( .A(n23055), .B(n23033), .Z(n23046) );
  XNOR U24420 ( .A(n23056), .B(n23057), .Z(n23033) );
  ANDN U24421 ( .B(n23058), .A(n23059), .Z(n23056) );
  XOR U24422 ( .A(n23060), .B(n23061), .Z(n23058) );
  IV U24423 ( .A(n23031), .Z(n23055) );
  XOR U24424 ( .A(n23029), .B(n23062), .Z(n23031) );
  XNOR U24425 ( .A(n23063), .B(n23064), .Z(n23062) );
  ANDN U24426 ( .B(n23065), .A(n23066), .Z(n23063) );
  XNOR U24427 ( .A(n23067), .B(n23068), .Z(n23065) );
  IV U24428 ( .A(n23032), .Z(n23029) );
  XOR U24429 ( .A(n23069), .B(n23070), .Z(n23032) );
  ANDN U24430 ( .B(n23071), .A(n23072), .Z(n23069) );
  XOR U24431 ( .A(n23070), .B(n23073), .Z(n23071) );
  XOR U24432 ( .A(n23074), .B(n23075), .Z(n23045) );
  XNOR U24433 ( .A(n23040), .B(n23076), .Z(n23075) );
  IV U24434 ( .A(n23043), .Z(n23076) );
  XOR U24435 ( .A(n23077), .B(n23078), .Z(n23043) );
  ANDN U24436 ( .B(n23079), .A(n23080), .Z(n23077) );
  XOR U24437 ( .A(n23078), .B(n23081), .Z(n23079) );
  XNOR U24438 ( .A(n23082), .B(n23083), .Z(n23040) );
  ANDN U24439 ( .B(n23084), .A(n23085), .Z(n23082) );
  XOR U24440 ( .A(n23083), .B(n23086), .Z(n23084) );
  IV U24441 ( .A(n23039), .Z(n23074) );
  XOR U24442 ( .A(n23037), .B(n23087), .Z(n23039) );
  XNOR U24443 ( .A(n23088), .B(n23089), .Z(n23087) );
  ANDN U24444 ( .B(n23090), .A(n23091), .Z(n23088) );
  XNOR U24445 ( .A(n23092), .B(n23093), .Z(n23090) );
  IV U24446 ( .A(n23041), .Z(n23037) );
  XOR U24447 ( .A(n23094), .B(n23095), .Z(n23041) );
  ANDN U24448 ( .B(n23096), .A(n23097), .Z(n23094) );
  XOR U24449 ( .A(n23098), .B(n23095), .Z(n23096) );
  XOR U24450 ( .A(n23052), .B(n22905), .Z(n23053) );
  XOR U24451 ( .A(n23099), .B(n23100), .Z(n22905) );
  AND U24452 ( .A(n232), .B(n23101), .Z(n23099) );
  XOR U24453 ( .A(n23102), .B(n23100), .Z(n23101) );
  XNOR U24454 ( .A(n23103), .B(n23104), .Z(n23052) );
  NAND U24455 ( .A(n23105), .B(n23106), .Z(n23104) );
  XOR U24456 ( .A(n23107), .B(n23004), .Z(n23106) );
  XOR U24457 ( .A(n23080), .B(n23081), .Z(n23004) );
  XOR U24458 ( .A(n23108), .B(n23073), .Z(n23081) );
  XOR U24459 ( .A(n23109), .B(n23061), .Z(n23073) );
  XOR U24460 ( .A(n23110), .B(n23111), .Z(n23061) );
  ANDN U24461 ( .B(n23112), .A(n23113), .Z(n23110) );
  XOR U24462 ( .A(n23111), .B(n23114), .Z(n23112) );
  IV U24463 ( .A(n23059), .Z(n23109) );
  XOR U24464 ( .A(n23057), .B(n23115), .Z(n23059) );
  XOR U24465 ( .A(n23116), .B(n23117), .Z(n23115) );
  ANDN U24466 ( .B(n23118), .A(n23119), .Z(n23116) );
  XOR U24467 ( .A(n23120), .B(n23117), .Z(n23118) );
  IV U24468 ( .A(n23060), .Z(n23057) );
  XOR U24469 ( .A(n23121), .B(n23122), .Z(n23060) );
  ANDN U24470 ( .B(n23123), .A(n23124), .Z(n23121) );
  XOR U24471 ( .A(n23122), .B(n23125), .Z(n23123) );
  IV U24472 ( .A(n23072), .Z(n23108) );
  XOR U24473 ( .A(n23126), .B(n23127), .Z(n23072) );
  XNOR U24474 ( .A(n23067), .B(n23128), .Z(n23127) );
  IV U24475 ( .A(n23070), .Z(n23128) );
  XOR U24476 ( .A(n23129), .B(n23130), .Z(n23070) );
  ANDN U24477 ( .B(n23131), .A(n23132), .Z(n23129) );
  XOR U24478 ( .A(n23130), .B(n23133), .Z(n23131) );
  XNOR U24479 ( .A(n23134), .B(n23135), .Z(n23067) );
  ANDN U24480 ( .B(n23136), .A(n23137), .Z(n23134) );
  XOR U24481 ( .A(n23135), .B(n23138), .Z(n23136) );
  IV U24482 ( .A(n23066), .Z(n23126) );
  XOR U24483 ( .A(n23064), .B(n23139), .Z(n23066) );
  XOR U24484 ( .A(n23140), .B(n23141), .Z(n23139) );
  ANDN U24485 ( .B(n23142), .A(n23143), .Z(n23140) );
  XOR U24486 ( .A(n23144), .B(n23141), .Z(n23142) );
  IV U24487 ( .A(n23068), .Z(n23064) );
  XOR U24488 ( .A(n23145), .B(n23146), .Z(n23068) );
  ANDN U24489 ( .B(n23147), .A(n23148), .Z(n23145) );
  XOR U24490 ( .A(n23149), .B(n23146), .Z(n23147) );
  XOR U24491 ( .A(n23150), .B(n23151), .Z(n23080) );
  XOR U24492 ( .A(n23098), .B(n23152), .Z(n23151) );
  IV U24493 ( .A(n23078), .Z(n23152) );
  XOR U24494 ( .A(n23153), .B(n23154), .Z(n23078) );
  ANDN U24495 ( .B(n23155), .A(n23156), .Z(n23153) );
  XOR U24496 ( .A(n23154), .B(n23157), .Z(n23155) );
  XOR U24497 ( .A(n23158), .B(n23086), .Z(n23098) );
  XOR U24498 ( .A(n23159), .B(n23160), .Z(n23086) );
  ANDN U24499 ( .B(n23161), .A(n23162), .Z(n23159) );
  XOR U24500 ( .A(n23160), .B(n23163), .Z(n23161) );
  IV U24501 ( .A(n23085), .Z(n23158) );
  XOR U24502 ( .A(n23164), .B(n23165), .Z(n23085) );
  XOR U24503 ( .A(n23166), .B(n23167), .Z(n23165) );
  ANDN U24504 ( .B(n23168), .A(n23169), .Z(n23166) );
  XOR U24505 ( .A(n23170), .B(n23167), .Z(n23168) );
  IV U24506 ( .A(n23083), .Z(n23164) );
  XOR U24507 ( .A(n23171), .B(n23172), .Z(n23083) );
  ANDN U24508 ( .B(n23173), .A(n23174), .Z(n23171) );
  XOR U24509 ( .A(n23172), .B(n23175), .Z(n23173) );
  IV U24510 ( .A(n23097), .Z(n23150) );
  XOR U24511 ( .A(n23176), .B(n23177), .Z(n23097) );
  XNOR U24512 ( .A(n23092), .B(n23178), .Z(n23177) );
  IV U24513 ( .A(n23095), .Z(n23178) );
  XOR U24514 ( .A(n23179), .B(n23180), .Z(n23095) );
  ANDN U24515 ( .B(n23181), .A(n23182), .Z(n23179) );
  XOR U24516 ( .A(n23183), .B(n23180), .Z(n23181) );
  XNOR U24517 ( .A(n23184), .B(n23185), .Z(n23092) );
  ANDN U24518 ( .B(n23186), .A(n23187), .Z(n23184) );
  XOR U24519 ( .A(n23185), .B(n23188), .Z(n23186) );
  IV U24520 ( .A(n23091), .Z(n23176) );
  XOR U24521 ( .A(n23089), .B(n23189), .Z(n23091) );
  XOR U24522 ( .A(n23190), .B(n23191), .Z(n23189) );
  ANDN U24523 ( .B(n23192), .A(n23193), .Z(n23190) );
  XOR U24524 ( .A(n23194), .B(n23191), .Z(n23192) );
  IV U24525 ( .A(n23093), .Z(n23089) );
  XOR U24526 ( .A(n23195), .B(n23196), .Z(n23093) );
  ANDN U24527 ( .B(n23197), .A(n23198), .Z(n23195) );
  XOR U24528 ( .A(n23199), .B(n23196), .Z(n23197) );
  IV U24529 ( .A(n23103), .Z(n23107) );
  XOR U24530 ( .A(n23103), .B(n23006), .Z(n23105) );
  XOR U24531 ( .A(n23200), .B(n23201), .Z(n23006) );
  AND U24532 ( .A(n232), .B(n23202), .Z(n23200) );
  XOR U24533 ( .A(n23203), .B(n23201), .Z(n23202) );
  NANDN U24534 ( .A(n23008), .B(n23010), .Z(n23103) );
  XOR U24535 ( .A(n23204), .B(n23205), .Z(n23010) );
  AND U24536 ( .A(n232), .B(n23206), .Z(n23204) );
  XOR U24537 ( .A(n23205), .B(n23207), .Z(n23206) );
  XNOR U24538 ( .A(n23208), .B(n23209), .Z(n232) );
  AND U24539 ( .A(n23210), .B(n23211), .Z(n23208) );
  XOR U24540 ( .A(n23209), .B(n23021), .Z(n23211) );
  XNOR U24541 ( .A(n23212), .B(n23213), .Z(n23021) );
  ANDN U24542 ( .B(n23214), .A(n23215), .Z(n23212) );
  XOR U24543 ( .A(n23213), .B(n23216), .Z(n23214) );
  XNOR U24544 ( .A(n23209), .B(n23023), .Z(n23210) );
  XOR U24545 ( .A(n23217), .B(n23218), .Z(n23023) );
  AND U24546 ( .A(n236), .B(n23219), .Z(n23217) );
  XOR U24547 ( .A(n23220), .B(n23218), .Z(n23219) );
  XOR U24548 ( .A(n23221), .B(n23222), .Z(n23209) );
  AND U24549 ( .A(n23223), .B(n23224), .Z(n23221) );
  XOR U24550 ( .A(n23222), .B(n23048), .Z(n23224) );
  XOR U24551 ( .A(n23215), .B(n23216), .Z(n23048) );
  XNOR U24552 ( .A(n23225), .B(n23226), .Z(n23216) );
  ANDN U24553 ( .B(n23227), .A(n23228), .Z(n23225) );
  XOR U24554 ( .A(n23229), .B(n23230), .Z(n23227) );
  XOR U24555 ( .A(n23231), .B(n23232), .Z(n23215) );
  XNOR U24556 ( .A(n23233), .B(n23234), .Z(n23232) );
  ANDN U24557 ( .B(n23235), .A(n23236), .Z(n23233) );
  XNOR U24558 ( .A(n23237), .B(n23238), .Z(n23235) );
  IV U24559 ( .A(n23213), .Z(n23231) );
  XOR U24560 ( .A(n23239), .B(n23240), .Z(n23213) );
  ANDN U24561 ( .B(n23241), .A(n23242), .Z(n23239) );
  XOR U24562 ( .A(n23240), .B(n23243), .Z(n23241) );
  XNOR U24563 ( .A(n23222), .B(n23050), .Z(n23223) );
  XOR U24564 ( .A(n23244), .B(n23245), .Z(n23050) );
  AND U24565 ( .A(n236), .B(n23246), .Z(n23244) );
  XOR U24566 ( .A(n23247), .B(n23245), .Z(n23246) );
  XNOR U24567 ( .A(n23248), .B(n23249), .Z(n23222) );
  AND U24568 ( .A(n23250), .B(n23251), .Z(n23248) );
  XNOR U24569 ( .A(n23249), .B(n23100), .Z(n23251) );
  XOR U24570 ( .A(n23242), .B(n23243), .Z(n23100) );
  XOR U24571 ( .A(n23252), .B(n23230), .Z(n23243) );
  XNOR U24572 ( .A(n23253), .B(n23254), .Z(n23230) );
  ANDN U24573 ( .B(n23255), .A(n23256), .Z(n23253) );
  XOR U24574 ( .A(n23257), .B(n23258), .Z(n23255) );
  IV U24575 ( .A(n23228), .Z(n23252) );
  XOR U24576 ( .A(n23226), .B(n23259), .Z(n23228) );
  XNOR U24577 ( .A(n23260), .B(n23261), .Z(n23259) );
  ANDN U24578 ( .B(n23262), .A(n23263), .Z(n23260) );
  XNOR U24579 ( .A(n23264), .B(n23265), .Z(n23262) );
  IV U24580 ( .A(n23229), .Z(n23226) );
  XOR U24581 ( .A(n23266), .B(n23267), .Z(n23229) );
  ANDN U24582 ( .B(n23268), .A(n23269), .Z(n23266) );
  XOR U24583 ( .A(n23267), .B(n23270), .Z(n23268) );
  XOR U24584 ( .A(n23271), .B(n23272), .Z(n23242) );
  XNOR U24585 ( .A(n23237), .B(n23273), .Z(n23272) );
  IV U24586 ( .A(n23240), .Z(n23273) );
  XOR U24587 ( .A(n23274), .B(n23275), .Z(n23240) );
  ANDN U24588 ( .B(n23276), .A(n23277), .Z(n23274) );
  XOR U24589 ( .A(n23275), .B(n23278), .Z(n23276) );
  XNOR U24590 ( .A(n23279), .B(n23280), .Z(n23237) );
  ANDN U24591 ( .B(n23281), .A(n23282), .Z(n23279) );
  XOR U24592 ( .A(n23280), .B(n23283), .Z(n23281) );
  IV U24593 ( .A(n23236), .Z(n23271) );
  XOR U24594 ( .A(n23234), .B(n23284), .Z(n23236) );
  XNOR U24595 ( .A(n23285), .B(n23286), .Z(n23284) );
  ANDN U24596 ( .B(n23287), .A(n23288), .Z(n23285) );
  XNOR U24597 ( .A(n23289), .B(n23290), .Z(n23287) );
  IV U24598 ( .A(n23238), .Z(n23234) );
  XOR U24599 ( .A(n23291), .B(n23292), .Z(n23238) );
  ANDN U24600 ( .B(n23293), .A(n23294), .Z(n23291) );
  XOR U24601 ( .A(n23295), .B(n23292), .Z(n23293) );
  XOR U24602 ( .A(n23249), .B(n23102), .Z(n23250) );
  XOR U24603 ( .A(n23296), .B(n23297), .Z(n23102) );
  AND U24604 ( .A(n236), .B(n23298), .Z(n23296) );
  XOR U24605 ( .A(n23299), .B(n23297), .Z(n23298) );
  XNOR U24606 ( .A(n23300), .B(n23301), .Z(n23249) );
  NAND U24607 ( .A(n23302), .B(n23303), .Z(n23301) );
  XOR U24608 ( .A(n23304), .B(n23201), .Z(n23303) );
  XOR U24609 ( .A(n23277), .B(n23278), .Z(n23201) );
  XOR U24610 ( .A(n23305), .B(n23270), .Z(n23278) );
  XOR U24611 ( .A(n23306), .B(n23258), .Z(n23270) );
  XOR U24612 ( .A(n23307), .B(n23308), .Z(n23258) );
  ANDN U24613 ( .B(n23309), .A(n23310), .Z(n23307) );
  XOR U24614 ( .A(n23308), .B(n23311), .Z(n23309) );
  IV U24615 ( .A(n23256), .Z(n23306) );
  XOR U24616 ( .A(n23254), .B(n23312), .Z(n23256) );
  XOR U24617 ( .A(n23313), .B(n23314), .Z(n23312) );
  ANDN U24618 ( .B(n23315), .A(n23316), .Z(n23313) );
  XOR U24619 ( .A(n23317), .B(n23314), .Z(n23315) );
  IV U24620 ( .A(n23257), .Z(n23254) );
  XOR U24621 ( .A(n23318), .B(n23319), .Z(n23257) );
  ANDN U24622 ( .B(n23320), .A(n23321), .Z(n23318) );
  XOR U24623 ( .A(n23319), .B(n23322), .Z(n23320) );
  IV U24624 ( .A(n23269), .Z(n23305) );
  XOR U24625 ( .A(n23323), .B(n23324), .Z(n23269) );
  XNOR U24626 ( .A(n23264), .B(n23325), .Z(n23324) );
  IV U24627 ( .A(n23267), .Z(n23325) );
  XOR U24628 ( .A(n23326), .B(n23327), .Z(n23267) );
  ANDN U24629 ( .B(n23328), .A(n23329), .Z(n23326) );
  XOR U24630 ( .A(n23327), .B(n23330), .Z(n23328) );
  XNOR U24631 ( .A(n23331), .B(n23332), .Z(n23264) );
  ANDN U24632 ( .B(n23333), .A(n23334), .Z(n23331) );
  XOR U24633 ( .A(n23332), .B(n23335), .Z(n23333) );
  IV U24634 ( .A(n23263), .Z(n23323) );
  XOR U24635 ( .A(n23261), .B(n23336), .Z(n23263) );
  XOR U24636 ( .A(n23337), .B(n23338), .Z(n23336) );
  ANDN U24637 ( .B(n23339), .A(n23340), .Z(n23337) );
  XOR U24638 ( .A(n23341), .B(n23338), .Z(n23339) );
  IV U24639 ( .A(n23265), .Z(n23261) );
  XOR U24640 ( .A(n23342), .B(n23343), .Z(n23265) );
  ANDN U24641 ( .B(n23344), .A(n23345), .Z(n23342) );
  XOR U24642 ( .A(n23346), .B(n23343), .Z(n23344) );
  XOR U24643 ( .A(n23347), .B(n23348), .Z(n23277) );
  XOR U24644 ( .A(n23295), .B(n23349), .Z(n23348) );
  IV U24645 ( .A(n23275), .Z(n23349) );
  XOR U24646 ( .A(n23350), .B(n23351), .Z(n23275) );
  ANDN U24647 ( .B(n23352), .A(n23353), .Z(n23350) );
  XOR U24648 ( .A(n23351), .B(n23354), .Z(n23352) );
  XOR U24649 ( .A(n23355), .B(n23283), .Z(n23295) );
  XOR U24650 ( .A(n23356), .B(n23357), .Z(n23283) );
  ANDN U24651 ( .B(n23358), .A(n23359), .Z(n23356) );
  XOR U24652 ( .A(n23357), .B(n23360), .Z(n23358) );
  IV U24653 ( .A(n23282), .Z(n23355) );
  XOR U24654 ( .A(n23361), .B(n23362), .Z(n23282) );
  XOR U24655 ( .A(n23363), .B(n23364), .Z(n23362) );
  ANDN U24656 ( .B(n23365), .A(n23366), .Z(n23363) );
  XOR U24657 ( .A(n23367), .B(n23364), .Z(n23365) );
  IV U24658 ( .A(n23280), .Z(n23361) );
  XOR U24659 ( .A(n23368), .B(n23369), .Z(n23280) );
  ANDN U24660 ( .B(n23370), .A(n23371), .Z(n23368) );
  XOR U24661 ( .A(n23369), .B(n23372), .Z(n23370) );
  IV U24662 ( .A(n23294), .Z(n23347) );
  XOR U24663 ( .A(n23373), .B(n23374), .Z(n23294) );
  XNOR U24664 ( .A(n23289), .B(n23375), .Z(n23374) );
  IV U24665 ( .A(n23292), .Z(n23375) );
  XOR U24666 ( .A(n23376), .B(n23377), .Z(n23292) );
  ANDN U24667 ( .B(n23378), .A(n23379), .Z(n23376) );
  XOR U24668 ( .A(n23380), .B(n23377), .Z(n23378) );
  XNOR U24669 ( .A(n23381), .B(n23382), .Z(n23289) );
  ANDN U24670 ( .B(n23383), .A(n23384), .Z(n23381) );
  XOR U24671 ( .A(n23382), .B(n23385), .Z(n23383) );
  IV U24672 ( .A(n23288), .Z(n23373) );
  XOR U24673 ( .A(n23286), .B(n23386), .Z(n23288) );
  XOR U24674 ( .A(n23387), .B(n23388), .Z(n23386) );
  ANDN U24675 ( .B(n23389), .A(n23390), .Z(n23387) );
  XOR U24676 ( .A(n23391), .B(n23388), .Z(n23389) );
  IV U24677 ( .A(n23290), .Z(n23286) );
  XOR U24678 ( .A(n23392), .B(n23393), .Z(n23290) );
  ANDN U24679 ( .B(n23394), .A(n23395), .Z(n23392) );
  XOR U24680 ( .A(n23396), .B(n23393), .Z(n23394) );
  IV U24681 ( .A(n23300), .Z(n23304) );
  XOR U24682 ( .A(n23300), .B(n23203), .Z(n23302) );
  XOR U24683 ( .A(n23397), .B(n23398), .Z(n23203) );
  AND U24684 ( .A(n236), .B(n23399), .Z(n23397) );
  XOR U24685 ( .A(n23400), .B(n23398), .Z(n23399) );
  NANDN U24686 ( .A(n23205), .B(n23207), .Z(n23300) );
  XOR U24687 ( .A(n23401), .B(n23402), .Z(n23207) );
  AND U24688 ( .A(n236), .B(n23403), .Z(n23401) );
  XOR U24689 ( .A(n23402), .B(n23404), .Z(n23403) );
  XNOR U24690 ( .A(n23405), .B(n23406), .Z(n236) );
  AND U24691 ( .A(n23407), .B(n23408), .Z(n23405) );
  XOR U24692 ( .A(n23406), .B(n23218), .Z(n23408) );
  XNOR U24693 ( .A(n23409), .B(n23410), .Z(n23218) );
  ANDN U24694 ( .B(n23411), .A(n23412), .Z(n23409) );
  XOR U24695 ( .A(n23410), .B(n23413), .Z(n23411) );
  XNOR U24696 ( .A(n23406), .B(n23220), .Z(n23407) );
  XOR U24697 ( .A(n23414), .B(n23415), .Z(n23220) );
  AND U24698 ( .A(n240), .B(n23416), .Z(n23414) );
  XOR U24699 ( .A(n23417), .B(n23415), .Z(n23416) );
  XOR U24700 ( .A(n23418), .B(n23419), .Z(n23406) );
  AND U24701 ( .A(n23420), .B(n23421), .Z(n23418) );
  XOR U24702 ( .A(n23419), .B(n23245), .Z(n23421) );
  XOR U24703 ( .A(n23412), .B(n23413), .Z(n23245) );
  XNOR U24704 ( .A(n23422), .B(n23423), .Z(n23413) );
  ANDN U24705 ( .B(n23424), .A(n23425), .Z(n23422) );
  XOR U24706 ( .A(n23426), .B(n23427), .Z(n23424) );
  XOR U24707 ( .A(n23428), .B(n23429), .Z(n23412) );
  XNOR U24708 ( .A(n23430), .B(n23431), .Z(n23429) );
  ANDN U24709 ( .B(n23432), .A(n23433), .Z(n23430) );
  XNOR U24710 ( .A(n23434), .B(n23435), .Z(n23432) );
  IV U24711 ( .A(n23410), .Z(n23428) );
  XOR U24712 ( .A(n23436), .B(n23437), .Z(n23410) );
  ANDN U24713 ( .B(n23438), .A(n23439), .Z(n23436) );
  XOR U24714 ( .A(n23437), .B(n23440), .Z(n23438) );
  XNOR U24715 ( .A(n23419), .B(n23247), .Z(n23420) );
  XOR U24716 ( .A(n23441), .B(n23442), .Z(n23247) );
  AND U24717 ( .A(n240), .B(n23443), .Z(n23441) );
  XOR U24718 ( .A(n23444), .B(n23442), .Z(n23443) );
  XNOR U24719 ( .A(n23445), .B(n23446), .Z(n23419) );
  AND U24720 ( .A(n23447), .B(n23448), .Z(n23445) );
  XNOR U24721 ( .A(n23446), .B(n23297), .Z(n23448) );
  XOR U24722 ( .A(n23439), .B(n23440), .Z(n23297) );
  XOR U24723 ( .A(n23449), .B(n23427), .Z(n23440) );
  XNOR U24724 ( .A(n23450), .B(n23451), .Z(n23427) );
  ANDN U24725 ( .B(n23452), .A(n23453), .Z(n23450) );
  XOR U24726 ( .A(n23454), .B(n23455), .Z(n23452) );
  IV U24727 ( .A(n23425), .Z(n23449) );
  XOR U24728 ( .A(n23423), .B(n23456), .Z(n23425) );
  XNOR U24729 ( .A(n23457), .B(n23458), .Z(n23456) );
  ANDN U24730 ( .B(n23459), .A(n23460), .Z(n23457) );
  XNOR U24731 ( .A(n23461), .B(n23462), .Z(n23459) );
  IV U24732 ( .A(n23426), .Z(n23423) );
  XOR U24733 ( .A(n23463), .B(n23464), .Z(n23426) );
  ANDN U24734 ( .B(n23465), .A(n23466), .Z(n23463) );
  XOR U24735 ( .A(n23464), .B(n23467), .Z(n23465) );
  XOR U24736 ( .A(n23468), .B(n23469), .Z(n23439) );
  XNOR U24737 ( .A(n23434), .B(n23470), .Z(n23469) );
  IV U24738 ( .A(n23437), .Z(n23470) );
  XOR U24739 ( .A(n23471), .B(n23472), .Z(n23437) );
  ANDN U24740 ( .B(n23473), .A(n23474), .Z(n23471) );
  XOR U24741 ( .A(n23472), .B(n23475), .Z(n23473) );
  XNOR U24742 ( .A(n23476), .B(n23477), .Z(n23434) );
  ANDN U24743 ( .B(n23478), .A(n23479), .Z(n23476) );
  XOR U24744 ( .A(n23477), .B(n23480), .Z(n23478) );
  IV U24745 ( .A(n23433), .Z(n23468) );
  XOR U24746 ( .A(n23431), .B(n23481), .Z(n23433) );
  XNOR U24747 ( .A(n23482), .B(n23483), .Z(n23481) );
  ANDN U24748 ( .B(n23484), .A(n23485), .Z(n23482) );
  XNOR U24749 ( .A(n23486), .B(n23487), .Z(n23484) );
  IV U24750 ( .A(n23435), .Z(n23431) );
  XOR U24751 ( .A(n23488), .B(n23489), .Z(n23435) );
  ANDN U24752 ( .B(n23490), .A(n23491), .Z(n23488) );
  XOR U24753 ( .A(n23492), .B(n23489), .Z(n23490) );
  XOR U24754 ( .A(n23446), .B(n23299), .Z(n23447) );
  XOR U24755 ( .A(n23493), .B(n23494), .Z(n23299) );
  AND U24756 ( .A(n240), .B(n23495), .Z(n23493) );
  XOR U24757 ( .A(n23496), .B(n23494), .Z(n23495) );
  XNOR U24758 ( .A(n23497), .B(n23498), .Z(n23446) );
  NAND U24759 ( .A(n23499), .B(n23500), .Z(n23498) );
  XOR U24760 ( .A(n23501), .B(n23398), .Z(n23500) );
  XOR U24761 ( .A(n23474), .B(n23475), .Z(n23398) );
  XOR U24762 ( .A(n23502), .B(n23467), .Z(n23475) );
  XOR U24763 ( .A(n23503), .B(n23455), .Z(n23467) );
  XOR U24764 ( .A(n23504), .B(n23505), .Z(n23455) );
  ANDN U24765 ( .B(n23506), .A(n23507), .Z(n23504) );
  XOR U24766 ( .A(n23505), .B(n23508), .Z(n23506) );
  IV U24767 ( .A(n23453), .Z(n23503) );
  XOR U24768 ( .A(n23451), .B(n23509), .Z(n23453) );
  XOR U24769 ( .A(n23510), .B(n23511), .Z(n23509) );
  ANDN U24770 ( .B(n23512), .A(n23513), .Z(n23510) );
  XOR U24771 ( .A(n23514), .B(n23511), .Z(n23512) );
  IV U24772 ( .A(n23454), .Z(n23451) );
  XOR U24773 ( .A(n23515), .B(n23516), .Z(n23454) );
  ANDN U24774 ( .B(n23517), .A(n23518), .Z(n23515) );
  XOR U24775 ( .A(n23516), .B(n23519), .Z(n23517) );
  IV U24776 ( .A(n23466), .Z(n23502) );
  XOR U24777 ( .A(n23520), .B(n23521), .Z(n23466) );
  XNOR U24778 ( .A(n23461), .B(n23522), .Z(n23521) );
  IV U24779 ( .A(n23464), .Z(n23522) );
  XOR U24780 ( .A(n23523), .B(n23524), .Z(n23464) );
  ANDN U24781 ( .B(n23525), .A(n23526), .Z(n23523) );
  XOR U24782 ( .A(n23524), .B(n23527), .Z(n23525) );
  XNOR U24783 ( .A(n23528), .B(n23529), .Z(n23461) );
  ANDN U24784 ( .B(n23530), .A(n23531), .Z(n23528) );
  XOR U24785 ( .A(n23529), .B(n23532), .Z(n23530) );
  IV U24786 ( .A(n23460), .Z(n23520) );
  XOR U24787 ( .A(n23458), .B(n23533), .Z(n23460) );
  XOR U24788 ( .A(n23534), .B(n23535), .Z(n23533) );
  ANDN U24789 ( .B(n23536), .A(n23537), .Z(n23534) );
  XOR U24790 ( .A(n23538), .B(n23535), .Z(n23536) );
  IV U24791 ( .A(n23462), .Z(n23458) );
  XOR U24792 ( .A(n23539), .B(n23540), .Z(n23462) );
  ANDN U24793 ( .B(n23541), .A(n23542), .Z(n23539) );
  XOR U24794 ( .A(n23543), .B(n23540), .Z(n23541) );
  XOR U24795 ( .A(n23544), .B(n23545), .Z(n23474) );
  XOR U24796 ( .A(n23492), .B(n23546), .Z(n23545) );
  IV U24797 ( .A(n23472), .Z(n23546) );
  XOR U24798 ( .A(n23547), .B(n23548), .Z(n23472) );
  ANDN U24799 ( .B(n23549), .A(n23550), .Z(n23547) );
  XOR U24800 ( .A(n23548), .B(n23551), .Z(n23549) );
  XOR U24801 ( .A(n23552), .B(n23480), .Z(n23492) );
  XOR U24802 ( .A(n23553), .B(n23554), .Z(n23480) );
  ANDN U24803 ( .B(n23555), .A(n23556), .Z(n23553) );
  XOR U24804 ( .A(n23554), .B(n23557), .Z(n23555) );
  IV U24805 ( .A(n23479), .Z(n23552) );
  XOR U24806 ( .A(n23558), .B(n23559), .Z(n23479) );
  XOR U24807 ( .A(n23560), .B(n23561), .Z(n23559) );
  ANDN U24808 ( .B(n23562), .A(n23563), .Z(n23560) );
  XOR U24809 ( .A(n23564), .B(n23561), .Z(n23562) );
  IV U24810 ( .A(n23477), .Z(n23558) );
  XOR U24811 ( .A(n23565), .B(n23566), .Z(n23477) );
  ANDN U24812 ( .B(n23567), .A(n23568), .Z(n23565) );
  XOR U24813 ( .A(n23566), .B(n23569), .Z(n23567) );
  IV U24814 ( .A(n23491), .Z(n23544) );
  XOR U24815 ( .A(n23570), .B(n23571), .Z(n23491) );
  XNOR U24816 ( .A(n23486), .B(n23572), .Z(n23571) );
  IV U24817 ( .A(n23489), .Z(n23572) );
  XOR U24818 ( .A(n23573), .B(n23574), .Z(n23489) );
  ANDN U24819 ( .B(n23575), .A(n23576), .Z(n23573) );
  XOR U24820 ( .A(n23577), .B(n23574), .Z(n23575) );
  XNOR U24821 ( .A(n23578), .B(n23579), .Z(n23486) );
  ANDN U24822 ( .B(n23580), .A(n23581), .Z(n23578) );
  XOR U24823 ( .A(n23579), .B(n23582), .Z(n23580) );
  IV U24824 ( .A(n23485), .Z(n23570) );
  XOR U24825 ( .A(n23483), .B(n23583), .Z(n23485) );
  XOR U24826 ( .A(n23584), .B(n23585), .Z(n23583) );
  ANDN U24827 ( .B(n23586), .A(n23587), .Z(n23584) );
  XOR U24828 ( .A(n23588), .B(n23585), .Z(n23586) );
  IV U24829 ( .A(n23487), .Z(n23483) );
  XOR U24830 ( .A(n23589), .B(n23590), .Z(n23487) );
  ANDN U24831 ( .B(n23591), .A(n23592), .Z(n23589) );
  XOR U24832 ( .A(n23593), .B(n23590), .Z(n23591) );
  IV U24833 ( .A(n23497), .Z(n23501) );
  XOR U24834 ( .A(n23497), .B(n23400), .Z(n23499) );
  XOR U24835 ( .A(n23594), .B(n23595), .Z(n23400) );
  AND U24836 ( .A(n240), .B(n23596), .Z(n23594) );
  XOR U24837 ( .A(n23597), .B(n23595), .Z(n23596) );
  NANDN U24838 ( .A(n23402), .B(n23404), .Z(n23497) );
  XOR U24839 ( .A(n23598), .B(n23599), .Z(n23404) );
  AND U24840 ( .A(n240), .B(n23600), .Z(n23598) );
  XOR U24841 ( .A(n23599), .B(n23601), .Z(n23600) );
  XNOR U24842 ( .A(n23602), .B(n23603), .Z(n240) );
  AND U24843 ( .A(n23604), .B(n23605), .Z(n23602) );
  XOR U24844 ( .A(n23603), .B(n23415), .Z(n23605) );
  XNOR U24845 ( .A(n23606), .B(n23607), .Z(n23415) );
  ANDN U24846 ( .B(n23608), .A(n23609), .Z(n23606) );
  XOR U24847 ( .A(n23607), .B(n23610), .Z(n23608) );
  XNOR U24848 ( .A(n23603), .B(n23417), .Z(n23604) );
  XOR U24849 ( .A(n23611), .B(n23612), .Z(n23417) );
  AND U24850 ( .A(n244), .B(n23613), .Z(n23611) );
  XOR U24851 ( .A(n23614), .B(n23612), .Z(n23613) );
  XOR U24852 ( .A(n23615), .B(n23616), .Z(n23603) );
  AND U24853 ( .A(n23617), .B(n23618), .Z(n23615) );
  XOR U24854 ( .A(n23616), .B(n23442), .Z(n23618) );
  XOR U24855 ( .A(n23609), .B(n23610), .Z(n23442) );
  XNOR U24856 ( .A(n23619), .B(n23620), .Z(n23610) );
  ANDN U24857 ( .B(n23621), .A(n23622), .Z(n23619) );
  XOR U24858 ( .A(n23623), .B(n23624), .Z(n23621) );
  XOR U24859 ( .A(n23625), .B(n23626), .Z(n23609) );
  XNOR U24860 ( .A(n23627), .B(n23628), .Z(n23626) );
  ANDN U24861 ( .B(n23629), .A(n23630), .Z(n23627) );
  XNOR U24862 ( .A(n23631), .B(n23632), .Z(n23629) );
  IV U24863 ( .A(n23607), .Z(n23625) );
  XOR U24864 ( .A(n23633), .B(n23634), .Z(n23607) );
  ANDN U24865 ( .B(n23635), .A(n23636), .Z(n23633) );
  XOR U24866 ( .A(n23634), .B(n23637), .Z(n23635) );
  XNOR U24867 ( .A(n23616), .B(n23444), .Z(n23617) );
  XOR U24868 ( .A(n23638), .B(n23639), .Z(n23444) );
  AND U24869 ( .A(n244), .B(n23640), .Z(n23638) );
  XOR U24870 ( .A(n23641), .B(n23639), .Z(n23640) );
  XNOR U24871 ( .A(n23642), .B(n23643), .Z(n23616) );
  AND U24872 ( .A(n23644), .B(n23645), .Z(n23642) );
  XNOR U24873 ( .A(n23643), .B(n23494), .Z(n23645) );
  XOR U24874 ( .A(n23636), .B(n23637), .Z(n23494) );
  XOR U24875 ( .A(n23646), .B(n23624), .Z(n23637) );
  XNOR U24876 ( .A(n23647), .B(n23648), .Z(n23624) );
  ANDN U24877 ( .B(n23649), .A(n23650), .Z(n23647) );
  XOR U24878 ( .A(n23651), .B(n23652), .Z(n23649) );
  IV U24879 ( .A(n23622), .Z(n23646) );
  XOR U24880 ( .A(n23620), .B(n23653), .Z(n23622) );
  XNOR U24881 ( .A(n23654), .B(n23655), .Z(n23653) );
  ANDN U24882 ( .B(n23656), .A(n23657), .Z(n23654) );
  XNOR U24883 ( .A(n23658), .B(n23659), .Z(n23656) );
  IV U24884 ( .A(n23623), .Z(n23620) );
  XOR U24885 ( .A(n23660), .B(n23661), .Z(n23623) );
  ANDN U24886 ( .B(n23662), .A(n23663), .Z(n23660) );
  XOR U24887 ( .A(n23661), .B(n23664), .Z(n23662) );
  XOR U24888 ( .A(n23665), .B(n23666), .Z(n23636) );
  XNOR U24889 ( .A(n23631), .B(n23667), .Z(n23666) );
  IV U24890 ( .A(n23634), .Z(n23667) );
  XOR U24891 ( .A(n23668), .B(n23669), .Z(n23634) );
  ANDN U24892 ( .B(n23670), .A(n23671), .Z(n23668) );
  XOR U24893 ( .A(n23669), .B(n23672), .Z(n23670) );
  XNOR U24894 ( .A(n23673), .B(n23674), .Z(n23631) );
  ANDN U24895 ( .B(n23675), .A(n23676), .Z(n23673) );
  XOR U24896 ( .A(n23674), .B(n23677), .Z(n23675) );
  IV U24897 ( .A(n23630), .Z(n23665) );
  XOR U24898 ( .A(n23628), .B(n23678), .Z(n23630) );
  XNOR U24899 ( .A(n23679), .B(n23680), .Z(n23678) );
  ANDN U24900 ( .B(n23681), .A(n23682), .Z(n23679) );
  XNOR U24901 ( .A(n23683), .B(n23684), .Z(n23681) );
  IV U24902 ( .A(n23632), .Z(n23628) );
  XOR U24903 ( .A(n23685), .B(n23686), .Z(n23632) );
  ANDN U24904 ( .B(n23687), .A(n23688), .Z(n23685) );
  XOR U24905 ( .A(n23689), .B(n23686), .Z(n23687) );
  XOR U24906 ( .A(n23643), .B(n23496), .Z(n23644) );
  XOR U24907 ( .A(n23690), .B(n23691), .Z(n23496) );
  AND U24908 ( .A(n244), .B(n23692), .Z(n23690) );
  XOR U24909 ( .A(n23693), .B(n23691), .Z(n23692) );
  XNOR U24910 ( .A(n23694), .B(n23695), .Z(n23643) );
  NAND U24911 ( .A(n23696), .B(n23697), .Z(n23695) );
  XOR U24912 ( .A(n23698), .B(n23595), .Z(n23697) );
  XOR U24913 ( .A(n23671), .B(n23672), .Z(n23595) );
  XOR U24914 ( .A(n23699), .B(n23664), .Z(n23672) );
  XOR U24915 ( .A(n23700), .B(n23652), .Z(n23664) );
  XOR U24916 ( .A(n23701), .B(n23702), .Z(n23652) );
  ANDN U24917 ( .B(n23703), .A(n23704), .Z(n23701) );
  XOR U24918 ( .A(n23702), .B(n23705), .Z(n23703) );
  IV U24919 ( .A(n23650), .Z(n23700) );
  XOR U24920 ( .A(n23648), .B(n23706), .Z(n23650) );
  XOR U24921 ( .A(n23707), .B(n23708), .Z(n23706) );
  ANDN U24922 ( .B(n23709), .A(n23710), .Z(n23707) );
  XOR U24923 ( .A(n23711), .B(n23708), .Z(n23709) );
  IV U24924 ( .A(n23651), .Z(n23648) );
  XOR U24925 ( .A(n23712), .B(n23713), .Z(n23651) );
  ANDN U24926 ( .B(n23714), .A(n23715), .Z(n23712) );
  XOR U24927 ( .A(n23713), .B(n23716), .Z(n23714) );
  IV U24928 ( .A(n23663), .Z(n23699) );
  XOR U24929 ( .A(n23717), .B(n23718), .Z(n23663) );
  XNOR U24930 ( .A(n23658), .B(n23719), .Z(n23718) );
  IV U24931 ( .A(n23661), .Z(n23719) );
  XOR U24932 ( .A(n23720), .B(n23721), .Z(n23661) );
  ANDN U24933 ( .B(n23722), .A(n23723), .Z(n23720) );
  XOR U24934 ( .A(n23721), .B(n23724), .Z(n23722) );
  XNOR U24935 ( .A(n23725), .B(n23726), .Z(n23658) );
  ANDN U24936 ( .B(n23727), .A(n23728), .Z(n23725) );
  XOR U24937 ( .A(n23726), .B(n23729), .Z(n23727) );
  IV U24938 ( .A(n23657), .Z(n23717) );
  XOR U24939 ( .A(n23655), .B(n23730), .Z(n23657) );
  XOR U24940 ( .A(n23731), .B(n23732), .Z(n23730) );
  ANDN U24941 ( .B(n23733), .A(n23734), .Z(n23731) );
  XOR U24942 ( .A(n23735), .B(n23732), .Z(n23733) );
  IV U24943 ( .A(n23659), .Z(n23655) );
  XOR U24944 ( .A(n23736), .B(n23737), .Z(n23659) );
  ANDN U24945 ( .B(n23738), .A(n23739), .Z(n23736) );
  XOR U24946 ( .A(n23740), .B(n23737), .Z(n23738) );
  XOR U24947 ( .A(n23741), .B(n23742), .Z(n23671) );
  XOR U24948 ( .A(n23689), .B(n23743), .Z(n23742) );
  IV U24949 ( .A(n23669), .Z(n23743) );
  XOR U24950 ( .A(n23744), .B(n23745), .Z(n23669) );
  ANDN U24951 ( .B(n23746), .A(n23747), .Z(n23744) );
  XOR U24952 ( .A(n23745), .B(n23748), .Z(n23746) );
  XOR U24953 ( .A(n23749), .B(n23677), .Z(n23689) );
  XOR U24954 ( .A(n23750), .B(n23751), .Z(n23677) );
  ANDN U24955 ( .B(n23752), .A(n23753), .Z(n23750) );
  XOR U24956 ( .A(n23751), .B(n23754), .Z(n23752) );
  IV U24957 ( .A(n23676), .Z(n23749) );
  XOR U24958 ( .A(n23755), .B(n23756), .Z(n23676) );
  XOR U24959 ( .A(n23757), .B(n23758), .Z(n23756) );
  ANDN U24960 ( .B(n23759), .A(n23760), .Z(n23757) );
  XOR U24961 ( .A(n23761), .B(n23758), .Z(n23759) );
  IV U24962 ( .A(n23674), .Z(n23755) );
  XOR U24963 ( .A(n23762), .B(n23763), .Z(n23674) );
  ANDN U24964 ( .B(n23764), .A(n23765), .Z(n23762) );
  XOR U24965 ( .A(n23763), .B(n23766), .Z(n23764) );
  IV U24966 ( .A(n23688), .Z(n23741) );
  XOR U24967 ( .A(n23767), .B(n23768), .Z(n23688) );
  XNOR U24968 ( .A(n23683), .B(n23769), .Z(n23768) );
  IV U24969 ( .A(n23686), .Z(n23769) );
  XOR U24970 ( .A(n23770), .B(n23771), .Z(n23686) );
  ANDN U24971 ( .B(n23772), .A(n23773), .Z(n23770) );
  XOR U24972 ( .A(n23774), .B(n23771), .Z(n23772) );
  XNOR U24973 ( .A(n23775), .B(n23776), .Z(n23683) );
  ANDN U24974 ( .B(n23777), .A(n23778), .Z(n23775) );
  XOR U24975 ( .A(n23776), .B(n23779), .Z(n23777) );
  IV U24976 ( .A(n23682), .Z(n23767) );
  XOR U24977 ( .A(n23680), .B(n23780), .Z(n23682) );
  XOR U24978 ( .A(n23781), .B(n23782), .Z(n23780) );
  ANDN U24979 ( .B(n23783), .A(n23784), .Z(n23781) );
  XOR U24980 ( .A(n23785), .B(n23782), .Z(n23783) );
  IV U24981 ( .A(n23684), .Z(n23680) );
  XOR U24982 ( .A(n23786), .B(n23787), .Z(n23684) );
  ANDN U24983 ( .B(n23788), .A(n23789), .Z(n23786) );
  XOR U24984 ( .A(n23790), .B(n23787), .Z(n23788) );
  IV U24985 ( .A(n23694), .Z(n23698) );
  XOR U24986 ( .A(n23694), .B(n23597), .Z(n23696) );
  XOR U24987 ( .A(n23791), .B(n23792), .Z(n23597) );
  AND U24988 ( .A(n244), .B(n23793), .Z(n23791) );
  XOR U24989 ( .A(n23794), .B(n23792), .Z(n23793) );
  NANDN U24990 ( .A(n23599), .B(n23601), .Z(n23694) );
  XOR U24991 ( .A(n23795), .B(n23796), .Z(n23601) );
  AND U24992 ( .A(n244), .B(n23797), .Z(n23795) );
  XOR U24993 ( .A(n23796), .B(n23798), .Z(n23797) );
  XNOR U24994 ( .A(n23799), .B(n23800), .Z(n244) );
  AND U24995 ( .A(n23801), .B(n23802), .Z(n23799) );
  XOR U24996 ( .A(n23800), .B(n23612), .Z(n23802) );
  XNOR U24997 ( .A(n23803), .B(n23804), .Z(n23612) );
  ANDN U24998 ( .B(n23805), .A(n23806), .Z(n23803) );
  XOR U24999 ( .A(n23804), .B(n23807), .Z(n23805) );
  XNOR U25000 ( .A(n23800), .B(n23614), .Z(n23801) );
  XOR U25001 ( .A(n23808), .B(n23809), .Z(n23614) );
  AND U25002 ( .A(n248), .B(n23810), .Z(n23808) );
  XOR U25003 ( .A(n23811), .B(n23809), .Z(n23810) );
  XOR U25004 ( .A(n23812), .B(n23813), .Z(n23800) );
  AND U25005 ( .A(n23814), .B(n23815), .Z(n23812) );
  XOR U25006 ( .A(n23813), .B(n23639), .Z(n23815) );
  XOR U25007 ( .A(n23806), .B(n23807), .Z(n23639) );
  XNOR U25008 ( .A(n23816), .B(n23817), .Z(n23807) );
  ANDN U25009 ( .B(n23818), .A(n23819), .Z(n23816) );
  XOR U25010 ( .A(n23820), .B(n23821), .Z(n23818) );
  XOR U25011 ( .A(n23822), .B(n23823), .Z(n23806) );
  XNOR U25012 ( .A(n23824), .B(n23825), .Z(n23823) );
  ANDN U25013 ( .B(n23826), .A(n23827), .Z(n23824) );
  XNOR U25014 ( .A(n23828), .B(n23829), .Z(n23826) );
  IV U25015 ( .A(n23804), .Z(n23822) );
  XOR U25016 ( .A(n23830), .B(n23831), .Z(n23804) );
  ANDN U25017 ( .B(n23832), .A(n23833), .Z(n23830) );
  XOR U25018 ( .A(n23831), .B(n23834), .Z(n23832) );
  XNOR U25019 ( .A(n23813), .B(n23641), .Z(n23814) );
  XOR U25020 ( .A(n23835), .B(n23836), .Z(n23641) );
  AND U25021 ( .A(n248), .B(n23837), .Z(n23835) );
  XOR U25022 ( .A(n23838), .B(n23836), .Z(n23837) );
  XNOR U25023 ( .A(n23839), .B(n23840), .Z(n23813) );
  AND U25024 ( .A(n23841), .B(n23842), .Z(n23839) );
  XNOR U25025 ( .A(n23840), .B(n23691), .Z(n23842) );
  XOR U25026 ( .A(n23833), .B(n23834), .Z(n23691) );
  XOR U25027 ( .A(n23843), .B(n23821), .Z(n23834) );
  XNOR U25028 ( .A(n23844), .B(n23845), .Z(n23821) );
  ANDN U25029 ( .B(n23846), .A(n23847), .Z(n23844) );
  XOR U25030 ( .A(n23848), .B(n23849), .Z(n23846) );
  IV U25031 ( .A(n23819), .Z(n23843) );
  XOR U25032 ( .A(n23817), .B(n23850), .Z(n23819) );
  XNOR U25033 ( .A(n23851), .B(n23852), .Z(n23850) );
  ANDN U25034 ( .B(n23853), .A(n23854), .Z(n23851) );
  XNOR U25035 ( .A(n23855), .B(n23856), .Z(n23853) );
  IV U25036 ( .A(n23820), .Z(n23817) );
  XOR U25037 ( .A(n23857), .B(n23858), .Z(n23820) );
  ANDN U25038 ( .B(n23859), .A(n23860), .Z(n23857) );
  XOR U25039 ( .A(n23858), .B(n23861), .Z(n23859) );
  XOR U25040 ( .A(n23862), .B(n23863), .Z(n23833) );
  XNOR U25041 ( .A(n23828), .B(n23864), .Z(n23863) );
  IV U25042 ( .A(n23831), .Z(n23864) );
  XOR U25043 ( .A(n23865), .B(n23866), .Z(n23831) );
  ANDN U25044 ( .B(n23867), .A(n23868), .Z(n23865) );
  XOR U25045 ( .A(n23866), .B(n23869), .Z(n23867) );
  XNOR U25046 ( .A(n23870), .B(n23871), .Z(n23828) );
  ANDN U25047 ( .B(n23872), .A(n23873), .Z(n23870) );
  XOR U25048 ( .A(n23871), .B(n23874), .Z(n23872) );
  IV U25049 ( .A(n23827), .Z(n23862) );
  XOR U25050 ( .A(n23825), .B(n23875), .Z(n23827) );
  XNOR U25051 ( .A(n23876), .B(n23877), .Z(n23875) );
  ANDN U25052 ( .B(n23878), .A(n23879), .Z(n23876) );
  XNOR U25053 ( .A(n23880), .B(n23881), .Z(n23878) );
  IV U25054 ( .A(n23829), .Z(n23825) );
  XOR U25055 ( .A(n23882), .B(n23883), .Z(n23829) );
  ANDN U25056 ( .B(n23884), .A(n23885), .Z(n23882) );
  XOR U25057 ( .A(n23886), .B(n23883), .Z(n23884) );
  XOR U25058 ( .A(n23840), .B(n23693), .Z(n23841) );
  XOR U25059 ( .A(n23887), .B(n23888), .Z(n23693) );
  AND U25060 ( .A(n248), .B(n23889), .Z(n23887) );
  XOR U25061 ( .A(n23890), .B(n23888), .Z(n23889) );
  XNOR U25062 ( .A(n23891), .B(n23892), .Z(n23840) );
  NAND U25063 ( .A(n23893), .B(n23894), .Z(n23892) );
  XOR U25064 ( .A(n23895), .B(n23792), .Z(n23894) );
  XOR U25065 ( .A(n23868), .B(n23869), .Z(n23792) );
  XOR U25066 ( .A(n23896), .B(n23861), .Z(n23869) );
  XOR U25067 ( .A(n23897), .B(n23849), .Z(n23861) );
  XOR U25068 ( .A(n23898), .B(n23899), .Z(n23849) );
  ANDN U25069 ( .B(n23900), .A(n23901), .Z(n23898) );
  XOR U25070 ( .A(n23899), .B(n23902), .Z(n23900) );
  IV U25071 ( .A(n23847), .Z(n23897) );
  XOR U25072 ( .A(n23845), .B(n23903), .Z(n23847) );
  XOR U25073 ( .A(n23904), .B(n23905), .Z(n23903) );
  ANDN U25074 ( .B(n23906), .A(n23907), .Z(n23904) );
  XOR U25075 ( .A(n23908), .B(n23905), .Z(n23906) );
  IV U25076 ( .A(n23848), .Z(n23845) );
  XOR U25077 ( .A(n23909), .B(n23910), .Z(n23848) );
  ANDN U25078 ( .B(n23911), .A(n23912), .Z(n23909) );
  XOR U25079 ( .A(n23910), .B(n23913), .Z(n23911) );
  IV U25080 ( .A(n23860), .Z(n23896) );
  XOR U25081 ( .A(n23914), .B(n23915), .Z(n23860) );
  XNOR U25082 ( .A(n23855), .B(n23916), .Z(n23915) );
  IV U25083 ( .A(n23858), .Z(n23916) );
  XOR U25084 ( .A(n23917), .B(n23918), .Z(n23858) );
  ANDN U25085 ( .B(n23919), .A(n23920), .Z(n23917) );
  XOR U25086 ( .A(n23918), .B(n23921), .Z(n23919) );
  XNOR U25087 ( .A(n23922), .B(n23923), .Z(n23855) );
  ANDN U25088 ( .B(n23924), .A(n23925), .Z(n23922) );
  XOR U25089 ( .A(n23923), .B(n23926), .Z(n23924) );
  IV U25090 ( .A(n23854), .Z(n23914) );
  XOR U25091 ( .A(n23852), .B(n23927), .Z(n23854) );
  XOR U25092 ( .A(n23928), .B(n23929), .Z(n23927) );
  ANDN U25093 ( .B(n23930), .A(n23931), .Z(n23928) );
  XOR U25094 ( .A(n23932), .B(n23929), .Z(n23930) );
  IV U25095 ( .A(n23856), .Z(n23852) );
  XOR U25096 ( .A(n23933), .B(n23934), .Z(n23856) );
  ANDN U25097 ( .B(n23935), .A(n23936), .Z(n23933) );
  XOR U25098 ( .A(n23937), .B(n23934), .Z(n23935) );
  XOR U25099 ( .A(n23938), .B(n23939), .Z(n23868) );
  XOR U25100 ( .A(n23886), .B(n23940), .Z(n23939) );
  IV U25101 ( .A(n23866), .Z(n23940) );
  XOR U25102 ( .A(n23941), .B(n23942), .Z(n23866) );
  ANDN U25103 ( .B(n23943), .A(n23944), .Z(n23941) );
  XOR U25104 ( .A(n23942), .B(n23945), .Z(n23943) );
  XOR U25105 ( .A(n23946), .B(n23874), .Z(n23886) );
  XOR U25106 ( .A(n23947), .B(n23948), .Z(n23874) );
  ANDN U25107 ( .B(n23949), .A(n23950), .Z(n23947) );
  XOR U25108 ( .A(n23948), .B(n23951), .Z(n23949) );
  IV U25109 ( .A(n23873), .Z(n23946) );
  XOR U25110 ( .A(n23952), .B(n23953), .Z(n23873) );
  XOR U25111 ( .A(n23954), .B(n23955), .Z(n23953) );
  ANDN U25112 ( .B(n23956), .A(n23957), .Z(n23954) );
  XOR U25113 ( .A(n23958), .B(n23955), .Z(n23956) );
  IV U25114 ( .A(n23871), .Z(n23952) );
  XOR U25115 ( .A(n23959), .B(n23960), .Z(n23871) );
  ANDN U25116 ( .B(n23961), .A(n23962), .Z(n23959) );
  XOR U25117 ( .A(n23960), .B(n23963), .Z(n23961) );
  IV U25118 ( .A(n23885), .Z(n23938) );
  XOR U25119 ( .A(n23964), .B(n23965), .Z(n23885) );
  XNOR U25120 ( .A(n23880), .B(n23966), .Z(n23965) );
  IV U25121 ( .A(n23883), .Z(n23966) );
  XOR U25122 ( .A(n23967), .B(n23968), .Z(n23883) );
  ANDN U25123 ( .B(n23969), .A(n23970), .Z(n23967) );
  XOR U25124 ( .A(n23971), .B(n23968), .Z(n23969) );
  XNOR U25125 ( .A(n23972), .B(n23973), .Z(n23880) );
  ANDN U25126 ( .B(n23974), .A(n23975), .Z(n23972) );
  XOR U25127 ( .A(n23973), .B(n23976), .Z(n23974) );
  IV U25128 ( .A(n23879), .Z(n23964) );
  XOR U25129 ( .A(n23877), .B(n23977), .Z(n23879) );
  XOR U25130 ( .A(n23978), .B(n23979), .Z(n23977) );
  ANDN U25131 ( .B(n23980), .A(n23981), .Z(n23978) );
  XOR U25132 ( .A(n23982), .B(n23979), .Z(n23980) );
  IV U25133 ( .A(n23881), .Z(n23877) );
  XOR U25134 ( .A(n23983), .B(n23984), .Z(n23881) );
  ANDN U25135 ( .B(n23985), .A(n23986), .Z(n23983) );
  XOR U25136 ( .A(n23987), .B(n23984), .Z(n23985) );
  IV U25137 ( .A(n23891), .Z(n23895) );
  XOR U25138 ( .A(n23891), .B(n23794), .Z(n23893) );
  XOR U25139 ( .A(n23988), .B(n23989), .Z(n23794) );
  AND U25140 ( .A(n248), .B(n23990), .Z(n23988) );
  XOR U25141 ( .A(n23991), .B(n23989), .Z(n23990) );
  NANDN U25142 ( .A(n23796), .B(n23798), .Z(n23891) );
  XOR U25143 ( .A(n23992), .B(n23993), .Z(n23798) );
  AND U25144 ( .A(n248), .B(n23994), .Z(n23992) );
  XOR U25145 ( .A(n23993), .B(n23995), .Z(n23994) );
  XNOR U25146 ( .A(n23996), .B(n23997), .Z(n248) );
  AND U25147 ( .A(n23998), .B(n23999), .Z(n23996) );
  XOR U25148 ( .A(n23997), .B(n23809), .Z(n23999) );
  XNOR U25149 ( .A(n24000), .B(n24001), .Z(n23809) );
  ANDN U25150 ( .B(n24002), .A(n24003), .Z(n24000) );
  XOR U25151 ( .A(n24001), .B(n24004), .Z(n24002) );
  XNOR U25152 ( .A(n23997), .B(n23811), .Z(n23998) );
  XOR U25153 ( .A(n24005), .B(n24006), .Z(n23811) );
  AND U25154 ( .A(n252), .B(n24007), .Z(n24005) );
  XOR U25155 ( .A(n24008), .B(n24006), .Z(n24007) );
  XOR U25156 ( .A(n24009), .B(n24010), .Z(n23997) );
  AND U25157 ( .A(n24011), .B(n24012), .Z(n24009) );
  XOR U25158 ( .A(n24010), .B(n23836), .Z(n24012) );
  XOR U25159 ( .A(n24003), .B(n24004), .Z(n23836) );
  XNOR U25160 ( .A(n24013), .B(n24014), .Z(n24004) );
  ANDN U25161 ( .B(n24015), .A(n24016), .Z(n24013) );
  XOR U25162 ( .A(n24017), .B(n24018), .Z(n24015) );
  XOR U25163 ( .A(n24019), .B(n24020), .Z(n24003) );
  XNOR U25164 ( .A(n24021), .B(n24022), .Z(n24020) );
  ANDN U25165 ( .B(n24023), .A(n24024), .Z(n24021) );
  XNOR U25166 ( .A(n24025), .B(n24026), .Z(n24023) );
  IV U25167 ( .A(n24001), .Z(n24019) );
  XOR U25168 ( .A(n24027), .B(n24028), .Z(n24001) );
  ANDN U25169 ( .B(n24029), .A(n24030), .Z(n24027) );
  XOR U25170 ( .A(n24028), .B(n24031), .Z(n24029) );
  XNOR U25171 ( .A(n24010), .B(n23838), .Z(n24011) );
  XOR U25172 ( .A(n24032), .B(n24033), .Z(n23838) );
  AND U25173 ( .A(n252), .B(n24034), .Z(n24032) );
  XOR U25174 ( .A(n24035), .B(n24033), .Z(n24034) );
  XNOR U25175 ( .A(n24036), .B(n24037), .Z(n24010) );
  AND U25176 ( .A(n24038), .B(n24039), .Z(n24036) );
  XNOR U25177 ( .A(n24037), .B(n23888), .Z(n24039) );
  XOR U25178 ( .A(n24030), .B(n24031), .Z(n23888) );
  XOR U25179 ( .A(n24040), .B(n24018), .Z(n24031) );
  XNOR U25180 ( .A(n24041), .B(n24042), .Z(n24018) );
  ANDN U25181 ( .B(n24043), .A(n24044), .Z(n24041) );
  XOR U25182 ( .A(n24045), .B(n24046), .Z(n24043) );
  IV U25183 ( .A(n24016), .Z(n24040) );
  XOR U25184 ( .A(n24014), .B(n24047), .Z(n24016) );
  XNOR U25185 ( .A(n24048), .B(n24049), .Z(n24047) );
  ANDN U25186 ( .B(n24050), .A(n24051), .Z(n24048) );
  XNOR U25187 ( .A(n24052), .B(n24053), .Z(n24050) );
  IV U25188 ( .A(n24017), .Z(n24014) );
  XOR U25189 ( .A(n24054), .B(n24055), .Z(n24017) );
  ANDN U25190 ( .B(n24056), .A(n24057), .Z(n24054) );
  XOR U25191 ( .A(n24055), .B(n24058), .Z(n24056) );
  XOR U25192 ( .A(n24059), .B(n24060), .Z(n24030) );
  XNOR U25193 ( .A(n24025), .B(n24061), .Z(n24060) );
  IV U25194 ( .A(n24028), .Z(n24061) );
  XOR U25195 ( .A(n24062), .B(n24063), .Z(n24028) );
  ANDN U25196 ( .B(n24064), .A(n24065), .Z(n24062) );
  XOR U25197 ( .A(n24063), .B(n24066), .Z(n24064) );
  XNOR U25198 ( .A(n24067), .B(n24068), .Z(n24025) );
  ANDN U25199 ( .B(n24069), .A(n24070), .Z(n24067) );
  XOR U25200 ( .A(n24068), .B(n24071), .Z(n24069) );
  IV U25201 ( .A(n24024), .Z(n24059) );
  XOR U25202 ( .A(n24022), .B(n24072), .Z(n24024) );
  XNOR U25203 ( .A(n24073), .B(n24074), .Z(n24072) );
  ANDN U25204 ( .B(n24075), .A(n24076), .Z(n24073) );
  XNOR U25205 ( .A(n24077), .B(n24078), .Z(n24075) );
  IV U25206 ( .A(n24026), .Z(n24022) );
  XOR U25207 ( .A(n24079), .B(n24080), .Z(n24026) );
  ANDN U25208 ( .B(n24081), .A(n24082), .Z(n24079) );
  XOR U25209 ( .A(n24083), .B(n24080), .Z(n24081) );
  XOR U25210 ( .A(n24037), .B(n23890), .Z(n24038) );
  XOR U25211 ( .A(n24084), .B(n24085), .Z(n23890) );
  AND U25212 ( .A(n252), .B(n24086), .Z(n24084) );
  XOR U25213 ( .A(n24087), .B(n24085), .Z(n24086) );
  XNOR U25214 ( .A(n24088), .B(n24089), .Z(n24037) );
  NAND U25215 ( .A(n24090), .B(n24091), .Z(n24089) );
  XOR U25216 ( .A(n24092), .B(n23989), .Z(n24091) );
  XOR U25217 ( .A(n24065), .B(n24066), .Z(n23989) );
  XOR U25218 ( .A(n24093), .B(n24058), .Z(n24066) );
  XOR U25219 ( .A(n24094), .B(n24046), .Z(n24058) );
  XOR U25220 ( .A(n24095), .B(n24096), .Z(n24046) );
  ANDN U25221 ( .B(n24097), .A(n24098), .Z(n24095) );
  XOR U25222 ( .A(n24096), .B(n24099), .Z(n24097) );
  IV U25223 ( .A(n24044), .Z(n24094) );
  XOR U25224 ( .A(n24042), .B(n24100), .Z(n24044) );
  XOR U25225 ( .A(n24101), .B(n24102), .Z(n24100) );
  ANDN U25226 ( .B(n24103), .A(n24104), .Z(n24101) );
  XOR U25227 ( .A(n24105), .B(n24102), .Z(n24103) );
  IV U25228 ( .A(n24045), .Z(n24042) );
  XOR U25229 ( .A(n24106), .B(n24107), .Z(n24045) );
  ANDN U25230 ( .B(n24108), .A(n24109), .Z(n24106) );
  XOR U25231 ( .A(n24107), .B(n24110), .Z(n24108) );
  IV U25232 ( .A(n24057), .Z(n24093) );
  XOR U25233 ( .A(n24111), .B(n24112), .Z(n24057) );
  XNOR U25234 ( .A(n24052), .B(n24113), .Z(n24112) );
  IV U25235 ( .A(n24055), .Z(n24113) );
  XOR U25236 ( .A(n24114), .B(n24115), .Z(n24055) );
  ANDN U25237 ( .B(n24116), .A(n24117), .Z(n24114) );
  XOR U25238 ( .A(n24115), .B(n24118), .Z(n24116) );
  XNOR U25239 ( .A(n24119), .B(n24120), .Z(n24052) );
  ANDN U25240 ( .B(n24121), .A(n24122), .Z(n24119) );
  XOR U25241 ( .A(n24120), .B(n24123), .Z(n24121) );
  IV U25242 ( .A(n24051), .Z(n24111) );
  XOR U25243 ( .A(n24049), .B(n24124), .Z(n24051) );
  XOR U25244 ( .A(n24125), .B(n24126), .Z(n24124) );
  ANDN U25245 ( .B(n24127), .A(n24128), .Z(n24125) );
  XOR U25246 ( .A(n24129), .B(n24126), .Z(n24127) );
  IV U25247 ( .A(n24053), .Z(n24049) );
  XOR U25248 ( .A(n24130), .B(n24131), .Z(n24053) );
  ANDN U25249 ( .B(n24132), .A(n24133), .Z(n24130) );
  XOR U25250 ( .A(n24134), .B(n24131), .Z(n24132) );
  XOR U25251 ( .A(n24135), .B(n24136), .Z(n24065) );
  XOR U25252 ( .A(n24083), .B(n24137), .Z(n24136) );
  IV U25253 ( .A(n24063), .Z(n24137) );
  XOR U25254 ( .A(n24138), .B(n24139), .Z(n24063) );
  ANDN U25255 ( .B(n24140), .A(n24141), .Z(n24138) );
  XOR U25256 ( .A(n24139), .B(n24142), .Z(n24140) );
  XOR U25257 ( .A(n24143), .B(n24071), .Z(n24083) );
  XOR U25258 ( .A(n24144), .B(n24145), .Z(n24071) );
  ANDN U25259 ( .B(n24146), .A(n24147), .Z(n24144) );
  XOR U25260 ( .A(n24145), .B(n24148), .Z(n24146) );
  IV U25261 ( .A(n24070), .Z(n24143) );
  XOR U25262 ( .A(n24149), .B(n24150), .Z(n24070) );
  XOR U25263 ( .A(n24151), .B(n24152), .Z(n24150) );
  ANDN U25264 ( .B(n24153), .A(n24154), .Z(n24151) );
  XOR U25265 ( .A(n24155), .B(n24152), .Z(n24153) );
  IV U25266 ( .A(n24068), .Z(n24149) );
  XOR U25267 ( .A(n24156), .B(n24157), .Z(n24068) );
  ANDN U25268 ( .B(n24158), .A(n24159), .Z(n24156) );
  XOR U25269 ( .A(n24157), .B(n24160), .Z(n24158) );
  IV U25270 ( .A(n24082), .Z(n24135) );
  XOR U25271 ( .A(n24161), .B(n24162), .Z(n24082) );
  XNOR U25272 ( .A(n24077), .B(n24163), .Z(n24162) );
  IV U25273 ( .A(n24080), .Z(n24163) );
  XOR U25274 ( .A(n24164), .B(n24165), .Z(n24080) );
  ANDN U25275 ( .B(n24166), .A(n24167), .Z(n24164) );
  XOR U25276 ( .A(n24168), .B(n24165), .Z(n24166) );
  XNOR U25277 ( .A(n24169), .B(n24170), .Z(n24077) );
  ANDN U25278 ( .B(n24171), .A(n24172), .Z(n24169) );
  XOR U25279 ( .A(n24170), .B(n24173), .Z(n24171) );
  IV U25280 ( .A(n24076), .Z(n24161) );
  XOR U25281 ( .A(n24074), .B(n24174), .Z(n24076) );
  XOR U25282 ( .A(n24175), .B(n24176), .Z(n24174) );
  ANDN U25283 ( .B(n24177), .A(n24178), .Z(n24175) );
  XOR U25284 ( .A(n24179), .B(n24176), .Z(n24177) );
  IV U25285 ( .A(n24078), .Z(n24074) );
  XOR U25286 ( .A(n24180), .B(n24181), .Z(n24078) );
  ANDN U25287 ( .B(n24182), .A(n24183), .Z(n24180) );
  XOR U25288 ( .A(n24184), .B(n24181), .Z(n24182) );
  IV U25289 ( .A(n24088), .Z(n24092) );
  XOR U25290 ( .A(n24088), .B(n23991), .Z(n24090) );
  XOR U25291 ( .A(n24185), .B(n24186), .Z(n23991) );
  AND U25292 ( .A(n252), .B(n24187), .Z(n24185) );
  XOR U25293 ( .A(n24188), .B(n24186), .Z(n24187) );
  NANDN U25294 ( .A(n23993), .B(n23995), .Z(n24088) );
  XOR U25295 ( .A(n24189), .B(n24190), .Z(n23995) );
  AND U25296 ( .A(n252), .B(n24191), .Z(n24189) );
  XOR U25297 ( .A(n24190), .B(n24192), .Z(n24191) );
  XNOR U25298 ( .A(n24193), .B(n24194), .Z(n252) );
  AND U25299 ( .A(n24195), .B(n24196), .Z(n24193) );
  XOR U25300 ( .A(n24194), .B(n24006), .Z(n24196) );
  XNOR U25301 ( .A(n24197), .B(n24198), .Z(n24006) );
  ANDN U25302 ( .B(n24199), .A(n24200), .Z(n24197) );
  XOR U25303 ( .A(n24198), .B(n24201), .Z(n24199) );
  XNOR U25304 ( .A(n24194), .B(n24008), .Z(n24195) );
  XOR U25305 ( .A(n24202), .B(n24203), .Z(n24008) );
  AND U25306 ( .A(n256), .B(n24204), .Z(n24202) );
  XOR U25307 ( .A(n24205), .B(n24203), .Z(n24204) );
  XOR U25308 ( .A(n24206), .B(n24207), .Z(n24194) );
  AND U25309 ( .A(n24208), .B(n24209), .Z(n24206) );
  XOR U25310 ( .A(n24207), .B(n24033), .Z(n24209) );
  XOR U25311 ( .A(n24200), .B(n24201), .Z(n24033) );
  XNOR U25312 ( .A(n24210), .B(n24211), .Z(n24201) );
  ANDN U25313 ( .B(n24212), .A(n24213), .Z(n24210) );
  XOR U25314 ( .A(n24214), .B(n24215), .Z(n24212) );
  XOR U25315 ( .A(n24216), .B(n24217), .Z(n24200) );
  XNOR U25316 ( .A(n24218), .B(n24219), .Z(n24217) );
  ANDN U25317 ( .B(n24220), .A(n24221), .Z(n24218) );
  XNOR U25318 ( .A(n24222), .B(n24223), .Z(n24220) );
  IV U25319 ( .A(n24198), .Z(n24216) );
  XOR U25320 ( .A(n24224), .B(n24225), .Z(n24198) );
  ANDN U25321 ( .B(n24226), .A(n24227), .Z(n24224) );
  XOR U25322 ( .A(n24225), .B(n24228), .Z(n24226) );
  XNOR U25323 ( .A(n24207), .B(n24035), .Z(n24208) );
  XOR U25324 ( .A(n24229), .B(n24230), .Z(n24035) );
  AND U25325 ( .A(n256), .B(n24231), .Z(n24229) );
  XOR U25326 ( .A(n24232), .B(n24230), .Z(n24231) );
  XNOR U25327 ( .A(n24233), .B(n24234), .Z(n24207) );
  AND U25328 ( .A(n24235), .B(n24236), .Z(n24233) );
  XNOR U25329 ( .A(n24234), .B(n24085), .Z(n24236) );
  XOR U25330 ( .A(n24227), .B(n24228), .Z(n24085) );
  XOR U25331 ( .A(n24237), .B(n24215), .Z(n24228) );
  XNOR U25332 ( .A(n24238), .B(n24239), .Z(n24215) );
  ANDN U25333 ( .B(n24240), .A(n24241), .Z(n24238) );
  XOR U25334 ( .A(n24242), .B(n24243), .Z(n24240) );
  IV U25335 ( .A(n24213), .Z(n24237) );
  XOR U25336 ( .A(n24211), .B(n24244), .Z(n24213) );
  XNOR U25337 ( .A(n24245), .B(n24246), .Z(n24244) );
  ANDN U25338 ( .B(n24247), .A(n24248), .Z(n24245) );
  XNOR U25339 ( .A(n24249), .B(n24250), .Z(n24247) );
  IV U25340 ( .A(n24214), .Z(n24211) );
  XOR U25341 ( .A(n24251), .B(n24252), .Z(n24214) );
  ANDN U25342 ( .B(n24253), .A(n24254), .Z(n24251) );
  XOR U25343 ( .A(n24252), .B(n24255), .Z(n24253) );
  XOR U25344 ( .A(n24256), .B(n24257), .Z(n24227) );
  XNOR U25345 ( .A(n24222), .B(n24258), .Z(n24257) );
  IV U25346 ( .A(n24225), .Z(n24258) );
  XOR U25347 ( .A(n24259), .B(n24260), .Z(n24225) );
  ANDN U25348 ( .B(n24261), .A(n24262), .Z(n24259) );
  XOR U25349 ( .A(n24260), .B(n24263), .Z(n24261) );
  XNOR U25350 ( .A(n24264), .B(n24265), .Z(n24222) );
  ANDN U25351 ( .B(n24266), .A(n24267), .Z(n24264) );
  XOR U25352 ( .A(n24265), .B(n24268), .Z(n24266) );
  IV U25353 ( .A(n24221), .Z(n24256) );
  XOR U25354 ( .A(n24219), .B(n24269), .Z(n24221) );
  XNOR U25355 ( .A(n24270), .B(n24271), .Z(n24269) );
  ANDN U25356 ( .B(n24272), .A(n24273), .Z(n24270) );
  XNOR U25357 ( .A(n24274), .B(n24275), .Z(n24272) );
  IV U25358 ( .A(n24223), .Z(n24219) );
  XOR U25359 ( .A(n24276), .B(n24277), .Z(n24223) );
  ANDN U25360 ( .B(n24278), .A(n24279), .Z(n24276) );
  XOR U25361 ( .A(n24280), .B(n24277), .Z(n24278) );
  XOR U25362 ( .A(n24234), .B(n24087), .Z(n24235) );
  XOR U25363 ( .A(n24281), .B(n24282), .Z(n24087) );
  AND U25364 ( .A(n256), .B(n24283), .Z(n24281) );
  XOR U25365 ( .A(n24284), .B(n24282), .Z(n24283) );
  XNOR U25366 ( .A(n24285), .B(n24286), .Z(n24234) );
  NAND U25367 ( .A(n24287), .B(n24288), .Z(n24286) );
  XOR U25368 ( .A(n24289), .B(n24186), .Z(n24288) );
  XOR U25369 ( .A(n24262), .B(n24263), .Z(n24186) );
  XOR U25370 ( .A(n24290), .B(n24255), .Z(n24263) );
  XOR U25371 ( .A(n24291), .B(n24243), .Z(n24255) );
  XOR U25372 ( .A(n24292), .B(n24293), .Z(n24243) );
  ANDN U25373 ( .B(n24294), .A(n24295), .Z(n24292) );
  XOR U25374 ( .A(n24293), .B(n24296), .Z(n24294) );
  IV U25375 ( .A(n24241), .Z(n24291) );
  XOR U25376 ( .A(n24239), .B(n24297), .Z(n24241) );
  XOR U25377 ( .A(n24298), .B(n24299), .Z(n24297) );
  ANDN U25378 ( .B(n24300), .A(n24301), .Z(n24298) );
  XOR U25379 ( .A(n24302), .B(n24299), .Z(n24300) );
  IV U25380 ( .A(n24242), .Z(n24239) );
  XOR U25381 ( .A(n24303), .B(n24304), .Z(n24242) );
  ANDN U25382 ( .B(n24305), .A(n24306), .Z(n24303) );
  XOR U25383 ( .A(n24304), .B(n24307), .Z(n24305) );
  IV U25384 ( .A(n24254), .Z(n24290) );
  XOR U25385 ( .A(n24308), .B(n24309), .Z(n24254) );
  XNOR U25386 ( .A(n24249), .B(n24310), .Z(n24309) );
  IV U25387 ( .A(n24252), .Z(n24310) );
  XOR U25388 ( .A(n24311), .B(n24312), .Z(n24252) );
  ANDN U25389 ( .B(n24313), .A(n24314), .Z(n24311) );
  XOR U25390 ( .A(n24312), .B(n24315), .Z(n24313) );
  XNOR U25391 ( .A(n24316), .B(n24317), .Z(n24249) );
  ANDN U25392 ( .B(n24318), .A(n24319), .Z(n24316) );
  XOR U25393 ( .A(n24317), .B(n24320), .Z(n24318) );
  IV U25394 ( .A(n24248), .Z(n24308) );
  XOR U25395 ( .A(n24246), .B(n24321), .Z(n24248) );
  XOR U25396 ( .A(n24322), .B(n24323), .Z(n24321) );
  ANDN U25397 ( .B(n24324), .A(n24325), .Z(n24322) );
  XOR U25398 ( .A(n24326), .B(n24323), .Z(n24324) );
  IV U25399 ( .A(n24250), .Z(n24246) );
  XOR U25400 ( .A(n24327), .B(n24328), .Z(n24250) );
  ANDN U25401 ( .B(n24329), .A(n24330), .Z(n24327) );
  XOR U25402 ( .A(n24331), .B(n24328), .Z(n24329) );
  XOR U25403 ( .A(n24332), .B(n24333), .Z(n24262) );
  XOR U25404 ( .A(n24280), .B(n24334), .Z(n24333) );
  IV U25405 ( .A(n24260), .Z(n24334) );
  XOR U25406 ( .A(n24335), .B(n24336), .Z(n24260) );
  ANDN U25407 ( .B(n24337), .A(n24338), .Z(n24335) );
  XOR U25408 ( .A(n24336), .B(n24339), .Z(n24337) );
  XOR U25409 ( .A(n24340), .B(n24268), .Z(n24280) );
  XOR U25410 ( .A(n24341), .B(n24342), .Z(n24268) );
  ANDN U25411 ( .B(n24343), .A(n24344), .Z(n24341) );
  XOR U25412 ( .A(n24342), .B(n24345), .Z(n24343) );
  IV U25413 ( .A(n24267), .Z(n24340) );
  XOR U25414 ( .A(n24346), .B(n24347), .Z(n24267) );
  XOR U25415 ( .A(n24348), .B(n24349), .Z(n24347) );
  ANDN U25416 ( .B(n24350), .A(n24351), .Z(n24348) );
  XOR U25417 ( .A(n24352), .B(n24349), .Z(n24350) );
  IV U25418 ( .A(n24265), .Z(n24346) );
  XOR U25419 ( .A(n24353), .B(n24354), .Z(n24265) );
  ANDN U25420 ( .B(n24355), .A(n24356), .Z(n24353) );
  XOR U25421 ( .A(n24354), .B(n24357), .Z(n24355) );
  IV U25422 ( .A(n24279), .Z(n24332) );
  XOR U25423 ( .A(n24358), .B(n24359), .Z(n24279) );
  XNOR U25424 ( .A(n24274), .B(n24360), .Z(n24359) );
  IV U25425 ( .A(n24277), .Z(n24360) );
  XOR U25426 ( .A(n24361), .B(n24362), .Z(n24277) );
  ANDN U25427 ( .B(n24363), .A(n24364), .Z(n24361) );
  XOR U25428 ( .A(n24365), .B(n24362), .Z(n24363) );
  XNOR U25429 ( .A(n24366), .B(n24367), .Z(n24274) );
  ANDN U25430 ( .B(n24368), .A(n24369), .Z(n24366) );
  XOR U25431 ( .A(n24367), .B(n24370), .Z(n24368) );
  IV U25432 ( .A(n24273), .Z(n24358) );
  XOR U25433 ( .A(n24271), .B(n24371), .Z(n24273) );
  XOR U25434 ( .A(n24372), .B(n24373), .Z(n24371) );
  ANDN U25435 ( .B(n24374), .A(n24375), .Z(n24372) );
  XOR U25436 ( .A(n24376), .B(n24373), .Z(n24374) );
  IV U25437 ( .A(n24275), .Z(n24271) );
  XOR U25438 ( .A(n24377), .B(n24378), .Z(n24275) );
  ANDN U25439 ( .B(n24379), .A(n24380), .Z(n24377) );
  XOR U25440 ( .A(n24381), .B(n24378), .Z(n24379) );
  IV U25441 ( .A(n24285), .Z(n24289) );
  XOR U25442 ( .A(n24285), .B(n24188), .Z(n24287) );
  XOR U25443 ( .A(n24382), .B(n24383), .Z(n24188) );
  AND U25444 ( .A(n256), .B(n24384), .Z(n24382) );
  XOR U25445 ( .A(n24385), .B(n24383), .Z(n24384) );
  NANDN U25446 ( .A(n24190), .B(n24192), .Z(n24285) );
  XOR U25447 ( .A(n24386), .B(n24387), .Z(n24192) );
  AND U25448 ( .A(n256), .B(n24388), .Z(n24386) );
  XOR U25449 ( .A(n24387), .B(n24389), .Z(n24388) );
  XNOR U25450 ( .A(n24390), .B(n24391), .Z(n256) );
  AND U25451 ( .A(n24392), .B(n24393), .Z(n24390) );
  XOR U25452 ( .A(n24391), .B(n24203), .Z(n24393) );
  XNOR U25453 ( .A(n24394), .B(n24395), .Z(n24203) );
  ANDN U25454 ( .B(n24396), .A(n24397), .Z(n24394) );
  XOR U25455 ( .A(n24395), .B(n24398), .Z(n24396) );
  XNOR U25456 ( .A(n24391), .B(n24205), .Z(n24392) );
  XOR U25457 ( .A(n24399), .B(n24400), .Z(n24205) );
  AND U25458 ( .A(n260), .B(n24401), .Z(n24399) );
  XOR U25459 ( .A(n24402), .B(n24400), .Z(n24401) );
  XOR U25460 ( .A(n24403), .B(n24404), .Z(n24391) );
  AND U25461 ( .A(n24405), .B(n24406), .Z(n24403) );
  XOR U25462 ( .A(n24404), .B(n24230), .Z(n24406) );
  XOR U25463 ( .A(n24397), .B(n24398), .Z(n24230) );
  XNOR U25464 ( .A(n24407), .B(n24408), .Z(n24398) );
  ANDN U25465 ( .B(n24409), .A(n24410), .Z(n24407) );
  XOR U25466 ( .A(n24411), .B(n24412), .Z(n24409) );
  XOR U25467 ( .A(n24413), .B(n24414), .Z(n24397) );
  XNOR U25468 ( .A(n24415), .B(n24416), .Z(n24414) );
  ANDN U25469 ( .B(n24417), .A(n24418), .Z(n24415) );
  XNOR U25470 ( .A(n24419), .B(n24420), .Z(n24417) );
  IV U25471 ( .A(n24395), .Z(n24413) );
  XOR U25472 ( .A(n24421), .B(n24422), .Z(n24395) );
  ANDN U25473 ( .B(n24423), .A(n24424), .Z(n24421) );
  XOR U25474 ( .A(n24422), .B(n24425), .Z(n24423) );
  XNOR U25475 ( .A(n24404), .B(n24232), .Z(n24405) );
  XOR U25476 ( .A(n24426), .B(n24427), .Z(n24232) );
  AND U25477 ( .A(n260), .B(n24428), .Z(n24426) );
  XOR U25478 ( .A(n24429), .B(n24427), .Z(n24428) );
  XNOR U25479 ( .A(n24430), .B(n24431), .Z(n24404) );
  AND U25480 ( .A(n24432), .B(n24433), .Z(n24430) );
  XNOR U25481 ( .A(n24431), .B(n24282), .Z(n24433) );
  XOR U25482 ( .A(n24424), .B(n24425), .Z(n24282) );
  XOR U25483 ( .A(n24434), .B(n24412), .Z(n24425) );
  XNOR U25484 ( .A(n24435), .B(n24436), .Z(n24412) );
  ANDN U25485 ( .B(n24437), .A(n24438), .Z(n24435) );
  XOR U25486 ( .A(n24439), .B(n24440), .Z(n24437) );
  IV U25487 ( .A(n24410), .Z(n24434) );
  XOR U25488 ( .A(n24408), .B(n24441), .Z(n24410) );
  XNOR U25489 ( .A(n24442), .B(n24443), .Z(n24441) );
  ANDN U25490 ( .B(n24444), .A(n24445), .Z(n24442) );
  XNOR U25491 ( .A(n24446), .B(n24447), .Z(n24444) );
  IV U25492 ( .A(n24411), .Z(n24408) );
  XOR U25493 ( .A(n24448), .B(n24449), .Z(n24411) );
  ANDN U25494 ( .B(n24450), .A(n24451), .Z(n24448) );
  XOR U25495 ( .A(n24449), .B(n24452), .Z(n24450) );
  XOR U25496 ( .A(n24453), .B(n24454), .Z(n24424) );
  XNOR U25497 ( .A(n24419), .B(n24455), .Z(n24454) );
  IV U25498 ( .A(n24422), .Z(n24455) );
  XOR U25499 ( .A(n24456), .B(n24457), .Z(n24422) );
  ANDN U25500 ( .B(n24458), .A(n24459), .Z(n24456) );
  XOR U25501 ( .A(n24457), .B(n24460), .Z(n24458) );
  XNOR U25502 ( .A(n24461), .B(n24462), .Z(n24419) );
  ANDN U25503 ( .B(n24463), .A(n24464), .Z(n24461) );
  XOR U25504 ( .A(n24462), .B(n24465), .Z(n24463) );
  IV U25505 ( .A(n24418), .Z(n24453) );
  XOR U25506 ( .A(n24416), .B(n24466), .Z(n24418) );
  XNOR U25507 ( .A(n24467), .B(n24468), .Z(n24466) );
  ANDN U25508 ( .B(n24469), .A(n24470), .Z(n24467) );
  XNOR U25509 ( .A(n24471), .B(n24472), .Z(n24469) );
  IV U25510 ( .A(n24420), .Z(n24416) );
  XOR U25511 ( .A(n24473), .B(n24474), .Z(n24420) );
  ANDN U25512 ( .B(n24475), .A(n24476), .Z(n24473) );
  XOR U25513 ( .A(n24477), .B(n24474), .Z(n24475) );
  XOR U25514 ( .A(n24431), .B(n24284), .Z(n24432) );
  XOR U25515 ( .A(n24478), .B(n24479), .Z(n24284) );
  AND U25516 ( .A(n260), .B(n24480), .Z(n24478) );
  XOR U25517 ( .A(n24481), .B(n24479), .Z(n24480) );
  XNOR U25518 ( .A(n24482), .B(n24483), .Z(n24431) );
  NAND U25519 ( .A(n24484), .B(n24485), .Z(n24483) );
  XOR U25520 ( .A(n24486), .B(n24383), .Z(n24485) );
  XOR U25521 ( .A(n24459), .B(n24460), .Z(n24383) );
  XOR U25522 ( .A(n24487), .B(n24452), .Z(n24460) );
  XOR U25523 ( .A(n24488), .B(n24440), .Z(n24452) );
  XOR U25524 ( .A(n24489), .B(n24490), .Z(n24440) );
  ANDN U25525 ( .B(n24491), .A(n24492), .Z(n24489) );
  XOR U25526 ( .A(n24490), .B(n24493), .Z(n24491) );
  IV U25527 ( .A(n24438), .Z(n24488) );
  XOR U25528 ( .A(n24436), .B(n24494), .Z(n24438) );
  XOR U25529 ( .A(n24495), .B(n24496), .Z(n24494) );
  ANDN U25530 ( .B(n24497), .A(n24498), .Z(n24495) );
  XOR U25531 ( .A(n24499), .B(n24496), .Z(n24497) );
  IV U25532 ( .A(n24439), .Z(n24436) );
  XOR U25533 ( .A(n24500), .B(n24501), .Z(n24439) );
  ANDN U25534 ( .B(n24502), .A(n24503), .Z(n24500) );
  XOR U25535 ( .A(n24501), .B(n24504), .Z(n24502) );
  IV U25536 ( .A(n24451), .Z(n24487) );
  XOR U25537 ( .A(n24505), .B(n24506), .Z(n24451) );
  XNOR U25538 ( .A(n24446), .B(n24507), .Z(n24506) );
  IV U25539 ( .A(n24449), .Z(n24507) );
  XOR U25540 ( .A(n24508), .B(n24509), .Z(n24449) );
  ANDN U25541 ( .B(n24510), .A(n24511), .Z(n24508) );
  XOR U25542 ( .A(n24509), .B(n24512), .Z(n24510) );
  XNOR U25543 ( .A(n24513), .B(n24514), .Z(n24446) );
  ANDN U25544 ( .B(n24515), .A(n24516), .Z(n24513) );
  XOR U25545 ( .A(n24514), .B(n24517), .Z(n24515) );
  IV U25546 ( .A(n24445), .Z(n24505) );
  XOR U25547 ( .A(n24443), .B(n24518), .Z(n24445) );
  XOR U25548 ( .A(n24519), .B(n24520), .Z(n24518) );
  ANDN U25549 ( .B(n24521), .A(n24522), .Z(n24519) );
  XOR U25550 ( .A(n24523), .B(n24520), .Z(n24521) );
  IV U25551 ( .A(n24447), .Z(n24443) );
  XOR U25552 ( .A(n24524), .B(n24525), .Z(n24447) );
  ANDN U25553 ( .B(n24526), .A(n24527), .Z(n24524) );
  XOR U25554 ( .A(n24528), .B(n24525), .Z(n24526) );
  XOR U25555 ( .A(n24529), .B(n24530), .Z(n24459) );
  XOR U25556 ( .A(n24477), .B(n24531), .Z(n24530) );
  IV U25557 ( .A(n24457), .Z(n24531) );
  XOR U25558 ( .A(n24532), .B(n24533), .Z(n24457) );
  ANDN U25559 ( .B(n24534), .A(n24535), .Z(n24532) );
  XOR U25560 ( .A(n24533), .B(n24536), .Z(n24534) );
  XOR U25561 ( .A(n24537), .B(n24465), .Z(n24477) );
  XOR U25562 ( .A(n24538), .B(n24539), .Z(n24465) );
  ANDN U25563 ( .B(n24540), .A(n24541), .Z(n24538) );
  XOR U25564 ( .A(n24539), .B(n24542), .Z(n24540) );
  IV U25565 ( .A(n24464), .Z(n24537) );
  XOR U25566 ( .A(n24543), .B(n24544), .Z(n24464) );
  XOR U25567 ( .A(n24545), .B(n24546), .Z(n24544) );
  ANDN U25568 ( .B(n24547), .A(n24548), .Z(n24545) );
  XOR U25569 ( .A(n24549), .B(n24546), .Z(n24547) );
  IV U25570 ( .A(n24462), .Z(n24543) );
  XOR U25571 ( .A(n24550), .B(n24551), .Z(n24462) );
  ANDN U25572 ( .B(n24552), .A(n24553), .Z(n24550) );
  XOR U25573 ( .A(n24551), .B(n24554), .Z(n24552) );
  IV U25574 ( .A(n24476), .Z(n24529) );
  XOR U25575 ( .A(n24555), .B(n24556), .Z(n24476) );
  XNOR U25576 ( .A(n24471), .B(n24557), .Z(n24556) );
  IV U25577 ( .A(n24474), .Z(n24557) );
  XOR U25578 ( .A(n24558), .B(n24559), .Z(n24474) );
  ANDN U25579 ( .B(n24560), .A(n24561), .Z(n24558) );
  XOR U25580 ( .A(n24562), .B(n24559), .Z(n24560) );
  XNOR U25581 ( .A(n24563), .B(n24564), .Z(n24471) );
  ANDN U25582 ( .B(n24565), .A(n24566), .Z(n24563) );
  XOR U25583 ( .A(n24564), .B(n24567), .Z(n24565) );
  IV U25584 ( .A(n24470), .Z(n24555) );
  XOR U25585 ( .A(n24468), .B(n24568), .Z(n24470) );
  XOR U25586 ( .A(n24569), .B(n24570), .Z(n24568) );
  ANDN U25587 ( .B(n24571), .A(n24572), .Z(n24569) );
  XOR U25588 ( .A(n24573), .B(n24570), .Z(n24571) );
  IV U25589 ( .A(n24472), .Z(n24468) );
  XOR U25590 ( .A(n24574), .B(n24575), .Z(n24472) );
  ANDN U25591 ( .B(n24576), .A(n24577), .Z(n24574) );
  XOR U25592 ( .A(n24578), .B(n24575), .Z(n24576) );
  IV U25593 ( .A(n24482), .Z(n24486) );
  XOR U25594 ( .A(n24482), .B(n24385), .Z(n24484) );
  XOR U25595 ( .A(n24579), .B(n24580), .Z(n24385) );
  AND U25596 ( .A(n260), .B(n24581), .Z(n24579) );
  XOR U25597 ( .A(n24582), .B(n24580), .Z(n24581) );
  NANDN U25598 ( .A(n24387), .B(n24389), .Z(n24482) );
  XOR U25599 ( .A(n24583), .B(n24584), .Z(n24389) );
  AND U25600 ( .A(n260), .B(n24585), .Z(n24583) );
  XOR U25601 ( .A(n24584), .B(n24586), .Z(n24585) );
  XNOR U25602 ( .A(n24587), .B(n24588), .Z(n260) );
  AND U25603 ( .A(n24589), .B(n24590), .Z(n24587) );
  XOR U25604 ( .A(n24588), .B(n24400), .Z(n24590) );
  XNOR U25605 ( .A(n24591), .B(n24592), .Z(n24400) );
  ANDN U25606 ( .B(n24593), .A(n24594), .Z(n24591) );
  XOR U25607 ( .A(n24592), .B(n24595), .Z(n24593) );
  XNOR U25608 ( .A(n24588), .B(n24402), .Z(n24589) );
  XOR U25609 ( .A(n24596), .B(n24597), .Z(n24402) );
  AND U25610 ( .A(n264), .B(n24598), .Z(n24596) );
  XOR U25611 ( .A(n24599), .B(n24597), .Z(n24598) );
  XOR U25612 ( .A(n24600), .B(n24601), .Z(n24588) );
  AND U25613 ( .A(n24602), .B(n24603), .Z(n24600) );
  XOR U25614 ( .A(n24601), .B(n24427), .Z(n24603) );
  XOR U25615 ( .A(n24594), .B(n24595), .Z(n24427) );
  XNOR U25616 ( .A(n24604), .B(n24605), .Z(n24595) );
  ANDN U25617 ( .B(n24606), .A(n24607), .Z(n24604) );
  XOR U25618 ( .A(n24608), .B(n24609), .Z(n24606) );
  XOR U25619 ( .A(n24610), .B(n24611), .Z(n24594) );
  XNOR U25620 ( .A(n24612), .B(n24613), .Z(n24611) );
  ANDN U25621 ( .B(n24614), .A(n24615), .Z(n24612) );
  XNOR U25622 ( .A(n24616), .B(n24617), .Z(n24614) );
  IV U25623 ( .A(n24592), .Z(n24610) );
  XOR U25624 ( .A(n24618), .B(n24619), .Z(n24592) );
  ANDN U25625 ( .B(n24620), .A(n24621), .Z(n24618) );
  XOR U25626 ( .A(n24619), .B(n24622), .Z(n24620) );
  XNOR U25627 ( .A(n24601), .B(n24429), .Z(n24602) );
  XOR U25628 ( .A(n24623), .B(n24624), .Z(n24429) );
  AND U25629 ( .A(n264), .B(n24625), .Z(n24623) );
  XOR U25630 ( .A(n24626), .B(n24624), .Z(n24625) );
  XNOR U25631 ( .A(n24627), .B(n24628), .Z(n24601) );
  AND U25632 ( .A(n24629), .B(n24630), .Z(n24627) );
  XNOR U25633 ( .A(n24628), .B(n24479), .Z(n24630) );
  XOR U25634 ( .A(n24621), .B(n24622), .Z(n24479) );
  XOR U25635 ( .A(n24631), .B(n24609), .Z(n24622) );
  XNOR U25636 ( .A(n24632), .B(n24633), .Z(n24609) );
  ANDN U25637 ( .B(n24634), .A(n24635), .Z(n24632) );
  XOR U25638 ( .A(n24636), .B(n24637), .Z(n24634) );
  IV U25639 ( .A(n24607), .Z(n24631) );
  XOR U25640 ( .A(n24605), .B(n24638), .Z(n24607) );
  XNOR U25641 ( .A(n24639), .B(n24640), .Z(n24638) );
  ANDN U25642 ( .B(n24641), .A(n24642), .Z(n24639) );
  XNOR U25643 ( .A(n24643), .B(n24644), .Z(n24641) );
  IV U25644 ( .A(n24608), .Z(n24605) );
  XOR U25645 ( .A(n24645), .B(n24646), .Z(n24608) );
  ANDN U25646 ( .B(n24647), .A(n24648), .Z(n24645) );
  XOR U25647 ( .A(n24646), .B(n24649), .Z(n24647) );
  XOR U25648 ( .A(n24650), .B(n24651), .Z(n24621) );
  XNOR U25649 ( .A(n24616), .B(n24652), .Z(n24651) );
  IV U25650 ( .A(n24619), .Z(n24652) );
  XOR U25651 ( .A(n24653), .B(n24654), .Z(n24619) );
  ANDN U25652 ( .B(n24655), .A(n24656), .Z(n24653) );
  XOR U25653 ( .A(n24654), .B(n24657), .Z(n24655) );
  XNOR U25654 ( .A(n24658), .B(n24659), .Z(n24616) );
  ANDN U25655 ( .B(n24660), .A(n24661), .Z(n24658) );
  XOR U25656 ( .A(n24659), .B(n24662), .Z(n24660) );
  IV U25657 ( .A(n24615), .Z(n24650) );
  XOR U25658 ( .A(n24613), .B(n24663), .Z(n24615) );
  XNOR U25659 ( .A(n24664), .B(n24665), .Z(n24663) );
  ANDN U25660 ( .B(n24666), .A(n24667), .Z(n24664) );
  XNOR U25661 ( .A(n24668), .B(n24669), .Z(n24666) );
  IV U25662 ( .A(n24617), .Z(n24613) );
  XOR U25663 ( .A(n24670), .B(n24671), .Z(n24617) );
  ANDN U25664 ( .B(n24672), .A(n24673), .Z(n24670) );
  XOR U25665 ( .A(n24674), .B(n24671), .Z(n24672) );
  XOR U25666 ( .A(n24628), .B(n24481), .Z(n24629) );
  XOR U25667 ( .A(n24675), .B(n24676), .Z(n24481) );
  AND U25668 ( .A(n264), .B(n24677), .Z(n24675) );
  XOR U25669 ( .A(n24678), .B(n24676), .Z(n24677) );
  XNOR U25670 ( .A(n24679), .B(n24680), .Z(n24628) );
  NAND U25671 ( .A(n24681), .B(n24682), .Z(n24680) );
  XOR U25672 ( .A(n24683), .B(n24580), .Z(n24682) );
  XOR U25673 ( .A(n24656), .B(n24657), .Z(n24580) );
  XOR U25674 ( .A(n24684), .B(n24649), .Z(n24657) );
  XOR U25675 ( .A(n24685), .B(n24637), .Z(n24649) );
  XOR U25676 ( .A(n24686), .B(n24687), .Z(n24637) );
  ANDN U25677 ( .B(n24688), .A(n24689), .Z(n24686) );
  XOR U25678 ( .A(n24687), .B(n24690), .Z(n24688) );
  IV U25679 ( .A(n24635), .Z(n24685) );
  XOR U25680 ( .A(n24633), .B(n24691), .Z(n24635) );
  XOR U25681 ( .A(n24692), .B(n24693), .Z(n24691) );
  ANDN U25682 ( .B(n24694), .A(n24695), .Z(n24692) );
  XOR U25683 ( .A(n24696), .B(n24693), .Z(n24694) );
  IV U25684 ( .A(n24636), .Z(n24633) );
  XOR U25685 ( .A(n24697), .B(n24698), .Z(n24636) );
  ANDN U25686 ( .B(n24699), .A(n24700), .Z(n24697) );
  XOR U25687 ( .A(n24698), .B(n24701), .Z(n24699) );
  IV U25688 ( .A(n24648), .Z(n24684) );
  XOR U25689 ( .A(n24702), .B(n24703), .Z(n24648) );
  XNOR U25690 ( .A(n24643), .B(n24704), .Z(n24703) );
  IV U25691 ( .A(n24646), .Z(n24704) );
  XOR U25692 ( .A(n24705), .B(n24706), .Z(n24646) );
  ANDN U25693 ( .B(n24707), .A(n24708), .Z(n24705) );
  XOR U25694 ( .A(n24706), .B(n24709), .Z(n24707) );
  XNOR U25695 ( .A(n24710), .B(n24711), .Z(n24643) );
  ANDN U25696 ( .B(n24712), .A(n24713), .Z(n24710) );
  XOR U25697 ( .A(n24711), .B(n24714), .Z(n24712) );
  IV U25698 ( .A(n24642), .Z(n24702) );
  XOR U25699 ( .A(n24640), .B(n24715), .Z(n24642) );
  XOR U25700 ( .A(n24716), .B(n24717), .Z(n24715) );
  ANDN U25701 ( .B(n24718), .A(n24719), .Z(n24716) );
  XOR U25702 ( .A(n24720), .B(n24717), .Z(n24718) );
  IV U25703 ( .A(n24644), .Z(n24640) );
  XOR U25704 ( .A(n24721), .B(n24722), .Z(n24644) );
  ANDN U25705 ( .B(n24723), .A(n24724), .Z(n24721) );
  XOR U25706 ( .A(n24725), .B(n24722), .Z(n24723) );
  XOR U25707 ( .A(n24726), .B(n24727), .Z(n24656) );
  XOR U25708 ( .A(n24674), .B(n24728), .Z(n24727) );
  IV U25709 ( .A(n24654), .Z(n24728) );
  XOR U25710 ( .A(n24729), .B(n24730), .Z(n24654) );
  ANDN U25711 ( .B(n24731), .A(n24732), .Z(n24729) );
  XOR U25712 ( .A(n24730), .B(n24733), .Z(n24731) );
  XOR U25713 ( .A(n24734), .B(n24662), .Z(n24674) );
  XOR U25714 ( .A(n24735), .B(n24736), .Z(n24662) );
  ANDN U25715 ( .B(n24737), .A(n24738), .Z(n24735) );
  XOR U25716 ( .A(n24736), .B(n24739), .Z(n24737) );
  IV U25717 ( .A(n24661), .Z(n24734) );
  XOR U25718 ( .A(n24740), .B(n24741), .Z(n24661) );
  XOR U25719 ( .A(n24742), .B(n24743), .Z(n24741) );
  ANDN U25720 ( .B(n24744), .A(n24745), .Z(n24742) );
  XOR U25721 ( .A(n24746), .B(n24743), .Z(n24744) );
  IV U25722 ( .A(n24659), .Z(n24740) );
  XOR U25723 ( .A(n24747), .B(n24748), .Z(n24659) );
  ANDN U25724 ( .B(n24749), .A(n24750), .Z(n24747) );
  XOR U25725 ( .A(n24748), .B(n24751), .Z(n24749) );
  IV U25726 ( .A(n24673), .Z(n24726) );
  XOR U25727 ( .A(n24752), .B(n24753), .Z(n24673) );
  XNOR U25728 ( .A(n24668), .B(n24754), .Z(n24753) );
  IV U25729 ( .A(n24671), .Z(n24754) );
  XOR U25730 ( .A(n24755), .B(n24756), .Z(n24671) );
  ANDN U25731 ( .B(n24757), .A(n24758), .Z(n24755) );
  XOR U25732 ( .A(n24759), .B(n24756), .Z(n24757) );
  XNOR U25733 ( .A(n24760), .B(n24761), .Z(n24668) );
  ANDN U25734 ( .B(n24762), .A(n24763), .Z(n24760) );
  XOR U25735 ( .A(n24761), .B(n24764), .Z(n24762) );
  IV U25736 ( .A(n24667), .Z(n24752) );
  XOR U25737 ( .A(n24665), .B(n24765), .Z(n24667) );
  XOR U25738 ( .A(n24766), .B(n24767), .Z(n24765) );
  ANDN U25739 ( .B(n24768), .A(n24769), .Z(n24766) );
  XOR U25740 ( .A(n24770), .B(n24767), .Z(n24768) );
  IV U25741 ( .A(n24669), .Z(n24665) );
  XOR U25742 ( .A(n24771), .B(n24772), .Z(n24669) );
  ANDN U25743 ( .B(n24773), .A(n24774), .Z(n24771) );
  XOR U25744 ( .A(n24775), .B(n24772), .Z(n24773) );
  IV U25745 ( .A(n24679), .Z(n24683) );
  XOR U25746 ( .A(n24679), .B(n24582), .Z(n24681) );
  XOR U25747 ( .A(n24776), .B(n24777), .Z(n24582) );
  AND U25748 ( .A(n264), .B(n24778), .Z(n24776) );
  XOR U25749 ( .A(n24779), .B(n24777), .Z(n24778) );
  NANDN U25750 ( .A(n24584), .B(n24586), .Z(n24679) );
  XOR U25751 ( .A(n24780), .B(n24781), .Z(n24586) );
  AND U25752 ( .A(n264), .B(n24782), .Z(n24780) );
  XOR U25753 ( .A(n24781), .B(n24783), .Z(n24782) );
  XNOR U25754 ( .A(n24784), .B(n24785), .Z(n264) );
  AND U25755 ( .A(n24786), .B(n24787), .Z(n24784) );
  XOR U25756 ( .A(n24785), .B(n24597), .Z(n24787) );
  XNOR U25757 ( .A(n24788), .B(n24789), .Z(n24597) );
  ANDN U25758 ( .B(n24790), .A(n24791), .Z(n24788) );
  XOR U25759 ( .A(n24789), .B(n24792), .Z(n24790) );
  XNOR U25760 ( .A(n24785), .B(n24599), .Z(n24786) );
  XOR U25761 ( .A(n24793), .B(n24794), .Z(n24599) );
  AND U25762 ( .A(n268), .B(n24795), .Z(n24793) );
  XOR U25763 ( .A(n24796), .B(n24794), .Z(n24795) );
  XOR U25764 ( .A(n24797), .B(n24798), .Z(n24785) );
  AND U25765 ( .A(n24799), .B(n24800), .Z(n24797) );
  XOR U25766 ( .A(n24798), .B(n24624), .Z(n24800) );
  XOR U25767 ( .A(n24791), .B(n24792), .Z(n24624) );
  XNOR U25768 ( .A(n24801), .B(n24802), .Z(n24792) );
  ANDN U25769 ( .B(n24803), .A(n24804), .Z(n24801) );
  XOR U25770 ( .A(n24805), .B(n24806), .Z(n24803) );
  XOR U25771 ( .A(n24807), .B(n24808), .Z(n24791) );
  XNOR U25772 ( .A(n24809), .B(n24810), .Z(n24808) );
  ANDN U25773 ( .B(n24811), .A(n24812), .Z(n24809) );
  XNOR U25774 ( .A(n24813), .B(n24814), .Z(n24811) );
  IV U25775 ( .A(n24789), .Z(n24807) );
  XOR U25776 ( .A(n24815), .B(n24816), .Z(n24789) );
  ANDN U25777 ( .B(n24817), .A(n24818), .Z(n24815) );
  XOR U25778 ( .A(n24816), .B(n24819), .Z(n24817) );
  XNOR U25779 ( .A(n24798), .B(n24626), .Z(n24799) );
  XOR U25780 ( .A(n24820), .B(n24821), .Z(n24626) );
  AND U25781 ( .A(n268), .B(n24822), .Z(n24820) );
  XOR U25782 ( .A(n24823), .B(n24821), .Z(n24822) );
  XNOR U25783 ( .A(n24824), .B(n24825), .Z(n24798) );
  AND U25784 ( .A(n24826), .B(n24827), .Z(n24824) );
  XNOR U25785 ( .A(n24825), .B(n24676), .Z(n24827) );
  XOR U25786 ( .A(n24818), .B(n24819), .Z(n24676) );
  XOR U25787 ( .A(n24828), .B(n24806), .Z(n24819) );
  XNOR U25788 ( .A(n24829), .B(n24830), .Z(n24806) );
  ANDN U25789 ( .B(n24831), .A(n24832), .Z(n24829) );
  XOR U25790 ( .A(n24833), .B(n24834), .Z(n24831) );
  IV U25791 ( .A(n24804), .Z(n24828) );
  XOR U25792 ( .A(n24802), .B(n24835), .Z(n24804) );
  XNOR U25793 ( .A(n24836), .B(n24837), .Z(n24835) );
  ANDN U25794 ( .B(n24838), .A(n24839), .Z(n24836) );
  XNOR U25795 ( .A(n24840), .B(n24841), .Z(n24838) );
  IV U25796 ( .A(n24805), .Z(n24802) );
  XOR U25797 ( .A(n24842), .B(n24843), .Z(n24805) );
  ANDN U25798 ( .B(n24844), .A(n24845), .Z(n24842) );
  XOR U25799 ( .A(n24843), .B(n24846), .Z(n24844) );
  XOR U25800 ( .A(n24847), .B(n24848), .Z(n24818) );
  XNOR U25801 ( .A(n24813), .B(n24849), .Z(n24848) );
  IV U25802 ( .A(n24816), .Z(n24849) );
  XOR U25803 ( .A(n24850), .B(n24851), .Z(n24816) );
  ANDN U25804 ( .B(n24852), .A(n24853), .Z(n24850) );
  XOR U25805 ( .A(n24851), .B(n24854), .Z(n24852) );
  XNOR U25806 ( .A(n24855), .B(n24856), .Z(n24813) );
  ANDN U25807 ( .B(n24857), .A(n24858), .Z(n24855) );
  XOR U25808 ( .A(n24856), .B(n24859), .Z(n24857) );
  IV U25809 ( .A(n24812), .Z(n24847) );
  XOR U25810 ( .A(n24810), .B(n24860), .Z(n24812) );
  XNOR U25811 ( .A(n24861), .B(n24862), .Z(n24860) );
  ANDN U25812 ( .B(n24863), .A(n24864), .Z(n24861) );
  XNOR U25813 ( .A(n24865), .B(n24866), .Z(n24863) );
  IV U25814 ( .A(n24814), .Z(n24810) );
  XOR U25815 ( .A(n24867), .B(n24868), .Z(n24814) );
  ANDN U25816 ( .B(n24869), .A(n24870), .Z(n24867) );
  XOR U25817 ( .A(n24871), .B(n24868), .Z(n24869) );
  XOR U25818 ( .A(n24825), .B(n24678), .Z(n24826) );
  XOR U25819 ( .A(n24872), .B(n24873), .Z(n24678) );
  AND U25820 ( .A(n268), .B(n24874), .Z(n24872) );
  XOR U25821 ( .A(n24875), .B(n24873), .Z(n24874) );
  XNOR U25822 ( .A(n24876), .B(n24877), .Z(n24825) );
  NAND U25823 ( .A(n24878), .B(n24879), .Z(n24877) );
  XOR U25824 ( .A(n24880), .B(n24777), .Z(n24879) );
  XOR U25825 ( .A(n24853), .B(n24854), .Z(n24777) );
  XOR U25826 ( .A(n24881), .B(n24846), .Z(n24854) );
  XOR U25827 ( .A(n24882), .B(n24834), .Z(n24846) );
  XOR U25828 ( .A(n24883), .B(n24884), .Z(n24834) );
  ANDN U25829 ( .B(n24885), .A(n24886), .Z(n24883) );
  XOR U25830 ( .A(n24884), .B(n24887), .Z(n24885) );
  IV U25831 ( .A(n24832), .Z(n24882) );
  XOR U25832 ( .A(n24830), .B(n24888), .Z(n24832) );
  XOR U25833 ( .A(n24889), .B(n24890), .Z(n24888) );
  ANDN U25834 ( .B(n24891), .A(n24892), .Z(n24889) );
  XOR U25835 ( .A(n24893), .B(n24890), .Z(n24891) );
  IV U25836 ( .A(n24833), .Z(n24830) );
  XOR U25837 ( .A(n24894), .B(n24895), .Z(n24833) );
  ANDN U25838 ( .B(n24896), .A(n24897), .Z(n24894) );
  XOR U25839 ( .A(n24895), .B(n24898), .Z(n24896) );
  IV U25840 ( .A(n24845), .Z(n24881) );
  XOR U25841 ( .A(n24899), .B(n24900), .Z(n24845) );
  XNOR U25842 ( .A(n24840), .B(n24901), .Z(n24900) );
  IV U25843 ( .A(n24843), .Z(n24901) );
  XOR U25844 ( .A(n24902), .B(n24903), .Z(n24843) );
  ANDN U25845 ( .B(n24904), .A(n24905), .Z(n24902) );
  XOR U25846 ( .A(n24903), .B(n24906), .Z(n24904) );
  XNOR U25847 ( .A(n24907), .B(n24908), .Z(n24840) );
  ANDN U25848 ( .B(n24909), .A(n24910), .Z(n24907) );
  XOR U25849 ( .A(n24908), .B(n24911), .Z(n24909) );
  IV U25850 ( .A(n24839), .Z(n24899) );
  XOR U25851 ( .A(n24837), .B(n24912), .Z(n24839) );
  XOR U25852 ( .A(n24913), .B(n24914), .Z(n24912) );
  ANDN U25853 ( .B(n24915), .A(n24916), .Z(n24913) );
  XOR U25854 ( .A(n24917), .B(n24914), .Z(n24915) );
  IV U25855 ( .A(n24841), .Z(n24837) );
  XOR U25856 ( .A(n24918), .B(n24919), .Z(n24841) );
  ANDN U25857 ( .B(n24920), .A(n24921), .Z(n24918) );
  XOR U25858 ( .A(n24922), .B(n24919), .Z(n24920) );
  XOR U25859 ( .A(n24923), .B(n24924), .Z(n24853) );
  XOR U25860 ( .A(n24871), .B(n24925), .Z(n24924) );
  IV U25861 ( .A(n24851), .Z(n24925) );
  XOR U25862 ( .A(n24926), .B(n24927), .Z(n24851) );
  ANDN U25863 ( .B(n24928), .A(n24929), .Z(n24926) );
  XOR U25864 ( .A(n24927), .B(n24930), .Z(n24928) );
  XOR U25865 ( .A(n24931), .B(n24859), .Z(n24871) );
  XOR U25866 ( .A(n24932), .B(n24933), .Z(n24859) );
  ANDN U25867 ( .B(n24934), .A(n24935), .Z(n24932) );
  XOR U25868 ( .A(n24933), .B(n24936), .Z(n24934) );
  IV U25869 ( .A(n24858), .Z(n24931) );
  XOR U25870 ( .A(n24937), .B(n24938), .Z(n24858) );
  XOR U25871 ( .A(n24939), .B(n24940), .Z(n24938) );
  ANDN U25872 ( .B(n24941), .A(n24942), .Z(n24939) );
  XOR U25873 ( .A(n24943), .B(n24940), .Z(n24941) );
  IV U25874 ( .A(n24856), .Z(n24937) );
  XOR U25875 ( .A(n24944), .B(n24945), .Z(n24856) );
  ANDN U25876 ( .B(n24946), .A(n24947), .Z(n24944) );
  XOR U25877 ( .A(n24945), .B(n24948), .Z(n24946) );
  IV U25878 ( .A(n24870), .Z(n24923) );
  XOR U25879 ( .A(n24949), .B(n24950), .Z(n24870) );
  XNOR U25880 ( .A(n24865), .B(n24951), .Z(n24950) );
  IV U25881 ( .A(n24868), .Z(n24951) );
  XOR U25882 ( .A(n24952), .B(n24953), .Z(n24868) );
  ANDN U25883 ( .B(n24954), .A(n24955), .Z(n24952) );
  XOR U25884 ( .A(n24956), .B(n24953), .Z(n24954) );
  XNOR U25885 ( .A(n24957), .B(n24958), .Z(n24865) );
  ANDN U25886 ( .B(n24959), .A(n24960), .Z(n24957) );
  XOR U25887 ( .A(n24958), .B(n24961), .Z(n24959) );
  IV U25888 ( .A(n24864), .Z(n24949) );
  XOR U25889 ( .A(n24862), .B(n24962), .Z(n24864) );
  XOR U25890 ( .A(n24963), .B(n24964), .Z(n24962) );
  ANDN U25891 ( .B(n24965), .A(n24966), .Z(n24963) );
  XOR U25892 ( .A(n24967), .B(n24964), .Z(n24965) );
  IV U25893 ( .A(n24866), .Z(n24862) );
  XOR U25894 ( .A(n24968), .B(n24969), .Z(n24866) );
  ANDN U25895 ( .B(n24970), .A(n24971), .Z(n24968) );
  XOR U25896 ( .A(n24972), .B(n24969), .Z(n24970) );
  IV U25897 ( .A(n24876), .Z(n24880) );
  XOR U25898 ( .A(n24876), .B(n24779), .Z(n24878) );
  XOR U25899 ( .A(n24973), .B(n24974), .Z(n24779) );
  AND U25900 ( .A(n268), .B(n24975), .Z(n24973) );
  XOR U25901 ( .A(n24976), .B(n24974), .Z(n24975) );
  NANDN U25902 ( .A(n24781), .B(n24783), .Z(n24876) );
  XOR U25903 ( .A(n24977), .B(n24978), .Z(n24783) );
  AND U25904 ( .A(n268), .B(n24979), .Z(n24977) );
  XOR U25905 ( .A(n24978), .B(n24980), .Z(n24979) );
  XNOR U25906 ( .A(n24981), .B(n24982), .Z(n268) );
  AND U25907 ( .A(n24983), .B(n24984), .Z(n24981) );
  XOR U25908 ( .A(n24982), .B(n24794), .Z(n24984) );
  XNOR U25909 ( .A(n24985), .B(n24986), .Z(n24794) );
  ANDN U25910 ( .B(n24987), .A(n24988), .Z(n24985) );
  XOR U25911 ( .A(n24986), .B(n24989), .Z(n24987) );
  XNOR U25912 ( .A(n24982), .B(n24796), .Z(n24983) );
  XOR U25913 ( .A(n24990), .B(n24991), .Z(n24796) );
  AND U25914 ( .A(n272), .B(n24992), .Z(n24990) );
  XOR U25915 ( .A(n24993), .B(n24991), .Z(n24992) );
  XOR U25916 ( .A(n24994), .B(n24995), .Z(n24982) );
  AND U25917 ( .A(n24996), .B(n24997), .Z(n24994) );
  XOR U25918 ( .A(n24995), .B(n24821), .Z(n24997) );
  XOR U25919 ( .A(n24988), .B(n24989), .Z(n24821) );
  XNOR U25920 ( .A(n24998), .B(n24999), .Z(n24989) );
  ANDN U25921 ( .B(n25000), .A(n25001), .Z(n24998) );
  XOR U25922 ( .A(n25002), .B(n25003), .Z(n25000) );
  XOR U25923 ( .A(n25004), .B(n25005), .Z(n24988) );
  XNOR U25924 ( .A(n25006), .B(n25007), .Z(n25005) );
  ANDN U25925 ( .B(n25008), .A(n25009), .Z(n25006) );
  XNOR U25926 ( .A(n25010), .B(n25011), .Z(n25008) );
  IV U25927 ( .A(n24986), .Z(n25004) );
  XOR U25928 ( .A(n25012), .B(n25013), .Z(n24986) );
  ANDN U25929 ( .B(n25014), .A(n25015), .Z(n25012) );
  XOR U25930 ( .A(n25013), .B(n25016), .Z(n25014) );
  XNOR U25931 ( .A(n24995), .B(n24823), .Z(n24996) );
  XOR U25932 ( .A(n25017), .B(n25018), .Z(n24823) );
  AND U25933 ( .A(n272), .B(n25019), .Z(n25017) );
  XOR U25934 ( .A(n25020), .B(n25018), .Z(n25019) );
  XNOR U25935 ( .A(n25021), .B(n25022), .Z(n24995) );
  AND U25936 ( .A(n25023), .B(n25024), .Z(n25021) );
  XNOR U25937 ( .A(n25022), .B(n24873), .Z(n25024) );
  XOR U25938 ( .A(n25015), .B(n25016), .Z(n24873) );
  XOR U25939 ( .A(n25025), .B(n25003), .Z(n25016) );
  XNOR U25940 ( .A(n25026), .B(n25027), .Z(n25003) );
  ANDN U25941 ( .B(n25028), .A(n25029), .Z(n25026) );
  XOR U25942 ( .A(n25030), .B(n25031), .Z(n25028) );
  IV U25943 ( .A(n25001), .Z(n25025) );
  XOR U25944 ( .A(n24999), .B(n25032), .Z(n25001) );
  XNOR U25945 ( .A(n25033), .B(n25034), .Z(n25032) );
  ANDN U25946 ( .B(n25035), .A(n25036), .Z(n25033) );
  XNOR U25947 ( .A(n25037), .B(n25038), .Z(n25035) );
  IV U25948 ( .A(n25002), .Z(n24999) );
  XOR U25949 ( .A(n25039), .B(n25040), .Z(n25002) );
  ANDN U25950 ( .B(n25041), .A(n25042), .Z(n25039) );
  XOR U25951 ( .A(n25040), .B(n25043), .Z(n25041) );
  XOR U25952 ( .A(n25044), .B(n25045), .Z(n25015) );
  XNOR U25953 ( .A(n25010), .B(n25046), .Z(n25045) );
  IV U25954 ( .A(n25013), .Z(n25046) );
  XOR U25955 ( .A(n25047), .B(n25048), .Z(n25013) );
  ANDN U25956 ( .B(n25049), .A(n25050), .Z(n25047) );
  XOR U25957 ( .A(n25048), .B(n25051), .Z(n25049) );
  XNOR U25958 ( .A(n25052), .B(n25053), .Z(n25010) );
  ANDN U25959 ( .B(n25054), .A(n25055), .Z(n25052) );
  XOR U25960 ( .A(n25053), .B(n25056), .Z(n25054) );
  IV U25961 ( .A(n25009), .Z(n25044) );
  XOR U25962 ( .A(n25007), .B(n25057), .Z(n25009) );
  XNOR U25963 ( .A(n25058), .B(n25059), .Z(n25057) );
  ANDN U25964 ( .B(n25060), .A(n25061), .Z(n25058) );
  XNOR U25965 ( .A(n25062), .B(n25063), .Z(n25060) );
  IV U25966 ( .A(n25011), .Z(n25007) );
  XOR U25967 ( .A(n25064), .B(n25065), .Z(n25011) );
  ANDN U25968 ( .B(n25066), .A(n25067), .Z(n25064) );
  XOR U25969 ( .A(n25068), .B(n25065), .Z(n25066) );
  XOR U25970 ( .A(n25022), .B(n24875), .Z(n25023) );
  XOR U25971 ( .A(n25069), .B(n25070), .Z(n24875) );
  AND U25972 ( .A(n272), .B(n25071), .Z(n25069) );
  XOR U25973 ( .A(n25072), .B(n25070), .Z(n25071) );
  XNOR U25974 ( .A(n25073), .B(n25074), .Z(n25022) );
  NAND U25975 ( .A(n25075), .B(n25076), .Z(n25074) );
  XOR U25976 ( .A(n25077), .B(n24974), .Z(n25076) );
  XOR U25977 ( .A(n25050), .B(n25051), .Z(n24974) );
  XOR U25978 ( .A(n25078), .B(n25043), .Z(n25051) );
  XOR U25979 ( .A(n25079), .B(n25031), .Z(n25043) );
  XOR U25980 ( .A(n25080), .B(n25081), .Z(n25031) );
  ANDN U25981 ( .B(n25082), .A(n25083), .Z(n25080) );
  XOR U25982 ( .A(n25081), .B(n25084), .Z(n25082) );
  IV U25983 ( .A(n25029), .Z(n25079) );
  XOR U25984 ( .A(n25027), .B(n25085), .Z(n25029) );
  XOR U25985 ( .A(n25086), .B(n25087), .Z(n25085) );
  ANDN U25986 ( .B(n25088), .A(n25089), .Z(n25086) );
  XOR U25987 ( .A(n25090), .B(n25087), .Z(n25088) );
  IV U25988 ( .A(n25030), .Z(n25027) );
  XOR U25989 ( .A(n25091), .B(n25092), .Z(n25030) );
  ANDN U25990 ( .B(n25093), .A(n25094), .Z(n25091) );
  XOR U25991 ( .A(n25092), .B(n25095), .Z(n25093) );
  IV U25992 ( .A(n25042), .Z(n25078) );
  XOR U25993 ( .A(n25096), .B(n25097), .Z(n25042) );
  XNOR U25994 ( .A(n25037), .B(n25098), .Z(n25097) );
  IV U25995 ( .A(n25040), .Z(n25098) );
  XOR U25996 ( .A(n25099), .B(n25100), .Z(n25040) );
  ANDN U25997 ( .B(n25101), .A(n25102), .Z(n25099) );
  XOR U25998 ( .A(n25100), .B(n25103), .Z(n25101) );
  XNOR U25999 ( .A(n25104), .B(n25105), .Z(n25037) );
  ANDN U26000 ( .B(n25106), .A(n25107), .Z(n25104) );
  XOR U26001 ( .A(n25105), .B(n25108), .Z(n25106) );
  IV U26002 ( .A(n25036), .Z(n25096) );
  XOR U26003 ( .A(n25034), .B(n25109), .Z(n25036) );
  XOR U26004 ( .A(n25110), .B(n25111), .Z(n25109) );
  ANDN U26005 ( .B(n25112), .A(n25113), .Z(n25110) );
  XOR U26006 ( .A(n25114), .B(n25111), .Z(n25112) );
  IV U26007 ( .A(n25038), .Z(n25034) );
  XOR U26008 ( .A(n25115), .B(n25116), .Z(n25038) );
  ANDN U26009 ( .B(n25117), .A(n25118), .Z(n25115) );
  XOR U26010 ( .A(n25119), .B(n25116), .Z(n25117) );
  XOR U26011 ( .A(n25120), .B(n25121), .Z(n25050) );
  XOR U26012 ( .A(n25068), .B(n25122), .Z(n25121) );
  IV U26013 ( .A(n25048), .Z(n25122) );
  XOR U26014 ( .A(n25123), .B(n25124), .Z(n25048) );
  ANDN U26015 ( .B(n25125), .A(n25126), .Z(n25123) );
  XOR U26016 ( .A(n25124), .B(n25127), .Z(n25125) );
  XOR U26017 ( .A(n25128), .B(n25056), .Z(n25068) );
  XOR U26018 ( .A(n25129), .B(n25130), .Z(n25056) );
  ANDN U26019 ( .B(n25131), .A(n25132), .Z(n25129) );
  XOR U26020 ( .A(n25130), .B(n25133), .Z(n25131) );
  IV U26021 ( .A(n25055), .Z(n25128) );
  XOR U26022 ( .A(n25134), .B(n25135), .Z(n25055) );
  XOR U26023 ( .A(n25136), .B(n25137), .Z(n25135) );
  ANDN U26024 ( .B(n25138), .A(n25139), .Z(n25136) );
  XOR U26025 ( .A(n25140), .B(n25137), .Z(n25138) );
  IV U26026 ( .A(n25053), .Z(n25134) );
  XOR U26027 ( .A(n25141), .B(n25142), .Z(n25053) );
  ANDN U26028 ( .B(n25143), .A(n25144), .Z(n25141) );
  XOR U26029 ( .A(n25142), .B(n25145), .Z(n25143) );
  IV U26030 ( .A(n25067), .Z(n25120) );
  XOR U26031 ( .A(n25146), .B(n25147), .Z(n25067) );
  XNOR U26032 ( .A(n25062), .B(n25148), .Z(n25147) );
  IV U26033 ( .A(n25065), .Z(n25148) );
  XOR U26034 ( .A(n25149), .B(n25150), .Z(n25065) );
  ANDN U26035 ( .B(n25151), .A(n25152), .Z(n25149) );
  XOR U26036 ( .A(n25153), .B(n25150), .Z(n25151) );
  XNOR U26037 ( .A(n25154), .B(n25155), .Z(n25062) );
  ANDN U26038 ( .B(n25156), .A(n25157), .Z(n25154) );
  XOR U26039 ( .A(n25155), .B(n25158), .Z(n25156) );
  IV U26040 ( .A(n25061), .Z(n25146) );
  XOR U26041 ( .A(n25059), .B(n25159), .Z(n25061) );
  XOR U26042 ( .A(n25160), .B(n25161), .Z(n25159) );
  ANDN U26043 ( .B(n25162), .A(n25163), .Z(n25160) );
  XOR U26044 ( .A(n25164), .B(n25161), .Z(n25162) );
  IV U26045 ( .A(n25063), .Z(n25059) );
  XOR U26046 ( .A(n25165), .B(n25166), .Z(n25063) );
  ANDN U26047 ( .B(n25167), .A(n25168), .Z(n25165) );
  XOR U26048 ( .A(n25169), .B(n25166), .Z(n25167) );
  IV U26049 ( .A(n25073), .Z(n25077) );
  XOR U26050 ( .A(n25073), .B(n24976), .Z(n25075) );
  XOR U26051 ( .A(n25170), .B(n25171), .Z(n24976) );
  AND U26052 ( .A(n272), .B(n25172), .Z(n25170) );
  XOR U26053 ( .A(n25173), .B(n25171), .Z(n25172) );
  NANDN U26054 ( .A(n24978), .B(n24980), .Z(n25073) );
  XOR U26055 ( .A(n25174), .B(n25175), .Z(n24980) );
  AND U26056 ( .A(n272), .B(n25176), .Z(n25174) );
  XOR U26057 ( .A(n25175), .B(n25177), .Z(n25176) );
  XNOR U26058 ( .A(n25178), .B(n25179), .Z(n272) );
  AND U26059 ( .A(n25180), .B(n25181), .Z(n25178) );
  XOR U26060 ( .A(n25179), .B(n24991), .Z(n25181) );
  XNOR U26061 ( .A(n25182), .B(n25183), .Z(n24991) );
  ANDN U26062 ( .B(n25184), .A(n25185), .Z(n25182) );
  XOR U26063 ( .A(n25183), .B(n25186), .Z(n25184) );
  XNOR U26064 ( .A(n25179), .B(n24993), .Z(n25180) );
  XOR U26065 ( .A(n25187), .B(n25188), .Z(n24993) );
  AND U26066 ( .A(n276), .B(n25189), .Z(n25187) );
  XOR U26067 ( .A(n25190), .B(n25188), .Z(n25189) );
  XOR U26068 ( .A(n25191), .B(n25192), .Z(n25179) );
  AND U26069 ( .A(n25193), .B(n25194), .Z(n25191) );
  XOR U26070 ( .A(n25192), .B(n25018), .Z(n25194) );
  XOR U26071 ( .A(n25185), .B(n25186), .Z(n25018) );
  XNOR U26072 ( .A(n25195), .B(n25196), .Z(n25186) );
  ANDN U26073 ( .B(n25197), .A(n25198), .Z(n25195) );
  XOR U26074 ( .A(n25199), .B(n25200), .Z(n25197) );
  XOR U26075 ( .A(n25201), .B(n25202), .Z(n25185) );
  XNOR U26076 ( .A(n25203), .B(n25204), .Z(n25202) );
  ANDN U26077 ( .B(n25205), .A(n25206), .Z(n25203) );
  XNOR U26078 ( .A(n25207), .B(n25208), .Z(n25205) );
  IV U26079 ( .A(n25183), .Z(n25201) );
  XOR U26080 ( .A(n25209), .B(n25210), .Z(n25183) );
  ANDN U26081 ( .B(n25211), .A(n25212), .Z(n25209) );
  XOR U26082 ( .A(n25210), .B(n25213), .Z(n25211) );
  XNOR U26083 ( .A(n25192), .B(n25020), .Z(n25193) );
  XOR U26084 ( .A(n25214), .B(n25215), .Z(n25020) );
  AND U26085 ( .A(n276), .B(n25216), .Z(n25214) );
  XOR U26086 ( .A(n25217), .B(n25215), .Z(n25216) );
  XNOR U26087 ( .A(n25218), .B(n25219), .Z(n25192) );
  AND U26088 ( .A(n25220), .B(n25221), .Z(n25218) );
  XNOR U26089 ( .A(n25219), .B(n25070), .Z(n25221) );
  XOR U26090 ( .A(n25212), .B(n25213), .Z(n25070) );
  XOR U26091 ( .A(n25222), .B(n25200), .Z(n25213) );
  XNOR U26092 ( .A(n25223), .B(n25224), .Z(n25200) );
  ANDN U26093 ( .B(n25225), .A(n25226), .Z(n25223) );
  XOR U26094 ( .A(n25227), .B(n25228), .Z(n25225) );
  IV U26095 ( .A(n25198), .Z(n25222) );
  XOR U26096 ( .A(n25196), .B(n25229), .Z(n25198) );
  XNOR U26097 ( .A(n25230), .B(n25231), .Z(n25229) );
  ANDN U26098 ( .B(n25232), .A(n25233), .Z(n25230) );
  XNOR U26099 ( .A(n25234), .B(n25235), .Z(n25232) );
  IV U26100 ( .A(n25199), .Z(n25196) );
  XOR U26101 ( .A(n25236), .B(n25237), .Z(n25199) );
  ANDN U26102 ( .B(n25238), .A(n25239), .Z(n25236) );
  XOR U26103 ( .A(n25237), .B(n25240), .Z(n25238) );
  XOR U26104 ( .A(n25241), .B(n25242), .Z(n25212) );
  XNOR U26105 ( .A(n25207), .B(n25243), .Z(n25242) );
  IV U26106 ( .A(n25210), .Z(n25243) );
  XOR U26107 ( .A(n25244), .B(n25245), .Z(n25210) );
  ANDN U26108 ( .B(n25246), .A(n25247), .Z(n25244) );
  XOR U26109 ( .A(n25245), .B(n25248), .Z(n25246) );
  XNOR U26110 ( .A(n25249), .B(n25250), .Z(n25207) );
  ANDN U26111 ( .B(n25251), .A(n25252), .Z(n25249) );
  XOR U26112 ( .A(n25250), .B(n25253), .Z(n25251) );
  IV U26113 ( .A(n25206), .Z(n25241) );
  XOR U26114 ( .A(n25204), .B(n25254), .Z(n25206) );
  XNOR U26115 ( .A(n25255), .B(n25256), .Z(n25254) );
  ANDN U26116 ( .B(n25257), .A(n25258), .Z(n25255) );
  XNOR U26117 ( .A(n25259), .B(n25260), .Z(n25257) );
  IV U26118 ( .A(n25208), .Z(n25204) );
  XOR U26119 ( .A(n25261), .B(n25262), .Z(n25208) );
  ANDN U26120 ( .B(n25263), .A(n25264), .Z(n25261) );
  XOR U26121 ( .A(n25265), .B(n25262), .Z(n25263) );
  XOR U26122 ( .A(n25219), .B(n25072), .Z(n25220) );
  XOR U26123 ( .A(n25266), .B(n25267), .Z(n25072) );
  AND U26124 ( .A(n276), .B(n25268), .Z(n25266) );
  XOR U26125 ( .A(n25269), .B(n25267), .Z(n25268) );
  XNOR U26126 ( .A(n25270), .B(n25271), .Z(n25219) );
  NAND U26127 ( .A(n25272), .B(n25273), .Z(n25271) );
  XOR U26128 ( .A(n25274), .B(n25171), .Z(n25273) );
  XOR U26129 ( .A(n25247), .B(n25248), .Z(n25171) );
  XOR U26130 ( .A(n25275), .B(n25240), .Z(n25248) );
  XOR U26131 ( .A(n25276), .B(n25228), .Z(n25240) );
  XOR U26132 ( .A(n25277), .B(n25278), .Z(n25228) );
  ANDN U26133 ( .B(n25279), .A(n25280), .Z(n25277) );
  XOR U26134 ( .A(n25278), .B(n25281), .Z(n25279) );
  IV U26135 ( .A(n25226), .Z(n25276) );
  XOR U26136 ( .A(n25224), .B(n25282), .Z(n25226) );
  XOR U26137 ( .A(n25283), .B(n25284), .Z(n25282) );
  ANDN U26138 ( .B(n25285), .A(n25286), .Z(n25283) );
  XOR U26139 ( .A(n25287), .B(n25284), .Z(n25285) );
  IV U26140 ( .A(n25227), .Z(n25224) );
  XOR U26141 ( .A(n25288), .B(n25289), .Z(n25227) );
  ANDN U26142 ( .B(n25290), .A(n25291), .Z(n25288) );
  XOR U26143 ( .A(n25289), .B(n25292), .Z(n25290) );
  IV U26144 ( .A(n25239), .Z(n25275) );
  XOR U26145 ( .A(n25293), .B(n25294), .Z(n25239) );
  XNOR U26146 ( .A(n25234), .B(n25295), .Z(n25294) );
  IV U26147 ( .A(n25237), .Z(n25295) );
  XOR U26148 ( .A(n25296), .B(n25297), .Z(n25237) );
  ANDN U26149 ( .B(n25298), .A(n25299), .Z(n25296) );
  XOR U26150 ( .A(n25297), .B(n25300), .Z(n25298) );
  XNOR U26151 ( .A(n25301), .B(n25302), .Z(n25234) );
  ANDN U26152 ( .B(n25303), .A(n25304), .Z(n25301) );
  XOR U26153 ( .A(n25302), .B(n25305), .Z(n25303) );
  IV U26154 ( .A(n25233), .Z(n25293) );
  XOR U26155 ( .A(n25231), .B(n25306), .Z(n25233) );
  XOR U26156 ( .A(n25307), .B(n25308), .Z(n25306) );
  ANDN U26157 ( .B(n25309), .A(n25310), .Z(n25307) );
  XOR U26158 ( .A(n25311), .B(n25308), .Z(n25309) );
  IV U26159 ( .A(n25235), .Z(n25231) );
  XOR U26160 ( .A(n25312), .B(n25313), .Z(n25235) );
  ANDN U26161 ( .B(n25314), .A(n25315), .Z(n25312) );
  XOR U26162 ( .A(n25316), .B(n25313), .Z(n25314) );
  XOR U26163 ( .A(n25317), .B(n25318), .Z(n25247) );
  XOR U26164 ( .A(n25265), .B(n25319), .Z(n25318) );
  IV U26165 ( .A(n25245), .Z(n25319) );
  XOR U26166 ( .A(n25320), .B(n25321), .Z(n25245) );
  ANDN U26167 ( .B(n25322), .A(n25323), .Z(n25320) );
  XOR U26168 ( .A(n25321), .B(n25324), .Z(n25322) );
  XOR U26169 ( .A(n25325), .B(n25253), .Z(n25265) );
  XOR U26170 ( .A(n25326), .B(n25327), .Z(n25253) );
  ANDN U26171 ( .B(n25328), .A(n25329), .Z(n25326) );
  XOR U26172 ( .A(n25327), .B(n25330), .Z(n25328) );
  IV U26173 ( .A(n25252), .Z(n25325) );
  XOR U26174 ( .A(n25331), .B(n25332), .Z(n25252) );
  XOR U26175 ( .A(n25333), .B(n25334), .Z(n25332) );
  ANDN U26176 ( .B(n25335), .A(n25336), .Z(n25333) );
  XOR U26177 ( .A(n25337), .B(n25334), .Z(n25335) );
  IV U26178 ( .A(n25250), .Z(n25331) );
  XOR U26179 ( .A(n25338), .B(n25339), .Z(n25250) );
  ANDN U26180 ( .B(n25340), .A(n25341), .Z(n25338) );
  XOR U26181 ( .A(n25339), .B(n25342), .Z(n25340) );
  IV U26182 ( .A(n25264), .Z(n25317) );
  XOR U26183 ( .A(n25343), .B(n25344), .Z(n25264) );
  XNOR U26184 ( .A(n25259), .B(n25345), .Z(n25344) );
  IV U26185 ( .A(n25262), .Z(n25345) );
  XOR U26186 ( .A(n25346), .B(n25347), .Z(n25262) );
  ANDN U26187 ( .B(n25348), .A(n25349), .Z(n25346) );
  XOR U26188 ( .A(n25350), .B(n25347), .Z(n25348) );
  XNOR U26189 ( .A(n25351), .B(n25352), .Z(n25259) );
  ANDN U26190 ( .B(n25353), .A(n25354), .Z(n25351) );
  XOR U26191 ( .A(n25352), .B(n25355), .Z(n25353) );
  IV U26192 ( .A(n25258), .Z(n25343) );
  XOR U26193 ( .A(n25256), .B(n25356), .Z(n25258) );
  XOR U26194 ( .A(n25357), .B(n25358), .Z(n25356) );
  ANDN U26195 ( .B(n25359), .A(n25360), .Z(n25357) );
  XOR U26196 ( .A(n25361), .B(n25358), .Z(n25359) );
  IV U26197 ( .A(n25260), .Z(n25256) );
  XOR U26198 ( .A(n25362), .B(n25363), .Z(n25260) );
  ANDN U26199 ( .B(n25364), .A(n25365), .Z(n25362) );
  XOR U26200 ( .A(n25366), .B(n25363), .Z(n25364) );
  IV U26201 ( .A(n25270), .Z(n25274) );
  XOR U26202 ( .A(n25270), .B(n25173), .Z(n25272) );
  XOR U26203 ( .A(n25367), .B(n25368), .Z(n25173) );
  AND U26204 ( .A(n276), .B(n25369), .Z(n25367) );
  XOR U26205 ( .A(n25370), .B(n25368), .Z(n25369) );
  NANDN U26206 ( .A(n25175), .B(n25177), .Z(n25270) );
  XOR U26207 ( .A(n25371), .B(n25372), .Z(n25177) );
  AND U26208 ( .A(n276), .B(n25373), .Z(n25371) );
  XOR U26209 ( .A(n25372), .B(n25374), .Z(n25373) );
  XNOR U26210 ( .A(n25375), .B(n25376), .Z(n276) );
  AND U26211 ( .A(n25377), .B(n25378), .Z(n25375) );
  XOR U26212 ( .A(n25376), .B(n25188), .Z(n25378) );
  XNOR U26213 ( .A(n25379), .B(n25380), .Z(n25188) );
  ANDN U26214 ( .B(n25381), .A(n25382), .Z(n25379) );
  XOR U26215 ( .A(n25380), .B(n25383), .Z(n25381) );
  XNOR U26216 ( .A(n25376), .B(n25190), .Z(n25377) );
  XOR U26217 ( .A(n25384), .B(n25385), .Z(n25190) );
  AND U26218 ( .A(n280), .B(n25386), .Z(n25384) );
  XOR U26219 ( .A(n25387), .B(n25385), .Z(n25386) );
  XOR U26220 ( .A(n25388), .B(n25389), .Z(n25376) );
  AND U26221 ( .A(n25390), .B(n25391), .Z(n25388) );
  XOR U26222 ( .A(n25389), .B(n25215), .Z(n25391) );
  XOR U26223 ( .A(n25382), .B(n25383), .Z(n25215) );
  XNOR U26224 ( .A(n25392), .B(n25393), .Z(n25383) );
  ANDN U26225 ( .B(n25394), .A(n25395), .Z(n25392) );
  XOR U26226 ( .A(n25396), .B(n25397), .Z(n25394) );
  XOR U26227 ( .A(n25398), .B(n25399), .Z(n25382) );
  XNOR U26228 ( .A(n25400), .B(n25401), .Z(n25399) );
  ANDN U26229 ( .B(n25402), .A(n25403), .Z(n25400) );
  XNOR U26230 ( .A(n25404), .B(n25405), .Z(n25402) );
  IV U26231 ( .A(n25380), .Z(n25398) );
  XOR U26232 ( .A(n25406), .B(n25407), .Z(n25380) );
  ANDN U26233 ( .B(n25408), .A(n25409), .Z(n25406) );
  XOR U26234 ( .A(n25407), .B(n25410), .Z(n25408) );
  XNOR U26235 ( .A(n25389), .B(n25217), .Z(n25390) );
  XOR U26236 ( .A(n25411), .B(n25412), .Z(n25217) );
  AND U26237 ( .A(n280), .B(n25413), .Z(n25411) );
  XOR U26238 ( .A(n25414), .B(n25412), .Z(n25413) );
  XNOR U26239 ( .A(n25415), .B(n25416), .Z(n25389) );
  AND U26240 ( .A(n25417), .B(n25418), .Z(n25415) );
  XNOR U26241 ( .A(n25416), .B(n25267), .Z(n25418) );
  XOR U26242 ( .A(n25409), .B(n25410), .Z(n25267) );
  XOR U26243 ( .A(n25419), .B(n25397), .Z(n25410) );
  XNOR U26244 ( .A(n25420), .B(n25421), .Z(n25397) );
  ANDN U26245 ( .B(n25422), .A(n25423), .Z(n25420) );
  XOR U26246 ( .A(n25424), .B(n25425), .Z(n25422) );
  IV U26247 ( .A(n25395), .Z(n25419) );
  XOR U26248 ( .A(n25393), .B(n25426), .Z(n25395) );
  XNOR U26249 ( .A(n25427), .B(n25428), .Z(n25426) );
  ANDN U26250 ( .B(n25429), .A(n25430), .Z(n25427) );
  XNOR U26251 ( .A(n25431), .B(n25432), .Z(n25429) );
  IV U26252 ( .A(n25396), .Z(n25393) );
  XOR U26253 ( .A(n25433), .B(n25434), .Z(n25396) );
  ANDN U26254 ( .B(n25435), .A(n25436), .Z(n25433) );
  XOR U26255 ( .A(n25434), .B(n25437), .Z(n25435) );
  XOR U26256 ( .A(n25438), .B(n25439), .Z(n25409) );
  XNOR U26257 ( .A(n25404), .B(n25440), .Z(n25439) );
  IV U26258 ( .A(n25407), .Z(n25440) );
  XOR U26259 ( .A(n25441), .B(n25442), .Z(n25407) );
  ANDN U26260 ( .B(n25443), .A(n25444), .Z(n25441) );
  XOR U26261 ( .A(n25442), .B(n25445), .Z(n25443) );
  XNOR U26262 ( .A(n25446), .B(n25447), .Z(n25404) );
  ANDN U26263 ( .B(n25448), .A(n25449), .Z(n25446) );
  XOR U26264 ( .A(n25447), .B(n25450), .Z(n25448) );
  IV U26265 ( .A(n25403), .Z(n25438) );
  XOR U26266 ( .A(n25401), .B(n25451), .Z(n25403) );
  XNOR U26267 ( .A(n25452), .B(n25453), .Z(n25451) );
  ANDN U26268 ( .B(n25454), .A(n25455), .Z(n25452) );
  XNOR U26269 ( .A(n25456), .B(n25457), .Z(n25454) );
  IV U26270 ( .A(n25405), .Z(n25401) );
  XOR U26271 ( .A(n25458), .B(n25459), .Z(n25405) );
  ANDN U26272 ( .B(n25460), .A(n25461), .Z(n25458) );
  XOR U26273 ( .A(n25462), .B(n25459), .Z(n25460) );
  XOR U26274 ( .A(n25416), .B(n25269), .Z(n25417) );
  XOR U26275 ( .A(n25463), .B(n25464), .Z(n25269) );
  AND U26276 ( .A(n280), .B(n25465), .Z(n25463) );
  XOR U26277 ( .A(n25466), .B(n25464), .Z(n25465) );
  XNOR U26278 ( .A(n25467), .B(n25468), .Z(n25416) );
  NAND U26279 ( .A(n25469), .B(n25470), .Z(n25468) );
  XOR U26280 ( .A(n25471), .B(n25368), .Z(n25470) );
  XOR U26281 ( .A(n25444), .B(n25445), .Z(n25368) );
  XOR U26282 ( .A(n25472), .B(n25437), .Z(n25445) );
  XOR U26283 ( .A(n25473), .B(n25425), .Z(n25437) );
  XOR U26284 ( .A(n25474), .B(n25475), .Z(n25425) );
  ANDN U26285 ( .B(n25476), .A(n25477), .Z(n25474) );
  XOR U26286 ( .A(n25475), .B(n25478), .Z(n25476) );
  IV U26287 ( .A(n25423), .Z(n25473) );
  XOR U26288 ( .A(n25421), .B(n25479), .Z(n25423) );
  XOR U26289 ( .A(n25480), .B(n25481), .Z(n25479) );
  ANDN U26290 ( .B(n25482), .A(n25483), .Z(n25480) );
  XOR U26291 ( .A(n25484), .B(n25481), .Z(n25482) );
  IV U26292 ( .A(n25424), .Z(n25421) );
  XOR U26293 ( .A(n25485), .B(n25486), .Z(n25424) );
  ANDN U26294 ( .B(n25487), .A(n25488), .Z(n25485) );
  XOR U26295 ( .A(n25486), .B(n25489), .Z(n25487) );
  IV U26296 ( .A(n25436), .Z(n25472) );
  XOR U26297 ( .A(n25490), .B(n25491), .Z(n25436) );
  XNOR U26298 ( .A(n25431), .B(n25492), .Z(n25491) );
  IV U26299 ( .A(n25434), .Z(n25492) );
  XOR U26300 ( .A(n25493), .B(n25494), .Z(n25434) );
  ANDN U26301 ( .B(n25495), .A(n25496), .Z(n25493) );
  XOR U26302 ( .A(n25494), .B(n25497), .Z(n25495) );
  XNOR U26303 ( .A(n25498), .B(n25499), .Z(n25431) );
  ANDN U26304 ( .B(n25500), .A(n25501), .Z(n25498) );
  XOR U26305 ( .A(n25499), .B(n25502), .Z(n25500) );
  IV U26306 ( .A(n25430), .Z(n25490) );
  XOR U26307 ( .A(n25428), .B(n25503), .Z(n25430) );
  XOR U26308 ( .A(n25504), .B(n25505), .Z(n25503) );
  ANDN U26309 ( .B(n25506), .A(n25507), .Z(n25504) );
  XOR U26310 ( .A(n25508), .B(n25505), .Z(n25506) );
  IV U26311 ( .A(n25432), .Z(n25428) );
  XOR U26312 ( .A(n25509), .B(n25510), .Z(n25432) );
  ANDN U26313 ( .B(n25511), .A(n25512), .Z(n25509) );
  XOR U26314 ( .A(n25513), .B(n25510), .Z(n25511) );
  XOR U26315 ( .A(n25514), .B(n25515), .Z(n25444) );
  XOR U26316 ( .A(n25462), .B(n25516), .Z(n25515) );
  IV U26317 ( .A(n25442), .Z(n25516) );
  XOR U26318 ( .A(n25517), .B(n25518), .Z(n25442) );
  ANDN U26319 ( .B(n25519), .A(n25520), .Z(n25517) );
  XOR U26320 ( .A(n25518), .B(n25521), .Z(n25519) );
  XOR U26321 ( .A(n25522), .B(n25450), .Z(n25462) );
  XOR U26322 ( .A(n25523), .B(n25524), .Z(n25450) );
  ANDN U26323 ( .B(n25525), .A(n25526), .Z(n25523) );
  XOR U26324 ( .A(n25524), .B(n25527), .Z(n25525) );
  IV U26325 ( .A(n25449), .Z(n25522) );
  XOR U26326 ( .A(n25528), .B(n25529), .Z(n25449) );
  XOR U26327 ( .A(n25530), .B(n25531), .Z(n25529) );
  ANDN U26328 ( .B(n25532), .A(n25533), .Z(n25530) );
  XOR U26329 ( .A(n25534), .B(n25531), .Z(n25532) );
  IV U26330 ( .A(n25447), .Z(n25528) );
  XOR U26331 ( .A(n25535), .B(n25536), .Z(n25447) );
  ANDN U26332 ( .B(n25537), .A(n25538), .Z(n25535) );
  XOR U26333 ( .A(n25536), .B(n25539), .Z(n25537) );
  IV U26334 ( .A(n25461), .Z(n25514) );
  XOR U26335 ( .A(n25540), .B(n25541), .Z(n25461) );
  XNOR U26336 ( .A(n25456), .B(n25542), .Z(n25541) );
  IV U26337 ( .A(n25459), .Z(n25542) );
  XOR U26338 ( .A(n25543), .B(n25544), .Z(n25459) );
  ANDN U26339 ( .B(n25545), .A(n25546), .Z(n25543) );
  XOR U26340 ( .A(n25547), .B(n25544), .Z(n25545) );
  XNOR U26341 ( .A(n25548), .B(n25549), .Z(n25456) );
  ANDN U26342 ( .B(n25550), .A(n25551), .Z(n25548) );
  XOR U26343 ( .A(n25549), .B(n25552), .Z(n25550) );
  IV U26344 ( .A(n25455), .Z(n25540) );
  XOR U26345 ( .A(n25453), .B(n25553), .Z(n25455) );
  XOR U26346 ( .A(n25554), .B(n25555), .Z(n25553) );
  ANDN U26347 ( .B(n25556), .A(n25557), .Z(n25554) );
  XOR U26348 ( .A(n25558), .B(n25555), .Z(n25556) );
  IV U26349 ( .A(n25457), .Z(n25453) );
  XOR U26350 ( .A(n25559), .B(n25560), .Z(n25457) );
  ANDN U26351 ( .B(n25561), .A(n25562), .Z(n25559) );
  XOR U26352 ( .A(n25563), .B(n25560), .Z(n25561) );
  IV U26353 ( .A(n25467), .Z(n25471) );
  XOR U26354 ( .A(n25467), .B(n25370), .Z(n25469) );
  XOR U26355 ( .A(n25564), .B(n25565), .Z(n25370) );
  AND U26356 ( .A(n280), .B(n25566), .Z(n25564) );
  XOR U26357 ( .A(n25567), .B(n25565), .Z(n25566) );
  NANDN U26358 ( .A(n25372), .B(n25374), .Z(n25467) );
  XOR U26359 ( .A(n25568), .B(n25569), .Z(n25374) );
  AND U26360 ( .A(n280), .B(n25570), .Z(n25568) );
  XOR U26361 ( .A(n25569), .B(n25571), .Z(n25570) );
  XNOR U26362 ( .A(n25572), .B(n25573), .Z(n280) );
  AND U26363 ( .A(n25574), .B(n25575), .Z(n25572) );
  XOR U26364 ( .A(n25573), .B(n25385), .Z(n25575) );
  XNOR U26365 ( .A(n25576), .B(n25577), .Z(n25385) );
  ANDN U26366 ( .B(n25578), .A(n25579), .Z(n25576) );
  XOR U26367 ( .A(n25577), .B(n25580), .Z(n25578) );
  XNOR U26368 ( .A(n25573), .B(n25387), .Z(n25574) );
  XOR U26369 ( .A(n25581), .B(n25582), .Z(n25387) );
  AND U26370 ( .A(n284), .B(n25583), .Z(n25581) );
  XOR U26371 ( .A(n25584), .B(n25582), .Z(n25583) );
  XOR U26372 ( .A(n25585), .B(n25586), .Z(n25573) );
  AND U26373 ( .A(n25587), .B(n25588), .Z(n25585) );
  XOR U26374 ( .A(n25586), .B(n25412), .Z(n25588) );
  XOR U26375 ( .A(n25579), .B(n25580), .Z(n25412) );
  XNOR U26376 ( .A(n25589), .B(n25590), .Z(n25580) );
  ANDN U26377 ( .B(n25591), .A(n25592), .Z(n25589) );
  XOR U26378 ( .A(n25593), .B(n25594), .Z(n25591) );
  XOR U26379 ( .A(n25595), .B(n25596), .Z(n25579) );
  XNOR U26380 ( .A(n25597), .B(n25598), .Z(n25596) );
  ANDN U26381 ( .B(n25599), .A(n25600), .Z(n25597) );
  XNOR U26382 ( .A(n25601), .B(n25602), .Z(n25599) );
  IV U26383 ( .A(n25577), .Z(n25595) );
  XOR U26384 ( .A(n25603), .B(n25604), .Z(n25577) );
  ANDN U26385 ( .B(n25605), .A(n25606), .Z(n25603) );
  XOR U26386 ( .A(n25604), .B(n25607), .Z(n25605) );
  XNOR U26387 ( .A(n25586), .B(n25414), .Z(n25587) );
  XOR U26388 ( .A(n25608), .B(n25609), .Z(n25414) );
  AND U26389 ( .A(n284), .B(n25610), .Z(n25608) );
  XOR U26390 ( .A(n25611), .B(n25609), .Z(n25610) );
  XNOR U26391 ( .A(n25612), .B(n25613), .Z(n25586) );
  AND U26392 ( .A(n25614), .B(n25615), .Z(n25612) );
  XNOR U26393 ( .A(n25613), .B(n25464), .Z(n25615) );
  XOR U26394 ( .A(n25606), .B(n25607), .Z(n25464) );
  XOR U26395 ( .A(n25616), .B(n25594), .Z(n25607) );
  XNOR U26396 ( .A(n25617), .B(n25618), .Z(n25594) );
  ANDN U26397 ( .B(n25619), .A(n25620), .Z(n25617) );
  XOR U26398 ( .A(n25621), .B(n25622), .Z(n25619) );
  IV U26399 ( .A(n25592), .Z(n25616) );
  XOR U26400 ( .A(n25590), .B(n25623), .Z(n25592) );
  XNOR U26401 ( .A(n25624), .B(n25625), .Z(n25623) );
  ANDN U26402 ( .B(n25626), .A(n25627), .Z(n25624) );
  XNOR U26403 ( .A(n25628), .B(n25629), .Z(n25626) );
  IV U26404 ( .A(n25593), .Z(n25590) );
  XOR U26405 ( .A(n25630), .B(n25631), .Z(n25593) );
  ANDN U26406 ( .B(n25632), .A(n25633), .Z(n25630) );
  XOR U26407 ( .A(n25631), .B(n25634), .Z(n25632) );
  XOR U26408 ( .A(n25635), .B(n25636), .Z(n25606) );
  XNOR U26409 ( .A(n25601), .B(n25637), .Z(n25636) );
  IV U26410 ( .A(n25604), .Z(n25637) );
  XOR U26411 ( .A(n25638), .B(n25639), .Z(n25604) );
  ANDN U26412 ( .B(n25640), .A(n25641), .Z(n25638) );
  XOR U26413 ( .A(n25639), .B(n25642), .Z(n25640) );
  XNOR U26414 ( .A(n25643), .B(n25644), .Z(n25601) );
  ANDN U26415 ( .B(n25645), .A(n25646), .Z(n25643) );
  XOR U26416 ( .A(n25644), .B(n25647), .Z(n25645) );
  IV U26417 ( .A(n25600), .Z(n25635) );
  XOR U26418 ( .A(n25598), .B(n25648), .Z(n25600) );
  XNOR U26419 ( .A(n25649), .B(n25650), .Z(n25648) );
  ANDN U26420 ( .B(n25651), .A(n25652), .Z(n25649) );
  XNOR U26421 ( .A(n25653), .B(n25654), .Z(n25651) );
  IV U26422 ( .A(n25602), .Z(n25598) );
  XOR U26423 ( .A(n25655), .B(n25656), .Z(n25602) );
  ANDN U26424 ( .B(n25657), .A(n25658), .Z(n25655) );
  XOR U26425 ( .A(n25659), .B(n25656), .Z(n25657) );
  XOR U26426 ( .A(n25613), .B(n25466), .Z(n25614) );
  XOR U26427 ( .A(n25660), .B(n25661), .Z(n25466) );
  AND U26428 ( .A(n284), .B(n25662), .Z(n25660) );
  XOR U26429 ( .A(n25663), .B(n25661), .Z(n25662) );
  XNOR U26430 ( .A(n25664), .B(n25665), .Z(n25613) );
  NAND U26431 ( .A(n25666), .B(n25667), .Z(n25665) );
  XOR U26432 ( .A(n25668), .B(n25565), .Z(n25667) );
  XOR U26433 ( .A(n25641), .B(n25642), .Z(n25565) );
  XOR U26434 ( .A(n25669), .B(n25634), .Z(n25642) );
  XOR U26435 ( .A(n25670), .B(n25622), .Z(n25634) );
  XOR U26436 ( .A(n25671), .B(n25672), .Z(n25622) );
  ANDN U26437 ( .B(n25673), .A(n25674), .Z(n25671) );
  XOR U26438 ( .A(n25672), .B(n25675), .Z(n25673) );
  IV U26439 ( .A(n25620), .Z(n25670) );
  XOR U26440 ( .A(n25618), .B(n25676), .Z(n25620) );
  XOR U26441 ( .A(n25677), .B(n25678), .Z(n25676) );
  ANDN U26442 ( .B(n25679), .A(n25680), .Z(n25677) );
  XOR U26443 ( .A(n25681), .B(n25678), .Z(n25679) );
  IV U26444 ( .A(n25621), .Z(n25618) );
  XOR U26445 ( .A(n25682), .B(n25683), .Z(n25621) );
  ANDN U26446 ( .B(n25684), .A(n25685), .Z(n25682) );
  XOR U26447 ( .A(n25683), .B(n25686), .Z(n25684) );
  IV U26448 ( .A(n25633), .Z(n25669) );
  XOR U26449 ( .A(n25687), .B(n25688), .Z(n25633) );
  XNOR U26450 ( .A(n25628), .B(n25689), .Z(n25688) );
  IV U26451 ( .A(n25631), .Z(n25689) );
  XOR U26452 ( .A(n25690), .B(n25691), .Z(n25631) );
  ANDN U26453 ( .B(n25692), .A(n25693), .Z(n25690) );
  XOR U26454 ( .A(n25691), .B(n25694), .Z(n25692) );
  XNOR U26455 ( .A(n25695), .B(n25696), .Z(n25628) );
  ANDN U26456 ( .B(n25697), .A(n25698), .Z(n25695) );
  XOR U26457 ( .A(n25696), .B(n25699), .Z(n25697) );
  IV U26458 ( .A(n25627), .Z(n25687) );
  XOR U26459 ( .A(n25625), .B(n25700), .Z(n25627) );
  XOR U26460 ( .A(n25701), .B(n25702), .Z(n25700) );
  ANDN U26461 ( .B(n25703), .A(n25704), .Z(n25701) );
  XOR U26462 ( .A(n25705), .B(n25702), .Z(n25703) );
  IV U26463 ( .A(n25629), .Z(n25625) );
  XOR U26464 ( .A(n25706), .B(n25707), .Z(n25629) );
  ANDN U26465 ( .B(n25708), .A(n25709), .Z(n25706) );
  XOR U26466 ( .A(n25710), .B(n25707), .Z(n25708) );
  XOR U26467 ( .A(n25711), .B(n25712), .Z(n25641) );
  XOR U26468 ( .A(n25659), .B(n25713), .Z(n25712) );
  IV U26469 ( .A(n25639), .Z(n25713) );
  XOR U26470 ( .A(n25714), .B(n25715), .Z(n25639) );
  ANDN U26471 ( .B(n25716), .A(n25717), .Z(n25714) );
  XOR U26472 ( .A(n25715), .B(n25718), .Z(n25716) );
  XOR U26473 ( .A(n25719), .B(n25647), .Z(n25659) );
  XOR U26474 ( .A(n25720), .B(n25721), .Z(n25647) );
  ANDN U26475 ( .B(n25722), .A(n25723), .Z(n25720) );
  XOR U26476 ( .A(n25721), .B(n25724), .Z(n25722) );
  IV U26477 ( .A(n25646), .Z(n25719) );
  XOR U26478 ( .A(n25725), .B(n25726), .Z(n25646) );
  XOR U26479 ( .A(n25727), .B(n25728), .Z(n25726) );
  ANDN U26480 ( .B(n25729), .A(n25730), .Z(n25727) );
  XOR U26481 ( .A(n25731), .B(n25728), .Z(n25729) );
  IV U26482 ( .A(n25644), .Z(n25725) );
  XOR U26483 ( .A(n25732), .B(n25733), .Z(n25644) );
  ANDN U26484 ( .B(n25734), .A(n25735), .Z(n25732) );
  XOR U26485 ( .A(n25733), .B(n25736), .Z(n25734) );
  IV U26486 ( .A(n25658), .Z(n25711) );
  XOR U26487 ( .A(n25737), .B(n25738), .Z(n25658) );
  XNOR U26488 ( .A(n25653), .B(n25739), .Z(n25738) );
  IV U26489 ( .A(n25656), .Z(n25739) );
  XOR U26490 ( .A(n25740), .B(n25741), .Z(n25656) );
  ANDN U26491 ( .B(n25742), .A(n25743), .Z(n25740) );
  XOR U26492 ( .A(n25744), .B(n25741), .Z(n25742) );
  XNOR U26493 ( .A(n25745), .B(n25746), .Z(n25653) );
  ANDN U26494 ( .B(n25747), .A(n25748), .Z(n25745) );
  XOR U26495 ( .A(n25746), .B(n25749), .Z(n25747) );
  IV U26496 ( .A(n25652), .Z(n25737) );
  XOR U26497 ( .A(n25650), .B(n25750), .Z(n25652) );
  XOR U26498 ( .A(n25751), .B(n25752), .Z(n25750) );
  ANDN U26499 ( .B(n25753), .A(n25754), .Z(n25751) );
  XOR U26500 ( .A(n25755), .B(n25752), .Z(n25753) );
  IV U26501 ( .A(n25654), .Z(n25650) );
  XOR U26502 ( .A(n25756), .B(n25757), .Z(n25654) );
  ANDN U26503 ( .B(n25758), .A(n25759), .Z(n25756) );
  XOR U26504 ( .A(n25760), .B(n25757), .Z(n25758) );
  IV U26505 ( .A(n25664), .Z(n25668) );
  XOR U26506 ( .A(n25664), .B(n25567), .Z(n25666) );
  XOR U26507 ( .A(n25761), .B(n25762), .Z(n25567) );
  AND U26508 ( .A(n284), .B(n25763), .Z(n25761) );
  XOR U26509 ( .A(n25764), .B(n25762), .Z(n25763) );
  NANDN U26510 ( .A(n25569), .B(n25571), .Z(n25664) );
  XOR U26511 ( .A(n25765), .B(n25766), .Z(n25571) );
  AND U26512 ( .A(n284), .B(n25767), .Z(n25765) );
  XOR U26513 ( .A(n25766), .B(n25768), .Z(n25767) );
  XNOR U26514 ( .A(n25769), .B(n25770), .Z(n284) );
  AND U26515 ( .A(n25771), .B(n25772), .Z(n25769) );
  XOR U26516 ( .A(n25770), .B(n25582), .Z(n25772) );
  XNOR U26517 ( .A(n25773), .B(n25774), .Z(n25582) );
  ANDN U26518 ( .B(n25775), .A(n25776), .Z(n25773) );
  XOR U26519 ( .A(n25774), .B(n25777), .Z(n25775) );
  XNOR U26520 ( .A(n25770), .B(n25584), .Z(n25771) );
  XOR U26521 ( .A(n25778), .B(n25779), .Z(n25584) );
  AND U26522 ( .A(n288), .B(n25780), .Z(n25778) );
  XOR U26523 ( .A(n25781), .B(n25779), .Z(n25780) );
  XOR U26524 ( .A(n25782), .B(n25783), .Z(n25770) );
  AND U26525 ( .A(n25784), .B(n25785), .Z(n25782) );
  XOR U26526 ( .A(n25783), .B(n25609), .Z(n25785) );
  XOR U26527 ( .A(n25776), .B(n25777), .Z(n25609) );
  XNOR U26528 ( .A(n25786), .B(n25787), .Z(n25777) );
  ANDN U26529 ( .B(n25788), .A(n25789), .Z(n25786) );
  XOR U26530 ( .A(n25790), .B(n25791), .Z(n25788) );
  XOR U26531 ( .A(n25792), .B(n25793), .Z(n25776) );
  XNOR U26532 ( .A(n25794), .B(n25795), .Z(n25793) );
  ANDN U26533 ( .B(n25796), .A(n25797), .Z(n25794) );
  XNOR U26534 ( .A(n25798), .B(n25799), .Z(n25796) );
  IV U26535 ( .A(n25774), .Z(n25792) );
  XOR U26536 ( .A(n25800), .B(n25801), .Z(n25774) );
  ANDN U26537 ( .B(n25802), .A(n25803), .Z(n25800) );
  XOR U26538 ( .A(n25801), .B(n25804), .Z(n25802) );
  XNOR U26539 ( .A(n25783), .B(n25611), .Z(n25784) );
  XOR U26540 ( .A(n25805), .B(n25806), .Z(n25611) );
  AND U26541 ( .A(n288), .B(n25807), .Z(n25805) );
  XOR U26542 ( .A(n25808), .B(n25806), .Z(n25807) );
  XNOR U26543 ( .A(n25809), .B(n25810), .Z(n25783) );
  AND U26544 ( .A(n25811), .B(n25812), .Z(n25809) );
  XNOR U26545 ( .A(n25810), .B(n25661), .Z(n25812) );
  XOR U26546 ( .A(n25803), .B(n25804), .Z(n25661) );
  XOR U26547 ( .A(n25813), .B(n25791), .Z(n25804) );
  XNOR U26548 ( .A(n25814), .B(n25815), .Z(n25791) );
  ANDN U26549 ( .B(n25816), .A(n25817), .Z(n25814) );
  XOR U26550 ( .A(n25818), .B(n25819), .Z(n25816) );
  IV U26551 ( .A(n25789), .Z(n25813) );
  XOR U26552 ( .A(n25787), .B(n25820), .Z(n25789) );
  XNOR U26553 ( .A(n25821), .B(n25822), .Z(n25820) );
  ANDN U26554 ( .B(n25823), .A(n25824), .Z(n25821) );
  XNOR U26555 ( .A(n25825), .B(n25826), .Z(n25823) );
  IV U26556 ( .A(n25790), .Z(n25787) );
  XOR U26557 ( .A(n25827), .B(n25828), .Z(n25790) );
  ANDN U26558 ( .B(n25829), .A(n25830), .Z(n25827) );
  XOR U26559 ( .A(n25828), .B(n25831), .Z(n25829) );
  XOR U26560 ( .A(n25832), .B(n25833), .Z(n25803) );
  XNOR U26561 ( .A(n25798), .B(n25834), .Z(n25833) );
  IV U26562 ( .A(n25801), .Z(n25834) );
  XOR U26563 ( .A(n25835), .B(n25836), .Z(n25801) );
  ANDN U26564 ( .B(n25837), .A(n25838), .Z(n25835) );
  XOR U26565 ( .A(n25836), .B(n25839), .Z(n25837) );
  XNOR U26566 ( .A(n25840), .B(n25841), .Z(n25798) );
  ANDN U26567 ( .B(n25842), .A(n25843), .Z(n25840) );
  XOR U26568 ( .A(n25841), .B(n25844), .Z(n25842) );
  IV U26569 ( .A(n25797), .Z(n25832) );
  XOR U26570 ( .A(n25795), .B(n25845), .Z(n25797) );
  XNOR U26571 ( .A(n25846), .B(n25847), .Z(n25845) );
  ANDN U26572 ( .B(n25848), .A(n25849), .Z(n25846) );
  XNOR U26573 ( .A(n25850), .B(n25851), .Z(n25848) );
  IV U26574 ( .A(n25799), .Z(n25795) );
  XOR U26575 ( .A(n25852), .B(n25853), .Z(n25799) );
  ANDN U26576 ( .B(n25854), .A(n25855), .Z(n25852) );
  XOR U26577 ( .A(n25856), .B(n25853), .Z(n25854) );
  XOR U26578 ( .A(n25810), .B(n25663), .Z(n25811) );
  XOR U26579 ( .A(n25857), .B(n25858), .Z(n25663) );
  AND U26580 ( .A(n288), .B(n25859), .Z(n25857) );
  XOR U26581 ( .A(n25860), .B(n25858), .Z(n25859) );
  XNOR U26582 ( .A(n25861), .B(n25862), .Z(n25810) );
  NAND U26583 ( .A(n25863), .B(n25864), .Z(n25862) );
  XOR U26584 ( .A(n25865), .B(n25762), .Z(n25864) );
  XOR U26585 ( .A(n25838), .B(n25839), .Z(n25762) );
  XOR U26586 ( .A(n25866), .B(n25831), .Z(n25839) );
  XOR U26587 ( .A(n25867), .B(n25819), .Z(n25831) );
  XOR U26588 ( .A(n25868), .B(n25869), .Z(n25819) );
  ANDN U26589 ( .B(n25870), .A(n25871), .Z(n25868) );
  XOR U26590 ( .A(n25869), .B(n25872), .Z(n25870) );
  IV U26591 ( .A(n25817), .Z(n25867) );
  XOR U26592 ( .A(n25815), .B(n25873), .Z(n25817) );
  XOR U26593 ( .A(n25874), .B(n25875), .Z(n25873) );
  ANDN U26594 ( .B(n25876), .A(n25877), .Z(n25874) );
  XOR U26595 ( .A(n25878), .B(n25875), .Z(n25876) );
  IV U26596 ( .A(n25818), .Z(n25815) );
  XOR U26597 ( .A(n25879), .B(n25880), .Z(n25818) );
  ANDN U26598 ( .B(n25881), .A(n25882), .Z(n25879) );
  XOR U26599 ( .A(n25880), .B(n25883), .Z(n25881) );
  IV U26600 ( .A(n25830), .Z(n25866) );
  XOR U26601 ( .A(n25884), .B(n25885), .Z(n25830) );
  XNOR U26602 ( .A(n25825), .B(n25886), .Z(n25885) );
  IV U26603 ( .A(n25828), .Z(n25886) );
  XOR U26604 ( .A(n25887), .B(n25888), .Z(n25828) );
  ANDN U26605 ( .B(n25889), .A(n25890), .Z(n25887) );
  XOR U26606 ( .A(n25888), .B(n25891), .Z(n25889) );
  XNOR U26607 ( .A(n25892), .B(n25893), .Z(n25825) );
  ANDN U26608 ( .B(n25894), .A(n25895), .Z(n25892) );
  XOR U26609 ( .A(n25893), .B(n25896), .Z(n25894) );
  IV U26610 ( .A(n25824), .Z(n25884) );
  XOR U26611 ( .A(n25822), .B(n25897), .Z(n25824) );
  XOR U26612 ( .A(n25898), .B(n25899), .Z(n25897) );
  ANDN U26613 ( .B(n25900), .A(n25901), .Z(n25898) );
  XOR U26614 ( .A(n25902), .B(n25899), .Z(n25900) );
  IV U26615 ( .A(n25826), .Z(n25822) );
  XOR U26616 ( .A(n25903), .B(n25904), .Z(n25826) );
  ANDN U26617 ( .B(n25905), .A(n25906), .Z(n25903) );
  XOR U26618 ( .A(n25907), .B(n25904), .Z(n25905) );
  XOR U26619 ( .A(n25908), .B(n25909), .Z(n25838) );
  XOR U26620 ( .A(n25856), .B(n25910), .Z(n25909) );
  IV U26621 ( .A(n25836), .Z(n25910) );
  XOR U26622 ( .A(n25911), .B(n25912), .Z(n25836) );
  ANDN U26623 ( .B(n25913), .A(n25914), .Z(n25911) );
  XOR U26624 ( .A(n25912), .B(n25915), .Z(n25913) );
  XOR U26625 ( .A(n25916), .B(n25844), .Z(n25856) );
  XOR U26626 ( .A(n25917), .B(n25918), .Z(n25844) );
  ANDN U26627 ( .B(n25919), .A(n25920), .Z(n25917) );
  XOR U26628 ( .A(n25918), .B(n25921), .Z(n25919) );
  IV U26629 ( .A(n25843), .Z(n25916) );
  XOR U26630 ( .A(n25922), .B(n25923), .Z(n25843) );
  XOR U26631 ( .A(n25924), .B(n25925), .Z(n25923) );
  ANDN U26632 ( .B(n25926), .A(n25927), .Z(n25924) );
  XOR U26633 ( .A(n25928), .B(n25925), .Z(n25926) );
  IV U26634 ( .A(n25841), .Z(n25922) );
  XOR U26635 ( .A(n25929), .B(n25930), .Z(n25841) );
  ANDN U26636 ( .B(n25931), .A(n25932), .Z(n25929) );
  XOR U26637 ( .A(n25930), .B(n25933), .Z(n25931) );
  IV U26638 ( .A(n25855), .Z(n25908) );
  XOR U26639 ( .A(n25934), .B(n25935), .Z(n25855) );
  XNOR U26640 ( .A(n25850), .B(n25936), .Z(n25935) );
  IV U26641 ( .A(n25853), .Z(n25936) );
  XOR U26642 ( .A(n25937), .B(n25938), .Z(n25853) );
  ANDN U26643 ( .B(n25939), .A(n25940), .Z(n25937) );
  XOR U26644 ( .A(n25941), .B(n25938), .Z(n25939) );
  XNOR U26645 ( .A(n25942), .B(n25943), .Z(n25850) );
  ANDN U26646 ( .B(n25944), .A(n25945), .Z(n25942) );
  XOR U26647 ( .A(n25943), .B(n25946), .Z(n25944) );
  IV U26648 ( .A(n25849), .Z(n25934) );
  XOR U26649 ( .A(n25847), .B(n25947), .Z(n25849) );
  XOR U26650 ( .A(n25948), .B(n25949), .Z(n25947) );
  ANDN U26651 ( .B(n25950), .A(n25951), .Z(n25948) );
  XOR U26652 ( .A(n25952), .B(n25949), .Z(n25950) );
  IV U26653 ( .A(n25851), .Z(n25847) );
  XOR U26654 ( .A(n25953), .B(n25954), .Z(n25851) );
  ANDN U26655 ( .B(n25955), .A(n25956), .Z(n25953) );
  XOR U26656 ( .A(n25957), .B(n25954), .Z(n25955) );
  IV U26657 ( .A(n25861), .Z(n25865) );
  XOR U26658 ( .A(n25861), .B(n25764), .Z(n25863) );
  XOR U26659 ( .A(n25958), .B(n25959), .Z(n25764) );
  AND U26660 ( .A(n288), .B(n25960), .Z(n25958) );
  XOR U26661 ( .A(n25961), .B(n25959), .Z(n25960) );
  NANDN U26662 ( .A(n25766), .B(n25768), .Z(n25861) );
  XOR U26663 ( .A(n25962), .B(n25963), .Z(n25768) );
  AND U26664 ( .A(n288), .B(n25964), .Z(n25962) );
  XOR U26665 ( .A(n25963), .B(n25965), .Z(n25964) );
  XNOR U26666 ( .A(n25966), .B(n25967), .Z(n288) );
  AND U26667 ( .A(n25968), .B(n25969), .Z(n25966) );
  XOR U26668 ( .A(n25967), .B(n25779), .Z(n25969) );
  XNOR U26669 ( .A(n25970), .B(n25971), .Z(n25779) );
  ANDN U26670 ( .B(n25972), .A(n25973), .Z(n25970) );
  XOR U26671 ( .A(n25971), .B(n25974), .Z(n25972) );
  XNOR U26672 ( .A(n25967), .B(n25781), .Z(n25968) );
  XOR U26673 ( .A(n25975), .B(n25976), .Z(n25781) );
  AND U26674 ( .A(n292), .B(n25977), .Z(n25975) );
  XOR U26675 ( .A(n25978), .B(n25976), .Z(n25977) );
  XOR U26676 ( .A(n25979), .B(n25980), .Z(n25967) );
  AND U26677 ( .A(n25981), .B(n25982), .Z(n25979) );
  XOR U26678 ( .A(n25980), .B(n25806), .Z(n25982) );
  XOR U26679 ( .A(n25973), .B(n25974), .Z(n25806) );
  XNOR U26680 ( .A(n25983), .B(n25984), .Z(n25974) );
  ANDN U26681 ( .B(n25985), .A(n25986), .Z(n25983) );
  XOR U26682 ( .A(n25987), .B(n25988), .Z(n25985) );
  XOR U26683 ( .A(n25989), .B(n25990), .Z(n25973) );
  XNOR U26684 ( .A(n25991), .B(n25992), .Z(n25990) );
  ANDN U26685 ( .B(n25993), .A(n25994), .Z(n25991) );
  XNOR U26686 ( .A(n25995), .B(n25996), .Z(n25993) );
  IV U26687 ( .A(n25971), .Z(n25989) );
  XOR U26688 ( .A(n25997), .B(n25998), .Z(n25971) );
  ANDN U26689 ( .B(n25999), .A(n26000), .Z(n25997) );
  XOR U26690 ( .A(n25998), .B(n26001), .Z(n25999) );
  XNOR U26691 ( .A(n25980), .B(n25808), .Z(n25981) );
  XOR U26692 ( .A(n26002), .B(n26003), .Z(n25808) );
  AND U26693 ( .A(n292), .B(n26004), .Z(n26002) );
  XOR U26694 ( .A(n26005), .B(n26003), .Z(n26004) );
  XNOR U26695 ( .A(n26006), .B(n26007), .Z(n25980) );
  AND U26696 ( .A(n26008), .B(n26009), .Z(n26006) );
  XNOR U26697 ( .A(n26007), .B(n25858), .Z(n26009) );
  XOR U26698 ( .A(n26000), .B(n26001), .Z(n25858) );
  XOR U26699 ( .A(n26010), .B(n25988), .Z(n26001) );
  XNOR U26700 ( .A(n26011), .B(n26012), .Z(n25988) );
  ANDN U26701 ( .B(n26013), .A(n26014), .Z(n26011) );
  XOR U26702 ( .A(n26015), .B(n26016), .Z(n26013) );
  IV U26703 ( .A(n25986), .Z(n26010) );
  XOR U26704 ( .A(n25984), .B(n26017), .Z(n25986) );
  XNOR U26705 ( .A(n26018), .B(n26019), .Z(n26017) );
  ANDN U26706 ( .B(n26020), .A(n26021), .Z(n26018) );
  XNOR U26707 ( .A(n26022), .B(n26023), .Z(n26020) );
  IV U26708 ( .A(n25987), .Z(n25984) );
  XOR U26709 ( .A(n26024), .B(n26025), .Z(n25987) );
  ANDN U26710 ( .B(n26026), .A(n26027), .Z(n26024) );
  XOR U26711 ( .A(n26025), .B(n26028), .Z(n26026) );
  XOR U26712 ( .A(n26029), .B(n26030), .Z(n26000) );
  XNOR U26713 ( .A(n25995), .B(n26031), .Z(n26030) );
  IV U26714 ( .A(n25998), .Z(n26031) );
  XOR U26715 ( .A(n26032), .B(n26033), .Z(n25998) );
  ANDN U26716 ( .B(n26034), .A(n26035), .Z(n26032) );
  XOR U26717 ( .A(n26033), .B(n26036), .Z(n26034) );
  XNOR U26718 ( .A(n26037), .B(n26038), .Z(n25995) );
  ANDN U26719 ( .B(n26039), .A(n26040), .Z(n26037) );
  XOR U26720 ( .A(n26038), .B(n26041), .Z(n26039) );
  IV U26721 ( .A(n25994), .Z(n26029) );
  XOR U26722 ( .A(n25992), .B(n26042), .Z(n25994) );
  XNOR U26723 ( .A(n26043), .B(n26044), .Z(n26042) );
  ANDN U26724 ( .B(n26045), .A(n26046), .Z(n26043) );
  XNOR U26725 ( .A(n26047), .B(n26048), .Z(n26045) );
  IV U26726 ( .A(n25996), .Z(n25992) );
  XOR U26727 ( .A(n26049), .B(n26050), .Z(n25996) );
  ANDN U26728 ( .B(n26051), .A(n26052), .Z(n26049) );
  XOR U26729 ( .A(n26053), .B(n26050), .Z(n26051) );
  XOR U26730 ( .A(n26007), .B(n25860), .Z(n26008) );
  XOR U26731 ( .A(n26054), .B(n26055), .Z(n25860) );
  AND U26732 ( .A(n292), .B(n26056), .Z(n26054) );
  XOR U26733 ( .A(n26057), .B(n26055), .Z(n26056) );
  XNOR U26734 ( .A(n26058), .B(n26059), .Z(n26007) );
  NAND U26735 ( .A(n26060), .B(n26061), .Z(n26059) );
  XOR U26736 ( .A(n26062), .B(n25959), .Z(n26061) );
  XOR U26737 ( .A(n26035), .B(n26036), .Z(n25959) );
  XOR U26738 ( .A(n26063), .B(n26028), .Z(n26036) );
  XOR U26739 ( .A(n26064), .B(n26016), .Z(n26028) );
  XOR U26740 ( .A(n26065), .B(n26066), .Z(n26016) );
  ANDN U26741 ( .B(n26067), .A(n26068), .Z(n26065) );
  XOR U26742 ( .A(n26066), .B(n26069), .Z(n26067) );
  IV U26743 ( .A(n26014), .Z(n26064) );
  XOR U26744 ( .A(n26012), .B(n26070), .Z(n26014) );
  XOR U26745 ( .A(n26071), .B(n26072), .Z(n26070) );
  ANDN U26746 ( .B(n26073), .A(n26074), .Z(n26071) );
  XOR U26747 ( .A(n26075), .B(n26072), .Z(n26073) );
  IV U26748 ( .A(n26015), .Z(n26012) );
  XOR U26749 ( .A(n26076), .B(n26077), .Z(n26015) );
  ANDN U26750 ( .B(n26078), .A(n26079), .Z(n26076) );
  XOR U26751 ( .A(n26077), .B(n26080), .Z(n26078) );
  IV U26752 ( .A(n26027), .Z(n26063) );
  XOR U26753 ( .A(n26081), .B(n26082), .Z(n26027) );
  XNOR U26754 ( .A(n26022), .B(n26083), .Z(n26082) );
  IV U26755 ( .A(n26025), .Z(n26083) );
  XOR U26756 ( .A(n26084), .B(n26085), .Z(n26025) );
  ANDN U26757 ( .B(n26086), .A(n26087), .Z(n26084) );
  XOR U26758 ( .A(n26085), .B(n26088), .Z(n26086) );
  XNOR U26759 ( .A(n26089), .B(n26090), .Z(n26022) );
  ANDN U26760 ( .B(n26091), .A(n26092), .Z(n26089) );
  XOR U26761 ( .A(n26090), .B(n26093), .Z(n26091) );
  IV U26762 ( .A(n26021), .Z(n26081) );
  XOR U26763 ( .A(n26019), .B(n26094), .Z(n26021) );
  XOR U26764 ( .A(n26095), .B(n26096), .Z(n26094) );
  ANDN U26765 ( .B(n26097), .A(n26098), .Z(n26095) );
  XOR U26766 ( .A(n26099), .B(n26096), .Z(n26097) );
  IV U26767 ( .A(n26023), .Z(n26019) );
  XOR U26768 ( .A(n26100), .B(n26101), .Z(n26023) );
  ANDN U26769 ( .B(n26102), .A(n26103), .Z(n26100) );
  XOR U26770 ( .A(n26104), .B(n26101), .Z(n26102) );
  XOR U26771 ( .A(n26105), .B(n26106), .Z(n26035) );
  XOR U26772 ( .A(n26053), .B(n26107), .Z(n26106) );
  IV U26773 ( .A(n26033), .Z(n26107) );
  XOR U26774 ( .A(n26108), .B(n26109), .Z(n26033) );
  ANDN U26775 ( .B(n26110), .A(n26111), .Z(n26108) );
  XOR U26776 ( .A(n26109), .B(n26112), .Z(n26110) );
  XOR U26777 ( .A(n26113), .B(n26041), .Z(n26053) );
  XOR U26778 ( .A(n26114), .B(n26115), .Z(n26041) );
  ANDN U26779 ( .B(n26116), .A(n26117), .Z(n26114) );
  XOR U26780 ( .A(n26115), .B(n26118), .Z(n26116) );
  IV U26781 ( .A(n26040), .Z(n26113) );
  XOR U26782 ( .A(n26119), .B(n26120), .Z(n26040) );
  XOR U26783 ( .A(n26121), .B(n26122), .Z(n26120) );
  ANDN U26784 ( .B(n26123), .A(n26124), .Z(n26121) );
  XOR U26785 ( .A(n26125), .B(n26122), .Z(n26123) );
  IV U26786 ( .A(n26038), .Z(n26119) );
  XOR U26787 ( .A(n26126), .B(n26127), .Z(n26038) );
  ANDN U26788 ( .B(n26128), .A(n26129), .Z(n26126) );
  XOR U26789 ( .A(n26127), .B(n26130), .Z(n26128) );
  IV U26790 ( .A(n26052), .Z(n26105) );
  XOR U26791 ( .A(n26131), .B(n26132), .Z(n26052) );
  XNOR U26792 ( .A(n26047), .B(n26133), .Z(n26132) );
  IV U26793 ( .A(n26050), .Z(n26133) );
  XOR U26794 ( .A(n26134), .B(n26135), .Z(n26050) );
  ANDN U26795 ( .B(n26136), .A(n26137), .Z(n26134) );
  XOR U26796 ( .A(n26138), .B(n26135), .Z(n26136) );
  XNOR U26797 ( .A(n26139), .B(n26140), .Z(n26047) );
  ANDN U26798 ( .B(n26141), .A(n26142), .Z(n26139) );
  XOR U26799 ( .A(n26140), .B(n26143), .Z(n26141) );
  IV U26800 ( .A(n26046), .Z(n26131) );
  XOR U26801 ( .A(n26044), .B(n26144), .Z(n26046) );
  XOR U26802 ( .A(n26145), .B(n26146), .Z(n26144) );
  ANDN U26803 ( .B(n26147), .A(n26148), .Z(n26145) );
  XOR U26804 ( .A(n26149), .B(n26146), .Z(n26147) );
  IV U26805 ( .A(n26048), .Z(n26044) );
  XOR U26806 ( .A(n26150), .B(n26151), .Z(n26048) );
  ANDN U26807 ( .B(n26152), .A(n26153), .Z(n26150) );
  XOR U26808 ( .A(n26154), .B(n26151), .Z(n26152) );
  IV U26809 ( .A(n26058), .Z(n26062) );
  XOR U26810 ( .A(n26058), .B(n25961), .Z(n26060) );
  XOR U26811 ( .A(n26155), .B(n26156), .Z(n25961) );
  AND U26812 ( .A(n292), .B(n26157), .Z(n26155) );
  XOR U26813 ( .A(n26158), .B(n26156), .Z(n26157) );
  NANDN U26814 ( .A(n25963), .B(n25965), .Z(n26058) );
  XOR U26815 ( .A(n26159), .B(n26160), .Z(n25965) );
  AND U26816 ( .A(n292), .B(n26161), .Z(n26159) );
  XOR U26817 ( .A(n26160), .B(n26162), .Z(n26161) );
  XNOR U26818 ( .A(n26163), .B(n26164), .Z(n292) );
  AND U26819 ( .A(n26165), .B(n26166), .Z(n26163) );
  XOR U26820 ( .A(n26164), .B(n25976), .Z(n26166) );
  XNOR U26821 ( .A(n26167), .B(n26168), .Z(n25976) );
  ANDN U26822 ( .B(n26169), .A(n26170), .Z(n26167) );
  XOR U26823 ( .A(n26168), .B(n26171), .Z(n26169) );
  XNOR U26824 ( .A(n26164), .B(n25978), .Z(n26165) );
  XOR U26825 ( .A(n26172), .B(n26173), .Z(n25978) );
  AND U26826 ( .A(n296), .B(n26174), .Z(n26172) );
  XOR U26827 ( .A(n26175), .B(n26173), .Z(n26174) );
  XOR U26828 ( .A(n26176), .B(n26177), .Z(n26164) );
  AND U26829 ( .A(n26178), .B(n26179), .Z(n26176) );
  XOR U26830 ( .A(n26177), .B(n26003), .Z(n26179) );
  XOR U26831 ( .A(n26170), .B(n26171), .Z(n26003) );
  XNOR U26832 ( .A(n26180), .B(n26181), .Z(n26171) );
  ANDN U26833 ( .B(n26182), .A(n26183), .Z(n26180) );
  XOR U26834 ( .A(n26184), .B(n26185), .Z(n26182) );
  XOR U26835 ( .A(n26186), .B(n26187), .Z(n26170) );
  XNOR U26836 ( .A(n26188), .B(n26189), .Z(n26187) );
  ANDN U26837 ( .B(n26190), .A(n26191), .Z(n26188) );
  XNOR U26838 ( .A(n26192), .B(n26193), .Z(n26190) );
  IV U26839 ( .A(n26168), .Z(n26186) );
  XOR U26840 ( .A(n26194), .B(n26195), .Z(n26168) );
  ANDN U26841 ( .B(n26196), .A(n26197), .Z(n26194) );
  XOR U26842 ( .A(n26195), .B(n26198), .Z(n26196) );
  XNOR U26843 ( .A(n26177), .B(n26005), .Z(n26178) );
  XOR U26844 ( .A(n26199), .B(n26200), .Z(n26005) );
  AND U26845 ( .A(n296), .B(n26201), .Z(n26199) );
  XOR U26846 ( .A(n26202), .B(n26200), .Z(n26201) );
  XNOR U26847 ( .A(n26203), .B(n26204), .Z(n26177) );
  AND U26848 ( .A(n26205), .B(n26206), .Z(n26203) );
  XNOR U26849 ( .A(n26204), .B(n26055), .Z(n26206) );
  XOR U26850 ( .A(n26197), .B(n26198), .Z(n26055) );
  XOR U26851 ( .A(n26207), .B(n26185), .Z(n26198) );
  XNOR U26852 ( .A(n26208), .B(n26209), .Z(n26185) );
  ANDN U26853 ( .B(n26210), .A(n26211), .Z(n26208) );
  XOR U26854 ( .A(n26212), .B(n26213), .Z(n26210) );
  IV U26855 ( .A(n26183), .Z(n26207) );
  XOR U26856 ( .A(n26181), .B(n26214), .Z(n26183) );
  XNOR U26857 ( .A(n26215), .B(n26216), .Z(n26214) );
  ANDN U26858 ( .B(n26217), .A(n26218), .Z(n26215) );
  XNOR U26859 ( .A(n26219), .B(n26220), .Z(n26217) );
  IV U26860 ( .A(n26184), .Z(n26181) );
  XOR U26861 ( .A(n26221), .B(n26222), .Z(n26184) );
  ANDN U26862 ( .B(n26223), .A(n26224), .Z(n26221) );
  XOR U26863 ( .A(n26222), .B(n26225), .Z(n26223) );
  XOR U26864 ( .A(n26226), .B(n26227), .Z(n26197) );
  XNOR U26865 ( .A(n26192), .B(n26228), .Z(n26227) );
  IV U26866 ( .A(n26195), .Z(n26228) );
  XOR U26867 ( .A(n26229), .B(n26230), .Z(n26195) );
  ANDN U26868 ( .B(n26231), .A(n26232), .Z(n26229) );
  XOR U26869 ( .A(n26230), .B(n26233), .Z(n26231) );
  XNOR U26870 ( .A(n26234), .B(n26235), .Z(n26192) );
  ANDN U26871 ( .B(n26236), .A(n26237), .Z(n26234) );
  XOR U26872 ( .A(n26235), .B(n26238), .Z(n26236) );
  IV U26873 ( .A(n26191), .Z(n26226) );
  XOR U26874 ( .A(n26189), .B(n26239), .Z(n26191) );
  XNOR U26875 ( .A(n26240), .B(n26241), .Z(n26239) );
  ANDN U26876 ( .B(n26242), .A(n26243), .Z(n26240) );
  XNOR U26877 ( .A(n26244), .B(n26245), .Z(n26242) );
  IV U26878 ( .A(n26193), .Z(n26189) );
  XOR U26879 ( .A(n26246), .B(n26247), .Z(n26193) );
  ANDN U26880 ( .B(n26248), .A(n26249), .Z(n26246) );
  XOR U26881 ( .A(n26250), .B(n26247), .Z(n26248) );
  XOR U26882 ( .A(n26204), .B(n26057), .Z(n26205) );
  XOR U26883 ( .A(n26251), .B(n26252), .Z(n26057) );
  AND U26884 ( .A(n296), .B(n26253), .Z(n26251) );
  XOR U26885 ( .A(n26254), .B(n26252), .Z(n26253) );
  XNOR U26886 ( .A(n26255), .B(n26256), .Z(n26204) );
  NAND U26887 ( .A(n26257), .B(n26258), .Z(n26256) );
  XOR U26888 ( .A(n26259), .B(n26156), .Z(n26258) );
  XOR U26889 ( .A(n26232), .B(n26233), .Z(n26156) );
  XOR U26890 ( .A(n26260), .B(n26225), .Z(n26233) );
  XOR U26891 ( .A(n26261), .B(n26213), .Z(n26225) );
  XOR U26892 ( .A(n26262), .B(n26263), .Z(n26213) );
  ANDN U26893 ( .B(n26264), .A(n26265), .Z(n26262) );
  XOR U26894 ( .A(n26263), .B(n26266), .Z(n26264) );
  IV U26895 ( .A(n26211), .Z(n26261) );
  XOR U26896 ( .A(n26209), .B(n26267), .Z(n26211) );
  XOR U26897 ( .A(n26268), .B(n26269), .Z(n26267) );
  ANDN U26898 ( .B(n26270), .A(n26271), .Z(n26268) );
  XOR U26899 ( .A(n26272), .B(n26269), .Z(n26270) );
  IV U26900 ( .A(n26212), .Z(n26209) );
  XOR U26901 ( .A(n26273), .B(n26274), .Z(n26212) );
  ANDN U26902 ( .B(n26275), .A(n26276), .Z(n26273) );
  XOR U26903 ( .A(n26274), .B(n26277), .Z(n26275) );
  IV U26904 ( .A(n26224), .Z(n26260) );
  XOR U26905 ( .A(n26278), .B(n26279), .Z(n26224) );
  XNOR U26906 ( .A(n26219), .B(n26280), .Z(n26279) );
  IV U26907 ( .A(n26222), .Z(n26280) );
  XOR U26908 ( .A(n26281), .B(n26282), .Z(n26222) );
  ANDN U26909 ( .B(n26283), .A(n26284), .Z(n26281) );
  XOR U26910 ( .A(n26282), .B(n26285), .Z(n26283) );
  XNOR U26911 ( .A(n26286), .B(n26287), .Z(n26219) );
  ANDN U26912 ( .B(n26288), .A(n26289), .Z(n26286) );
  XOR U26913 ( .A(n26287), .B(n26290), .Z(n26288) );
  IV U26914 ( .A(n26218), .Z(n26278) );
  XOR U26915 ( .A(n26216), .B(n26291), .Z(n26218) );
  XOR U26916 ( .A(n26292), .B(n26293), .Z(n26291) );
  ANDN U26917 ( .B(n26294), .A(n26295), .Z(n26292) );
  XOR U26918 ( .A(n26296), .B(n26293), .Z(n26294) );
  IV U26919 ( .A(n26220), .Z(n26216) );
  XOR U26920 ( .A(n26297), .B(n26298), .Z(n26220) );
  ANDN U26921 ( .B(n26299), .A(n26300), .Z(n26297) );
  XOR U26922 ( .A(n26301), .B(n26298), .Z(n26299) );
  XOR U26923 ( .A(n26302), .B(n26303), .Z(n26232) );
  XOR U26924 ( .A(n26250), .B(n26304), .Z(n26303) );
  IV U26925 ( .A(n26230), .Z(n26304) );
  XOR U26926 ( .A(n26305), .B(n26306), .Z(n26230) );
  ANDN U26927 ( .B(n26307), .A(n26308), .Z(n26305) );
  XOR U26928 ( .A(n26306), .B(n26309), .Z(n26307) );
  XOR U26929 ( .A(n26310), .B(n26238), .Z(n26250) );
  XOR U26930 ( .A(n26311), .B(n26312), .Z(n26238) );
  ANDN U26931 ( .B(n26313), .A(n26314), .Z(n26311) );
  XOR U26932 ( .A(n26312), .B(n26315), .Z(n26313) );
  IV U26933 ( .A(n26237), .Z(n26310) );
  XOR U26934 ( .A(n26316), .B(n26317), .Z(n26237) );
  XOR U26935 ( .A(n26318), .B(n26319), .Z(n26317) );
  ANDN U26936 ( .B(n26320), .A(n26321), .Z(n26318) );
  XOR U26937 ( .A(n26322), .B(n26319), .Z(n26320) );
  IV U26938 ( .A(n26235), .Z(n26316) );
  XOR U26939 ( .A(n26323), .B(n26324), .Z(n26235) );
  ANDN U26940 ( .B(n26325), .A(n26326), .Z(n26323) );
  XOR U26941 ( .A(n26324), .B(n26327), .Z(n26325) );
  IV U26942 ( .A(n26249), .Z(n26302) );
  XOR U26943 ( .A(n26328), .B(n26329), .Z(n26249) );
  XNOR U26944 ( .A(n26244), .B(n26330), .Z(n26329) );
  IV U26945 ( .A(n26247), .Z(n26330) );
  XOR U26946 ( .A(n26331), .B(n26332), .Z(n26247) );
  ANDN U26947 ( .B(n26333), .A(n26334), .Z(n26331) );
  XOR U26948 ( .A(n26335), .B(n26332), .Z(n26333) );
  XNOR U26949 ( .A(n26336), .B(n26337), .Z(n26244) );
  ANDN U26950 ( .B(n26338), .A(n26339), .Z(n26336) );
  XOR U26951 ( .A(n26337), .B(n26340), .Z(n26338) );
  IV U26952 ( .A(n26243), .Z(n26328) );
  XOR U26953 ( .A(n26241), .B(n26341), .Z(n26243) );
  XOR U26954 ( .A(n26342), .B(n26343), .Z(n26341) );
  ANDN U26955 ( .B(n26344), .A(n26345), .Z(n26342) );
  XOR U26956 ( .A(n26346), .B(n26343), .Z(n26344) );
  IV U26957 ( .A(n26245), .Z(n26241) );
  XOR U26958 ( .A(n26347), .B(n26348), .Z(n26245) );
  ANDN U26959 ( .B(n26349), .A(n26350), .Z(n26347) );
  XOR U26960 ( .A(n26351), .B(n26348), .Z(n26349) );
  IV U26961 ( .A(n26255), .Z(n26259) );
  XOR U26962 ( .A(n26255), .B(n26158), .Z(n26257) );
  XOR U26963 ( .A(n26352), .B(n26353), .Z(n26158) );
  AND U26964 ( .A(n296), .B(n26354), .Z(n26352) );
  XOR U26965 ( .A(n26355), .B(n26353), .Z(n26354) );
  NANDN U26966 ( .A(n26160), .B(n26162), .Z(n26255) );
  XOR U26967 ( .A(n26356), .B(n26357), .Z(n26162) );
  AND U26968 ( .A(n296), .B(n26358), .Z(n26356) );
  XOR U26969 ( .A(n26357), .B(n26359), .Z(n26358) );
  XNOR U26970 ( .A(n26360), .B(n26361), .Z(n296) );
  AND U26971 ( .A(n26362), .B(n26363), .Z(n26360) );
  XOR U26972 ( .A(n26361), .B(n26173), .Z(n26363) );
  XNOR U26973 ( .A(n26364), .B(n26365), .Z(n26173) );
  ANDN U26974 ( .B(n26366), .A(n26367), .Z(n26364) );
  XOR U26975 ( .A(n26365), .B(n26368), .Z(n26366) );
  XNOR U26976 ( .A(n26361), .B(n26175), .Z(n26362) );
  XOR U26977 ( .A(n26369), .B(n26370), .Z(n26175) );
  AND U26978 ( .A(n300), .B(n26371), .Z(n26369) );
  XOR U26979 ( .A(n26372), .B(n26370), .Z(n26371) );
  XOR U26980 ( .A(n26373), .B(n26374), .Z(n26361) );
  AND U26981 ( .A(n26375), .B(n26376), .Z(n26373) );
  XOR U26982 ( .A(n26374), .B(n26200), .Z(n26376) );
  XOR U26983 ( .A(n26367), .B(n26368), .Z(n26200) );
  XNOR U26984 ( .A(n26377), .B(n26378), .Z(n26368) );
  ANDN U26985 ( .B(n26379), .A(n26380), .Z(n26377) );
  XOR U26986 ( .A(n26381), .B(n26382), .Z(n26379) );
  XOR U26987 ( .A(n26383), .B(n26384), .Z(n26367) );
  XNOR U26988 ( .A(n26385), .B(n26386), .Z(n26384) );
  ANDN U26989 ( .B(n26387), .A(n26388), .Z(n26385) );
  XNOR U26990 ( .A(n26389), .B(n26390), .Z(n26387) );
  IV U26991 ( .A(n26365), .Z(n26383) );
  XOR U26992 ( .A(n26391), .B(n26392), .Z(n26365) );
  ANDN U26993 ( .B(n26393), .A(n26394), .Z(n26391) );
  XOR U26994 ( .A(n26392), .B(n26395), .Z(n26393) );
  XNOR U26995 ( .A(n26374), .B(n26202), .Z(n26375) );
  XOR U26996 ( .A(n26396), .B(n26397), .Z(n26202) );
  AND U26997 ( .A(n300), .B(n26398), .Z(n26396) );
  XOR U26998 ( .A(n26399), .B(n26397), .Z(n26398) );
  XNOR U26999 ( .A(n26400), .B(n26401), .Z(n26374) );
  AND U27000 ( .A(n26402), .B(n26403), .Z(n26400) );
  XNOR U27001 ( .A(n26401), .B(n26252), .Z(n26403) );
  XOR U27002 ( .A(n26394), .B(n26395), .Z(n26252) );
  XOR U27003 ( .A(n26404), .B(n26382), .Z(n26395) );
  XNOR U27004 ( .A(n26405), .B(n26406), .Z(n26382) );
  ANDN U27005 ( .B(n26407), .A(n26408), .Z(n26405) );
  XOR U27006 ( .A(n26409), .B(n26410), .Z(n26407) );
  IV U27007 ( .A(n26380), .Z(n26404) );
  XOR U27008 ( .A(n26378), .B(n26411), .Z(n26380) );
  XNOR U27009 ( .A(n26412), .B(n26413), .Z(n26411) );
  ANDN U27010 ( .B(n26414), .A(n26415), .Z(n26412) );
  XNOR U27011 ( .A(n26416), .B(n26417), .Z(n26414) );
  IV U27012 ( .A(n26381), .Z(n26378) );
  XOR U27013 ( .A(n26418), .B(n26419), .Z(n26381) );
  ANDN U27014 ( .B(n26420), .A(n26421), .Z(n26418) );
  XOR U27015 ( .A(n26419), .B(n26422), .Z(n26420) );
  XOR U27016 ( .A(n26423), .B(n26424), .Z(n26394) );
  XNOR U27017 ( .A(n26389), .B(n26425), .Z(n26424) );
  IV U27018 ( .A(n26392), .Z(n26425) );
  XOR U27019 ( .A(n26426), .B(n26427), .Z(n26392) );
  ANDN U27020 ( .B(n26428), .A(n26429), .Z(n26426) );
  XOR U27021 ( .A(n26427), .B(n26430), .Z(n26428) );
  XNOR U27022 ( .A(n26431), .B(n26432), .Z(n26389) );
  ANDN U27023 ( .B(n26433), .A(n26434), .Z(n26431) );
  XOR U27024 ( .A(n26432), .B(n26435), .Z(n26433) );
  IV U27025 ( .A(n26388), .Z(n26423) );
  XOR U27026 ( .A(n26386), .B(n26436), .Z(n26388) );
  XNOR U27027 ( .A(n26437), .B(n26438), .Z(n26436) );
  ANDN U27028 ( .B(n26439), .A(n26440), .Z(n26437) );
  XNOR U27029 ( .A(n26441), .B(n26442), .Z(n26439) );
  IV U27030 ( .A(n26390), .Z(n26386) );
  XOR U27031 ( .A(n26443), .B(n26444), .Z(n26390) );
  ANDN U27032 ( .B(n26445), .A(n26446), .Z(n26443) );
  XOR U27033 ( .A(n26447), .B(n26444), .Z(n26445) );
  XOR U27034 ( .A(n26401), .B(n26254), .Z(n26402) );
  XOR U27035 ( .A(n26448), .B(n26449), .Z(n26254) );
  AND U27036 ( .A(n300), .B(n26450), .Z(n26448) );
  XOR U27037 ( .A(n26451), .B(n26449), .Z(n26450) );
  XNOR U27038 ( .A(n26452), .B(n26453), .Z(n26401) );
  NAND U27039 ( .A(n26454), .B(n26455), .Z(n26453) );
  XOR U27040 ( .A(n26456), .B(n26353), .Z(n26455) );
  XOR U27041 ( .A(n26429), .B(n26430), .Z(n26353) );
  XOR U27042 ( .A(n26457), .B(n26422), .Z(n26430) );
  XOR U27043 ( .A(n26458), .B(n26410), .Z(n26422) );
  XOR U27044 ( .A(n26459), .B(n26460), .Z(n26410) );
  ANDN U27045 ( .B(n26461), .A(n26462), .Z(n26459) );
  XOR U27046 ( .A(n26460), .B(n26463), .Z(n26461) );
  IV U27047 ( .A(n26408), .Z(n26458) );
  XOR U27048 ( .A(n26406), .B(n26464), .Z(n26408) );
  XOR U27049 ( .A(n26465), .B(n26466), .Z(n26464) );
  ANDN U27050 ( .B(n26467), .A(n26468), .Z(n26465) );
  XOR U27051 ( .A(n26469), .B(n26466), .Z(n26467) );
  IV U27052 ( .A(n26409), .Z(n26406) );
  XOR U27053 ( .A(n26470), .B(n26471), .Z(n26409) );
  ANDN U27054 ( .B(n26472), .A(n26473), .Z(n26470) );
  XOR U27055 ( .A(n26471), .B(n26474), .Z(n26472) );
  IV U27056 ( .A(n26421), .Z(n26457) );
  XOR U27057 ( .A(n26475), .B(n26476), .Z(n26421) );
  XNOR U27058 ( .A(n26416), .B(n26477), .Z(n26476) );
  IV U27059 ( .A(n26419), .Z(n26477) );
  XOR U27060 ( .A(n26478), .B(n26479), .Z(n26419) );
  ANDN U27061 ( .B(n26480), .A(n26481), .Z(n26478) );
  XOR U27062 ( .A(n26479), .B(n26482), .Z(n26480) );
  XNOR U27063 ( .A(n26483), .B(n26484), .Z(n26416) );
  ANDN U27064 ( .B(n26485), .A(n26486), .Z(n26483) );
  XOR U27065 ( .A(n26484), .B(n26487), .Z(n26485) );
  IV U27066 ( .A(n26415), .Z(n26475) );
  XOR U27067 ( .A(n26413), .B(n26488), .Z(n26415) );
  XOR U27068 ( .A(n26489), .B(n26490), .Z(n26488) );
  ANDN U27069 ( .B(n26491), .A(n26492), .Z(n26489) );
  XOR U27070 ( .A(n26493), .B(n26490), .Z(n26491) );
  IV U27071 ( .A(n26417), .Z(n26413) );
  XOR U27072 ( .A(n26494), .B(n26495), .Z(n26417) );
  ANDN U27073 ( .B(n26496), .A(n26497), .Z(n26494) );
  XOR U27074 ( .A(n26498), .B(n26495), .Z(n26496) );
  XOR U27075 ( .A(n26499), .B(n26500), .Z(n26429) );
  XOR U27076 ( .A(n26447), .B(n26501), .Z(n26500) );
  IV U27077 ( .A(n26427), .Z(n26501) );
  XOR U27078 ( .A(n26502), .B(n26503), .Z(n26427) );
  ANDN U27079 ( .B(n26504), .A(n26505), .Z(n26502) );
  XOR U27080 ( .A(n26503), .B(n26506), .Z(n26504) );
  XOR U27081 ( .A(n26507), .B(n26435), .Z(n26447) );
  XOR U27082 ( .A(n26508), .B(n26509), .Z(n26435) );
  ANDN U27083 ( .B(n26510), .A(n26511), .Z(n26508) );
  XOR U27084 ( .A(n26509), .B(n26512), .Z(n26510) );
  IV U27085 ( .A(n26434), .Z(n26507) );
  XOR U27086 ( .A(n26513), .B(n26514), .Z(n26434) );
  XOR U27087 ( .A(n26515), .B(n26516), .Z(n26514) );
  ANDN U27088 ( .B(n26517), .A(n26518), .Z(n26515) );
  XOR U27089 ( .A(n26519), .B(n26516), .Z(n26517) );
  IV U27090 ( .A(n26432), .Z(n26513) );
  XOR U27091 ( .A(n26520), .B(n26521), .Z(n26432) );
  ANDN U27092 ( .B(n26522), .A(n26523), .Z(n26520) );
  XOR U27093 ( .A(n26521), .B(n26524), .Z(n26522) );
  IV U27094 ( .A(n26446), .Z(n26499) );
  XOR U27095 ( .A(n26525), .B(n26526), .Z(n26446) );
  XNOR U27096 ( .A(n26441), .B(n26527), .Z(n26526) );
  IV U27097 ( .A(n26444), .Z(n26527) );
  XOR U27098 ( .A(n26528), .B(n26529), .Z(n26444) );
  ANDN U27099 ( .B(n26530), .A(n26531), .Z(n26528) );
  XOR U27100 ( .A(n26532), .B(n26529), .Z(n26530) );
  XNOR U27101 ( .A(n26533), .B(n26534), .Z(n26441) );
  ANDN U27102 ( .B(n26535), .A(n26536), .Z(n26533) );
  XOR U27103 ( .A(n26534), .B(n26537), .Z(n26535) );
  IV U27104 ( .A(n26440), .Z(n26525) );
  XOR U27105 ( .A(n26438), .B(n26538), .Z(n26440) );
  XOR U27106 ( .A(n26539), .B(n26540), .Z(n26538) );
  ANDN U27107 ( .B(n26541), .A(n26542), .Z(n26539) );
  XOR U27108 ( .A(n26543), .B(n26540), .Z(n26541) );
  IV U27109 ( .A(n26442), .Z(n26438) );
  XOR U27110 ( .A(n26544), .B(n26545), .Z(n26442) );
  ANDN U27111 ( .B(n26546), .A(n26547), .Z(n26544) );
  XOR U27112 ( .A(n26548), .B(n26545), .Z(n26546) );
  IV U27113 ( .A(n26452), .Z(n26456) );
  XOR U27114 ( .A(n26452), .B(n26355), .Z(n26454) );
  XOR U27115 ( .A(n26549), .B(n26550), .Z(n26355) );
  AND U27116 ( .A(n300), .B(n26551), .Z(n26549) );
  XOR U27117 ( .A(n26552), .B(n26550), .Z(n26551) );
  NANDN U27118 ( .A(n26357), .B(n26359), .Z(n26452) );
  XOR U27119 ( .A(n26553), .B(n26554), .Z(n26359) );
  AND U27120 ( .A(n300), .B(n26555), .Z(n26553) );
  XOR U27121 ( .A(n26554), .B(n26556), .Z(n26555) );
  XNOR U27122 ( .A(n26557), .B(n26558), .Z(n300) );
  AND U27123 ( .A(n26559), .B(n26560), .Z(n26557) );
  XOR U27124 ( .A(n26558), .B(n26370), .Z(n26560) );
  XNOR U27125 ( .A(n26561), .B(n26562), .Z(n26370) );
  ANDN U27126 ( .B(n26563), .A(n26564), .Z(n26561) );
  XOR U27127 ( .A(n26562), .B(n26565), .Z(n26563) );
  XNOR U27128 ( .A(n26558), .B(n26372), .Z(n26559) );
  XOR U27129 ( .A(n26566), .B(n26567), .Z(n26372) );
  AND U27130 ( .A(n304), .B(n26568), .Z(n26566) );
  XOR U27131 ( .A(n26569), .B(n26567), .Z(n26568) );
  XOR U27132 ( .A(n26570), .B(n26571), .Z(n26558) );
  AND U27133 ( .A(n26572), .B(n26573), .Z(n26570) );
  XOR U27134 ( .A(n26571), .B(n26397), .Z(n26573) );
  XOR U27135 ( .A(n26564), .B(n26565), .Z(n26397) );
  XNOR U27136 ( .A(n26574), .B(n26575), .Z(n26565) );
  ANDN U27137 ( .B(n26576), .A(n26577), .Z(n26574) );
  XOR U27138 ( .A(n26578), .B(n26579), .Z(n26576) );
  XOR U27139 ( .A(n26580), .B(n26581), .Z(n26564) );
  XNOR U27140 ( .A(n26582), .B(n26583), .Z(n26581) );
  ANDN U27141 ( .B(n26584), .A(n26585), .Z(n26582) );
  XNOR U27142 ( .A(n26586), .B(n26587), .Z(n26584) );
  IV U27143 ( .A(n26562), .Z(n26580) );
  XOR U27144 ( .A(n26588), .B(n26589), .Z(n26562) );
  ANDN U27145 ( .B(n26590), .A(n26591), .Z(n26588) );
  XOR U27146 ( .A(n26589), .B(n26592), .Z(n26590) );
  XNOR U27147 ( .A(n26571), .B(n26399), .Z(n26572) );
  XOR U27148 ( .A(n26593), .B(n26594), .Z(n26399) );
  AND U27149 ( .A(n304), .B(n26595), .Z(n26593) );
  XOR U27150 ( .A(n26596), .B(n26594), .Z(n26595) );
  XNOR U27151 ( .A(n26597), .B(n26598), .Z(n26571) );
  AND U27152 ( .A(n26599), .B(n26600), .Z(n26597) );
  XNOR U27153 ( .A(n26598), .B(n26449), .Z(n26600) );
  XOR U27154 ( .A(n26591), .B(n26592), .Z(n26449) );
  XOR U27155 ( .A(n26601), .B(n26579), .Z(n26592) );
  XNOR U27156 ( .A(n26602), .B(n26603), .Z(n26579) );
  ANDN U27157 ( .B(n26604), .A(n26605), .Z(n26602) );
  XOR U27158 ( .A(n26606), .B(n26607), .Z(n26604) );
  IV U27159 ( .A(n26577), .Z(n26601) );
  XOR U27160 ( .A(n26575), .B(n26608), .Z(n26577) );
  XNOR U27161 ( .A(n26609), .B(n26610), .Z(n26608) );
  ANDN U27162 ( .B(n26611), .A(n26612), .Z(n26609) );
  XNOR U27163 ( .A(n26613), .B(n26614), .Z(n26611) );
  IV U27164 ( .A(n26578), .Z(n26575) );
  XOR U27165 ( .A(n26615), .B(n26616), .Z(n26578) );
  ANDN U27166 ( .B(n26617), .A(n26618), .Z(n26615) );
  XOR U27167 ( .A(n26616), .B(n26619), .Z(n26617) );
  XOR U27168 ( .A(n26620), .B(n26621), .Z(n26591) );
  XNOR U27169 ( .A(n26586), .B(n26622), .Z(n26621) );
  IV U27170 ( .A(n26589), .Z(n26622) );
  XOR U27171 ( .A(n26623), .B(n26624), .Z(n26589) );
  ANDN U27172 ( .B(n26625), .A(n26626), .Z(n26623) );
  XOR U27173 ( .A(n26624), .B(n26627), .Z(n26625) );
  XNOR U27174 ( .A(n26628), .B(n26629), .Z(n26586) );
  ANDN U27175 ( .B(n26630), .A(n26631), .Z(n26628) );
  XOR U27176 ( .A(n26629), .B(n26632), .Z(n26630) );
  IV U27177 ( .A(n26585), .Z(n26620) );
  XOR U27178 ( .A(n26583), .B(n26633), .Z(n26585) );
  XNOR U27179 ( .A(n26634), .B(n26635), .Z(n26633) );
  ANDN U27180 ( .B(n26636), .A(n26637), .Z(n26634) );
  XNOR U27181 ( .A(n26638), .B(n26639), .Z(n26636) );
  IV U27182 ( .A(n26587), .Z(n26583) );
  XOR U27183 ( .A(n26640), .B(n26641), .Z(n26587) );
  ANDN U27184 ( .B(n26642), .A(n26643), .Z(n26640) );
  XOR U27185 ( .A(n26644), .B(n26641), .Z(n26642) );
  XOR U27186 ( .A(n26598), .B(n26451), .Z(n26599) );
  XOR U27187 ( .A(n26645), .B(n26646), .Z(n26451) );
  AND U27188 ( .A(n304), .B(n26647), .Z(n26645) );
  XOR U27189 ( .A(n26648), .B(n26646), .Z(n26647) );
  XNOR U27190 ( .A(n26649), .B(n26650), .Z(n26598) );
  NAND U27191 ( .A(n26651), .B(n26652), .Z(n26650) );
  XOR U27192 ( .A(n26653), .B(n26550), .Z(n26652) );
  XOR U27193 ( .A(n26626), .B(n26627), .Z(n26550) );
  XOR U27194 ( .A(n26654), .B(n26619), .Z(n26627) );
  XOR U27195 ( .A(n26655), .B(n26607), .Z(n26619) );
  XOR U27196 ( .A(n26656), .B(n26657), .Z(n26607) );
  ANDN U27197 ( .B(n26658), .A(n26659), .Z(n26656) );
  XOR U27198 ( .A(n26657), .B(n26660), .Z(n26658) );
  IV U27199 ( .A(n26605), .Z(n26655) );
  XOR U27200 ( .A(n26603), .B(n26661), .Z(n26605) );
  XOR U27201 ( .A(n26662), .B(n26663), .Z(n26661) );
  ANDN U27202 ( .B(n26664), .A(n26665), .Z(n26662) );
  XOR U27203 ( .A(n26666), .B(n26663), .Z(n26664) );
  IV U27204 ( .A(n26606), .Z(n26603) );
  XOR U27205 ( .A(n26667), .B(n26668), .Z(n26606) );
  ANDN U27206 ( .B(n26669), .A(n26670), .Z(n26667) );
  XOR U27207 ( .A(n26668), .B(n26671), .Z(n26669) );
  IV U27208 ( .A(n26618), .Z(n26654) );
  XOR U27209 ( .A(n26672), .B(n26673), .Z(n26618) );
  XNOR U27210 ( .A(n26613), .B(n26674), .Z(n26673) );
  IV U27211 ( .A(n26616), .Z(n26674) );
  XOR U27212 ( .A(n26675), .B(n26676), .Z(n26616) );
  ANDN U27213 ( .B(n26677), .A(n26678), .Z(n26675) );
  XOR U27214 ( .A(n26676), .B(n26679), .Z(n26677) );
  XNOR U27215 ( .A(n26680), .B(n26681), .Z(n26613) );
  ANDN U27216 ( .B(n26682), .A(n26683), .Z(n26680) );
  XOR U27217 ( .A(n26681), .B(n26684), .Z(n26682) );
  IV U27218 ( .A(n26612), .Z(n26672) );
  XOR U27219 ( .A(n26610), .B(n26685), .Z(n26612) );
  XOR U27220 ( .A(n26686), .B(n26687), .Z(n26685) );
  ANDN U27221 ( .B(n26688), .A(n26689), .Z(n26686) );
  XOR U27222 ( .A(n26690), .B(n26687), .Z(n26688) );
  IV U27223 ( .A(n26614), .Z(n26610) );
  XOR U27224 ( .A(n26691), .B(n26692), .Z(n26614) );
  ANDN U27225 ( .B(n26693), .A(n26694), .Z(n26691) );
  XOR U27226 ( .A(n26695), .B(n26692), .Z(n26693) );
  XOR U27227 ( .A(n26696), .B(n26697), .Z(n26626) );
  XOR U27228 ( .A(n26644), .B(n26698), .Z(n26697) );
  IV U27229 ( .A(n26624), .Z(n26698) );
  XOR U27230 ( .A(n26699), .B(n26700), .Z(n26624) );
  ANDN U27231 ( .B(n26701), .A(n26702), .Z(n26699) );
  XOR U27232 ( .A(n26700), .B(n26703), .Z(n26701) );
  XOR U27233 ( .A(n26704), .B(n26632), .Z(n26644) );
  XOR U27234 ( .A(n26705), .B(n26706), .Z(n26632) );
  ANDN U27235 ( .B(n26707), .A(n26708), .Z(n26705) );
  XOR U27236 ( .A(n26706), .B(n26709), .Z(n26707) );
  IV U27237 ( .A(n26631), .Z(n26704) );
  XOR U27238 ( .A(n26710), .B(n26711), .Z(n26631) );
  XOR U27239 ( .A(n26712), .B(n26713), .Z(n26711) );
  ANDN U27240 ( .B(n26714), .A(n26715), .Z(n26712) );
  XOR U27241 ( .A(n26716), .B(n26713), .Z(n26714) );
  IV U27242 ( .A(n26629), .Z(n26710) );
  XOR U27243 ( .A(n26717), .B(n26718), .Z(n26629) );
  ANDN U27244 ( .B(n26719), .A(n26720), .Z(n26717) );
  XOR U27245 ( .A(n26718), .B(n26721), .Z(n26719) );
  IV U27246 ( .A(n26643), .Z(n26696) );
  XOR U27247 ( .A(n26722), .B(n26723), .Z(n26643) );
  XNOR U27248 ( .A(n26638), .B(n26724), .Z(n26723) );
  IV U27249 ( .A(n26641), .Z(n26724) );
  XOR U27250 ( .A(n26725), .B(n26726), .Z(n26641) );
  ANDN U27251 ( .B(n26727), .A(n26728), .Z(n26725) );
  XOR U27252 ( .A(n26729), .B(n26726), .Z(n26727) );
  XNOR U27253 ( .A(n26730), .B(n26731), .Z(n26638) );
  ANDN U27254 ( .B(n26732), .A(n26733), .Z(n26730) );
  XOR U27255 ( .A(n26731), .B(n26734), .Z(n26732) );
  IV U27256 ( .A(n26637), .Z(n26722) );
  XOR U27257 ( .A(n26635), .B(n26735), .Z(n26637) );
  XOR U27258 ( .A(n26736), .B(n26737), .Z(n26735) );
  ANDN U27259 ( .B(n26738), .A(n26739), .Z(n26736) );
  XOR U27260 ( .A(n26740), .B(n26737), .Z(n26738) );
  IV U27261 ( .A(n26639), .Z(n26635) );
  XOR U27262 ( .A(n26741), .B(n26742), .Z(n26639) );
  ANDN U27263 ( .B(n26743), .A(n26744), .Z(n26741) );
  XOR U27264 ( .A(n26745), .B(n26742), .Z(n26743) );
  IV U27265 ( .A(n26649), .Z(n26653) );
  XOR U27266 ( .A(n26649), .B(n26552), .Z(n26651) );
  XOR U27267 ( .A(n26746), .B(n26747), .Z(n26552) );
  AND U27268 ( .A(n304), .B(n26748), .Z(n26746) );
  XOR U27269 ( .A(n26749), .B(n26747), .Z(n26748) );
  NANDN U27270 ( .A(n26554), .B(n26556), .Z(n26649) );
  XOR U27271 ( .A(n26750), .B(n26751), .Z(n26556) );
  AND U27272 ( .A(n304), .B(n26752), .Z(n26750) );
  XOR U27273 ( .A(n26751), .B(n26753), .Z(n26752) );
  XNOR U27274 ( .A(n26754), .B(n26755), .Z(n304) );
  AND U27275 ( .A(n26756), .B(n26757), .Z(n26754) );
  XOR U27276 ( .A(n26755), .B(n26567), .Z(n26757) );
  XNOR U27277 ( .A(n26758), .B(n26759), .Z(n26567) );
  ANDN U27278 ( .B(n26760), .A(n26761), .Z(n26758) );
  XOR U27279 ( .A(n26759), .B(n26762), .Z(n26760) );
  XNOR U27280 ( .A(n26755), .B(n26569), .Z(n26756) );
  XOR U27281 ( .A(n26763), .B(n26764), .Z(n26569) );
  AND U27282 ( .A(n308), .B(n26765), .Z(n26763) );
  XOR U27283 ( .A(n26766), .B(n26764), .Z(n26765) );
  XOR U27284 ( .A(n26767), .B(n26768), .Z(n26755) );
  AND U27285 ( .A(n26769), .B(n26770), .Z(n26767) );
  XOR U27286 ( .A(n26768), .B(n26594), .Z(n26770) );
  XOR U27287 ( .A(n26761), .B(n26762), .Z(n26594) );
  XNOR U27288 ( .A(n26771), .B(n26772), .Z(n26762) );
  ANDN U27289 ( .B(n26773), .A(n26774), .Z(n26771) );
  XOR U27290 ( .A(n26775), .B(n26776), .Z(n26773) );
  XOR U27291 ( .A(n26777), .B(n26778), .Z(n26761) );
  XNOR U27292 ( .A(n26779), .B(n26780), .Z(n26778) );
  ANDN U27293 ( .B(n26781), .A(n26782), .Z(n26779) );
  XNOR U27294 ( .A(n26783), .B(n26784), .Z(n26781) );
  IV U27295 ( .A(n26759), .Z(n26777) );
  XOR U27296 ( .A(n26785), .B(n26786), .Z(n26759) );
  ANDN U27297 ( .B(n26787), .A(n26788), .Z(n26785) );
  XOR U27298 ( .A(n26786), .B(n26789), .Z(n26787) );
  XNOR U27299 ( .A(n26768), .B(n26596), .Z(n26769) );
  XOR U27300 ( .A(n26790), .B(n26791), .Z(n26596) );
  AND U27301 ( .A(n308), .B(n26792), .Z(n26790) );
  XOR U27302 ( .A(n26793), .B(n26791), .Z(n26792) );
  XNOR U27303 ( .A(n26794), .B(n26795), .Z(n26768) );
  AND U27304 ( .A(n26796), .B(n26797), .Z(n26794) );
  XNOR U27305 ( .A(n26795), .B(n26646), .Z(n26797) );
  XOR U27306 ( .A(n26788), .B(n26789), .Z(n26646) );
  XOR U27307 ( .A(n26798), .B(n26776), .Z(n26789) );
  XNOR U27308 ( .A(n26799), .B(n26800), .Z(n26776) );
  ANDN U27309 ( .B(n26801), .A(n26802), .Z(n26799) );
  XOR U27310 ( .A(n26803), .B(n26804), .Z(n26801) );
  IV U27311 ( .A(n26774), .Z(n26798) );
  XOR U27312 ( .A(n26772), .B(n26805), .Z(n26774) );
  XNOR U27313 ( .A(n26806), .B(n26807), .Z(n26805) );
  ANDN U27314 ( .B(n26808), .A(n26809), .Z(n26806) );
  XNOR U27315 ( .A(n26810), .B(n26811), .Z(n26808) );
  IV U27316 ( .A(n26775), .Z(n26772) );
  XOR U27317 ( .A(n26812), .B(n26813), .Z(n26775) );
  ANDN U27318 ( .B(n26814), .A(n26815), .Z(n26812) );
  XOR U27319 ( .A(n26813), .B(n26816), .Z(n26814) );
  XOR U27320 ( .A(n26817), .B(n26818), .Z(n26788) );
  XNOR U27321 ( .A(n26783), .B(n26819), .Z(n26818) );
  IV U27322 ( .A(n26786), .Z(n26819) );
  XOR U27323 ( .A(n26820), .B(n26821), .Z(n26786) );
  ANDN U27324 ( .B(n26822), .A(n26823), .Z(n26820) );
  XOR U27325 ( .A(n26821), .B(n26824), .Z(n26822) );
  XNOR U27326 ( .A(n26825), .B(n26826), .Z(n26783) );
  ANDN U27327 ( .B(n26827), .A(n26828), .Z(n26825) );
  XOR U27328 ( .A(n26826), .B(n26829), .Z(n26827) );
  IV U27329 ( .A(n26782), .Z(n26817) );
  XOR U27330 ( .A(n26780), .B(n26830), .Z(n26782) );
  XNOR U27331 ( .A(n26831), .B(n26832), .Z(n26830) );
  ANDN U27332 ( .B(n26833), .A(n26834), .Z(n26831) );
  XNOR U27333 ( .A(n26835), .B(n26836), .Z(n26833) );
  IV U27334 ( .A(n26784), .Z(n26780) );
  XOR U27335 ( .A(n26837), .B(n26838), .Z(n26784) );
  ANDN U27336 ( .B(n26839), .A(n26840), .Z(n26837) );
  XOR U27337 ( .A(n26841), .B(n26838), .Z(n26839) );
  XOR U27338 ( .A(n26795), .B(n26648), .Z(n26796) );
  XOR U27339 ( .A(n26842), .B(n26843), .Z(n26648) );
  AND U27340 ( .A(n308), .B(n26844), .Z(n26842) );
  XOR U27341 ( .A(n26845), .B(n26843), .Z(n26844) );
  XNOR U27342 ( .A(n26846), .B(n26847), .Z(n26795) );
  NAND U27343 ( .A(n26848), .B(n26849), .Z(n26847) );
  XOR U27344 ( .A(n26850), .B(n26747), .Z(n26849) );
  XOR U27345 ( .A(n26823), .B(n26824), .Z(n26747) );
  XOR U27346 ( .A(n26851), .B(n26816), .Z(n26824) );
  XOR U27347 ( .A(n26852), .B(n26804), .Z(n26816) );
  XOR U27348 ( .A(n26853), .B(n26854), .Z(n26804) );
  ANDN U27349 ( .B(n26855), .A(n26856), .Z(n26853) );
  XOR U27350 ( .A(n26854), .B(n26857), .Z(n26855) );
  IV U27351 ( .A(n26802), .Z(n26852) );
  XOR U27352 ( .A(n26800), .B(n26858), .Z(n26802) );
  XOR U27353 ( .A(n26859), .B(n26860), .Z(n26858) );
  ANDN U27354 ( .B(n26861), .A(n26862), .Z(n26859) );
  XOR U27355 ( .A(n26863), .B(n26860), .Z(n26861) );
  IV U27356 ( .A(n26803), .Z(n26800) );
  XOR U27357 ( .A(n26864), .B(n26865), .Z(n26803) );
  ANDN U27358 ( .B(n26866), .A(n26867), .Z(n26864) );
  XOR U27359 ( .A(n26865), .B(n26868), .Z(n26866) );
  IV U27360 ( .A(n26815), .Z(n26851) );
  XOR U27361 ( .A(n26869), .B(n26870), .Z(n26815) );
  XNOR U27362 ( .A(n26810), .B(n26871), .Z(n26870) );
  IV U27363 ( .A(n26813), .Z(n26871) );
  XOR U27364 ( .A(n26872), .B(n26873), .Z(n26813) );
  ANDN U27365 ( .B(n26874), .A(n26875), .Z(n26872) );
  XOR U27366 ( .A(n26873), .B(n26876), .Z(n26874) );
  XNOR U27367 ( .A(n26877), .B(n26878), .Z(n26810) );
  ANDN U27368 ( .B(n26879), .A(n26880), .Z(n26877) );
  XOR U27369 ( .A(n26878), .B(n26881), .Z(n26879) );
  IV U27370 ( .A(n26809), .Z(n26869) );
  XOR U27371 ( .A(n26807), .B(n26882), .Z(n26809) );
  XOR U27372 ( .A(n26883), .B(n26884), .Z(n26882) );
  ANDN U27373 ( .B(n26885), .A(n26886), .Z(n26883) );
  XOR U27374 ( .A(n26887), .B(n26884), .Z(n26885) );
  IV U27375 ( .A(n26811), .Z(n26807) );
  XOR U27376 ( .A(n26888), .B(n26889), .Z(n26811) );
  ANDN U27377 ( .B(n26890), .A(n26891), .Z(n26888) );
  XOR U27378 ( .A(n26892), .B(n26889), .Z(n26890) );
  XOR U27379 ( .A(n26893), .B(n26894), .Z(n26823) );
  XOR U27380 ( .A(n26841), .B(n26895), .Z(n26894) );
  IV U27381 ( .A(n26821), .Z(n26895) );
  XOR U27382 ( .A(n26896), .B(n26897), .Z(n26821) );
  ANDN U27383 ( .B(n26898), .A(n26899), .Z(n26896) );
  XOR U27384 ( .A(n26897), .B(n26900), .Z(n26898) );
  XOR U27385 ( .A(n26901), .B(n26829), .Z(n26841) );
  XOR U27386 ( .A(n26902), .B(n26903), .Z(n26829) );
  ANDN U27387 ( .B(n26904), .A(n26905), .Z(n26902) );
  XOR U27388 ( .A(n26903), .B(n26906), .Z(n26904) );
  IV U27389 ( .A(n26828), .Z(n26901) );
  XOR U27390 ( .A(n26907), .B(n26908), .Z(n26828) );
  XOR U27391 ( .A(n26909), .B(n26910), .Z(n26908) );
  ANDN U27392 ( .B(n26911), .A(n26912), .Z(n26909) );
  XOR U27393 ( .A(n26913), .B(n26910), .Z(n26911) );
  IV U27394 ( .A(n26826), .Z(n26907) );
  XOR U27395 ( .A(n26914), .B(n26915), .Z(n26826) );
  ANDN U27396 ( .B(n26916), .A(n26917), .Z(n26914) );
  XOR U27397 ( .A(n26915), .B(n26918), .Z(n26916) );
  IV U27398 ( .A(n26840), .Z(n26893) );
  XOR U27399 ( .A(n26919), .B(n26920), .Z(n26840) );
  XNOR U27400 ( .A(n26835), .B(n26921), .Z(n26920) );
  IV U27401 ( .A(n26838), .Z(n26921) );
  XOR U27402 ( .A(n26922), .B(n26923), .Z(n26838) );
  ANDN U27403 ( .B(n26924), .A(n26925), .Z(n26922) );
  XOR U27404 ( .A(n26926), .B(n26923), .Z(n26924) );
  XNOR U27405 ( .A(n26927), .B(n26928), .Z(n26835) );
  ANDN U27406 ( .B(n26929), .A(n26930), .Z(n26927) );
  XOR U27407 ( .A(n26928), .B(n26931), .Z(n26929) );
  IV U27408 ( .A(n26834), .Z(n26919) );
  XOR U27409 ( .A(n26832), .B(n26932), .Z(n26834) );
  XOR U27410 ( .A(n26933), .B(n26934), .Z(n26932) );
  ANDN U27411 ( .B(n26935), .A(n26936), .Z(n26933) );
  XOR U27412 ( .A(n26937), .B(n26934), .Z(n26935) );
  IV U27413 ( .A(n26836), .Z(n26832) );
  XOR U27414 ( .A(n26938), .B(n26939), .Z(n26836) );
  ANDN U27415 ( .B(n26940), .A(n26941), .Z(n26938) );
  XOR U27416 ( .A(n26942), .B(n26939), .Z(n26940) );
  IV U27417 ( .A(n26846), .Z(n26850) );
  XOR U27418 ( .A(n26846), .B(n26749), .Z(n26848) );
  XOR U27419 ( .A(n26943), .B(n26944), .Z(n26749) );
  AND U27420 ( .A(n308), .B(n26945), .Z(n26943) );
  XOR U27421 ( .A(n26946), .B(n26944), .Z(n26945) );
  NANDN U27422 ( .A(n26751), .B(n26753), .Z(n26846) );
  XOR U27423 ( .A(n26947), .B(n26948), .Z(n26753) );
  AND U27424 ( .A(n308), .B(n26949), .Z(n26947) );
  XOR U27425 ( .A(n26948), .B(n26950), .Z(n26949) );
  XNOR U27426 ( .A(n26951), .B(n26952), .Z(n308) );
  AND U27427 ( .A(n26953), .B(n26954), .Z(n26951) );
  XOR U27428 ( .A(n26952), .B(n26764), .Z(n26954) );
  XNOR U27429 ( .A(n26955), .B(n26956), .Z(n26764) );
  ANDN U27430 ( .B(n26957), .A(n26958), .Z(n26955) );
  XOR U27431 ( .A(n26956), .B(n26959), .Z(n26957) );
  XNOR U27432 ( .A(n26952), .B(n26766), .Z(n26953) );
  XOR U27433 ( .A(n26960), .B(n26961), .Z(n26766) );
  AND U27434 ( .A(n312), .B(n26962), .Z(n26960) );
  XOR U27435 ( .A(n26963), .B(n26961), .Z(n26962) );
  XOR U27436 ( .A(n26964), .B(n26965), .Z(n26952) );
  AND U27437 ( .A(n26966), .B(n26967), .Z(n26964) );
  XOR U27438 ( .A(n26965), .B(n26791), .Z(n26967) );
  XOR U27439 ( .A(n26958), .B(n26959), .Z(n26791) );
  XNOR U27440 ( .A(n26968), .B(n26969), .Z(n26959) );
  ANDN U27441 ( .B(n26970), .A(n26971), .Z(n26968) );
  XOR U27442 ( .A(n26972), .B(n26973), .Z(n26970) );
  XOR U27443 ( .A(n26974), .B(n26975), .Z(n26958) );
  XNOR U27444 ( .A(n26976), .B(n26977), .Z(n26975) );
  ANDN U27445 ( .B(n26978), .A(n26979), .Z(n26976) );
  XNOR U27446 ( .A(n26980), .B(n26981), .Z(n26978) );
  IV U27447 ( .A(n26956), .Z(n26974) );
  XOR U27448 ( .A(n26982), .B(n26983), .Z(n26956) );
  ANDN U27449 ( .B(n26984), .A(n26985), .Z(n26982) );
  XOR U27450 ( .A(n26983), .B(n26986), .Z(n26984) );
  XNOR U27451 ( .A(n26965), .B(n26793), .Z(n26966) );
  XOR U27452 ( .A(n26987), .B(n26988), .Z(n26793) );
  AND U27453 ( .A(n312), .B(n26989), .Z(n26987) );
  XOR U27454 ( .A(n26990), .B(n26988), .Z(n26989) );
  XNOR U27455 ( .A(n26991), .B(n26992), .Z(n26965) );
  AND U27456 ( .A(n26993), .B(n26994), .Z(n26991) );
  XNOR U27457 ( .A(n26992), .B(n26843), .Z(n26994) );
  XOR U27458 ( .A(n26985), .B(n26986), .Z(n26843) );
  XOR U27459 ( .A(n26995), .B(n26973), .Z(n26986) );
  XNOR U27460 ( .A(n26996), .B(n26997), .Z(n26973) );
  ANDN U27461 ( .B(n26998), .A(n26999), .Z(n26996) );
  XOR U27462 ( .A(n27000), .B(n27001), .Z(n26998) );
  IV U27463 ( .A(n26971), .Z(n26995) );
  XOR U27464 ( .A(n26969), .B(n27002), .Z(n26971) );
  XNOR U27465 ( .A(n27003), .B(n27004), .Z(n27002) );
  ANDN U27466 ( .B(n27005), .A(n27006), .Z(n27003) );
  XNOR U27467 ( .A(n27007), .B(n27008), .Z(n27005) );
  IV U27468 ( .A(n26972), .Z(n26969) );
  XOR U27469 ( .A(n27009), .B(n27010), .Z(n26972) );
  ANDN U27470 ( .B(n27011), .A(n27012), .Z(n27009) );
  XOR U27471 ( .A(n27010), .B(n27013), .Z(n27011) );
  XOR U27472 ( .A(n27014), .B(n27015), .Z(n26985) );
  XNOR U27473 ( .A(n26980), .B(n27016), .Z(n27015) );
  IV U27474 ( .A(n26983), .Z(n27016) );
  XOR U27475 ( .A(n27017), .B(n27018), .Z(n26983) );
  ANDN U27476 ( .B(n27019), .A(n27020), .Z(n27017) );
  XOR U27477 ( .A(n27018), .B(n27021), .Z(n27019) );
  XNOR U27478 ( .A(n27022), .B(n27023), .Z(n26980) );
  ANDN U27479 ( .B(n27024), .A(n27025), .Z(n27022) );
  XOR U27480 ( .A(n27023), .B(n27026), .Z(n27024) );
  IV U27481 ( .A(n26979), .Z(n27014) );
  XOR U27482 ( .A(n26977), .B(n27027), .Z(n26979) );
  XNOR U27483 ( .A(n27028), .B(n27029), .Z(n27027) );
  ANDN U27484 ( .B(n27030), .A(n27031), .Z(n27028) );
  XNOR U27485 ( .A(n27032), .B(n27033), .Z(n27030) );
  IV U27486 ( .A(n26981), .Z(n26977) );
  XOR U27487 ( .A(n27034), .B(n27035), .Z(n26981) );
  ANDN U27488 ( .B(n27036), .A(n27037), .Z(n27034) );
  XOR U27489 ( .A(n27038), .B(n27035), .Z(n27036) );
  XOR U27490 ( .A(n26992), .B(n26845), .Z(n26993) );
  XOR U27491 ( .A(n27039), .B(n27040), .Z(n26845) );
  AND U27492 ( .A(n312), .B(n27041), .Z(n27039) );
  XOR U27493 ( .A(n27042), .B(n27040), .Z(n27041) );
  XNOR U27494 ( .A(n27043), .B(n27044), .Z(n26992) );
  NAND U27495 ( .A(n27045), .B(n27046), .Z(n27044) );
  XOR U27496 ( .A(n27047), .B(n26944), .Z(n27046) );
  XOR U27497 ( .A(n27020), .B(n27021), .Z(n26944) );
  XOR U27498 ( .A(n27048), .B(n27013), .Z(n27021) );
  XOR U27499 ( .A(n27049), .B(n27001), .Z(n27013) );
  XOR U27500 ( .A(n27050), .B(n27051), .Z(n27001) );
  ANDN U27501 ( .B(n27052), .A(n27053), .Z(n27050) );
  XOR U27502 ( .A(n27051), .B(n27054), .Z(n27052) );
  IV U27503 ( .A(n26999), .Z(n27049) );
  XOR U27504 ( .A(n26997), .B(n27055), .Z(n26999) );
  XOR U27505 ( .A(n27056), .B(n27057), .Z(n27055) );
  ANDN U27506 ( .B(n27058), .A(n27059), .Z(n27056) );
  XOR U27507 ( .A(n27060), .B(n27057), .Z(n27058) );
  IV U27508 ( .A(n27000), .Z(n26997) );
  XOR U27509 ( .A(n27061), .B(n27062), .Z(n27000) );
  ANDN U27510 ( .B(n27063), .A(n27064), .Z(n27061) );
  XOR U27511 ( .A(n27062), .B(n27065), .Z(n27063) );
  IV U27512 ( .A(n27012), .Z(n27048) );
  XOR U27513 ( .A(n27066), .B(n27067), .Z(n27012) );
  XNOR U27514 ( .A(n27007), .B(n27068), .Z(n27067) );
  IV U27515 ( .A(n27010), .Z(n27068) );
  XOR U27516 ( .A(n27069), .B(n27070), .Z(n27010) );
  ANDN U27517 ( .B(n27071), .A(n27072), .Z(n27069) );
  XOR U27518 ( .A(n27070), .B(n27073), .Z(n27071) );
  XNOR U27519 ( .A(n27074), .B(n27075), .Z(n27007) );
  ANDN U27520 ( .B(n27076), .A(n27077), .Z(n27074) );
  XOR U27521 ( .A(n27075), .B(n27078), .Z(n27076) );
  IV U27522 ( .A(n27006), .Z(n27066) );
  XOR U27523 ( .A(n27004), .B(n27079), .Z(n27006) );
  XOR U27524 ( .A(n27080), .B(n27081), .Z(n27079) );
  ANDN U27525 ( .B(n27082), .A(n27083), .Z(n27080) );
  XOR U27526 ( .A(n27084), .B(n27081), .Z(n27082) );
  IV U27527 ( .A(n27008), .Z(n27004) );
  XOR U27528 ( .A(n27085), .B(n27086), .Z(n27008) );
  ANDN U27529 ( .B(n27087), .A(n27088), .Z(n27085) );
  XOR U27530 ( .A(n27089), .B(n27086), .Z(n27087) );
  XOR U27531 ( .A(n27090), .B(n27091), .Z(n27020) );
  XOR U27532 ( .A(n27038), .B(n27092), .Z(n27091) );
  IV U27533 ( .A(n27018), .Z(n27092) );
  XOR U27534 ( .A(n27093), .B(n27094), .Z(n27018) );
  ANDN U27535 ( .B(n27095), .A(n27096), .Z(n27093) );
  XOR U27536 ( .A(n27094), .B(n27097), .Z(n27095) );
  XOR U27537 ( .A(n27098), .B(n27026), .Z(n27038) );
  XOR U27538 ( .A(n27099), .B(n27100), .Z(n27026) );
  ANDN U27539 ( .B(n27101), .A(n27102), .Z(n27099) );
  XOR U27540 ( .A(n27100), .B(n27103), .Z(n27101) );
  IV U27541 ( .A(n27025), .Z(n27098) );
  XOR U27542 ( .A(n27104), .B(n27105), .Z(n27025) );
  XOR U27543 ( .A(n27106), .B(n27107), .Z(n27105) );
  ANDN U27544 ( .B(n27108), .A(n27109), .Z(n27106) );
  XOR U27545 ( .A(n27110), .B(n27107), .Z(n27108) );
  IV U27546 ( .A(n27023), .Z(n27104) );
  XOR U27547 ( .A(n27111), .B(n27112), .Z(n27023) );
  ANDN U27548 ( .B(n27113), .A(n27114), .Z(n27111) );
  XOR U27549 ( .A(n27112), .B(n27115), .Z(n27113) );
  IV U27550 ( .A(n27037), .Z(n27090) );
  XOR U27551 ( .A(n27116), .B(n27117), .Z(n27037) );
  XNOR U27552 ( .A(n27032), .B(n27118), .Z(n27117) );
  IV U27553 ( .A(n27035), .Z(n27118) );
  XOR U27554 ( .A(n27119), .B(n27120), .Z(n27035) );
  ANDN U27555 ( .B(n27121), .A(n27122), .Z(n27119) );
  XOR U27556 ( .A(n27123), .B(n27120), .Z(n27121) );
  XNOR U27557 ( .A(n27124), .B(n27125), .Z(n27032) );
  ANDN U27558 ( .B(n27126), .A(n27127), .Z(n27124) );
  XOR U27559 ( .A(n27125), .B(n27128), .Z(n27126) );
  IV U27560 ( .A(n27031), .Z(n27116) );
  XOR U27561 ( .A(n27029), .B(n27129), .Z(n27031) );
  XOR U27562 ( .A(n27130), .B(n27131), .Z(n27129) );
  ANDN U27563 ( .B(n27132), .A(n27133), .Z(n27130) );
  XOR U27564 ( .A(n27134), .B(n27131), .Z(n27132) );
  IV U27565 ( .A(n27033), .Z(n27029) );
  XOR U27566 ( .A(n27135), .B(n27136), .Z(n27033) );
  ANDN U27567 ( .B(n27137), .A(n27138), .Z(n27135) );
  XOR U27568 ( .A(n27139), .B(n27136), .Z(n27137) );
  IV U27569 ( .A(n27043), .Z(n27047) );
  XOR U27570 ( .A(n27043), .B(n26946), .Z(n27045) );
  XOR U27571 ( .A(n27140), .B(n27141), .Z(n26946) );
  AND U27572 ( .A(n312), .B(n27142), .Z(n27140) );
  XOR U27573 ( .A(n27143), .B(n27141), .Z(n27142) );
  NANDN U27574 ( .A(n26948), .B(n26950), .Z(n27043) );
  XOR U27575 ( .A(n27144), .B(n27145), .Z(n26950) );
  AND U27576 ( .A(n312), .B(n27146), .Z(n27144) );
  XOR U27577 ( .A(n27145), .B(n27147), .Z(n27146) );
  XNOR U27578 ( .A(n27148), .B(n27149), .Z(n312) );
  AND U27579 ( .A(n27150), .B(n27151), .Z(n27148) );
  XOR U27580 ( .A(n27149), .B(n26961), .Z(n27151) );
  XNOR U27581 ( .A(n27152), .B(n27153), .Z(n26961) );
  ANDN U27582 ( .B(n27154), .A(n27155), .Z(n27152) );
  XOR U27583 ( .A(n27153), .B(n27156), .Z(n27154) );
  XNOR U27584 ( .A(n27149), .B(n26963), .Z(n27150) );
  XOR U27585 ( .A(n27157), .B(n27158), .Z(n26963) );
  AND U27586 ( .A(n316), .B(n27159), .Z(n27157) );
  XOR U27587 ( .A(n27160), .B(n27158), .Z(n27159) );
  XOR U27588 ( .A(n27161), .B(n27162), .Z(n27149) );
  AND U27589 ( .A(n27163), .B(n27164), .Z(n27161) );
  XOR U27590 ( .A(n27162), .B(n26988), .Z(n27164) );
  XOR U27591 ( .A(n27155), .B(n27156), .Z(n26988) );
  XNOR U27592 ( .A(n27165), .B(n27166), .Z(n27156) );
  ANDN U27593 ( .B(n27167), .A(n27168), .Z(n27165) );
  XOR U27594 ( .A(n27169), .B(n27170), .Z(n27167) );
  XOR U27595 ( .A(n27171), .B(n27172), .Z(n27155) );
  XNOR U27596 ( .A(n27173), .B(n27174), .Z(n27172) );
  ANDN U27597 ( .B(n27175), .A(n27176), .Z(n27173) );
  XNOR U27598 ( .A(n27177), .B(n27178), .Z(n27175) );
  IV U27599 ( .A(n27153), .Z(n27171) );
  XOR U27600 ( .A(n27179), .B(n27180), .Z(n27153) );
  ANDN U27601 ( .B(n27181), .A(n27182), .Z(n27179) );
  XOR U27602 ( .A(n27180), .B(n27183), .Z(n27181) );
  XNOR U27603 ( .A(n27162), .B(n26990), .Z(n27163) );
  XOR U27604 ( .A(n27184), .B(n27185), .Z(n26990) );
  AND U27605 ( .A(n316), .B(n27186), .Z(n27184) );
  XOR U27606 ( .A(n27187), .B(n27185), .Z(n27186) );
  XNOR U27607 ( .A(n27188), .B(n27189), .Z(n27162) );
  AND U27608 ( .A(n27190), .B(n27191), .Z(n27188) );
  XNOR U27609 ( .A(n27189), .B(n27040), .Z(n27191) );
  XOR U27610 ( .A(n27182), .B(n27183), .Z(n27040) );
  XOR U27611 ( .A(n27192), .B(n27170), .Z(n27183) );
  XNOR U27612 ( .A(n27193), .B(n27194), .Z(n27170) );
  ANDN U27613 ( .B(n27195), .A(n27196), .Z(n27193) );
  XOR U27614 ( .A(n27197), .B(n27198), .Z(n27195) );
  IV U27615 ( .A(n27168), .Z(n27192) );
  XOR U27616 ( .A(n27166), .B(n27199), .Z(n27168) );
  XNOR U27617 ( .A(n27200), .B(n27201), .Z(n27199) );
  ANDN U27618 ( .B(n27202), .A(n27203), .Z(n27200) );
  XNOR U27619 ( .A(n27204), .B(n27205), .Z(n27202) );
  IV U27620 ( .A(n27169), .Z(n27166) );
  XOR U27621 ( .A(n27206), .B(n27207), .Z(n27169) );
  ANDN U27622 ( .B(n27208), .A(n27209), .Z(n27206) );
  XOR U27623 ( .A(n27207), .B(n27210), .Z(n27208) );
  XOR U27624 ( .A(n27211), .B(n27212), .Z(n27182) );
  XNOR U27625 ( .A(n27177), .B(n27213), .Z(n27212) );
  IV U27626 ( .A(n27180), .Z(n27213) );
  XOR U27627 ( .A(n27214), .B(n27215), .Z(n27180) );
  ANDN U27628 ( .B(n27216), .A(n27217), .Z(n27214) );
  XOR U27629 ( .A(n27215), .B(n27218), .Z(n27216) );
  XNOR U27630 ( .A(n27219), .B(n27220), .Z(n27177) );
  ANDN U27631 ( .B(n27221), .A(n27222), .Z(n27219) );
  XOR U27632 ( .A(n27220), .B(n27223), .Z(n27221) );
  IV U27633 ( .A(n27176), .Z(n27211) );
  XOR U27634 ( .A(n27174), .B(n27224), .Z(n27176) );
  XNOR U27635 ( .A(n27225), .B(n27226), .Z(n27224) );
  ANDN U27636 ( .B(n27227), .A(n27228), .Z(n27225) );
  XNOR U27637 ( .A(n27229), .B(n27230), .Z(n27227) );
  IV U27638 ( .A(n27178), .Z(n27174) );
  XOR U27639 ( .A(n27231), .B(n27232), .Z(n27178) );
  ANDN U27640 ( .B(n27233), .A(n27234), .Z(n27231) );
  XOR U27641 ( .A(n27235), .B(n27232), .Z(n27233) );
  XOR U27642 ( .A(n27189), .B(n27042), .Z(n27190) );
  XOR U27643 ( .A(n27236), .B(n27237), .Z(n27042) );
  AND U27644 ( .A(n316), .B(n27238), .Z(n27236) );
  XOR U27645 ( .A(n27239), .B(n27237), .Z(n27238) );
  XNOR U27646 ( .A(n27240), .B(n27241), .Z(n27189) );
  NAND U27647 ( .A(n27242), .B(n27243), .Z(n27241) );
  XOR U27648 ( .A(n27244), .B(n27141), .Z(n27243) );
  XOR U27649 ( .A(n27217), .B(n27218), .Z(n27141) );
  XOR U27650 ( .A(n27245), .B(n27210), .Z(n27218) );
  XOR U27651 ( .A(n27246), .B(n27198), .Z(n27210) );
  XOR U27652 ( .A(n27247), .B(n27248), .Z(n27198) );
  ANDN U27653 ( .B(n27249), .A(n27250), .Z(n27247) );
  XOR U27654 ( .A(n27248), .B(n27251), .Z(n27249) );
  IV U27655 ( .A(n27196), .Z(n27246) );
  XOR U27656 ( .A(n27194), .B(n27252), .Z(n27196) );
  XOR U27657 ( .A(n27253), .B(n27254), .Z(n27252) );
  ANDN U27658 ( .B(n27255), .A(n27256), .Z(n27253) );
  XOR U27659 ( .A(n27257), .B(n27254), .Z(n27255) );
  IV U27660 ( .A(n27197), .Z(n27194) );
  XOR U27661 ( .A(n27258), .B(n27259), .Z(n27197) );
  ANDN U27662 ( .B(n27260), .A(n27261), .Z(n27258) );
  XOR U27663 ( .A(n27259), .B(n27262), .Z(n27260) );
  IV U27664 ( .A(n27209), .Z(n27245) );
  XOR U27665 ( .A(n27263), .B(n27264), .Z(n27209) );
  XNOR U27666 ( .A(n27204), .B(n27265), .Z(n27264) );
  IV U27667 ( .A(n27207), .Z(n27265) );
  XOR U27668 ( .A(n27266), .B(n27267), .Z(n27207) );
  ANDN U27669 ( .B(n27268), .A(n27269), .Z(n27266) );
  XOR U27670 ( .A(n27267), .B(n27270), .Z(n27268) );
  XNOR U27671 ( .A(n27271), .B(n27272), .Z(n27204) );
  ANDN U27672 ( .B(n27273), .A(n27274), .Z(n27271) );
  XOR U27673 ( .A(n27272), .B(n27275), .Z(n27273) );
  IV U27674 ( .A(n27203), .Z(n27263) );
  XOR U27675 ( .A(n27201), .B(n27276), .Z(n27203) );
  XOR U27676 ( .A(n27277), .B(n27278), .Z(n27276) );
  ANDN U27677 ( .B(n27279), .A(n27280), .Z(n27277) );
  XOR U27678 ( .A(n27281), .B(n27278), .Z(n27279) );
  IV U27679 ( .A(n27205), .Z(n27201) );
  XOR U27680 ( .A(n27282), .B(n27283), .Z(n27205) );
  ANDN U27681 ( .B(n27284), .A(n27285), .Z(n27282) );
  XOR U27682 ( .A(n27286), .B(n27283), .Z(n27284) );
  XOR U27683 ( .A(n27287), .B(n27288), .Z(n27217) );
  XOR U27684 ( .A(n27235), .B(n27289), .Z(n27288) );
  IV U27685 ( .A(n27215), .Z(n27289) );
  XOR U27686 ( .A(n27290), .B(n27291), .Z(n27215) );
  ANDN U27687 ( .B(n27292), .A(n27293), .Z(n27290) );
  XOR U27688 ( .A(n27291), .B(n27294), .Z(n27292) );
  XOR U27689 ( .A(n27295), .B(n27223), .Z(n27235) );
  XOR U27690 ( .A(n27296), .B(n27297), .Z(n27223) );
  ANDN U27691 ( .B(n27298), .A(n27299), .Z(n27296) );
  XOR U27692 ( .A(n27297), .B(n27300), .Z(n27298) );
  IV U27693 ( .A(n27222), .Z(n27295) );
  XOR U27694 ( .A(n27301), .B(n27302), .Z(n27222) );
  XOR U27695 ( .A(n27303), .B(n27304), .Z(n27302) );
  ANDN U27696 ( .B(n27305), .A(n27306), .Z(n27303) );
  XOR U27697 ( .A(n27307), .B(n27304), .Z(n27305) );
  IV U27698 ( .A(n27220), .Z(n27301) );
  XOR U27699 ( .A(n27308), .B(n27309), .Z(n27220) );
  ANDN U27700 ( .B(n27310), .A(n27311), .Z(n27308) );
  XOR U27701 ( .A(n27309), .B(n27312), .Z(n27310) );
  IV U27702 ( .A(n27234), .Z(n27287) );
  XOR U27703 ( .A(n27313), .B(n27314), .Z(n27234) );
  XNOR U27704 ( .A(n27229), .B(n27315), .Z(n27314) );
  IV U27705 ( .A(n27232), .Z(n27315) );
  XOR U27706 ( .A(n27316), .B(n27317), .Z(n27232) );
  ANDN U27707 ( .B(n27318), .A(n27319), .Z(n27316) );
  XOR U27708 ( .A(n27320), .B(n27317), .Z(n27318) );
  XNOR U27709 ( .A(n27321), .B(n27322), .Z(n27229) );
  ANDN U27710 ( .B(n27323), .A(n27324), .Z(n27321) );
  XOR U27711 ( .A(n27322), .B(n27325), .Z(n27323) );
  IV U27712 ( .A(n27228), .Z(n27313) );
  XOR U27713 ( .A(n27226), .B(n27326), .Z(n27228) );
  XOR U27714 ( .A(n27327), .B(n27328), .Z(n27326) );
  ANDN U27715 ( .B(n27329), .A(n27330), .Z(n27327) );
  XOR U27716 ( .A(n27331), .B(n27328), .Z(n27329) );
  IV U27717 ( .A(n27230), .Z(n27226) );
  XOR U27718 ( .A(n27332), .B(n27333), .Z(n27230) );
  ANDN U27719 ( .B(n27334), .A(n27335), .Z(n27332) );
  XOR U27720 ( .A(n27336), .B(n27333), .Z(n27334) );
  IV U27721 ( .A(n27240), .Z(n27244) );
  XOR U27722 ( .A(n27240), .B(n27143), .Z(n27242) );
  XOR U27723 ( .A(n27337), .B(n27338), .Z(n27143) );
  AND U27724 ( .A(n316), .B(n27339), .Z(n27337) );
  XOR U27725 ( .A(n27340), .B(n27338), .Z(n27339) );
  NANDN U27726 ( .A(n27145), .B(n27147), .Z(n27240) );
  XOR U27727 ( .A(n27341), .B(n27342), .Z(n27147) );
  AND U27728 ( .A(n316), .B(n27343), .Z(n27341) );
  XOR U27729 ( .A(n27342), .B(n27344), .Z(n27343) );
  XNOR U27730 ( .A(n27345), .B(n27346), .Z(n316) );
  AND U27731 ( .A(n27347), .B(n27348), .Z(n27345) );
  XOR U27732 ( .A(n27346), .B(n27158), .Z(n27348) );
  XNOR U27733 ( .A(n27349), .B(n27350), .Z(n27158) );
  ANDN U27734 ( .B(n27351), .A(n27352), .Z(n27349) );
  XOR U27735 ( .A(n27350), .B(n27353), .Z(n27351) );
  XNOR U27736 ( .A(n27346), .B(n27160), .Z(n27347) );
  XOR U27737 ( .A(n27354), .B(n27355), .Z(n27160) );
  AND U27738 ( .A(n320), .B(n27356), .Z(n27354) );
  XOR U27739 ( .A(n27357), .B(n27355), .Z(n27356) );
  XOR U27740 ( .A(n27358), .B(n27359), .Z(n27346) );
  AND U27741 ( .A(n27360), .B(n27361), .Z(n27358) );
  XOR U27742 ( .A(n27359), .B(n27185), .Z(n27361) );
  XOR U27743 ( .A(n27352), .B(n27353), .Z(n27185) );
  XNOR U27744 ( .A(n27362), .B(n27363), .Z(n27353) );
  ANDN U27745 ( .B(n27364), .A(n27365), .Z(n27362) );
  XOR U27746 ( .A(n27366), .B(n27367), .Z(n27364) );
  XOR U27747 ( .A(n27368), .B(n27369), .Z(n27352) );
  XNOR U27748 ( .A(n27370), .B(n27371), .Z(n27369) );
  ANDN U27749 ( .B(n27372), .A(n27373), .Z(n27370) );
  XNOR U27750 ( .A(n27374), .B(n27375), .Z(n27372) );
  IV U27751 ( .A(n27350), .Z(n27368) );
  XOR U27752 ( .A(n27376), .B(n27377), .Z(n27350) );
  ANDN U27753 ( .B(n27378), .A(n27379), .Z(n27376) );
  XOR U27754 ( .A(n27377), .B(n27380), .Z(n27378) );
  XNOR U27755 ( .A(n27359), .B(n27187), .Z(n27360) );
  XOR U27756 ( .A(n27381), .B(n27382), .Z(n27187) );
  AND U27757 ( .A(n320), .B(n27383), .Z(n27381) );
  XOR U27758 ( .A(n27384), .B(n27382), .Z(n27383) );
  XNOR U27759 ( .A(n27385), .B(n27386), .Z(n27359) );
  AND U27760 ( .A(n27387), .B(n27388), .Z(n27385) );
  XNOR U27761 ( .A(n27386), .B(n27237), .Z(n27388) );
  XOR U27762 ( .A(n27379), .B(n27380), .Z(n27237) );
  XOR U27763 ( .A(n27389), .B(n27367), .Z(n27380) );
  XNOR U27764 ( .A(n27390), .B(n27391), .Z(n27367) );
  ANDN U27765 ( .B(n27392), .A(n27393), .Z(n27390) );
  XOR U27766 ( .A(n27394), .B(n27395), .Z(n27392) );
  IV U27767 ( .A(n27365), .Z(n27389) );
  XOR U27768 ( .A(n27363), .B(n27396), .Z(n27365) );
  XNOR U27769 ( .A(n27397), .B(n27398), .Z(n27396) );
  ANDN U27770 ( .B(n27399), .A(n27400), .Z(n27397) );
  XNOR U27771 ( .A(n27401), .B(n27402), .Z(n27399) );
  IV U27772 ( .A(n27366), .Z(n27363) );
  XOR U27773 ( .A(n27403), .B(n27404), .Z(n27366) );
  ANDN U27774 ( .B(n27405), .A(n27406), .Z(n27403) );
  XOR U27775 ( .A(n27404), .B(n27407), .Z(n27405) );
  XOR U27776 ( .A(n27408), .B(n27409), .Z(n27379) );
  XNOR U27777 ( .A(n27374), .B(n27410), .Z(n27409) );
  IV U27778 ( .A(n27377), .Z(n27410) );
  XOR U27779 ( .A(n27411), .B(n27412), .Z(n27377) );
  ANDN U27780 ( .B(n27413), .A(n27414), .Z(n27411) );
  XOR U27781 ( .A(n27412), .B(n27415), .Z(n27413) );
  XNOR U27782 ( .A(n27416), .B(n27417), .Z(n27374) );
  ANDN U27783 ( .B(n27418), .A(n27419), .Z(n27416) );
  XOR U27784 ( .A(n27417), .B(n27420), .Z(n27418) );
  IV U27785 ( .A(n27373), .Z(n27408) );
  XOR U27786 ( .A(n27371), .B(n27421), .Z(n27373) );
  XNOR U27787 ( .A(n27422), .B(n27423), .Z(n27421) );
  ANDN U27788 ( .B(n27424), .A(n27425), .Z(n27422) );
  XNOR U27789 ( .A(n27426), .B(n27427), .Z(n27424) );
  IV U27790 ( .A(n27375), .Z(n27371) );
  XOR U27791 ( .A(n27428), .B(n27429), .Z(n27375) );
  ANDN U27792 ( .B(n27430), .A(n27431), .Z(n27428) );
  XOR U27793 ( .A(n27432), .B(n27429), .Z(n27430) );
  XOR U27794 ( .A(n27386), .B(n27239), .Z(n27387) );
  XOR U27795 ( .A(n27433), .B(n27434), .Z(n27239) );
  AND U27796 ( .A(n320), .B(n27435), .Z(n27433) );
  XOR U27797 ( .A(n27436), .B(n27434), .Z(n27435) );
  XNOR U27798 ( .A(n27437), .B(n27438), .Z(n27386) );
  NAND U27799 ( .A(n27439), .B(n27440), .Z(n27438) );
  XOR U27800 ( .A(n27441), .B(n27338), .Z(n27440) );
  XOR U27801 ( .A(n27414), .B(n27415), .Z(n27338) );
  XOR U27802 ( .A(n27442), .B(n27407), .Z(n27415) );
  XOR U27803 ( .A(n27443), .B(n27395), .Z(n27407) );
  XOR U27804 ( .A(n27444), .B(n27445), .Z(n27395) );
  ANDN U27805 ( .B(n27446), .A(n27447), .Z(n27444) );
  XOR U27806 ( .A(n27445), .B(n27448), .Z(n27446) );
  IV U27807 ( .A(n27393), .Z(n27443) );
  XOR U27808 ( .A(n27391), .B(n27449), .Z(n27393) );
  XOR U27809 ( .A(n27450), .B(n27451), .Z(n27449) );
  ANDN U27810 ( .B(n27452), .A(n27453), .Z(n27450) );
  XOR U27811 ( .A(n27454), .B(n27451), .Z(n27452) );
  IV U27812 ( .A(n27394), .Z(n27391) );
  XOR U27813 ( .A(n27455), .B(n27456), .Z(n27394) );
  ANDN U27814 ( .B(n27457), .A(n27458), .Z(n27455) );
  XOR U27815 ( .A(n27456), .B(n27459), .Z(n27457) );
  IV U27816 ( .A(n27406), .Z(n27442) );
  XOR U27817 ( .A(n27460), .B(n27461), .Z(n27406) );
  XNOR U27818 ( .A(n27401), .B(n27462), .Z(n27461) );
  IV U27819 ( .A(n27404), .Z(n27462) );
  XOR U27820 ( .A(n27463), .B(n27464), .Z(n27404) );
  ANDN U27821 ( .B(n27465), .A(n27466), .Z(n27463) );
  XOR U27822 ( .A(n27464), .B(n27467), .Z(n27465) );
  XNOR U27823 ( .A(n27468), .B(n27469), .Z(n27401) );
  ANDN U27824 ( .B(n27470), .A(n27471), .Z(n27468) );
  XOR U27825 ( .A(n27469), .B(n27472), .Z(n27470) );
  IV U27826 ( .A(n27400), .Z(n27460) );
  XOR U27827 ( .A(n27398), .B(n27473), .Z(n27400) );
  XOR U27828 ( .A(n27474), .B(n27475), .Z(n27473) );
  ANDN U27829 ( .B(n27476), .A(n27477), .Z(n27474) );
  XOR U27830 ( .A(n27478), .B(n27475), .Z(n27476) );
  IV U27831 ( .A(n27402), .Z(n27398) );
  XOR U27832 ( .A(n27479), .B(n27480), .Z(n27402) );
  ANDN U27833 ( .B(n27481), .A(n27482), .Z(n27479) );
  XOR U27834 ( .A(n27483), .B(n27480), .Z(n27481) );
  XOR U27835 ( .A(n27484), .B(n27485), .Z(n27414) );
  XOR U27836 ( .A(n27432), .B(n27486), .Z(n27485) );
  IV U27837 ( .A(n27412), .Z(n27486) );
  XOR U27838 ( .A(n27487), .B(n27488), .Z(n27412) );
  ANDN U27839 ( .B(n27489), .A(n27490), .Z(n27487) );
  XOR U27840 ( .A(n27488), .B(n27491), .Z(n27489) );
  XOR U27841 ( .A(n27492), .B(n27420), .Z(n27432) );
  XOR U27842 ( .A(n27493), .B(n27494), .Z(n27420) );
  ANDN U27843 ( .B(n27495), .A(n27496), .Z(n27493) );
  XOR U27844 ( .A(n27494), .B(n27497), .Z(n27495) );
  IV U27845 ( .A(n27419), .Z(n27492) );
  XOR U27846 ( .A(n27498), .B(n27499), .Z(n27419) );
  XOR U27847 ( .A(n27500), .B(n27501), .Z(n27499) );
  ANDN U27848 ( .B(n27502), .A(n27503), .Z(n27500) );
  XOR U27849 ( .A(n27504), .B(n27501), .Z(n27502) );
  IV U27850 ( .A(n27417), .Z(n27498) );
  XOR U27851 ( .A(n27505), .B(n27506), .Z(n27417) );
  ANDN U27852 ( .B(n27507), .A(n27508), .Z(n27505) );
  XOR U27853 ( .A(n27506), .B(n27509), .Z(n27507) );
  IV U27854 ( .A(n27431), .Z(n27484) );
  XOR U27855 ( .A(n27510), .B(n27511), .Z(n27431) );
  XNOR U27856 ( .A(n27426), .B(n27512), .Z(n27511) );
  IV U27857 ( .A(n27429), .Z(n27512) );
  XOR U27858 ( .A(n27513), .B(n27514), .Z(n27429) );
  ANDN U27859 ( .B(n27515), .A(n27516), .Z(n27513) );
  XOR U27860 ( .A(n27517), .B(n27514), .Z(n27515) );
  XNOR U27861 ( .A(n27518), .B(n27519), .Z(n27426) );
  ANDN U27862 ( .B(n27520), .A(n27521), .Z(n27518) );
  XOR U27863 ( .A(n27519), .B(n27522), .Z(n27520) );
  IV U27864 ( .A(n27425), .Z(n27510) );
  XOR U27865 ( .A(n27423), .B(n27523), .Z(n27425) );
  XOR U27866 ( .A(n27524), .B(n27525), .Z(n27523) );
  ANDN U27867 ( .B(n27526), .A(n27527), .Z(n27524) );
  XOR U27868 ( .A(n27528), .B(n27525), .Z(n27526) );
  IV U27869 ( .A(n27427), .Z(n27423) );
  XOR U27870 ( .A(n27529), .B(n27530), .Z(n27427) );
  ANDN U27871 ( .B(n27531), .A(n27532), .Z(n27529) );
  XOR U27872 ( .A(n27533), .B(n27530), .Z(n27531) );
  IV U27873 ( .A(n27437), .Z(n27441) );
  XOR U27874 ( .A(n27437), .B(n27340), .Z(n27439) );
  XOR U27875 ( .A(n27534), .B(n27535), .Z(n27340) );
  AND U27876 ( .A(n320), .B(n27536), .Z(n27534) );
  XOR U27877 ( .A(n27537), .B(n27535), .Z(n27536) );
  NANDN U27878 ( .A(n27342), .B(n27344), .Z(n27437) );
  XOR U27879 ( .A(n27538), .B(n27539), .Z(n27344) );
  AND U27880 ( .A(n320), .B(n27540), .Z(n27538) );
  XOR U27881 ( .A(n27539), .B(n27541), .Z(n27540) );
  XNOR U27882 ( .A(n27542), .B(n27543), .Z(n320) );
  AND U27883 ( .A(n27544), .B(n27545), .Z(n27542) );
  XOR U27884 ( .A(n27543), .B(n27355), .Z(n27545) );
  XNOR U27885 ( .A(n27546), .B(n27547), .Z(n27355) );
  ANDN U27886 ( .B(n27548), .A(n27549), .Z(n27546) );
  XOR U27887 ( .A(n27547), .B(n27550), .Z(n27548) );
  XNOR U27888 ( .A(n27543), .B(n27357), .Z(n27544) );
  XOR U27889 ( .A(n27551), .B(n27552), .Z(n27357) );
  AND U27890 ( .A(n324), .B(n27553), .Z(n27551) );
  XOR U27891 ( .A(n27554), .B(n27552), .Z(n27553) );
  XOR U27892 ( .A(n27555), .B(n27556), .Z(n27543) );
  AND U27893 ( .A(n27557), .B(n27558), .Z(n27555) );
  XOR U27894 ( .A(n27556), .B(n27382), .Z(n27558) );
  XOR U27895 ( .A(n27549), .B(n27550), .Z(n27382) );
  XNOR U27896 ( .A(n27559), .B(n27560), .Z(n27550) );
  ANDN U27897 ( .B(n27561), .A(n27562), .Z(n27559) );
  XOR U27898 ( .A(n27563), .B(n27564), .Z(n27561) );
  XOR U27899 ( .A(n27565), .B(n27566), .Z(n27549) );
  XNOR U27900 ( .A(n27567), .B(n27568), .Z(n27566) );
  ANDN U27901 ( .B(n27569), .A(n27570), .Z(n27567) );
  XNOR U27902 ( .A(n27571), .B(n27572), .Z(n27569) );
  IV U27903 ( .A(n27547), .Z(n27565) );
  XOR U27904 ( .A(n27573), .B(n27574), .Z(n27547) );
  ANDN U27905 ( .B(n27575), .A(n27576), .Z(n27573) );
  XOR U27906 ( .A(n27574), .B(n27577), .Z(n27575) );
  XNOR U27907 ( .A(n27556), .B(n27384), .Z(n27557) );
  XOR U27908 ( .A(n27578), .B(n27579), .Z(n27384) );
  AND U27909 ( .A(n324), .B(n27580), .Z(n27578) );
  XOR U27910 ( .A(n27581), .B(n27579), .Z(n27580) );
  XNOR U27911 ( .A(n27582), .B(n27583), .Z(n27556) );
  AND U27912 ( .A(n27584), .B(n27585), .Z(n27582) );
  XNOR U27913 ( .A(n27583), .B(n27434), .Z(n27585) );
  XOR U27914 ( .A(n27576), .B(n27577), .Z(n27434) );
  XOR U27915 ( .A(n27586), .B(n27564), .Z(n27577) );
  XNOR U27916 ( .A(n27587), .B(n27588), .Z(n27564) );
  ANDN U27917 ( .B(n27589), .A(n27590), .Z(n27587) );
  XOR U27918 ( .A(n27591), .B(n27592), .Z(n27589) );
  IV U27919 ( .A(n27562), .Z(n27586) );
  XOR U27920 ( .A(n27560), .B(n27593), .Z(n27562) );
  XNOR U27921 ( .A(n27594), .B(n27595), .Z(n27593) );
  ANDN U27922 ( .B(n27596), .A(n27597), .Z(n27594) );
  XNOR U27923 ( .A(n27598), .B(n27599), .Z(n27596) );
  IV U27924 ( .A(n27563), .Z(n27560) );
  XOR U27925 ( .A(n27600), .B(n27601), .Z(n27563) );
  ANDN U27926 ( .B(n27602), .A(n27603), .Z(n27600) );
  XOR U27927 ( .A(n27601), .B(n27604), .Z(n27602) );
  XOR U27928 ( .A(n27605), .B(n27606), .Z(n27576) );
  XNOR U27929 ( .A(n27571), .B(n27607), .Z(n27606) );
  IV U27930 ( .A(n27574), .Z(n27607) );
  XOR U27931 ( .A(n27608), .B(n27609), .Z(n27574) );
  ANDN U27932 ( .B(n27610), .A(n27611), .Z(n27608) );
  XOR U27933 ( .A(n27609), .B(n27612), .Z(n27610) );
  XNOR U27934 ( .A(n27613), .B(n27614), .Z(n27571) );
  ANDN U27935 ( .B(n27615), .A(n27616), .Z(n27613) );
  XOR U27936 ( .A(n27614), .B(n27617), .Z(n27615) );
  IV U27937 ( .A(n27570), .Z(n27605) );
  XOR U27938 ( .A(n27568), .B(n27618), .Z(n27570) );
  XNOR U27939 ( .A(n27619), .B(n27620), .Z(n27618) );
  ANDN U27940 ( .B(n27621), .A(n27622), .Z(n27619) );
  XNOR U27941 ( .A(n27623), .B(n27624), .Z(n27621) );
  IV U27942 ( .A(n27572), .Z(n27568) );
  XOR U27943 ( .A(n27625), .B(n27626), .Z(n27572) );
  ANDN U27944 ( .B(n27627), .A(n27628), .Z(n27625) );
  XOR U27945 ( .A(n27629), .B(n27626), .Z(n27627) );
  XOR U27946 ( .A(n27583), .B(n27436), .Z(n27584) );
  XOR U27947 ( .A(n27630), .B(n27631), .Z(n27436) );
  AND U27948 ( .A(n324), .B(n27632), .Z(n27630) );
  XOR U27949 ( .A(n27633), .B(n27631), .Z(n27632) );
  XNOR U27950 ( .A(n27634), .B(n27635), .Z(n27583) );
  NAND U27951 ( .A(n27636), .B(n27637), .Z(n27635) );
  XOR U27952 ( .A(n27638), .B(n27535), .Z(n27637) );
  XOR U27953 ( .A(n27611), .B(n27612), .Z(n27535) );
  XOR U27954 ( .A(n27639), .B(n27604), .Z(n27612) );
  XOR U27955 ( .A(n27640), .B(n27592), .Z(n27604) );
  XOR U27956 ( .A(n27641), .B(n27642), .Z(n27592) );
  ANDN U27957 ( .B(n27643), .A(n27644), .Z(n27641) );
  XOR U27958 ( .A(n27642), .B(n27645), .Z(n27643) );
  IV U27959 ( .A(n27590), .Z(n27640) );
  XOR U27960 ( .A(n27588), .B(n27646), .Z(n27590) );
  XOR U27961 ( .A(n27647), .B(n27648), .Z(n27646) );
  ANDN U27962 ( .B(n27649), .A(n27650), .Z(n27647) );
  XOR U27963 ( .A(n27651), .B(n27648), .Z(n27649) );
  IV U27964 ( .A(n27591), .Z(n27588) );
  XOR U27965 ( .A(n27652), .B(n27653), .Z(n27591) );
  ANDN U27966 ( .B(n27654), .A(n27655), .Z(n27652) );
  XOR U27967 ( .A(n27653), .B(n27656), .Z(n27654) );
  IV U27968 ( .A(n27603), .Z(n27639) );
  XOR U27969 ( .A(n27657), .B(n27658), .Z(n27603) );
  XNOR U27970 ( .A(n27598), .B(n27659), .Z(n27658) );
  IV U27971 ( .A(n27601), .Z(n27659) );
  XOR U27972 ( .A(n27660), .B(n27661), .Z(n27601) );
  ANDN U27973 ( .B(n27662), .A(n27663), .Z(n27660) );
  XOR U27974 ( .A(n27661), .B(n27664), .Z(n27662) );
  XNOR U27975 ( .A(n27665), .B(n27666), .Z(n27598) );
  ANDN U27976 ( .B(n27667), .A(n27668), .Z(n27665) );
  XOR U27977 ( .A(n27666), .B(n27669), .Z(n27667) );
  IV U27978 ( .A(n27597), .Z(n27657) );
  XOR U27979 ( .A(n27595), .B(n27670), .Z(n27597) );
  XOR U27980 ( .A(n27671), .B(n27672), .Z(n27670) );
  ANDN U27981 ( .B(n27673), .A(n27674), .Z(n27671) );
  XOR U27982 ( .A(n27675), .B(n27672), .Z(n27673) );
  IV U27983 ( .A(n27599), .Z(n27595) );
  XOR U27984 ( .A(n27676), .B(n27677), .Z(n27599) );
  ANDN U27985 ( .B(n27678), .A(n27679), .Z(n27676) );
  XOR U27986 ( .A(n27680), .B(n27677), .Z(n27678) );
  XOR U27987 ( .A(n27681), .B(n27682), .Z(n27611) );
  XOR U27988 ( .A(n27629), .B(n27683), .Z(n27682) );
  IV U27989 ( .A(n27609), .Z(n27683) );
  XOR U27990 ( .A(n27684), .B(n27685), .Z(n27609) );
  ANDN U27991 ( .B(n27686), .A(n27687), .Z(n27684) );
  XOR U27992 ( .A(n27685), .B(n27688), .Z(n27686) );
  XOR U27993 ( .A(n27689), .B(n27617), .Z(n27629) );
  XOR U27994 ( .A(n27690), .B(n27691), .Z(n27617) );
  ANDN U27995 ( .B(n27692), .A(n27693), .Z(n27690) );
  XOR U27996 ( .A(n27691), .B(n27694), .Z(n27692) );
  IV U27997 ( .A(n27616), .Z(n27689) );
  XOR U27998 ( .A(n27695), .B(n27696), .Z(n27616) );
  XOR U27999 ( .A(n27697), .B(n27698), .Z(n27696) );
  ANDN U28000 ( .B(n27699), .A(n27700), .Z(n27697) );
  XOR U28001 ( .A(n27701), .B(n27698), .Z(n27699) );
  IV U28002 ( .A(n27614), .Z(n27695) );
  XOR U28003 ( .A(n27702), .B(n27703), .Z(n27614) );
  ANDN U28004 ( .B(n27704), .A(n27705), .Z(n27702) );
  XOR U28005 ( .A(n27703), .B(n27706), .Z(n27704) );
  IV U28006 ( .A(n27628), .Z(n27681) );
  XOR U28007 ( .A(n27707), .B(n27708), .Z(n27628) );
  XNOR U28008 ( .A(n27623), .B(n27709), .Z(n27708) );
  IV U28009 ( .A(n27626), .Z(n27709) );
  XOR U28010 ( .A(n27710), .B(n27711), .Z(n27626) );
  ANDN U28011 ( .B(n27712), .A(n27713), .Z(n27710) );
  XOR U28012 ( .A(n27714), .B(n27711), .Z(n27712) );
  XNOR U28013 ( .A(n27715), .B(n27716), .Z(n27623) );
  ANDN U28014 ( .B(n27717), .A(n27718), .Z(n27715) );
  XOR U28015 ( .A(n27716), .B(n27719), .Z(n27717) );
  IV U28016 ( .A(n27622), .Z(n27707) );
  XOR U28017 ( .A(n27620), .B(n27720), .Z(n27622) );
  XOR U28018 ( .A(n27721), .B(n27722), .Z(n27720) );
  ANDN U28019 ( .B(n27723), .A(n27724), .Z(n27721) );
  XOR U28020 ( .A(n27725), .B(n27722), .Z(n27723) );
  IV U28021 ( .A(n27624), .Z(n27620) );
  XOR U28022 ( .A(n27726), .B(n27727), .Z(n27624) );
  ANDN U28023 ( .B(n27728), .A(n27729), .Z(n27726) );
  XOR U28024 ( .A(n27730), .B(n27727), .Z(n27728) );
  IV U28025 ( .A(n27634), .Z(n27638) );
  XOR U28026 ( .A(n27634), .B(n27537), .Z(n27636) );
  XOR U28027 ( .A(n27731), .B(n27732), .Z(n27537) );
  AND U28028 ( .A(n324), .B(n27733), .Z(n27731) );
  XOR U28029 ( .A(n27734), .B(n27732), .Z(n27733) );
  NANDN U28030 ( .A(n27539), .B(n27541), .Z(n27634) );
  XOR U28031 ( .A(n27735), .B(n27736), .Z(n27541) );
  AND U28032 ( .A(n324), .B(n27737), .Z(n27735) );
  XOR U28033 ( .A(n27736), .B(n27738), .Z(n27737) );
  XNOR U28034 ( .A(n27739), .B(n27740), .Z(n324) );
  AND U28035 ( .A(n27741), .B(n27742), .Z(n27739) );
  XOR U28036 ( .A(n27740), .B(n27552), .Z(n27742) );
  XNOR U28037 ( .A(n27743), .B(n27744), .Z(n27552) );
  ANDN U28038 ( .B(n27745), .A(n27746), .Z(n27743) );
  XOR U28039 ( .A(n27744), .B(n27747), .Z(n27745) );
  XNOR U28040 ( .A(n27740), .B(n27554), .Z(n27741) );
  XOR U28041 ( .A(n27748), .B(n27749), .Z(n27554) );
  AND U28042 ( .A(n328), .B(n27750), .Z(n27748) );
  XOR U28043 ( .A(n27751), .B(n27749), .Z(n27750) );
  XOR U28044 ( .A(n27752), .B(n27753), .Z(n27740) );
  AND U28045 ( .A(n27754), .B(n27755), .Z(n27752) );
  XOR U28046 ( .A(n27753), .B(n27579), .Z(n27755) );
  XOR U28047 ( .A(n27746), .B(n27747), .Z(n27579) );
  XNOR U28048 ( .A(n27756), .B(n27757), .Z(n27747) );
  ANDN U28049 ( .B(n27758), .A(n27759), .Z(n27756) );
  XOR U28050 ( .A(n27760), .B(n27761), .Z(n27758) );
  XOR U28051 ( .A(n27762), .B(n27763), .Z(n27746) );
  XNOR U28052 ( .A(n27764), .B(n27765), .Z(n27763) );
  ANDN U28053 ( .B(n27766), .A(n27767), .Z(n27764) );
  XNOR U28054 ( .A(n27768), .B(n27769), .Z(n27766) );
  IV U28055 ( .A(n27744), .Z(n27762) );
  XOR U28056 ( .A(n27770), .B(n27771), .Z(n27744) );
  ANDN U28057 ( .B(n27772), .A(n27773), .Z(n27770) );
  XOR U28058 ( .A(n27771), .B(n27774), .Z(n27772) );
  XNOR U28059 ( .A(n27753), .B(n27581), .Z(n27754) );
  XOR U28060 ( .A(n27775), .B(n27776), .Z(n27581) );
  AND U28061 ( .A(n328), .B(n27777), .Z(n27775) );
  XOR U28062 ( .A(n27778), .B(n27776), .Z(n27777) );
  XNOR U28063 ( .A(n27779), .B(n27780), .Z(n27753) );
  AND U28064 ( .A(n27781), .B(n27782), .Z(n27779) );
  XNOR U28065 ( .A(n27780), .B(n27631), .Z(n27782) );
  XOR U28066 ( .A(n27773), .B(n27774), .Z(n27631) );
  XOR U28067 ( .A(n27783), .B(n27761), .Z(n27774) );
  XNOR U28068 ( .A(n27784), .B(n27785), .Z(n27761) );
  ANDN U28069 ( .B(n27786), .A(n27787), .Z(n27784) );
  XOR U28070 ( .A(n27788), .B(n27789), .Z(n27786) );
  IV U28071 ( .A(n27759), .Z(n27783) );
  XOR U28072 ( .A(n27757), .B(n27790), .Z(n27759) );
  XNOR U28073 ( .A(n27791), .B(n27792), .Z(n27790) );
  ANDN U28074 ( .B(n27793), .A(n27794), .Z(n27791) );
  XNOR U28075 ( .A(n27795), .B(n27796), .Z(n27793) );
  IV U28076 ( .A(n27760), .Z(n27757) );
  XOR U28077 ( .A(n27797), .B(n27798), .Z(n27760) );
  ANDN U28078 ( .B(n27799), .A(n27800), .Z(n27797) );
  XOR U28079 ( .A(n27798), .B(n27801), .Z(n27799) );
  XOR U28080 ( .A(n27802), .B(n27803), .Z(n27773) );
  XNOR U28081 ( .A(n27768), .B(n27804), .Z(n27803) );
  IV U28082 ( .A(n27771), .Z(n27804) );
  XOR U28083 ( .A(n27805), .B(n27806), .Z(n27771) );
  ANDN U28084 ( .B(n27807), .A(n27808), .Z(n27805) );
  XOR U28085 ( .A(n27806), .B(n27809), .Z(n27807) );
  XNOR U28086 ( .A(n27810), .B(n27811), .Z(n27768) );
  ANDN U28087 ( .B(n27812), .A(n27813), .Z(n27810) );
  XOR U28088 ( .A(n27811), .B(n27814), .Z(n27812) );
  IV U28089 ( .A(n27767), .Z(n27802) );
  XOR U28090 ( .A(n27765), .B(n27815), .Z(n27767) );
  XNOR U28091 ( .A(n27816), .B(n27817), .Z(n27815) );
  ANDN U28092 ( .B(n27818), .A(n27819), .Z(n27816) );
  XNOR U28093 ( .A(n27820), .B(n27821), .Z(n27818) );
  IV U28094 ( .A(n27769), .Z(n27765) );
  XOR U28095 ( .A(n27822), .B(n27823), .Z(n27769) );
  ANDN U28096 ( .B(n27824), .A(n27825), .Z(n27822) );
  XOR U28097 ( .A(n27826), .B(n27823), .Z(n27824) );
  XOR U28098 ( .A(n27780), .B(n27633), .Z(n27781) );
  XOR U28099 ( .A(n27827), .B(n27828), .Z(n27633) );
  AND U28100 ( .A(n328), .B(n27829), .Z(n27827) );
  XOR U28101 ( .A(n27830), .B(n27828), .Z(n27829) );
  XNOR U28102 ( .A(n27831), .B(n27832), .Z(n27780) );
  NAND U28103 ( .A(n27833), .B(n27834), .Z(n27832) );
  XOR U28104 ( .A(n27835), .B(n27732), .Z(n27834) );
  XOR U28105 ( .A(n27808), .B(n27809), .Z(n27732) );
  XOR U28106 ( .A(n27836), .B(n27801), .Z(n27809) );
  XOR U28107 ( .A(n27837), .B(n27789), .Z(n27801) );
  XOR U28108 ( .A(n27838), .B(n27839), .Z(n27789) );
  ANDN U28109 ( .B(n27840), .A(n27841), .Z(n27838) );
  XOR U28110 ( .A(n27839), .B(n27842), .Z(n27840) );
  IV U28111 ( .A(n27787), .Z(n27837) );
  XOR U28112 ( .A(n27785), .B(n27843), .Z(n27787) );
  XOR U28113 ( .A(n27844), .B(n27845), .Z(n27843) );
  ANDN U28114 ( .B(n27846), .A(n27847), .Z(n27844) );
  XOR U28115 ( .A(n27848), .B(n27845), .Z(n27846) );
  IV U28116 ( .A(n27788), .Z(n27785) );
  XOR U28117 ( .A(n27849), .B(n27850), .Z(n27788) );
  ANDN U28118 ( .B(n27851), .A(n27852), .Z(n27849) );
  XOR U28119 ( .A(n27850), .B(n27853), .Z(n27851) );
  IV U28120 ( .A(n27800), .Z(n27836) );
  XOR U28121 ( .A(n27854), .B(n27855), .Z(n27800) );
  XNOR U28122 ( .A(n27795), .B(n27856), .Z(n27855) );
  IV U28123 ( .A(n27798), .Z(n27856) );
  XOR U28124 ( .A(n27857), .B(n27858), .Z(n27798) );
  ANDN U28125 ( .B(n27859), .A(n27860), .Z(n27857) );
  XOR U28126 ( .A(n27858), .B(n27861), .Z(n27859) );
  XNOR U28127 ( .A(n27862), .B(n27863), .Z(n27795) );
  ANDN U28128 ( .B(n27864), .A(n27865), .Z(n27862) );
  XOR U28129 ( .A(n27863), .B(n27866), .Z(n27864) );
  IV U28130 ( .A(n27794), .Z(n27854) );
  XOR U28131 ( .A(n27792), .B(n27867), .Z(n27794) );
  XOR U28132 ( .A(n27868), .B(n27869), .Z(n27867) );
  ANDN U28133 ( .B(n27870), .A(n27871), .Z(n27868) );
  XOR U28134 ( .A(n27872), .B(n27869), .Z(n27870) );
  IV U28135 ( .A(n27796), .Z(n27792) );
  XOR U28136 ( .A(n27873), .B(n27874), .Z(n27796) );
  ANDN U28137 ( .B(n27875), .A(n27876), .Z(n27873) );
  XOR U28138 ( .A(n27877), .B(n27874), .Z(n27875) );
  XOR U28139 ( .A(n27878), .B(n27879), .Z(n27808) );
  XOR U28140 ( .A(n27826), .B(n27880), .Z(n27879) );
  IV U28141 ( .A(n27806), .Z(n27880) );
  XOR U28142 ( .A(n27881), .B(n27882), .Z(n27806) );
  ANDN U28143 ( .B(n27883), .A(n27884), .Z(n27881) );
  XOR U28144 ( .A(n27882), .B(n27885), .Z(n27883) );
  XOR U28145 ( .A(n27886), .B(n27814), .Z(n27826) );
  XOR U28146 ( .A(n27887), .B(n27888), .Z(n27814) );
  ANDN U28147 ( .B(n27889), .A(n27890), .Z(n27887) );
  XOR U28148 ( .A(n27888), .B(n27891), .Z(n27889) );
  IV U28149 ( .A(n27813), .Z(n27886) );
  XOR U28150 ( .A(n27892), .B(n27893), .Z(n27813) );
  XOR U28151 ( .A(n27894), .B(n27895), .Z(n27893) );
  ANDN U28152 ( .B(n27896), .A(n27897), .Z(n27894) );
  XOR U28153 ( .A(n27898), .B(n27895), .Z(n27896) );
  IV U28154 ( .A(n27811), .Z(n27892) );
  XOR U28155 ( .A(n27899), .B(n27900), .Z(n27811) );
  ANDN U28156 ( .B(n27901), .A(n27902), .Z(n27899) );
  XOR U28157 ( .A(n27900), .B(n27903), .Z(n27901) );
  IV U28158 ( .A(n27825), .Z(n27878) );
  XOR U28159 ( .A(n27904), .B(n27905), .Z(n27825) );
  XNOR U28160 ( .A(n27820), .B(n27906), .Z(n27905) );
  IV U28161 ( .A(n27823), .Z(n27906) );
  XOR U28162 ( .A(n27907), .B(n27908), .Z(n27823) );
  ANDN U28163 ( .B(n27909), .A(n27910), .Z(n27907) );
  XOR U28164 ( .A(n27911), .B(n27908), .Z(n27909) );
  XNOR U28165 ( .A(n27912), .B(n27913), .Z(n27820) );
  ANDN U28166 ( .B(n27914), .A(n27915), .Z(n27912) );
  XOR U28167 ( .A(n27913), .B(n27916), .Z(n27914) );
  IV U28168 ( .A(n27819), .Z(n27904) );
  XOR U28169 ( .A(n27817), .B(n27917), .Z(n27819) );
  XOR U28170 ( .A(n27918), .B(n27919), .Z(n27917) );
  ANDN U28171 ( .B(n27920), .A(n27921), .Z(n27918) );
  XOR U28172 ( .A(n27922), .B(n27919), .Z(n27920) );
  IV U28173 ( .A(n27821), .Z(n27817) );
  XOR U28174 ( .A(n27923), .B(n27924), .Z(n27821) );
  ANDN U28175 ( .B(n27925), .A(n27926), .Z(n27923) );
  XOR U28176 ( .A(n27927), .B(n27924), .Z(n27925) );
  IV U28177 ( .A(n27831), .Z(n27835) );
  XOR U28178 ( .A(n27831), .B(n27734), .Z(n27833) );
  XOR U28179 ( .A(n27928), .B(n27929), .Z(n27734) );
  AND U28180 ( .A(n328), .B(n27930), .Z(n27928) );
  XOR U28181 ( .A(n27931), .B(n27929), .Z(n27930) );
  NANDN U28182 ( .A(n27736), .B(n27738), .Z(n27831) );
  XOR U28183 ( .A(n27932), .B(n27933), .Z(n27738) );
  AND U28184 ( .A(n328), .B(n27934), .Z(n27932) );
  XOR U28185 ( .A(n27933), .B(n27935), .Z(n27934) );
  XNOR U28186 ( .A(n27936), .B(n27937), .Z(n328) );
  AND U28187 ( .A(n27938), .B(n27939), .Z(n27936) );
  XOR U28188 ( .A(n27937), .B(n27749), .Z(n27939) );
  XNOR U28189 ( .A(n27940), .B(n27941), .Z(n27749) );
  ANDN U28190 ( .B(n27942), .A(n27943), .Z(n27940) );
  XOR U28191 ( .A(n27941), .B(n27944), .Z(n27942) );
  XNOR U28192 ( .A(n27937), .B(n27751), .Z(n27938) );
  XOR U28193 ( .A(n27945), .B(n27946), .Z(n27751) );
  AND U28194 ( .A(n332), .B(n27947), .Z(n27945) );
  XOR U28195 ( .A(n27948), .B(n27946), .Z(n27947) );
  XOR U28196 ( .A(n27949), .B(n27950), .Z(n27937) );
  AND U28197 ( .A(n27951), .B(n27952), .Z(n27949) );
  XOR U28198 ( .A(n27950), .B(n27776), .Z(n27952) );
  XOR U28199 ( .A(n27943), .B(n27944), .Z(n27776) );
  XNOR U28200 ( .A(n27953), .B(n27954), .Z(n27944) );
  ANDN U28201 ( .B(n27955), .A(n27956), .Z(n27953) );
  XOR U28202 ( .A(n27957), .B(n27958), .Z(n27955) );
  XOR U28203 ( .A(n27959), .B(n27960), .Z(n27943) );
  XNOR U28204 ( .A(n27961), .B(n27962), .Z(n27960) );
  ANDN U28205 ( .B(n27963), .A(n27964), .Z(n27961) );
  XNOR U28206 ( .A(n27965), .B(n27966), .Z(n27963) );
  IV U28207 ( .A(n27941), .Z(n27959) );
  XOR U28208 ( .A(n27967), .B(n27968), .Z(n27941) );
  ANDN U28209 ( .B(n27969), .A(n27970), .Z(n27967) );
  XOR U28210 ( .A(n27968), .B(n27971), .Z(n27969) );
  XNOR U28211 ( .A(n27950), .B(n27778), .Z(n27951) );
  XOR U28212 ( .A(n27972), .B(n27973), .Z(n27778) );
  AND U28213 ( .A(n332), .B(n27974), .Z(n27972) );
  XOR U28214 ( .A(n27975), .B(n27973), .Z(n27974) );
  XNOR U28215 ( .A(n27976), .B(n27977), .Z(n27950) );
  AND U28216 ( .A(n27978), .B(n27979), .Z(n27976) );
  XNOR U28217 ( .A(n27977), .B(n27828), .Z(n27979) );
  XOR U28218 ( .A(n27970), .B(n27971), .Z(n27828) );
  XOR U28219 ( .A(n27980), .B(n27958), .Z(n27971) );
  XNOR U28220 ( .A(n27981), .B(n27982), .Z(n27958) );
  ANDN U28221 ( .B(n27983), .A(n27984), .Z(n27981) );
  XOR U28222 ( .A(n27985), .B(n27986), .Z(n27983) );
  IV U28223 ( .A(n27956), .Z(n27980) );
  XOR U28224 ( .A(n27954), .B(n27987), .Z(n27956) );
  XNOR U28225 ( .A(n27988), .B(n27989), .Z(n27987) );
  ANDN U28226 ( .B(n27990), .A(n27991), .Z(n27988) );
  XNOR U28227 ( .A(n27992), .B(n27993), .Z(n27990) );
  IV U28228 ( .A(n27957), .Z(n27954) );
  XOR U28229 ( .A(n27994), .B(n27995), .Z(n27957) );
  ANDN U28230 ( .B(n27996), .A(n27997), .Z(n27994) );
  XOR U28231 ( .A(n27995), .B(n27998), .Z(n27996) );
  XOR U28232 ( .A(n27999), .B(n28000), .Z(n27970) );
  XNOR U28233 ( .A(n27965), .B(n28001), .Z(n28000) );
  IV U28234 ( .A(n27968), .Z(n28001) );
  XOR U28235 ( .A(n28002), .B(n28003), .Z(n27968) );
  ANDN U28236 ( .B(n28004), .A(n28005), .Z(n28002) );
  XOR U28237 ( .A(n28003), .B(n28006), .Z(n28004) );
  XNOR U28238 ( .A(n28007), .B(n28008), .Z(n27965) );
  ANDN U28239 ( .B(n28009), .A(n28010), .Z(n28007) );
  XOR U28240 ( .A(n28008), .B(n28011), .Z(n28009) );
  IV U28241 ( .A(n27964), .Z(n27999) );
  XOR U28242 ( .A(n27962), .B(n28012), .Z(n27964) );
  XNOR U28243 ( .A(n28013), .B(n28014), .Z(n28012) );
  ANDN U28244 ( .B(n28015), .A(n28016), .Z(n28013) );
  XNOR U28245 ( .A(n28017), .B(n28018), .Z(n28015) );
  IV U28246 ( .A(n27966), .Z(n27962) );
  XOR U28247 ( .A(n28019), .B(n28020), .Z(n27966) );
  ANDN U28248 ( .B(n28021), .A(n28022), .Z(n28019) );
  XOR U28249 ( .A(n28023), .B(n28020), .Z(n28021) );
  XOR U28250 ( .A(n27977), .B(n27830), .Z(n27978) );
  XOR U28251 ( .A(n28024), .B(n28025), .Z(n27830) );
  AND U28252 ( .A(n332), .B(n28026), .Z(n28024) );
  XOR U28253 ( .A(n28027), .B(n28025), .Z(n28026) );
  XNOR U28254 ( .A(n28028), .B(n28029), .Z(n27977) );
  NAND U28255 ( .A(n28030), .B(n28031), .Z(n28029) );
  XOR U28256 ( .A(n28032), .B(n27929), .Z(n28031) );
  XOR U28257 ( .A(n28005), .B(n28006), .Z(n27929) );
  XOR U28258 ( .A(n28033), .B(n27998), .Z(n28006) );
  XOR U28259 ( .A(n28034), .B(n27986), .Z(n27998) );
  XOR U28260 ( .A(n28035), .B(n28036), .Z(n27986) );
  ANDN U28261 ( .B(n28037), .A(n28038), .Z(n28035) );
  XOR U28262 ( .A(n28036), .B(n28039), .Z(n28037) );
  IV U28263 ( .A(n27984), .Z(n28034) );
  XOR U28264 ( .A(n27982), .B(n28040), .Z(n27984) );
  XOR U28265 ( .A(n28041), .B(n28042), .Z(n28040) );
  ANDN U28266 ( .B(n28043), .A(n28044), .Z(n28041) );
  XOR U28267 ( .A(n28045), .B(n28042), .Z(n28043) );
  IV U28268 ( .A(n27985), .Z(n27982) );
  XOR U28269 ( .A(n28046), .B(n28047), .Z(n27985) );
  ANDN U28270 ( .B(n28048), .A(n28049), .Z(n28046) );
  XOR U28271 ( .A(n28047), .B(n28050), .Z(n28048) );
  IV U28272 ( .A(n27997), .Z(n28033) );
  XOR U28273 ( .A(n28051), .B(n28052), .Z(n27997) );
  XNOR U28274 ( .A(n27992), .B(n28053), .Z(n28052) );
  IV U28275 ( .A(n27995), .Z(n28053) );
  XOR U28276 ( .A(n28054), .B(n28055), .Z(n27995) );
  ANDN U28277 ( .B(n28056), .A(n28057), .Z(n28054) );
  XOR U28278 ( .A(n28055), .B(n28058), .Z(n28056) );
  XNOR U28279 ( .A(n28059), .B(n28060), .Z(n27992) );
  ANDN U28280 ( .B(n28061), .A(n28062), .Z(n28059) );
  XOR U28281 ( .A(n28060), .B(n28063), .Z(n28061) );
  IV U28282 ( .A(n27991), .Z(n28051) );
  XOR U28283 ( .A(n27989), .B(n28064), .Z(n27991) );
  XOR U28284 ( .A(n28065), .B(n28066), .Z(n28064) );
  ANDN U28285 ( .B(n28067), .A(n28068), .Z(n28065) );
  XOR U28286 ( .A(n28069), .B(n28066), .Z(n28067) );
  IV U28287 ( .A(n27993), .Z(n27989) );
  XOR U28288 ( .A(n28070), .B(n28071), .Z(n27993) );
  ANDN U28289 ( .B(n28072), .A(n28073), .Z(n28070) );
  XOR U28290 ( .A(n28074), .B(n28071), .Z(n28072) );
  XOR U28291 ( .A(n28075), .B(n28076), .Z(n28005) );
  XOR U28292 ( .A(n28023), .B(n28077), .Z(n28076) );
  IV U28293 ( .A(n28003), .Z(n28077) );
  XOR U28294 ( .A(n28078), .B(n28079), .Z(n28003) );
  ANDN U28295 ( .B(n28080), .A(n28081), .Z(n28078) );
  XOR U28296 ( .A(n28079), .B(n28082), .Z(n28080) );
  XOR U28297 ( .A(n28083), .B(n28011), .Z(n28023) );
  XOR U28298 ( .A(n28084), .B(n28085), .Z(n28011) );
  ANDN U28299 ( .B(n28086), .A(n28087), .Z(n28084) );
  XOR U28300 ( .A(n28085), .B(n28088), .Z(n28086) );
  IV U28301 ( .A(n28010), .Z(n28083) );
  XOR U28302 ( .A(n28089), .B(n28090), .Z(n28010) );
  XOR U28303 ( .A(n28091), .B(n28092), .Z(n28090) );
  ANDN U28304 ( .B(n28093), .A(n28094), .Z(n28091) );
  XOR U28305 ( .A(n28095), .B(n28092), .Z(n28093) );
  IV U28306 ( .A(n28008), .Z(n28089) );
  XOR U28307 ( .A(n28096), .B(n28097), .Z(n28008) );
  ANDN U28308 ( .B(n28098), .A(n28099), .Z(n28096) );
  XOR U28309 ( .A(n28097), .B(n28100), .Z(n28098) );
  IV U28310 ( .A(n28022), .Z(n28075) );
  XOR U28311 ( .A(n28101), .B(n28102), .Z(n28022) );
  XNOR U28312 ( .A(n28017), .B(n28103), .Z(n28102) );
  IV U28313 ( .A(n28020), .Z(n28103) );
  XOR U28314 ( .A(n28104), .B(n28105), .Z(n28020) );
  ANDN U28315 ( .B(n28106), .A(n28107), .Z(n28104) );
  XOR U28316 ( .A(n28108), .B(n28105), .Z(n28106) );
  XNOR U28317 ( .A(n28109), .B(n28110), .Z(n28017) );
  ANDN U28318 ( .B(n28111), .A(n28112), .Z(n28109) );
  XOR U28319 ( .A(n28110), .B(n28113), .Z(n28111) );
  IV U28320 ( .A(n28016), .Z(n28101) );
  XOR U28321 ( .A(n28014), .B(n28114), .Z(n28016) );
  XOR U28322 ( .A(n28115), .B(n28116), .Z(n28114) );
  ANDN U28323 ( .B(n28117), .A(n28118), .Z(n28115) );
  XOR U28324 ( .A(n28119), .B(n28116), .Z(n28117) );
  IV U28325 ( .A(n28018), .Z(n28014) );
  XOR U28326 ( .A(n28120), .B(n28121), .Z(n28018) );
  ANDN U28327 ( .B(n28122), .A(n28123), .Z(n28120) );
  XOR U28328 ( .A(n28124), .B(n28121), .Z(n28122) );
  IV U28329 ( .A(n28028), .Z(n28032) );
  XOR U28330 ( .A(n28028), .B(n27931), .Z(n28030) );
  XOR U28331 ( .A(n28125), .B(n28126), .Z(n27931) );
  AND U28332 ( .A(n332), .B(n28127), .Z(n28125) );
  XOR U28333 ( .A(n28128), .B(n28126), .Z(n28127) );
  NANDN U28334 ( .A(n27933), .B(n27935), .Z(n28028) );
  XOR U28335 ( .A(n28129), .B(n28130), .Z(n27935) );
  AND U28336 ( .A(n332), .B(n28131), .Z(n28129) );
  XOR U28337 ( .A(n28130), .B(n28132), .Z(n28131) );
  XNOR U28338 ( .A(n28133), .B(n28134), .Z(n332) );
  AND U28339 ( .A(n28135), .B(n28136), .Z(n28133) );
  XOR U28340 ( .A(n28134), .B(n27946), .Z(n28136) );
  XNOR U28341 ( .A(n28137), .B(n28138), .Z(n27946) );
  ANDN U28342 ( .B(n28139), .A(n28140), .Z(n28137) );
  XOR U28343 ( .A(n28138), .B(n28141), .Z(n28139) );
  XNOR U28344 ( .A(n28134), .B(n27948), .Z(n28135) );
  XOR U28345 ( .A(n28142), .B(n28143), .Z(n27948) );
  AND U28346 ( .A(n336), .B(n28144), .Z(n28142) );
  XOR U28347 ( .A(n28145), .B(n28143), .Z(n28144) );
  XOR U28348 ( .A(n28146), .B(n28147), .Z(n28134) );
  AND U28349 ( .A(n28148), .B(n28149), .Z(n28146) );
  XOR U28350 ( .A(n28147), .B(n27973), .Z(n28149) );
  XOR U28351 ( .A(n28140), .B(n28141), .Z(n27973) );
  XNOR U28352 ( .A(n28150), .B(n28151), .Z(n28141) );
  ANDN U28353 ( .B(n28152), .A(n28153), .Z(n28150) );
  XOR U28354 ( .A(n28154), .B(n28155), .Z(n28152) );
  XOR U28355 ( .A(n28156), .B(n28157), .Z(n28140) );
  XNOR U28356 ( .A(n28158), .B(n28159), .Z(n28157) );
  ANDN U28357 ( .B(n28160), .A(n28161), .Z(n28158) );
  XNOR U28358 ( .A(n28162), .B(n28163), .Z(n28160) );
  IV U28359 ( .A(n28138), .Z(n28156) );
  XOR U28360 ( .A(n28164), .B(n28165), .Z(n28138) );
  ANDN U28361 ( .B(n28166), .A(n28167), .Z(n28164) );
  XOR U28362 ( .A(n28165), .B(n28168), .Z(n28166) );
  XNOR U28363 ( .A(n28147), .B(n27975), .Z(n28148) );
  XOR U28364 ( .A(n28169), .B(n28170), .Z(n27975) );
  AND U28365 ( .A(n336), .B(n28171), .Z(n28169) );
  XOR U28366 ( .A(n28172), .B(n28170), .Z(n28171) );
  XNOR U28367 ( .A(n28173), .B(n28174), .Z(n28147) );
  AND U28368 ( .A(n28175), .B(n28176), .Z(n28173) );
  XNOR U28369 ( .A(n28174), .B(n28025), .Z(n28176) );
  XOR U28370 ( .A(n28167), .B(n28168), .Z(n28025) );
  XOR U28371 ( .A(n28177), .B(n28155), .Z(n28168) );
  XNOR U28372 ( .A(n28178), .B(n28179), .Z(n28155) );
  ANDN U28373 ( .B(n28180), .A(n28181), .Z(n28178) );
  XOR U28374 ( .A(n28182), .B(n28183), .Z(n28180) );
  IV U28375 ( .A(n28153), .Z(n28177) );
  XOR U28376 ( .A(n28151), .B(n28184), .Z(n28153) );
  XNOR U28377 ( .A(n28185), .B(n28186), .Z(n28184) );
  ANDN U28378 ( .B(n28187), .A(n28188), .Z(n28185) );
  XNOR U28379 ( .A(n28189), .B(n28190), .Z(n28187) );
  IV U28380 ( .A(n28154), .Z(n28151) );
  XOR U28381 ( .A(n28191), .B(n28192), .Z(n28154) );
  ANDN U28382 ( .B(n28193), .A(n28194), .Z(n28191) );
  XOR U28383 ( .A(n28192), .B(n28195), .Z(n28193) );
  XOR U28384 ( .A(n28196), .B(n28197), .Z(n28167) );
  XNOR U28385 ( .A(n28162), .B(n28198), .Z(n28197) );
  IV U28386 ( .A(n28165), .Z(n28198) );
  XOR U28387 ( .A(n28199), .B(n28200), .Z(n28165) );
  ANDN U28388 ( .B(n28201), .A(n28202), .Z(n28199) );
  XOR U28389 ( .A(n28200), .B(n28203), .Z(n28201) );
  XNOR U28390 ( .A(n28204), .B(n28205), .Z(n28162) );
  ANDN U28391 ( .B(n28206), .A(n28207), .Z(n28204) );
  XOR U28392 ( .A(n28205), .B(n28208), .Z(n28206) );
  IV U28393 ( .A(n28161), .Z(n28196) );
  XOR U28394 ( .A(n28159), .B(n28209), .Z(n28161) );
  XNOR U28395 ( .A(n28210), .B(n28211), .Z(n28209) );
  ANDN U28396 ( .B(n28212), .A(n28213), .Z(n28210) );
  XNOR U28397 ( .A(n28214), .B(n28215), .Z(n28212) );
  IV U28398 ( .A(n28163), .Z(n28159) );
  XOR U28399 ( .A(n28216), .B(n28217), .Z(n28163) );
  ANDN U28400 ( .B(n28218), .A(n28219), .Z(n28216) );
  XOR U28401 ( .A(n28220), .B(n28217), .Z(n28218) );
  XOR U28402 ( .A(n28174), .B(n28027), .Z(n28175) );
  XOR U28403 ( .A(n28221), .B(n28222), .Z(n28027) );
  AND U28404 ( .A(n336), .B(n28223), .Z(n28221) );
  XOR U28405 ( .A(n28224), .B(n28222), .Z(n28223) );
  XNOR U28406 ( .A(n28225), .B(n28226), .Z(n28174) );
  NAND U28407 ( .A(n28227), .B(n28228), .Z(n28226) );
  XOR U28408 ( .A(n28229), .B(n28126), .Z(n28228) );
  XOR U28409 ( .A(n28202), .B(n28203), .Z(n28126) );
  XOR U28410 ( .A(n28230), .B(n28195), .Z(n28203) );
  XOR U28411 ( .A(n28231), .B(n28183), .Z(n28195) );
  XOR U28412 ( .A(n28232), .B(n28233), .Z(n28183) );
  ANDN U28413 ( .B(n28234), .A(n28235), .Z(n28232) );
  XOR U28414 ( .A(n28233), .B(n28236), .Z(n28234) );
  IV U28415 ( .A(n28181), .Z(n28231) );
  XOR U28416 ( .A(n28179), .B(n28237), .Z(n28181) );
  XOR U28417 ( .A(n28238), .B(n28239), .Z(n28237) );
  ANDN U28418 ( .B(n28240), .A(n28241), .Z(n28238) );
  XOR U28419 ( .A(n28242), .B(n28239), .Z(n28240) );
  IV U28420 ( .A(n28182), .Z(n28179) );
  XOR U28421 ( .A(n28243), .B(n28244), .Z(n28182) );
  ANDN U28422 ( .B(n28245), .A(n28246), .Z(n28243) );
  XOR U28423 ( .A(n28244), .B(n28247), .Z(n28245) );
  IV U28424 ( .A(n28194), .Z(n28230) );
  XOR U28425 ( .A(n28248), .B(n28249), .Z(n28194) );
  XNOR U28426 ( .A(n28189), .B(n28250), .Z(n28249) );
  IV U28427 ( .A(n28192), .Z(n28250) );
  XOR U28428 ( .A(n28251), .B(n28252), .Z(n28192) );
  ANDN U28429 ( .B(n28253), .A(n28254), .Z(n28251) );
  XOR U28430 ( .A(n28252), .B(n28255), .Z(n28253) );
  XNOR U28431 ( .A(n28256), .B(n28257), .Z(n28189) );
  ANDN U28432 ( .B(n28258), .A(n28259), .Z(n28256) );
  XOR U28433 ( .A(n28257), .B(n28260), .Z(n28258) );
  IV U28434 ( .A(n28188), .Z(n28248) );
  XOR U28435 ( .A(n28186), .B(n28261), .Z(n28188) );
  XOR U28436 ( .A(n28262), .B(n28263), .Z(n28261) );
  ANDN U28437 ( .B(n28264), .A(n28265), .Z(n28262) );
  XOR U28438 ( .A(n28266), .B(n28263), .Z(n28264) );
  IV U28439 ( .A(n28190), .Z(n28186) );
  XOR U28440 ( .A(n28267), .B(n28268), .Z(n28190) );
  ANDN U28441 ( .B(n28269), .A(n28270), .Z(n28267) );
  XOR U28442 ( .A(n28271), .B(n28268), .Z(n28269) );
  XOR U28443 ( .A(n28272), .B(n28273), .Z(n28202) );
  XOR U28444 ( .A(n28220), .B(n28274), .Z(n28273) );
  IV U28445 ( .A(n28200), .Z(n28274) );
  XOR U28446 ( .A(n28275), .B(n28276), .Z(n28200) );
  ANDN U28447 ( .B(n28277), .A(n28278), .Z(n28275) );
  XOR U28448 ( .A(n28276), .B(n28279), .Z(n28277) );
  XOR U28449 ( .A(n28280), .B(n28208), .Z(n28220) );
  XOR U28450 ( .A(n28281), .B(n28282), .Z(n28208) );
  ANDN U28451 ( .B(n28283), .A(n28284), .Z(n28281) );
  XOR U28452 ( .A(n28282), .B(n28285), .Z(n28283) );
  IV U28453 ( .A(n28207), .Z(n28280) );
  XOR U28454 ( .A(n28286), .B(n28287), .Z(n28207) );
  XOR U28455 ( .A(n28288), .B(n28289), .Z(n28287) );
  ANDN U28456 ( .B(n28290), .A(n28291), .Z(n28288) );
  XOR U28457 ( .A(n28292), .B(n28289), .Z(n28290) );
  IV U28458 ( .A(n28205), .Z(n28286) );
  XOR U28459 ( .A(n28293), .B(n28294), .Z(n28205) );
  ANDN U28460 ( .B(n28295), .A(n28296), .Z(n28293) );
  XOR U28461 ( .A(n28294), .B(n28297), .Z(n28295) );
  IV U28462 ( .A(n28219), .Z(n28272) );
  XOR U28463 ( .A(n28298), .B(n28299), .Z(n28219) );
  XNOR U28464 ( .A(n28214), .B(n28300), .Z(n28299) );
  IV U28465 ( .A(n28217), .Z(n28300) );
  XOR U28466 ( .A(n28301), .B(n28302), .Z(n28217) );
  ANDN U28467 ( .B(n28303), .A(n28304), .Z(n28301) );
  XOR U28468 ( .A(n28305), .B(n28302), .Z(n28303) );
  XNOR U28469 ( .A(n28306), .B(n28307), .Z(n28214) );
  ANDN U28470 ( .B(n28308), .A(n28309), .Z(n28306) );
  XOR U28471 ( .A(n28307), .B(n28310), .Z(n28308) );
  IV U28472 ( .A(n28213), .Z(n28298) );
  XOR U28473 ( .A(n28211), .B(n28311), .Z(n28213) );
  XOR U28474 ( .A(n28312), .B(n28313), .Z(n28311) );
  ANDN U28475 ( .B(n28314), .A(n28315), .Z(n28312) );
  XOR U28476 ( .A(n28316), .B(n28313), .Z(n28314) );
  IV U28477 ( .A(n28215), .Z(n28211) );
  XOR U28478 ( .A(n28317), .B(n28318), .Z(n28215) );
  ANDN U28479 ( .B(n28319), .A(n28320), .Z(n28317) );
  XOR U28480 ( .A(n28321), .B(n28318), .Z(n28319) );
  IV U28481 ( .A(n28225), .Z(n28229) );
  XOR U28482 ( .A(n28225), .B(n28128), .Z(n28227) );
  XOR U28483 ( .A(n28322), .B(n28323), .Z(n28128) );
  AND U28484 ( .A(n336), .B(n28324), .Z(n28322) );
  XOR U28485 ( .A(n28325), .B(n28323), .Z(n28324) );
  NANDN U28486 ( .A(n28130), .B(n28132), .Z(n28225) );
  XOR U28487 ( .A(n28326), .B(n28327), .Z(n28132) );
  AND U28488 ( .A(n336), .B(n28328), .Z(n28326) );
  XOR U28489 ( .A(n28327), .B(n28329), .Z(n28328) );
  XNOR U28490 ( .A(n28330), .B(n28331), .Z(n336) );
  AND U28491 ( .A(n28332), .B(n28333), .Z(n28330) );
  XOR U28492 ( .A(n28331), .B(n28143), .Z(n28333) );
  XNOR U28493 ( .A(n28334), .B(n28335), .Z(n28143) );
  ANDN U28494 ( .B(n28336), .A(n28337), .Z(n28334) );
  XOR U28495 ( .A(n28335), .B(n28338), .Z(n28336) );
  XNOR U28496 ( .A(n28331), .B(n28145), .Z(n28332) );
  XOR U28497 ( .A(n28339), .B(n28340), .Z(n28145) );
  AND U28498 ( .A(n340), .B(n28341), .Z(n28339) );
  XOR U28499 ( .A(n28342), .B(n28340), .Z(n28341) );
  XOR U28500 ( .A(n28343), .B(n28344), .Z(n28331) );
  AND U28501 ( .A(n28345), .B(n28346), .Z(n28343) );
  XOR U28502 ( .A(n28344), .B(n28170), .Z(n28346) );
  XOR U28503 ( .A(n28337), .B(n28338), .Z(n28170) );
  XNOR U28504 ( .A(n28347), .B(n28348), .Z(n28338) );
  ANDN U28505 ( .B(n28349), .A(n28350), .Z(n28347) );
  XOR U28506 ( .A(n28351), .B(n28352), .Z(n28349) );
  XOR U28507 ( .A(n28353), .B(n28354), .Z(n28337) );
  XNOR U28508 ( .A(n28355), .B(n28356), .Z(n28354) );
  ANDN U28509 ( .B(n28357), .A(n28358), .Z(n28355) );
  XNOR U28510 ( .A(n28359), .B(n28360), .Z(n28357) );
  IV U28511 ( .A(n28335), .Z(n28353) );
  XOR U28512 ( .A(n28361), .B(n28362), .Z(n28335) );
  ANDN U28513 ( .B(n28363), .A(n28364), .Z(n28361) );
  XOR U28514 ( .A(n28362), .B(n28365), .Z(n28363) );
  XNOR U28515 ( .A(n28344), .B(n28172), .Z(n28345) );
  XOR U28516 ( .A(n28366), .B(n28367), .Z(n28172) );
  AND U28517 ( .A(n340), .B(n28368), .Z(n28366) );
  XOR U28518 ( .A(n28369), .B(n28367), .Z(n28368) );
  XNOR U28519 ( .A(n28370), .B(n28371), .Z(n28344) );
  AND U28520 ( .A(n28372), .B(n28373), .Z(n28370) );
  XNOR U28521 ( .A(n28371), .B(n28222), .Z(n28373) );
  XOR U28522 ( .A(n28364), .B(n28365), .Z(n28222) );
  XOR U28523 ( .A(n28374), .B(n28352), .Z(n28365) );
  XNOR U28524 ( .A(n28375), .B(n28376), .Z(n28352) );
  ANDN U28525 ( .B(n28377), .A(n28378), .Z(n28375) );
  XOR U28526 ( .A(n28379), .B(n28380), .Z(n28377) );
  IV U28527 ( .A(n28350), .Z(n28374) );
  XOR U28528 ( .A(n28348), .B(n28381), .Z(n28350) );
  XNOR U28529 ( .A(n28382), .B(n28383), .Z(n28381) );
  ANDN U28530 ( .B(n28384), .A(n28385), .Z(n28382) );
  XNOR U28531 ( .A(n28386), .B(n28387), .Z(n28384) );
  IV U28532 ( .A(n28351), .Z(n28348) );
  XOR U28533 ( .A(n28388), .B(n28389), .Z(n28351) );
  ANDN U28534 ( .B(n28390), .A(n28391), .Z(n28388) );
  XOR U28535 ( .A(n28389), .B(n28392), .Z(n28390) );
  XOR U28536 ( .A(n28393), .B(n28394), .Z(n28364) );
  XNOR U28537 ( .A(n28359), .B(n28395), .Z(n28394) );
  IV U28538 ( .A(n28362), .Z(n28395) );
  XOR U28539 ( .A(n28396), .B(n28397), .Z(n28362) );
  ANDN U28540 ( .B(n28398), .A(n28399), .Z(n28396) );
  XOR U28541 ( .A(n28397), .B(n28400), .Z(n28398) );
  XNOR U28542 ( .A(n28401), .B(n28402), .Z(n28359) );
  ANDN U28543 ( .B(n28403), .A(n28404), .Z(n28401) );
  XOR U28544 ( .A(n28402), .B(n28405), .Z(n28403) );
  IV U28545 ( .A(n28358), .Z(n28393) );
  XOR U28546 ( .A(n28356), .B(n28406), .Z(n28358) );
  XNOR U28547 ( .A(n28407), .B(n28408), .Z(n28406) );
  ANDN U28548 ( .B(n28409), .A(n28410), .Z(n28407) );
  XNOR U28549 ( .A(n28411), .B(n28412), .Z(n28409) );
  IV U28550 ( .A(n28360), .Z(n28356) );
  XOR U28551 ( .A(n28413), .B(n28414), .Z(n28360) );
  ANDN U28552 ( .B(n28415), .A(n28416), .Z(n28413) );
  XOR U28553 ( .A(n28417), .B(n28414), .Z(n28415) );
  XOR U28554 ( .A(n28371), .B(n28224), .Z(n28372) );
  XOR U28555 ( .A(n28418), .B(n28419), .Z(n28224) );
  AND U28556 ( .A(n340), .B(n28420), .Z(n28418) );
  XOR U28557 ( .A(n28421), .B(n28419), .Z(n28420) );
  XNOR U28558 ( .A(n28422), .B(n28423), .Z(n28371) );
  NAND U28559 ( .A(n28424), .B(n28425), .Z(n28423) );
  XOR U28560 ( .A(n28426), .B(n28323), .Z(n28425) );
  XOR U28561 ( .A(n28399), .B(n28400), .Z(n28323) );
  XOR U28562 ( .A(n28427), .B(n28392), .Z(n28400) );
  XOR U28563 ( .A(n28428), .B(n28380), .Z(n28392) );
  XOR U28564 ( .A(n28429), .B(n28430), .Z(n28380) );
  ANDN U28565 ( .B(n28431), .A(n28432), .Z(n28429) );
  XOR U28566 ( .A(n28430), .B(n28433), .Z(n28431) );
  IV U28567 ( .A(n28378), .Z(n28428) );
  XOR U28568 ( .A(n28376), .B(n28434), .Z(n28378) );
  XOR U28569 ( .A(n28435), .B(n28436), .Z(n28434) );
  ANDN U28570 ( .B(n28437), .A(n28438), .Z(n28435) );
  XOR U28571 ( .A(n28439), .B(n28436), .Z(n28437) );
  IV U28572 ( .A(n28379), .Z(n28376) );
  XOR U28573 ( .A(n28440), .B(n28441), .Z(n28379) );
  ANDN U28574 ( .B(n28442), .A(n28443), .Z(n28440) );
  XOR U28575 ( .A(n28441), .B(n28444), .Z(n28442) );
  IV U28576 ( .A(n28391), .Z(n28427) );
  XOR U28577 ( .A(n28445), .B(n28446), .Z(n28391) );
  XNOR U28578 ( .A(n28386), .B(n28447), .Z(n28446) );
  IV U28579 ( .A(n28389), .Z(n28447) );
  XOR U28580 ( .A(n28448), .B(n28449), .Z(n28389) );
  ANDN U28581 ( .B(n28450), .A(n28451), .Z(n28448) );
  XOR U28582 ( .A(n28449), .B(n28452), .Z(n28450) );
  XNOR U28583 ( .A(n28453), .B(n28454), .Z(n28386) );
  ANDN U28584 ( .B(n28455), .A(n28456), .Z(n28453) );
  XOR U28585 ( .A(n28454), .B(n28457), .Z(n28455) );
  IV U28586 ( .A(n28385), .Z(n28445) );
  XOR U28587 ( .A(n28383), .B(n28458), .Z(n28385) );
  XOR U28588 ( .A(n28459), .B(n28460), .Z(n28458) );
  ANDN U28589 ( .B(n28461), .A(n28462), .Z(n28459) );
  XOR U28590 ( .A(n28463), .B(n28460), .Z(n28461) );
  IV U28591 ( .A(n28387), .Z(n28383) );
  XOR U28592 ( .A(n28464), .B(n28465), .Z(n28387) );
  ANDN U28593 ( .B(n28466), .A(n28467), .Z(n28464) );
  XOR U28594 ( .A(n28468), .B(n28465), .Z(n28466) );
  XOR U28595 ( .A(n28469), .B(n28470), .Z(n28399) );
  XOR U28596 ( .A(n28417), .B(n28471), .Z(n28470) );
  IV U28597 ( .A(n28397), .Z(n28471) );
  XOR U28598 ( .A(n28472), .B(n28473), .Z(n28397) );
  ANDN U28599 ( .B(n28474), .A(n28475), .Z(n28472) );
  XOR U28600 ( .A(n28473), .B(n28476), .Z(n28474) );
  XOR U28601 ( .A(n28477), .B(n28405), .Z(n28417) );
  XOR U28602 ( .A(n28478), .B(n28479), .Z(n28405) );
  ANDN U28603 ( .B(n28480), .A(n28481), .Z(n28478) );
  XOR U28604 ( .A(n28479), .B(n28482), .Z(n28480) );
  IV U28605 ( .A(n28404), .Z(n28477) );
  XOR U28606 ( .A(n28483), .B(n28484), .Z(n28404) );
  XOR U28607 ( .A(n28485), .B(n28486), .Z(n28484) );
  ANDN U28608 ( .B(n28487), .A(n28488), .Z(n28485) );
  XOR U28609 ( .A(n28489), .B(n28486), .Z(n28487) );
  IV U28610 ( .A(n28402), .Z(n28483) );
  XOR U28611 ( .A(n28490), .B(n28491), .Z(n28402) );
  ANDN U28612 ( .B(n28492), .A(n28493), .Z(n28490) );
  XOR U28613 ( .A(n28491), .B(n28494), .Z(n28492) );
  IV U28614 ( .A(n28416), .Z(n28469) );
  XOR U28615 ( .A(n28495), .B(n28496), .Z(n28416) );
  XNOR U28616 ( .A(n28411), .B(n28497), .Z(n28496) );
  IV U28617 ( .A(n28414), .Z(n28497) );
  XOR U28618 ( .A(n28498), .B(n28499), .Z(n28414) );
  ANDN U28619 ( .B(n28500), .A(n28501), .Z(n28498) );
  XOR U28620 ( .A(n28502), .B(n28499), .Z(n28500) );
  XNOR U28621 ( .A(n28503), .B(n28504), .Z(n28411) );
  ANDN U28622 ( .B(n28505), .A(n28506), .Z(n28503) );
  XOR U28623 ( .A(n28504), .B(n28507), .Z(n28505) );
  IV U28624 ( .A(n28410), .Z(n28495) );
  XOR U28625 ( .A(n28408), .B(n28508), .Z(n28410) );
  XOR U28626 ( .A(n28509), .B(n28510), .Z(n28508) );
  ANDN U28627 ( .B(n28511), .A(n28512), .Z(n28509) );
  XOR U28628 ( .A(n28513), .B(n28510), .Z(n28511) );
  IV U28629 ( .A(n28412), .Z(n28408) );
  XOR U28630 ( .A(n28514), .B(n28515), .Z(n28412) );
  ANDN U28631 ( .B(n28516), .A(n28517), .Z(n28514) );
  XOR U28632 ( .A(n28518), .B(n28515), .Z(n28516) );
  IV U28633 ( .A(n28422), .Z(n28426) );
  XOR U28634 ( .A(n28422), .B(n28325), .Z(n28424) );
  XOR U28635 ( .A(n28519), .B(n28520), .Z(n28325) );
  AND U28636 ( .A(n340), .B(n28521), .Z(n28519) );
  XOR U28637 ( .A(n28522), .B(n28520), .Z(n28521) );
  NANDN U28638 ( .A(n28327), .B(n28329), .Z(n28422) );
  XOR U28639 ( .A(n28523), .B(n28524), .Z(n28329) );
  AND U28640 ( .A(n340), .B(n28525), .Z(n28523) );
  XOR U28641 ( .A(n28524), .B(n28526), .Z(n28525) );
  XNOR U28642 ( .A(n28527), .B(n28528), .Z(n340) );
  AND U28643 ( .A(n28529), .B(n28530), .Z(n28527) );
  XOR U28644 ( .A(n28528), .B(n28340), .Z(n28530) );
  XNOR U28645 ( .A(n28531), .B(n28532), .Z(n28340) );
  ANDN U28646 ( .B(n28533), .A(n28534), .Z(n28531) );
  XOR U28647 ( .A(n28532), .B(n28535), .Z(n28533) );
  XNOR U28648 ( .A(n28528), .B(n28342), .Z(n28529) );
  XOR U28649 ( .A(n28536), .B(n28537), .Z(n28342) );
  AND U28650 ( .A(n344), .B(n28538), .Z(n28536) );
  XOR U28651 ( .A(n28539), .B(n28537), .Z(n28538) );
  XOR U28652 ( .A(n28540), .B(n28541), .Z(n28528) );
  AND U28653 ( .A(n28542), .B(n28543), .Z(n28540) );
  XOR U28654 ( .A(n28541), .B(n28367), .Z(n28543) );
  XOR U28655 ( .A(n28534), .B(n28535), .Z(n28367) );
  XNOR U28656 ( .A(n28544), .B(n28545), .Z(n28535) );
  ANDN U28657 ( .B(n28546), .A(n28547), .Z(n28544) );
  XOR U28658 ( .A(n28548), .B(n28549), .Z(n28546) );
  XOR U28659 ( .A(n28550), .B(n28551), .Z(n28534) );
  XNOR U28660 ( .A(n28552), .B(n28553), .Z(n28551) );
  ANDN U28661 ( .B(n28554), .A(n28555), .Z(n28552) );
  XNOR U28662 ( .A(n28556), .B(n28557), .Z(n28554) );
  IV U28663 ( .A(n28532), .Z(n28550) );
  XOR U28664 ( .A(n28558), .B(n28559), .Z(n28532) );
  ANDN U28665 ( .B(n28560), .A(n28561), .Z(n28558) );
  XOR U28666 ( .A(n28559), .B(n28562), .Z(n28560) );
  XNOR U28667 ( .A(n28541), .B(n28369), .Z(n28542) );
  XOR U28668 ( .A(n28563), .B(n28564), .Z(n28369) );
  AND U28669 ( .A(n344), .B(n28565), .Z(n28563) );
  XOR U28670 ( .A(n28566), .B(n28564), .Z(n28565) );
  XNOR U28671 ( .A(n28567), .B(n28568), .Z(n28541) );
  AND U28672 ( .A(n28569), .B(n28570), .Z(n28567) );
  XNOR U28673 ( .A(n28568), .B(n28419), .Z(n28570) );
  XOR U28674 ( .A(n28561), .B(n28562), .Z(n28419) );
  XOR U28675 ( .A(n28571), .B(n28549), .Z(n28562) );
  XNOR U28676 ( .A(n28572), .B(n28573), .Z(n28549) );
  ANDN U28677 ( .B(n28574), .A(n28575), .Z(n28572) );
  XOR U28678 ( .A(n28576), .B(n28577), .Z(n28574) );
  IV U28679 ( .A(n28547), .Z(n28571) );
  XOR U28680 ( .A(n28545), .B(n28578), .Z(n28547) );
  XNOR U28681 ( .A(n28579), .B(n28580), .Z(n28578) );
  ANDN U28682 ( .B(n28581), .A(n28582), .Z(n28579) );
  XNOR U28683 ( .A(n28583), .B(n28584), .Z(n28581) );
  IV U28684 ( .A(n28548), .Z(n28545) );
  XOR U28685 ( .A(n28585), .B(n28586), .Z(n28548) );
  ANDN U28686 ( .B(n28587), .A(n28588), .Z(n28585) );
  XOR U28687 ( .A(n28586), .B(n28589), .Z(n28587) );
  XOR U28688 ( .A(n28590), .B(n28591), .Z(n28561) );
  XNOR U28689 ( .A(n28556), .B(n28592), .Z(n28591) );
  IV U28690 ( .A(n28559), .Z(n28592) );
  XOR U28691 ( .A(n28593), .B(n28594), .Z(n28559) );
  ANDN U28692 ( .B(n28595), .A(n28596), .Z(n28593) );
  XOR U28693 ( .A(n28594), .B(n28597), .Z(n28595) );
  XNOR U28694 ( .A(n28598), .B(n28599), .Z(n28556) );
  ANDN U28695 ( .B(n28600), .A(n28601), .Z(n28598) );
  XOR U28696 ( .A(n28599), .B(n28602), .Z(n28600) );
  IV U28697 ( .A(n28555), .Z(n28590) );
  XOR U28698 ( .A(n28553), .B(n28603), .Z(n28555) );
  XNOR U28699 ( .A(n28604), .B(n28605), .Z(n28603) );
  ANDN U28700 ( .B(n28606), .A(n28607), .Z(n28604) );
  XNOR U28701 ( .A(n28608), .B(n28609), .Z(n28606) );
  IV U28702 ( .A(n28557), .Z(n28553) );
  XOR U28703 ( .A(n28610), .B(n28611), .Z(n28557) );
  ANDN U28704 ( .B(n28612), .A(n28613), .Z(n28610) );
  XOR U28705 ( .A(n28614), .B(n28611), .Z(n28612) );
  XOR U28706 ( .A(n28568), .B(n28421), .Z(n28569) );
  XOR U28707 ( .A(n28615), .B(n28616), .Z(n28421) );
  AND U28708 ( .A(n344), .B(n28617), .Z(n28615) );
  XOR U28709 ( .A(n28618), .B(n28616), .Z(n28617) );
  XNOR U28710 ( .A(n28619), .B(n28620), .Z(n28568) );
  NAND U28711 ( .A(n28621), .B(n28622), .Z(n28620) );
  XOR U28712 ( .A(n28623), .B(n28520), .Z(n28622) );
  XOR U28713 ( .A(n28596), .B(n28597), .Z(n28520) );
  XOR U28714 ( .A(n28624), .B(n28589), .Z(n28597) );
  XOR U28715 ( .A(n28625), .B(n28577), .Z(n28589) );
  XOR U28716 ( .A(n28626), .B(n28627), .Z(n28577) );
  ANDN U28717 ( .B(n28628), .A(n28629), .Z(n28626) );
  XOR U28718 ( .A(n28627), .B(n28630), .Z(n28628) );
  IV U28719 ( .A(n28575), .Z(n28625) );
  XOR U28720 ( .A(n28573), .B(n28631), .Z(n28575) );
  XOR U28721 ( .A(n28632), .B(n28633), .Z(n28631) );
  ANDN U28722 ( .B(n28634), .A(n28635), .Z(n28632) );
  XOR U28723 ( .A(n28636), .B(n28633), .Z(n28634) );
  IV U28724 ( .A(n28576), .Z(n28573) );
  XOR U28725 ( .A(n28637), .B(n28638), .Z(n28576) );
  ANDN U28726 ( .B(n28639), .A(n28640), .Z(n28637) );
  XOR U28727 ( .A(n28638), .B(n28641), .Z(n28639) );
  IV U28728 ( .A(n28588), .Z(n28624) );
  XOR U28729 ( .A(n28642), .B(n28643), .Z(n28588) );
  XNOR U28730 ( .A(n28583), .B(n28644), .Z(n28643) );
  IV U28731 ( .A(n28586), .Z(n28644) );
  XOR U28732 ( .A(n28645), .B(n28646), .Z(n28586) );
  ANDN U28733 ( .B(n28647), .A(n28648), .Z(n28645) );
  XOR U28734 ( .A(n28646), .B(n28649), .Z(n28647) );
  XNOR U28735 ( .A(n28650), .B(n28651), .Z(n28583) );
  ANDN U28736 ( .B(n28652), .A(n28653), .Z(n28650) );
  XOR U28737 ( .A(n28651), .B(n28654), .Z(n28652) );
  IV U28738 ( .A(n28582), .Z(n28642) );
  XOR U28739 ( .A(n28580), .B(n28655), .Z(n28582) );
  XOR U28740 ( .A(n28656), .B(n28657), .Z(n28655) );
  ANDN U28741 ( .B(n28658), .A(n28659), .Z(n28656) );
  XOR U28742 ( .A(n28660), .B(n28657), .Z(n28658) );
  IV U28743 ( .A(n28584), .Z(n28580) );
  XOR U28744 ( .A(n28661), .B(n28662), .Z(n28584) );
  ANDN U28745 ( .B(n28663), .A(n28664), .Z(n28661) );
  XOR U28746 ( .A(n28665), .B(n28662), .Z(n28663) );
  XOR U28747 ( .A(n28666), .B(n28667), .Z(n28596) );
  XOR U28748 ( .A(n28614), .B(n28668), .Z(n28667) );
  IV U28749 ( .A(n28594), .Z(n28668) );
  XOR U28750 ( .A(n28669), .B(n28670), .Z(n28594) );
  ANDN U28751 ( .B(n28671), .A(n28672), .Z(n28669) );
  XOR U28752 ( .A(n28670), .B(n28673), .Z(n28671) );
  XOR U28753 ( .A(n28674), .B(n28602), .Z(n28614) );
  XOR U28754 ( .A(n28675), .B(n28676), .Z(n28602) );
  ANDN U28755 ( .B(n28677), .A(n28678), .Z(n28675) );
  XOR U28756 ( .A(n28676), .B(n28679), .Z(n28677) );
  IV U28757 ( .A(n28601), .Z(n28674) );
  XOR U28758 ( .A(n28680), .B(n28681), .Z(n28601) );
  XOR U28759 ( .A(n28682), .B(n28683), .Z(n28681) );
  ANDN U28760 ( .B(n28684), .A(n28685), .Z(n28682) );
  XOR U28761 ( .A(n28686), .B(n28683), .Z(n28684) );
  IV U28762 ( .A(n28599), .Z(n28680) );
  XOR U28763 ( .A(n28687), .B(n28688), .Z(n28599) );
  ANDN U28764 ( .B(n28689), .A(n28690), .Z(n28687) );
  XOR U28765 ( .A(n28688), .B(n28691), .Z(n28689) );
  IV U28766 ( .A(n28613), .Z(n28666) );
  XOR U28767 ( .A(n28692), .B(n28693), .Z(n28613) );
  XNOR U28768 ( .A(n28608), .B(n28694), .Z(n28693) );
  IV U28769 ( .A(n28611), .Z(n28694) );
  XOR U28770 ( .A(n28695), .B(n28696), .Z(n28611) );
  ANDN U28771 ( .B(n28697), .A(n28698), .Z(n28695) );
  XOR U28772 ( .A(n28699), .B(n28696), .Z(n28697) );
  XNOR U28773 ( .A(n28700), .B(n28701), .Z(n28608) );
  ANDN U28774 ( .B(n28702), .A(n28703), .Z(n28700) );
  XOR U28775 ( .A(n28701), .B(n28704), .Z(n28702) );
  IV U28776 ( .A(n28607), .Z(n28692) );
  XOR U28777 ( .A(n28605), .B(n28705), .Z(n28607) );
  XOR U28778 ( .A(n28706), .B(n28707), .Z(n28705) );
  ANDN U28779 ( .B(n28708), .A(n28709), .Z(n28706) );
  XOR U28780 ( .A(n28710), .B(n28707), .Z(n28708) );
  IV U28781 ( .A(n28609), .Z(n28605) );
  XOR U28782 ( .A(n28711), .B(n28712), .Z(n28609) );
  ANDN U28783 ( .B(n28713), .A(n28714), .Z(n28711) );
  XOR U28784 ( .A(n28715), .B(n28712), .Z(n28713) );
  IV U28785 ( .A(n28619), .Z(n28623) );
  XOR U28786 ( .A(n28619), .B(n28522), .Z(n28621) );
  XOR U28787 ( .A(n28716), .B(n28717), .Z(n28522) );
  AND U28788 ( .A(n344), .B(n28718), .Z(n28716) );
  XOR U28789 ( .A(n28719), .B(n28717), .Z(n28718) );
  NANDN U28790 ( .A(n28524), .B(n28526), .Z(n28619) );
  XOR U28791 ( .A(n28720), .B(n28721), .Z(n28526) );
  AND U28792 ( .A(n344), .B(n28722), .Z(n28720) );
  XOR U28793 ( .A(n28721), .B(n28723), .Z(n28722) );
  XNOR U28794 ( .A(n28724), .B(n28725), .Z(n344) );
  AND U28795 ( .A(n28726), .B(n28727), .Z(n28724) );
  XOR U28796 ( .A(n28725), .B(n28537), .Z(n28727) );
  XNOR U28797 ( .A(n28728), .B(n28729), .Z(n28537) );
  ANDN U28798 ( .B(n28730), .A(n28731), .Z(n28728) );
  XOR U28799 ( .A(n28729), .B(n28732), .Z(n28730) );
  XNOR U28800 ( .A(n28725), .B(n28539), .Z(n28726) );
  XOR U28801 ( .A(n28733), .B(n28734), .Z(n28539) );
  AND U28802 ( .A(n348), .B(n28735), .Z(n28733) );
  XOR U28803 ( .A(n28736), .B(n28734), .Z(n28735) );
  XOR U28804 ( .A(n28737), .B(n28738), .Z(n28725) );
  AND U28805 ( .A(n28739), .B(n28740), .Z(n28737) );
  XOR U28806 ( .A(n28738), .B(n28564), .Z(n28740) );
  XOR U28807 ( .A(n28731), .B(n28732), .Z(n28564) );
  XNOR U28808 ( .A(n28741), .B(n28742), .Z(n28732) );
  ANDN U28809 ( .B(n28743), .A(n28744), .Z(n28741) );
  XOR U28810 ( .A(n28745), .B(n28746), .Z(n28743) );
  XOR U28811 ( .A(n28747), .B(n28748), .Z(n28731) );
  XNOR U28812 ( .A(n28749), .B(n28750), .Z(n28748) );
  ANDN U28813 ( .B(n28751), .A(n28752), .Z(n28749) );
  XNOR U28814 ( .A(n28753), .B(n28754), .Z(n28751) );
  IV U28815 ( .A(n28729), .Z(n28747) );
  XOR U28816 ( .A(n28755), .B(n28756), .Z(n28729) );
  ANDN U28817 ( .B(n28757), .A(n28758), .Z(n28755) );
  XOR U28818 ( .A(n28756), .B(n28759), .Z(n28757) );
  XNOR U28819 ( .A(n28738), .B(n28566), .Z(n28739) );
  XOR U28820 ( .A(n28760), .B(n28761), .Z(n28566) );
  AND U28821 ( .A(n348), .B(n28762), .Z(n28760) );
  XOR U28822 ( .A(n28763), .B(n28761), .Z(n28762) );
  XNOR U28823 ( .A(n28764), .B(n28765), .Z(n28738) );
  AND U28824 ( .A(n28766), .B(n28767), .Z(n28764) );
  XNOR U28825 ( .A(n28765), .B(n28616), .Z(n28767) );
  XOR U28826 ( .A(n28758), .B(n28759), .Z(n28616) );
  XOR U28827 ( .A(n28768), .B(n28746), .Z(n28759) );
  XNOR U28828 ( .A(n28769), .B(n28770), .Z(n28746) );
  ANDN U28829 ( .B(n28771), .A(n28772), .Z(n28769) );
  XOR U28830 ( .A(n28773), .B(n28774), .Z(n28771) );
  IV U28831 ( .A(n28744), .Z(n28768) );
  XOR U28832 ( .A(n28742), .B(n28775), .Z(n28744) );
  XNOR U28833 ( .A(n28776), .B(n28777), .Z(n28775) );
  ANDN U28834 ( .B(n28778), .A(n28779), .Z(n28776) );
  XNOR U28835 ( .A(n28780), .B(n28781), .Z(n28778) );
  IV U28836 ( .A(n28745), .Z(n28742) );
  XOR U28837 ( .A(n28782), .B(n28783), .Z(n28745) );
  ANDN U28838 ( .B(n28784), .A(n28785), .Z(n28782) );
  XOR U28839 ( .A(n28783), .B(n28786), .Z(n28784) );
  XOR U28840 ( .A(n28787), .B(n28788), .Z(n28758) );
  XNOR U28841 ( .A(n28753), .B(n28789), .Z(n28788) );
  IV U28842 ( .A(n28756), .Z(n28789) );
  XOR U28843 ( .A(n28790), .B(n28791), .Z(n28756) );
  ANDN U28844 ( .B(n28792), .A(n28793), .Z(n28790) );
  XOR U28845 ( .A(n28791), .B(n28794), .Z(n28792) );
  XNOR U28846 ( .A(n28795), .B(n28796), .Z(n28753) );
  ANDN U28847 ( .B(n28797), .A(n28798), .Z(n28795) );
  XOR U28848 ( .A(n28796), .B(n28799), .Z(n28797) );
  IV U28849 ( .A(n28752), .Z(n28787) );
  XOR U28850 ( .A(n28750), .B(n28800), .Z(n28752) );
  XNOR U28851 ( .A(n28801), .B(n28802), .Z(n28800) );
  ANDN U28852 ( .B(n28803), .A(n28804), .Z(n28801) );
  XNOR U28853 ( .A(n28805), .B(n28806), .Z(n28803) );
  IV U28854 ( .A(n28754), .Z(n28750) );
  XOR U28855 ( .A(n28807), .B(n28808), .Z(n28754) );
  ANDN U28856 ( .B(n28809), .A(n28810), .Z(n28807) );
  XOR U28857 ( .A(n28811), .B(n28808), .Z(n28809) );
  XOR U28858 ( .A(n28765), .B(n28618), .Z(n28766) );
  XOR U28859 ( .A(n28812), .B(n28813), .Z(n28618) );
  AND U28860 ( .A(n348), .B(n28814), .Z(n28812) );
  XOR U28861 ( .A(n28815), .B(n28813), .Z(n28814) );
  XNOR U28862 ( .A(n28816), .B(n28817), .Z(n28765) );
  NAND U28863 ( .A(n28818), .B(n28819), .Z(n28817) );
  XOR U28864 ( .A(n28820), .B(n28717), .Z(n28819) );
  XOR U28865 ( .A(n28793), .B(n28794), .Z(n28717) );
  XOR U28866 ( .A(n28821), .B(n28786), .Z(n28794) );
  XOR U28867 ( .A(n28822), .B(n28774), .Z(n28786) );
  XOR U28868 ( .A(n28823), .B(n28824), .Z(n28774) );
  ANDN U28869 ( .B(n28825), .A(n28826), .Z(n28823) );
  XOR U28870 ( .A(n28824), .B(n28827), .Z(n28825) );
  IV U28871 ( .A(n28772), .Z(n28822) );
  XOR U28872 ( .A(n28770), .B(n28828), .Z(n28772) );
  XOR U28873 ( .A(n28829), .B(n28830), .Z(n28828) );
  ANDN U28874 ( .B(n28831), .A(n28832), .Z(n28829) );
  XOR U28875 ( .A(n28833), .B(n28830), .Z(n28831) );
  IV U28876 ( .A(n28773), .Z(n28770) );
  XOR U28877 ( .A(n28834), .B(n28835), .Z(n28773) );
  ANDN U28878 ( .B(n28836), .A(n28837), .Z(n28834) );
  XOR U28879 ( .A(n28835), .B(n28838), .Z(n28836) );
  IV U28880 ( .A(n28785), .Z(n28821) );
  XOR U28881 ( .A(n28839), .B(n28840), .Z(n28785) );
  XNOR U28882 ( .A(n28780), .B(n28841), .Z(n28840) );
  IV U28883 ( .A(n28783), .Z(n28841) );
  XOR U28884 ( .A(n28842), .B(n28843), .Z(n28783) );
  ANDN U28885 ( .B(n28844), .A(n28845), .Z(n28842) );
  XOR U28886 ( .A(n28843), .B(n28846), .Z(n28844) );
  XNOR U28887 ( .A(n28847), .B(n28848), .Z(n28780) );
  ANDN U28888 ( .B(n28849), .A(n28850), .Z(n28847) );
  XOR U28889 ( .A(n28848), .B(n28851), .Z(n28849) );
  IV U28890 ( .A(n28779), .Z(n28839) );
  XOR U28891 ( .A(n28777), .B(n28852), .Z(n28779) );
  XOR U28892 ( .A(n28853), .B(n28854), .Z(n28852) );
  ANDN U28893 ( .B(n28855), .A(n28856), .Z(n28853) );
  XOR U28894 ( .A(n28857), .B(n28854), .Z(n28855) );
  IV U28895 ( .A(n28781), .Z(n28777) );
  XOR U28896 ( .A(n28858), .B(n28859), .Z(n28781) );
  ANDN U28897 ( .B(n28860), .A(n28861), .Z(n28858) );
  XOR U28898 ( .A(n28862), .B(n28859), .Z(n28860) );
  XOR U28899 ( .A(n28863), .B(n28864), .Z(n28793) );
  XOR U28900 ( .A(n28811), .B(n28865), .Z(n28864) );
  IV U28901 ( .A(n28791), .Z(n28865) );
  XOR U28902 ( .A(n28866), .B(n28867), .Z(n28791) );
  ANDN U28903 ( .B(n28868), .A(n28869), .Z(n28866) );
  XOR U28904 ( .A(n28867), .B(n28870), .Z(n28868) );
  XOR U28905 ( .A(n28871), .B(n28799), .Z(n28811) );
  XOR U28906 ( .A(n28872), .B(n28873), .Z(n28799) );
  ANDN U28907 ( .B(n28874), .A(n28875), .Z(n28872) );
  XOR U28908 ( .A(n28873), .B(n28876), .Z(n28874) );
  IV U28909 ( .A(n28798), .Z(n28871) );
  XOR U28910 ( .A(n28877), .B(n28878), .Z(n28798) );
  XOR U28911 ( .A(n28879), .B(n28880), .Z(n28878) );
  ANDN U28912 ( .B(n28881), .A(n28882), .Z(n28879) );
  XOR U28913 ( .A(n28883), .B(n28880), .Z(n28881) );
  IV U28914 ( .A(n28796), .Z(n28877) );
  XOR U28915 ( .A(n28884), .B(n28885), .Z(n28796) );
  ANDN U28916 ( .B(n28886), .A(n28887), .Z(n28884) );
  XOR U28917 ( .A(n28885), .B(n28888), .Z(n28886) );
  IV U28918 ( .A(n28810), .Z(n28863) );
  XOR U28919 ( .A(n28889), .B(n28890), .Z(n28810) );
  XNOR U28920 ( .A(n28805), .B(n28891), .Z(n28890) );
  IV U28921 ( .A(n28808), .Z(n28891) );
  XOR U28922 ( .A(n28892), .B(n28893), .Z(n28808) );
  ANDN U28923 ( .B(n28894), .A(n28895), .Z(n28892) );
  XOR U28924 ( .A(n28896), .B(n28893), .Z(n28894) );
  XNOR U28925 ( .A(n28897), .B(n28898), .Z(n28805) );
  ANDN U28926 ( .B(n28899), .A(n28900), .Z(n28897) );
  XOR U28927 ( .A(n28898), .B(n28901), .Z(n28899) );
  IV U28928 ( .A(n28804), .Z(n28889) );
  XOR U28929 ( .A(n28802), .B(n28902), .Z(n28804) );
  XOR U28930 ( .A(n28903), .B(n28904), .Z(n28902) );
  ANDN U28931 ( .B(n28905), .A(n28906), .Z(n28903) );
  XOR U28932 ( .A(n28907), .B(n28904), .Z(n28905) );
  IV U28933 ( .A(n28806), .Z(n28802) );
  XOR U28934 ( .A(n28908), .B(n28909), .Z(n28806) );
  ANDN U28935 ( .B(n28910), .A(n28911), .Z(n28908) );
  XOR U28936 ( .A(n28912), .B(n28909), .Z(n28910) );
  IV U28937 ( .A(n28816), .Z(n28820) );
  XOR U28938 ( .A(n28816), .B(n28719), .Z(n28818) );
  XOR U28939 ( .A(n28913), .B(n28914), .Z(n28719) );
  AND U28940 ( .A(n348), .B(n28915), .Z(n28913) );
  XOR U28941 ( .A(n28916), .B(n28914), .Z(n28915) );
  NANDN U28942 ( .A(n28721), .B(n28723), .Z(n28816) );
  XOR U28943 ( .A(n28917), .B(n28918), .Z(n28723) );
  AND U28944 ( .A(n348), .B(n28919), .Z(n28917) );
  XOR U28945 ( .A(n28918), .B(n28920), .Z(n28919) );
  XNOR U28946 ( .A(n28921), .B(n28922), .Z(n348) );
  AND U28947 ( .A(n28923), .B(n28924), .Z(n28921) );
  XOR U28948 ( .A(n28922), .B(n28734), .Z(n28924) );
  XNOR U28949 ( .A(n28925), .B(n28926), .Z(n28734) );
  ANDN U28950 ( .B(n28927), .A(n28928), .Z(n28925) );
  XOR U28951 ( .A(n28926), .B(n28929), .Z(n28927) );
  XNOR U28952 ( .A(n28922), .B(n28736), .Z(n28923) );
  XOR U28953 ( .A(n28930), .B(n28931), .Z(n28736) );
  AND U28954 ( .A(n352), .B(n28932), .Z(n28930) );
  XOR U28955 ( .A(n28933), .B(n28931), .Z(n28932) );
  XOR U28956 ( .A(n28934), .B(n28935), .Z(n28922) );
  AND U28957 ( .A(n28936), .B(n28937), .Z(n28934) );
  XOR U28958 ( .A(n28935), .B(n28761), .Z(n28937) );
  XOR U28959 ( .A(n28928), .B(n28929), .Z(n28761) );
  XNOR U28960 ( .A(n28938), .B(n28939), .Z(n28929) );
  ANDN U28961 ( .B(n28940), .A(n28941), .Z(n28938) );
  XOR U28962 ( .A(n28942), .B(n28943), .Z(n28940) );
  XOR U28963 ( .A(n28944), .B(n28945), .Z(n28928) );
  XNOR U28964 ( .A(n28946), .B(n28947), .Z(n28945) );
  ANDN U28965 ( .B(n28948), .A(n28949), .Z(n28946) );
  XNOR U28966 ( .A(n28950), .B(n28951), .Z(n28948) );
  IV U28967 ( .A(n28926), .Z(n28944) );
  XOR U28968 ( .A(n28952), .B(n28953), .Z(n28926) );
  ANDN U28969 ( .B(n28954), .A(n28955), .Z(n28952) );
  XOR U28970 ( .A(n28953), .B(n28956), .Z(n28954) );
  XNOR U28971 ( .A(n28935), .B(n28763), .Z(n28936) );
  XOR U28972 ( .A(n28957), .B(n28958), .Z(n28763) );
  AND U28973 ( .A(n352), .B(n28959), .Z(n28957) );
  XOR U28974 ( .A(n28960), .B(n28958), .Z(n28959) );
  XNOR U28975 ( .A(n28961), .B(n28962), .Z(n28935) );
  AND U28976 ( .A(n28963), .B(n28964), .Z(n28961) );
  XNOR U28977 ( .A(n28962), .B(n28813), .Z(n28964) );
  XOR U28978 ( .A(n28955), .B(n28956), .Z(n28813) );
  XOR U28979 ( .A(n28965), .B(n28943), .Z(n28956) );
  XNOR U28980 ( .A(n28966), .B(n28967), .Z(n28943) );
  ANDN U28981 ( .B(n28968), .A(n28969), .Z(n28966) );
  XOR U28982 ( .A(n28970), .B(n28971), .Z(n28968) );
  IV U28983 ( .A(n28941), .Z(n28965) );
  XOR U28984 ( .A(n28939), .B(n28972), .Z(n28941) );
  XNOR U28985 ( .A(n28973), .B(n28974), .Z(n28972) );
  ANDN U28986 ( .B(n28975), .A(n28976), .Z(n28973) );
  XNOR U28987 ( .A(n28977), .B(n28978), .Z(n28975) );
  IV U28988 ( .A(n28942), .Z(n28939) );
  XOR U28989 ( .A(n28979), .B(n28980), .Z(n28942) );
  ANDN U28990 ( .B(n28981), .A(n28982), .Z(n28979) );
  XOR U28991 ( .A(n28980), .B(n28983), .Z(n28981) );
  XOR U28992 ( .A(n28984), .B(n28985), .Z(n28955) );
  XNOR U28993 ( .A(n28950), .B(n28986), .Z(n28985) );
  IV U28994 ( .A(n28953), .Z(n28986) );
  XOR U28995 ( .A(n28987), .B(n28988), .Z(n28953) );
  ANDN U28996 ( .B(n28989), .A(n28990), .Z(n28987) );
  XOR U28997 ( .A(n28988), .B(n28991), .Z(n28989) );
  XNOR U28998 ( .A(n28992), .B(n28993), .Z(n28950) );
  ANDN U28999 ( .B(n28994), .A(n28995), .Z(n28992) );
  XOR U29000 ( .A(n28993), .B(n28996), .Z(n28994) );
  IV U29001 ( .A(n28949), .Z(n28984) );
  XOR U29002 ( .A(n28947), .B(n28997), .Z(n28949) );
  XNOR U29003 ( .A(n28998), .B(n28999), .Z(n28997) );
  ANDN U29004 ( .B(n29000), .A(n29001), .Z(n28998) );
  XNOR U29005 ( .A(n29002), .B(n29003), .Z(n29000) );
  IV U29006 ( .A(n28951), .Z(n28947) );
  XOR U29007 ( .A(n29004), .B(n29005), .Z(n28951) );
  ANDN U29008 ( .B(n29006), .A(n29007), .Z(n29004) );
  XOR U29009 ( .A(n29008), .B(n29005), .Z(n29006) );
  XOR U29010 ( .A(n28962), .B(n28815), .Z(n28963) );
  XOR U29011 ( .A(n29009), .B(n29010), .Z(n28815) );
  AND U29012 ( .A(n352), .B(n29011), .Z(n29009) );
  XOR U29013 ( .A(n29012), .B(n29010), .Z(n29011) );
  XNOR U29014 ( .A(n29013), .B(n29014), .Z(n28962) );
  NAND U29015 ( .A(n29015), .B(n29016), .Z(n29014) );
  XOR U29016 ( .A(n29017), .B(n28914), .Z(n29016) );
  XOR U29017 ( .A(n28990), .B(n28991), .Z(n28914) );
  XOR U29018 ( .A(n29018), .B(n28983), .Z(n28991) );
  XOR U29019 ( .A(n29019), .B(n28971), .Z(n28983) );
  XOR U29020 ( .A(n29020), .B(n29021), .Z(n28971) );
  ANDN U29021 ( .B(n29022), .A(n29023), .Z(n29020) );
  XOR U29022 ( .A(n29021), .B(n29024), .Z(n29022) );
  IV U29023 ( .A(n28969), .Z(n29019) );
  XOR U29024 ( .A(n28967), .B(n29025), .Z(n28969) );
  XOR U29025 ( .A(n29026), .B(n29027), .Z(n29025) );
  ANDN U29026 ( .B(n29028), .A(n29029), .Z(n29026) );
  XOR U29027 ( .A(n29030), .B(n29027), .Z(n29028) );
  IV U29028 ( .A(n28970), .Z(n28967) );
  XOR U29029 ( .A(n29031), .B(n29032), .Z(n28970) );
  ANDN U29030 ( .B(n29033), .A(n29034), .Z(n29031) );
  XOR U29031 ( .A(n29032), .B(n29035), .Z(n29033) );
  IV U29032 ( .A(n28982), .Z(n29018) );
  XOR U29033 ( .A(n29036), .B(n29037), .Z(n28982) );
  XNOR U29034 ( .A(n28977), .B(n29038), .Z(n29037) );
  IV U29035 ( .A(n28980), .Z(n29038) );
  XOR U29036 ( .A(n29039), .B(n29040), .Z(n28980) );
  ANDN U29037 ( .B(n29041), .A(n29042), .Z(n29039) );
  XOR U29038 ( .A(n29040), .B(n29043), .Z(n29041) );
  XNOR U29039 ( .A(n29044), .B(n29045), .Z(n28977) );
  ANDN U29040 ( .B(n29046), .A(n29047), .Z(n29044) );
  XOR U29041 ( .A(n29045), .B(n29048), .Z(n29046) );
  IV U29042 ( .A(n28976), .Z(n29036) );
  XOR U29043 ( .A(n28974), .B(n29049), .Z(n28976) );
  XOR U29044 ( .A(n29050), .B(n29051), .Z(n29049) );
  ANDN U29045 ( .B(n29052), .A(n29053), .Z(n29050) );
  XOR U29046 ( .A(n29054), .B(n29051), .Z(n29052) );
  IV U29047 ( .A(n28978), .Z(n28974) );
  XOR U29048 ( .A(n29055), .B(n29056), .Z(n28978) );
  ANDN U29049 ( .B(n29057), .A(n29058), .Z(n29055) );
  XOR U29050 ( .A(n29059), .B(n29056), .Z(n29057) );
  XOR U29051 ( .A(n29060), .B(n29061), .Z(n28990) );
  XOR U29052 ( .A(n29008), .B(n29062), .Z(n29061) );
  IV U29053 ( .A(n28988), .Z(n29062) );
  XOR U29054 ( .A(n29063), .B(n29064), .Z(n28988) );
  ANDN U29055 ( .B(n29065), .A(n29066), .Z(n29063) );
  XOR U29056 ( .A(n29064), .B(n29067), .Z(n29065) );
  XOR U29057 ( .A(n29068), .B(n28996), .Z(n29008) );
  XOR U29058 ( .A(n29069), .B(n29070), .Z(n28996) );
  ANDN U29059 ( .B(n29071), .A(n29072), .Z(n29069) );
  XOR U29060 ( .A(n29070), .B(n29073), .Z(n29071) );
  IV U29061 ( .A(n28995), .Z(n29068) );
  XOR U29062 ( .A(n29074), .B(n29075), .Z(n28995) );
  XOR U29063 ( .A(n29076), .B(n29077), .Z(n29075) );
  ANDN U29064 ( .B(n29078), .A(n29079), .Z(n29076) );
  XOR U29065 ( .A(n29080), .B(n29077), .Z(n29078) );
  IV U29066 ( .A(n28993), .Z(n29074) );
  XOR U29067 ( .A(n29081), .B(n29082), .Z(n28993) );
  ANDN U29068 ( .B(n29083), .A(n29084), .Z(n29081) );
  XOR U29069 ( .A(n29082), .B(n29085), .Z(n29083) );
  IV U29070 ( .A(n29007), .Z(n29060) );
  XOR U29071 ( .A(n29086), .B(n29087), .Z(n29007) );
  XNOR U29072 ( .A(n29002), .B(n29088), .Z(n29087) );
  IV U29073 ( .A(n29005), .Z(n29088) );
  XOR U29074 ( .A(n29089), .B(n29090), .Z(n29005) );
  ANDN U29075 ( .B(n29091), .A(n29092), .Z(n29089) );
  XOR U29076 ( .A(n29093), .B(n29090), .Z(n29091) );
  XNOR U29077 ( .A(n29094), .B(n29095), .Z(n29002) );
  ANDN U29078 ( .B(n29096), .A(n29097), .Z(n29094) );
  XOR U29079 ( .A(n29095), .B(n29098), .Z(n29096) );
  IV U29080 ( .A(n29001), .Z(n29086) );
  XOR U29081 ( .A(n28999), .B(n29099), .Z(n29001) );
  XOR U29082 ( .A(n29100), .B(n29101), .Z(n29099) );
  ANDN U29083 ( .B(n29102), .A(n29103), .Z(n29100) );
  XOR U29084 ( .A(n29104), .B(n29101), .Z(n29102) );
  IV U29085 ( .A(n29003), .Z(n28999) );
  XOR U29086 ( .A(n29105), .B(n29106), .Z(n29003) );
  ANDN U29087 ( .B(n29107), .A(n29108), .Z(n29105) );
  XOR U29088 ( .A(n29109), .B(n29106), .Z(n29107) );
  IV U29089 ( .A(n29013), .Z(n29017) );
  XOR U29090 ( .A(n29013), .B(n28916), .Z(n29015) );
  XOR U29091 ( .A(n29110), .B(n29111), .Z(n28916) );
  AND U29092 ( .A(n352), .B(n29112), .Z(n29110) );
  XOR U29093 ( .A(n29113), .B(n29111), .Z(n29112) );
  NANDN U29094 ( .A(n28918), .B(n28920), .Z(n29013) );
  XOR U29095 ( .A(n29114), .B(n29115), .Z(n28920) );
  AND U29096 ( .A(n352), .B(n29116), .Z(n29114) );
  XOR U29097 ( .A(n29115), .B(n29117), .Z(n29116) );
  XNOR U29098 ( .A(n29118), .B(n29119), .Z(n352) );
  AND U29099 ( .A(n29120), .B(n29121), .Z(n29118) );
  XOR U29100 ( .A(n29119), .B(n28931), .Z(n29121) );
  XNOR U29101 ( .A(n29122), .B(n29123), .Z(n28931) );
  ANDN U29102 ( .B(n29124), .A(n29125), .Z(n29122) );
  XOR U29103 ( .A(n29123), .B(n29126), .Z(n29124) );
  XNOR U29104 ( .A(n29119), .B(n28933), .Z(n29120) );
  XOR U29105 ( .A(n29127), .B(n29128), .Z(n28933) );
  AND U29106 ( .A(n356), .B(n29129), .Z(n29127) );
  XOR U29107 ( .A(n29130), .B(n29128), .Z(n29129) );
  XOR U29108 ( .A(n29131), .B(n29132), .Z(n29119) );
  AND U29109 ( .A(n29133), .B(n29134), .Z(n29131) );
  XOR U29110 ( .A(n29132), .B(n28958), .Z(n29134) );
  XOR U29111 ( .A(n29125), .B(n29126), .Z(n28958) );
  XNOR U29112 ( .A(n29135), .B(n29136), .Z(n29126) );
  ANDN U29113 ( .B(n29137), .A(n29138), .Z(n29135) );
  XOR U29114 ( .A(n29139), .B(n29140), .Z(n29137) );
  XOR U29115 ( .A(n29141), .B(n29142), .Z(n29125) );
  XNOR U29116 ( .A(n29143), .B(n29144), .Z(n29142) );
  ANDN U29117 ( .B(n29145), .A(n29146), .Z(n29143) );
  XNOR U29118 ( .A(n29147), .B(n29148), .Z(n29145) );
  IV U29119 ( .A(n29123), .Z(n29141) );
  XOR U29120 ( .A(n29149), .B(n29150), .Z(n29123) );
  ANDN U29121 ( .B(n29151), .A(n29152), .Z(n29149) );
  XOR U29122 ( .A(n29150), .B(n29153), .Z(n29151) );
  XNOR U29123 ( .A(n29132), .B(n28960), .Z(n29133) );
  XOR U29124 ( .A(n29154), .B(n29155), .Z(n28960) );
  AND U29125 ( .A(n356), .B(n29156), .Z(n29154) );
  XOR U29126 ( .A(n29157), .B(n29155), .Z(n29156) );
  XNOR U29127 ( .A(n29158), .B(n29159), .Z(n29132) );
  AND U29128 ( .A(n29160), .B(n29161), .Z(n29158) );
  XNOR U29129 ( .A(n29159), .B(n29010), .Z(n29161) );
  XOR U29130 ( .A(n29152), .B(n29153), .Z(n29010) );
  XOR U29131 ( .A(n29162), .B(n29140), .Z(n29153) );
  XNOR U29132 ( .A(n29163), .B(n29164), .Z(n29140) );
  ANDN U29133 ( .B(n29165), .A(n29166), .Z(n29163) );
  XOR U29134 ( .A(n29167), .B(n29168), .Z(n29165) );
  IV U29135 ( .A(n29138), .Z(n29162) );
  XOR U29136 ( .A(n29136), .B(n29169), .Z(n29138) );
  XNOR U29137 ( .A(n29170), .B(n29171), .Z(n29169) );
  ANDN U29138 ( .B(n29172), .A(n29173), .Z(n29170) );
  XNOR U29139 ( .A(n29174), .B(n29175), .Z(n29172) );
  IV U29140 ( .A(n29139), .Z(n29136) );
  XOR U29141 ( .A(n29176), .B(n29177), .Z(n29139) );
  ANDN U29142 ( .B(n29178), .A(n29179), .Z(n29176) );
  XOR U29143 ( .A(n29177), .B(n29180), .Z(n29178) );
  XOR U29144 ( .A(n29181), .B(n29182), .Z(n29152) );
  XNOR U29145 ( .A(n29147), .B(n29183), .Z(n29182) );
  IV U29146 ( .A(n29150), .Z(n29183) );
  XOR U29147 ( .A(n29184), .B(n29185), .Z(n29150) );
  ANDN U29148 ( .B(n29186), .A(n29187), .Z(n29184) );
  XOR U29149 ( .A(n29185), .B(n29188), .Z(n29186) );
  XNOR U29150 ( .A(n29189), .B(n29190), .Z(n29147) );
  ANDN U29151 ( .B(n29191), .A(n29192), .Z(n29189) );
  XOR U29152 ( .A(n29190), .B(n29193), .Z(n29191) );
  IV U29153 ( .A(n29146), .Z(n29181) );
  XOR U29154 ( .A(n29144), .B(n29194), .Z(n29146) );
  XNOR U29155 ( .A(n29195), .B(n29196), .Z(n29194) );
  ANDN U29156 ( .B(n29197), .A(n29198), .Z(n29195) );
  XNOR U29157 ( .A(n29199), .B(n29200), .Z(n29197) );
  IV U29158 ( .A(n29148), .Z(n29144) );
  XOR U29159 ( .A(n29201), .B(n29202), .Z(n29148) );
  ANDN U29160 ( .B(n29203), .A(n29204), .Z(n29201) );
  XOR U29161 ( .A(n29205), .B(n29202), .Z(n29203) );
  XOR U29162 ( .A(n29159), .B(n29012), .Z(n29160) );
  XOR U29163 ( .A(n29206), .B(n29207), .Z(n29012) );
  AND U29164 ( .A(n356), .B(n29208), .Z(n29206) );
  XOR U29165 ( .A(n29209), .B(n29207), .Z(n29208) );
  XNOR U29166 ( .A(n29210), .B(n29211), .Z(n29159) );
  NAND U29167 ( .A(n29212), .B(n29213), .Z(n29211) );
  XOR U29168 ( .A(n29214), .B(n29111), .Z(n29213) );
  XOR U29169 ( .A(n29187), .B(n29188), .Z(n29111) );
  XOR U29170 ( .A(n29215), .B(n29180), .Z(n29188) );
  XOR U29171 ( .A(n29216), .B(n29168), .Z(n29180) );
  XOR U29172 ( .A(n29217), .B(n29218), .Z(n29168) );
  ANDN U29173 ( .B(n29219), .A(n29220), .Z(n29217) );
  XOR U29174 ( .A(n29218), .B(n29221), .Z(n29219) );
  IV U29175 ( .A(n29166), .Z(n29216) );
  XOR U29176 ( .A(n29164), .B(n29222), .Z(n29166) );
  XOR U29177 ( .A(n29223), .B(n29224), .Z(n29222) );
  ANDN U29178 ( .B(n29225), .A(n29226), .Z(n29223) );
  XOR U29179 ( .A(n29227), .B(n29224), .Z(n29225) );
  IV U29180 ( .A(n29167), .Z(n29164) );
  XOR U29181 ( .A(n29228), .B(n29229), .Z(n29167) );
  ANDN U29182 ( .B(n29230), .A(n29231), .Z(n29228) );
  XOR U29183 ( .A(n29229), .B(n29232), .Z(n29230) );
  IV U29184 ( .A(n29179), .Z(n29215) );
  XOR U29185 ( .A(n29233), .B(n29234), .Z(n29179) );
  XNOR U29186 ( .A(n29174), .B(n29235), .Z(n29234) );
  IV U29187 ( .A(n29177), .Z(n29235) );
  XOR U29188 ( .A(n29236), .B(n29237), .Z(n29177) );
  ANDN U29189 ( .B(n29238), .A(n29239), .Z(n29236) );
  XOR U29190 ( .A(n29237), .B(n29240), .Z(n29238) );
  XNOR U29191 ( .A(n29241), .B(n29242), .Z(n29174) );
  ANDN U29192 ( .B(n29243), .A(n29244), .Z(n29241) );
  XOR U29193 ( .A(n29242), .B(n29245), .Z(n29243) );
  IV U29194 ( .A(n29173), .Z(n29233) );
  XOR U29195 ( .A(n29171), .B(n29246), .Z(n29173) );
  XOR U29196 ( .A(n29247), .B(n29248), .Z(n29246) );
  ANDN U29197 ( .B(n29249), .A(n29250), .Z(n29247) );
  XOR U29198 ( .A(n29251), .B(n29248), .Z(n29249) );
  IV U29199 ( .A(n29175), .Z(n29171) );
  XOR U29200 ( .A(n29252), .B(n29253), .Z(n29175) );
  ANDN U29201 ( .B(n29254), .A(n29255), .Z(n29252) );
  XOR U29202 ( .A(n29256), .B(n29253), .Z(n29254) );
  XOR U29203 ( .A(n29257), .B(n29258), .Z(n29187) );
  XOR U29204 ( .A(n29205), .B(n29259), .Z(n29258) );
  IV U29205 ( .A(n29185), .Z(n29259) );
  XOR U29206 ( .A(n29260), .B(n29261), .Z(n29185) );
  ANDN U29207 ( .B(n29262), .A(n29263), .Z(n29260) );
  XOR U29208 ( .A(n29261), .B(n29264), .Z(n29262) );
  XOR U29209 ( .A(n29265), .B(n29193), .Z(n29205) );
  XOR U29210 ( .A(n29266), .B(n29267), .Z(n29193) );
  ANDN U29211 ( .B(n29268), .A(n29269), .Z(n29266) );
  XOR U29212 ( .A(n29267), .B(n29270), .Z(n29268) );
  IV U29213 ( .A(n29192), .Z(n29265) );
  XOR U29214 ( .A(n29271), .B(n29272), .Z(n29192) );
  XOR U29215 ( .A(n29273), .B(n29274), .Z(n29272) );
  ANDN U29216 ( .B(n29275), .A(n29276), .Z(n29273) );
  XOR U29217 ( .A(n29277), .B(n29274), .Z(n29275) );
  IV U29218 ( .A(n29190), .Z(n29271) );
  XOR U29219 ( .A(n29278), .B(n29279), .Z(n29190) );
  ANDN U29220 ( .B(n29280), .A(n29281), .Z(n29278) );
  XOR U29221 ( .A(n29279), .B(n29282), .Z(n29280) );
  IV U29222 ( .A(n29204), .Z(n29257) );
  XOR U29223 ( .A(n29283), .B(n29284), .Z(n29204) );
  XNOR U29224 ( .A(n29199), .B(n29285), .Z(n29284) );
  IV U29225 ( .A(n29202), .Z(n29285) );
  XOR U29226 ( .A(n29286), .B(n29287), .Z(n29202) );
  ANDN U29227 ( .B(n29288), .A(n29289), .Z(n29286) );
  XOR U29228 ( .A(n29290), .B(n29287), .Z(n29288) );
  XNOR U29229 ( .A(n29291), .B(n29292), .Z(n29199) );
  ANDN U29230 ( .B(n29293), .A(n29294), .Z(n29291) );
  XOR U29231 ( .A(n29292), .B(n29295), .Z(n29293) );
  IV U29232 ( .A(n29198), .Z(n29283) );
  XOR U29233 ( .A(n29196), .B(n29296), .Z(n29198) );
  XOR U29234 ( .A(n29297), .B(n29298), .Z(n29296) );
  ANDN U29235 ( .B(n29299), .A(n29300), .Z(n29297) );
  XOR U29236 ( .A(n29301), .B(n29298), .Z(n29299) );
  IV U29237 ( .A(n29200), .Z(n29196) );
  XOR U29238 ( .A(n29302), .B(n29303), .Z(n29200) );
  ANDN U29239 ( .B(n29304), .A(n29305), .Z(n29302) );
  XOR U29240 ( .A(n29306), .B(n29303), .Z(n29304) );
  IV U29241 ( .A(n29210), .Z(n29214) );
  XOR U29242 ( .A(n29210), .B(n29113), .Z(n29212) );
  XOR U29243 ( .A(n29307), .B(n29308), .Z(n29113) );
  AND U29244 ( .A(n356), .B(n29309), .Z(n29307) );
  XOR U29245 ( .A(n29310), .B(n29308), .Z(n29309) );
  NANDN U29246 ( .A(n29115), .B(n29117), .Z(n29210) );
  XOR U29247 ( .A(n29311), .B(n29312), .Z(n29117) );
  AND U29248 ( .A(n356), .B(n29313), .Z(n29311) );
  XOR U29249 ( .A(n29312), .B(n29314), .Z(n29313) );
  XNOR U29250 ( .A(n29315), .B(n29316), .Z(n356) );
  AND U29251 ( .A(n29317), .B(n29318), .Z(n29315) );
  XOR U29252 ( .A(n29316), .B(n29128), .Z(n29318) );
  XNOR U29253 ( .A(n29319), .B(n29320), .Z(n29128) );
  ANDN U29254 ( .B(n29321), .A(n29322), .Z(n29319) );
  XOR U29255 ( .A(n29320), .B(n29323), .Z(n29321) );
  XNOR U29256 ( .A(n29316), .B(n29130), .Z(n29317) );
  XOR U29257 ( .A(n29324), .B(n29325), .Z(n29130) );
  AND U29258 ( .A(n360), .B(n29326), .Z(n29324) );
  XOR U29259 ( .A(n29327), .B(n29325), .Z(n29326) );
  XOR U29260 ( .A(n29328), .B(n29329), .Z(n29316) );
  AND U29261 ( .A(n29330), .B(n29331), .Z(n29328) );
  XOR U29262 ( .A(n29329), .B(n29155), .Z(n29331) );
  XOR U29263 ( .A(n29322), .B(n29323), .Z(n29155) );
  XNOR U29264 ( .A(n29332), .B(n29333), .Z(n29323) );
  ANDN U29265 ( .B(n29334), .A(n29335), .Z(n29332) );
  XOR U29266 ( .A(n29336), .B(n29337), .Z(n29334) );
  XOR U29267 ( .A(n29338), .B(n29339), .Z(n29322) );
  XNOR U29268 ( .A(n29340), .B(n29341), .Z(n29339) );
  ANDN U29269 ( .B(n29342), .A(n29343), .Z(n29340) );
  XNOR U29270 ( .A(n29344), .B(n29345), .Z(n29342) );
  IV U29271 ( .A(n29320), .Z(n29338) );
  XOR U29272 ( .A(n29346), .B(n29347), .Z(n29320) );
  ANDN U29273 ( .B(n29348), .A(n29349), .Z(n29346) );
  XOR U29274 ( .A(n29347), .B(n29350), .Z(n29348) );
  XNOR U29275 ( .A(n29329), .B(n29157), .Z(n29330) );
  XOR U29276 ( .A(n29351), .B(n29352), .Z(n29157) );
  AND U29277 ( .A(n360), .B(n29353), .Z(n29351) );
  XOR U29278 ( .A(n29354), .B(n29352), .Z(n29353) );
  XNOR U29279 ( .A(n29355), .B(n29356), .Z(n29329) );
  AND U29280 ( .A(n29357), .B(n29358), .Z(n29355) );
  XNOR U29281 ( .A(n29356), .B(n29207), .Z(n29358) );
  XOR U29282 ( .A(n29349), .B(n29350), .Z(n29207) );
  XOR U29283 ( .A(n29359), .B(n29337), .Z(n29350) );
  XNOR U29284 ( .A(n29360), .B(n29361), .Z(n29337) );
  ANDN U29285 ( .B(n29362), .A(n29363), .Z(n29360) );
  XOR U29286 ( .A(n29364), .B(n29365), .Z(n29362) );
  IV U29287 ( .A(n29335), .Z(n29359) );
  XOR U29288 ( .A(n29333), .B(n29366), .Z(n29335) );
  XNOR U29289 ( .A(n29367), .B(n29368), .Z(n29366) );
  ANDN U29290 ( .B(n29369), .A(n29370), .Z(n29367) );
  XNOR U29291 ( .A(n29371), .B(n29372), .Z(n29369) );
  IV U29292 ( .A(n29336), .Z(n29333) );
  XOR U29293 ( .A(n29373), .B(n29374), .Z(n29336) );
  ANDN U29294 ( .B(n29375), .A(n29376), .Z(n29373) );
  XOR U29295 ( .A(n29374), .B(n29377), .Z(n29375) );
  XOR U29296 ( .A(n29378), .B(n29379), .Z(n29349) );
  XNOR U29297 ( .A(n29344), .B(n29380), .Z(n29379) );
  IV U29298 ( .A(n29347), .Z(n29380) );
  XOR U29299 ( .A(n29381), .B(n29382), .Z(n29347) );
  ANDN U29300 ( .B(n29383), .A(n29384), .Z(n29381) );
  XOR U29301 ( .A(n29382), .B(n29385), .Z(n29383) );
  XNOR U29302 ( .A(n29386), .B(n29387), .Z(n29344) );
  ANDN U29303 ( .B(n29388), .A(n29389), .Z(n29386) );
  XOR U29304 ( .A(n29387), .B(n29390), .Z(n29388) );
  IV U29305 ( .A(n29343), .Z(n29378) );
  XOR U29306 ( .A(n29341), .B(n29391), .Z(n29343) );
  XNOR U29307 ( .A(n29392), .B(n29393), .Z(n29391) );
  ANDN U29308 ( .B(n29394), .A(n29395), .Z(n29392) );
  XNOR U29309 ( .A(n29396), .B(n29397), .Z(n29394) );
  IV U29310 ( .A(n29345), .Z(n29341) );
  XOR U29311 ( .A(n29398), .B(n29399), .Z(n29345) );
  ANDN U29312 ( .B(n29400), .A(n29401), .Z(n29398) );
  XOR U29313 ( .A(n29402), .B(n29399), .Z(n29400) );
  XOR U29314 ( .A(n29356), .B(n29209), .Z(n29357) );
  XOR U29315 ( .A(n29403), .B(n29404), .Z(n29209) );
  AND U29316 ( .A(n360), .B(n29405), .Z(n29403) );
  XOR U29317 ( .A(n29406), .B(n29404), .Z(n29405) );
  XNOR U29318 ( .A(n29407), .B(n29408), .Z(n29356) );
  NAND U29319 ( .A(n29409), .B(n29410), .Z(n29408) );
  XOR U29320 ( .A(n29411), .B(n29308), .Z(n29410) );
  XOR U29321 ( .A(n29384), .B(n29385), .Z(n29308) );
  XOR U29322 ( .A(n29412), .B(n29377), .Z(n29385) );
  XOR U29323 ( .A(n29413), .B(n29365), .Z(n29377) );
  XOR U29324 ( .A(n29414), .B(n29415), .Z(n29365) );
  ANDN U29325 ( .B(n29416), .A(n29417), .Z(n29414) );
  XOR U29326 ( .A(n29415), .B(n29418), .Z(n29416) );
  IV U29327 ( .A(n29363), .Z(n29413) );
  XOR U29328 ( .A(n29361), .B(n29419), .Z(n29363) );
  XOR U29329 ( .A(n29420), .B(n29421), .Z(n29419) );
  ANDN U29330 ( .B(n29422), .A(n29423), .Z(n29420) );
  XOR U29331 ( .A(n29424), .B(n29421), .Z(n29422) );
  IV U29332 ( .A(n29364), .Z(n29361) );
  XOR U29333 ( .A(n29425), .B(n29426), .Z(n29364) );
  ANDN U29334 ( .B(n29427), .A(n29428), .Z(n29425) );
  XOR U29335 ( .A(n29426), .B(n29429), .Z(n29427) );
  IV U29336 ( .A(n29376), .Z(n29412) );
  XOR U29337 ( .A(n29430), .B(n29431), .Z(n29376) );
  XNOR U29338 ( .A(n29371), .B(n29432), .Z(n29431) );
  IV U29339 ( .A(n29374), .Z(n29432) );
  XOR U29340 ( .A(n29433), .B(n29434), .Z(n29374) );
  ANDN U29341 ( .B(n29435), .A(n29436), .Z(n29433) );
  XOR U29342 ( .A(n29434), .B(n29437), .Z(n29435) );
  XNOR U29343 ( .A(n29438), .B(n29439), .Z(n29371) );
  ANDN U29344 ( .B(n29440), .A(n29441), .Z(n29438) );
  XOR U29345 ( .A(n29439), .B(n29442), .Z(n29440) );
  IV U29346 ( .A(n29370), .Z(n29430) );
  XOR U29347 ( .A(n29368), .B(n29443), .Z(n29370) );
  XOR U29348 ( .A(n29444), .B(n29445), .Z(n29443) );
  ANDN U29349 ( .B(n29446), .A(n29447), .Z(n29444) );
  XOR U29350 ( .A(n29448), .B(n29445), .Z(n29446) );
  IV U29351 ( .A(n29372), .Z(n29368) );
  XOR U29352 ( .A(n29449), .B(n29450), .Z(n29372) );
  ANDN U29353 ( .B(n29451), .A(n29452), .Z(n29449) );
  XOR U29354 ( .A(n29453), .B(n29450), .Z(n29451) );
  XOR U29355 ( .A(n29454), .B(n29455), .Z(n29384) );
  XOR U29356 ( .A(n29402), .B(n29456), .Z(n29455) );
  IV U29357 ( .A(n29382), .Z(n29456) );
  XOR U29358 ( .A(n29457), .B(n29458), .Z(n29382) );
  ANDN U29359 ( .B(n29459), .A(n29460), .Z(n29457) );
  XOR U29360 ( .A(n29458), .B(n29461), .Z(n29459) );
  XOR U29361 ( .A(n29462), .B(n29390), .Z(n29402) );
  XOR U29362 ( .A(n29463), .B(n29464), .Z(n29390) );
  ANDN U29363 ( .B(n29465), .A(n29466), .Z(n29463) );
  XOR U29364 ( .A(n29464), .B(n29467), .Z(n29465) );
  IV U29365 ( .A(n29389), .Z(n29462) );
  XOR U29366 ( .A(n29468), .B(n29469), .Z(n29389) );
  XOR U29367 ( .A(n29470), .B(n29471), .Z(n29469) );
  ANDN U29368 ( .B(n29472), .A(n29473), .Z(n29470) );
  XOR U29369 ( .A(n29474), .B(n29471), .Z(n29472) );
  IV U29370 ( .A(n29387), .Z(n29468) );
  XOR U29371 ( .A(n29475), .B(n29476), .Z(n29387) );
  ANDN U29372 ( .B(n29477), .A(n29478), .Z(n29475) );
  XOR U29373 ( .A(n29476), .B(n29479), .Z(n29477) );
  IV U29374 ( .A(n29401), .Z(n29454) );
  XOR U29375 ( .A(n29480), .B(n29481), .Z(n29401) );
  XNOR U29376 ( .A(n29396), .B(n29482), .Z(n29481) );
  IV U29377 ( .A(n29399), .Z(n29482) );
  XOR U29378 ( .A(n29483), .B(n29484), .Z(n29399) );
  ANDN U29379 ( .B(n29485), .A(n29486), .Z(n29483) );
  XOR U29380 ( .A(n29487), .B(n29484), .Z(n29485) );
  XNOR U29381 ( .A(n29488), .B(n29489), .Z(n29396) );
  ANDN U29382 ( .B(n29490), .A(n29491), .Z(n29488) );
  XOR U29383 ( .A(n29489), .B(n29492), .Z(n29490) );
  IV U29384 ( .A(n29395), .Z(n29480) );
  XOR U29385 ( .A(n29393), .B(n29493), .Z(n29395) );
  XOR U29386 ( .A(n29494), .B(n29495), .Z(n29493) );
  ANDN U29387 ( .B(n29496), .A(n29497), .Z(n29494) );
  XOR U29388 ( .A(n29498), .B(n29495), .Z(n29496) );
  IV U29389 ( .A(n29397), .Z(n29393) );
  XOR U29390 ( .A(n29499), .B(n29500), .Z(n29397) );
  ANDN U29391 ( .B(n29501), .A(n29502), .Z(n29499) );
  XOR U29392 ( .A(n29503), .B(n29500), .Z(n29501) );
  IV U29393 ( .A(n29407), .Z(n29411) );
  XOR U29394 ( .A(n29407), .B(n29310), .Z(n29409) );
  XOR U29395 ( .A(n29504), .B(n29505), .Z(n29310) );
  AND U29396 ( .A(n360), .B(n29506), .Z(n29504) );
  XOR U29397 ( .A(n29507), .B(n29505), .Z(n29506) );
  NANDN U29398 ( .A(n29312), .B(n29314), .Z(n29407) );
  XOR U29399 ( .A(n29508), .B(n29509), .Z(n29314) );
  AND U29400 ( .A(n360), .B(n29510), .Z(n29508) );
  XOR U29401 ( .A(n29509), .B(n29511), .Z(n29510) );
  XNOR U29402 ( .A(n29512), .B(n29513), .Z(n360) );
  AND U29403 ( .A(n29514), .B(n29515), .Z(n29512) );
  XOR U29404 ( .A(n29513), .B(n29325), .Z(n29515) );
  XNOR U29405 ( .A(n29516), .B(n29517), .Z(n29325) );
  ANDN U29406 ( .B(n29518), .A(n29519), .Z(n29516) );
  XOR U29407 ( .A(n29517), .B(n29520), .Z(n29518) );
  XNOR U29408 ( .A(n29513), .B(n29327), .Z(n29514) );
  XOR U29409 ( .A(n29521), .B(n29522), .Z(n29327) );
  AND U29410 ( .A(n364), .B(n29523), .Z(n29521) );
  XOR U29411 ( .A(n29524), .B(n29522), .Z(n29523) );
  XOR U29412 ( .A(n29525), .B(n29526), .Z(n29513) );
  AND U29413 ( .A(n29527), .B(n29528), .Z(n29525) );
  XOR U29414 ( .A(n29526), .B(n29352), .Z(n29528) );
  XOR U29415 ( .A(n29519), .B(n29520), .Z(n29352) );
  XNOR U29416 ( .A(n29529), .B(n29530), .Z(n29520) );
  ANDN U29417 ( .B(n29531), .A(n29532), .Z(n29529) );
  XOR U29418 ( .A(n29533), .B(n29534), .Z(n29531) );
  XOR U29419 ( .A(n29535), .B(n29536), .Z(n29519) );
  XNOR U29420 ( .A(n29537), .B(n29538), .Z(n29536) );
  ANDN U29421 ( .B(n29539), .A(n29540), .Z(n29537) );
  XNOR U29422 ( .A(n29541), .B(n29542), .Z(n29539) );
  IV U29423 ( .A(n29517), .Z(n29535) );
  XOR U29424 ( .A(n29543), .B(n29544), .Z(n29517) );
  ANDN U29425 ( .B(n29545), .A(n29546), .Z(n29543) );
  XOR U29426 ( .A(n29544), .B(n29547), .Z(n29545) );
  XNOR U29427 ( .A(n29526), .B(n29354), .Z(n29527) );
  XOR U29428 ( .A(n29548), .B(n29549), .Z(n29354) );
  AND U29429 ( .A(n364), .B(n29550), .Z(n29548) );
  XOR U29430 ( .A(n29551), .B(n29549), .Z(n29550) );
  XNOR U29431 ( .A(n29552), .B(n29553), .Z(n29526) );
  AND U29432 ( .A(n29554), .B(n29555), .Z(n29552) );
  XNOR U29433 ( .A(n29553), .B(n29404), .Z(n29555) );
  XOR U29434 ( .A(n29546), .B(n29547), .Z(n29404) );
  XOR U29435 ( .A(n29556), .B(n29534), .Z(n29547) );
  XNOR U29436 ( .A(n29557), .B(n29558), .Z(n29534) );
  ANDN U29437 ( .B(n29559), .A(n29560), .Z(n29557) );
  XOR U29438 ( .A(n29561), .B(n29562), .Z(n29559) );
  IV U29439 ( .A(n29532), .Z(n29556) );
  XOR U29440 ( .A(n29530), .B(n29563), .Z(n29532) );
  XNOR U29441 ( .A(n29564), .B(n29565), .Z(n29563) );
  ANDN U29442 ( .B(n29566), .A(n29567), .Z(n29564) );
  XNOR U29443 ( .A(n29568), .B(n29569), .Z(n29566) );
  IV U29444 ( .A(n29533), .Z(n29530) );
  XOR U29445 ( .A(n29570), .B(n29571), .Z(n29533) );
  ANDN U29446 ( .B(n29572), .A(n29573), .Z(n29570) );
  XOR U29447 ( .A(n29571), .B(n29574), .Z(n29572) );
  XOR U29448 ( .A(n29575), .B(n29576), .Z(n29546) );
  XNOR U29449 ( .A(n29541), .B(n29577), .Z(n29576) );
  IV U29450 ( .A(n29544), .Z(n29577) );
  XOR U29451 ( .A(n29578), .B(n29579), .Z(n29544) );
  ANDN U29452 ( .B(n29580), .A(n29581), .Z(n29578) );
  XOR U29453 ( .A(n29579), .B(n29582), .Z(n29580) );
  XNOR U29454 ( .A(n29583), .B(n29584), .Z(n29541) );
  ANDN U29455 ( .B(n29585), .A(n29586), .Z(n29583) );
  XOR U29456 ( .A(n29584), .B(n29587), .Z(n29585) );
  IV U29457 ( .A(n29540), .Z(n29575) );
  XOR U29458 ( .A(n29538), .B(n29588), .Z(n29540) );
  XNOR U29459 ( .A(n29589), .B(n29590), .Z(n29588) );
  ANDN U29460 ( .B(n29591), .A(n29592), .Z(n29589) );
  XNOR U29461 ( .A(n29593), .B(n29594), .Z(n29591) );
  IV U29462 ( .A(n29542), .Z(n29538) );
  XOR U29463 ( .A(n29595), .B(n29596), .Z(n29542) );
  ANDN U29464 ( .B(n29597), .A(n29598), .Z(n29595) );
  XOR U29465 ( .A(n29599), .B(n29596), .Z(n29597) );
  XOR U29466 ( .A(n29553), .B(n29406), .Z(n29554) );
  XOR U29467 ( .A(n29600), .B(n29601), .Z(n29406) );
  AND U29468 ( .A(n364), .B(n29602), .Z(n29600) );
  XOR U29469 ( .A(n29603), .B(n29601), .Z(n29602) );
  XNOR U29470 ( .A(n29604), .B(n29605), .Z(n29553) );
  NAND U29471 ( .A(n29606), .B(n29607), .Z(n29605) );
  XOR U29472 ( .A(n29608), .B(n29505), .Z(n29607) );
  XOR U29473 ( .A(n29581), .B(n29582), .Z(n29505) );
  XOR U29474 ( .A(n29609), .B(n29574), .Z(n29582) );
  XOR U29475 ( .A(n29610), .B(n29562), .Z(n29574) );
  XOR U29476 ( .A(n29611), .B(n29612), .Z(n29562) );
  ANDN U29477 ( .B(n29613), .A(n29614), .Z(n29611) );
  XOR U29478 ( .A(n29612), .B(n29615), .Z(n29613) );
  IV U29479 ( .A(n29560), .Z(n29610) );
  XOR U29480 ( .A(n29558), .B(n29616), .Z(n29560) );
  XOR U29481 ( .A(n29617), .B(n29618), .Z(n29616) );
  ANDN U29482 ( .B(n29619), .A(n29620), .Z(n29617) );
  XOR U29483 ( .A(n29621), .B(n29618), .Z(n29619) );
  IV U29484 ( .A(n29561), .Z(n29558) );
  XOR U29485 ( .A(n29622), .B(n29623), .Z(n29561) );
  ANDN U29486 ( .B(n29624), .A(n29625), .Z(n29622) );
  XOR U29487 ( .A(n29623), .B(n29626), .Z(n29624) );
  IV U29488 ( .A(n29573), .Z(n29609) );
  XOR U29489 ( .A(n29627), .B(n29628), .Z(n29573) );
  XNOR U29490 ( .A(n29568), .B(n29629), .Z(n29628) );
  IV U29491 ( .A(n29571), .Z(n29629) );
  XOR U29492 ( .A(n29630), .B(n29631), .Z(n29571) );
  ANDN U29493 ( .B(n29632), .A(n29633), .Z(n29630) );
  XOR U29494 ( .A(n29631), .B(n29634), .Z(n29632) );
  XNOR U29495 ( .A(n29635), .B(n29636), .Z(n29568) );
  ANDN U29496 ( .B(n29637), .A(n29638), .Z(n29635) );
  XOR U29497 ( .A(n29636), .B(n29639), .Z(n29637) );
  IV U29498 ( .A(n29567), .Z(n29627) );
  XOR U29499 ( .A(n29565), .B(n29640), .Z(n29567) );
  XOR U29500 ( .A(n29641), .B(n29642), .Z(n29640) );
  ANDN U29501 ( .B(n29643), .A(n29644), .Z(n29641) );
  XOR U29502 ( .A(n29645), .B(n29642), .Z(n29643) );
  IV U29503 ( .A(n29569), .Z(n29565) );
  XOR U29504 ( .A(n29646), .B(n29647), .Z(n29569) );
  ANDN U29505 ( .B(n29648), .A(n29649), .Z(n29646) );
  XOR U29506 ( .A(n29650), .B(n29647), .Z(n29648) );
  XOR U29507 ( .A(n29651), .B(n29652), .Z(n29581) );
  XOR U29508 ( .A(n29599), .B(n29653), .Z(n29652) );
  IV U29509 ( .A(n29579), .Z(n29653) );
  XOR U29510 ( .A(n29654), .B(n29655), .Z(n29579) );
  ANDN U29511 ( .B(n29656), .A(n29657), .Z(n29654) );
  XOR U29512 ( .A(n29655), .B(n29658), .Z(n29656) );
  XOR U29513 ( .A(n29659), .B(n29587), .Z(n29599) );
  XOR U29514 ( .A(n29660), .B(n29661), .Z(n29587) );
  ANDN U29515 ( .B(n29662), .A(n29663), .Z(n29660) );
  XOR U29516 ( .A(n29661), .B(n29664), .Z(n29662) );
  IV U29517 ( .A(n29586), .Z(n29659) );
  XOR U29518 ( .A(n29665), .B(n29666), .Z(n29586) );
  XOR U29519 ( .A(n29667), .B(n29668), .Z(n29666) );
  ANDN U29520 ( .B(n29669), .A(n29670), .Z(n29667) );
  XOR U29521 ( .A(n29671), .B(n29668), .Z(n29669) );
  IV U29522 ( .A(n29584), .Z(n29665) );
  XOR U29523 ( .A(n29672), .B(n29673), .Z(n29584) );
  ANDN U29524 ( .B(n29674), .A(n29675), .Z(n29672) );
  XOR U29525 ( .A(n29673), .B(n29676), .Z(n29674) );
  IV U29526 ( .A(n29598), .Z(n29651) );
  XOR U29527 ( .A(n29677), .B(n29678), .Z(n29598) );
  XNOR U29528 ( .A(n29593), .B(n29679), .Z(n29678) );
  IV U29529 ( .A(n29596), .Z(n29679) );
  XOR U29530 ( .A(n29680), .B(n29681), .Z(n29596) );
  ANDN U29531 ( .B(n29682), .A(n29683), .Z(n29680) );
  XOR U29532 ( .A(n29684), .B(n29681), .Z(n29682) );
  XNOR U29533 ( .A(n29685), .B(n29686), .Z(n29593) );
  ANDN U29534 ( .B(n29687), .A(n29688), .Z(n29685) );
  XOR U29535 ( .A(n29686), .B(n29689), .Z(n29687) );
  IV U29536 ( .A(n29592), .Z(n29677) );
  XOR U29537 ( .A(n29590), .B(n29690), .Z(n29592) );
  XOR U29538 ( .A(n29691), .B(n29692), .Z(n29690) );
  ANDN U29539 ( .B(n29693), .A(n29694), .Z(n29691) );
  XOR U29540 ( .A(n29695), .B(n29692), .Z(n29693) );
  IV U29541 ( .A(n29594), .Z(n29590) );
  XOR U29542 ( .A(n29696), .B(n29697), .Z(n29594) );
  ANDN U29543 ( .B(n29698), .A(n29699), .Z(n29696) );
  XOR U29544 ( .A(n29700), .B(n29697), .Z(n29698) );
  IV U29545 ( .A(n29604), .Z(n29608) );
  XOR U29546 ( .A(n29604), .B(n29507), .Z(n29606) );
  XOR U29547 ( .A(n29701), .B(n29702), .Z(n29507) );
  AND U29548 ( .A(n364), .B(n29703), .Z(n29701) );
  XOR U29549 ( .A(n29704), .B(n29702), .Z(n29703) );
  NANDN U29550 ( .A(n29509), .B(n29511), .Z(n29604) );
  XOR U29551 ( .A(n29705), .B(n29706), .Z(n29511) );
  AND U29552 ( .A(n364), .B(n29707), .Z(n29705) );
  XOR U29553 ( .A(n29706), .B(n29708), .Z(n29707) );
  XNOR U29554 ( .A(n29709), .B(n29710), .Z(n364) );
  AND U29555 ( .A(n29711), .B(n29712), .Z(n29709) );
  XOR U29556 ( .A(n29710), .B(n29522), .Z(n29712) );
  XNOR U29557 ( .A(n29713), .B(n29714), .Z(n29522) );
  ANDN U29558 ( .B(n29715), .A(n29716), .Z(n29713) );
  XOR U29559 ( .A(n29714), .B(n29717), .Z(n29715) );
  XNOR U29560 ( .A(n29710), .B(n29524), .Z(n29711) );
  XOR U29561 ( .A(n29718), .B(n29719), .Z(n29524) );
  AND U29562 ( .A(n368), .B(n29720), .Z(n29718) );
  XOR U29563 ( .A(n29721), .B(n29719), .Z(n29720) );
  XOR U29564 ( .A(n29722), .B(n29723), .Z(n29710) );
  AND U29565 ( .A(n29724), .B(n29725), .Z(n29722) );
  XOR U29566 ( .A(n29723), .B(n29549), .Z(n29725) );
  XOR U29567 ( .A(n29716), .B(n29717), .Z(n29549) );
  XNOR U29568 ( .A(n29726), .B(n29727), .Z(n29717) );
  ANDN U29569 ( .B(n29728), .A(n29729), .Z(n29726) );
  XOR U29570 ( .A(n29730), .B(n29731), .Z(n29728) );
  XOR U29571 ( .A(n29732), .B(n29733), .Z(n29716) );
  XNOR U29572 ( .A(n29734), .B(n29735), .Z(n29733) );
  ANDN U29573 ( .B(n29736), .A(n29737), .Z(n29734) );
  XNOR U29574 ( .A(n29738), .B(n29739), .Z(n29736) );
  IV U29575 ( .A(n29714), .Z(n29732) );
  XOR U29576 ( .A(n29740), .B(n29741), .Z(n29714) );
  ANDN U29577 ( .B(n29742), .A(n29743), .Z(n29740) );
  XOR U29578 ( .A(n29741), .B(n29744), .Z(n29742) );
  XNOR U29579 ( .A(n29723), .B(n29551), .Z(n29724) );
  XOR U29580 ( .A(n29745), .B(n29746), .Z(n29551) );
  AND U29581 ( .A(n368), .B(n29747), .Z(n29745) );
  XOR U29582 ( .A(n29748), .B(n29746), .Z(n29747) );
  XNOR U29583 ( .A(n29749), .B(n29750), .Z(n29723) );
  AND U29584 ( .A(n29751), .B(n29752), .Z(n29749) );
  XNOR U29585 ( .A(n29750), .B(n29601), .Z(n29752) );
  XOR U29586 ( .A(n29743), .B(n29744), .Z(n29601) );
  XOR U29587 ( .A(n29753), .B(n29731), .Z(n29744) );
  XNOR U29588 ( .A(n29754), .B(n29755), .Z(n29731) );
  ANDN U29589 ( .B(n29756), .A(n29757), .Z(n29754) );
  XOR U29590 ( .A(n29758), .B(n29759), .Z(n29756) );
  IV U29591 ( .A(n29729), .Z(n29753) );
  XOR U29592 ( .A(n29727), .B(n29760), .Z(n29729) );
  XNOR U29593 ( .A(n29761), .B(n29762), .Z(n29760) );
  ANDN U29594 ( .B(n29763), .A(n29764), .Z(n29761) );
  XNOR U29595 ( .A(n29765), .B(n29766), .Z(n29763) );
  IV U29596 ( .A(n29730), .Z(n29727) );
  XOR U29597 ( .A(n29767), .B(n29768), .Z(n29730) );
  ANDN U29598 ( .B(n29769), .A(n29770), .Z(n29767) );
  XOR U29599 ( .A(n29768), .B(n29771), .Z(n29769) );
  XOR U29600 ( .A(n29772), .B(n29773), .Z(n29743) );
  XNOR U29601 ( .A(n29738), .B(n29774), .Z(n29773) );
  IV U29602 ( .A(n29741), .Z(n29774) );
  XOR U29603 ( .A(n29775), .B(n29776), .Z(n29741) );
  ANDN U29604 ( .B(n29777), .A(n29778), .Z(n29775) );
  XOR U29605 ( .A(n29776), .B(n29779), .Z(n29777) );
  XNOR U29606 ( .A(n29780), .B(n29781), .Z(n29738) );
  ANDN U29607 ( .B(n29782), .A(n29783), .Z(n29780) );
  XOR U29608 ( .A(n29781), .B(n29784), .Z(n29782) );
  IV U29609 ( .A(n29737), .Z(n29772) );
  XOR U29610 ( .A(n29735), .B(n29785), .Z(n29737) );
  XNOR U29611 ( .A(n29786), .B(n29787), .Z(n29785) );
  ANDN U29612 ( .B(n29788), .A(n29789), .Z(n29786) );
  XNOR U29613 ( .A(n29790), .B(n29791), .Z(n29788) );
  IV U29614 ( .A(n29739), .Z(n29735) );
  XOR U29615 ( .A(n29792), .B(n29793), .Z(n29739) );
  ANDN U29616 ( .B(n29794), .A(n29795), .Z(n29792) );
  XOR U29617 ( .A(n29796), .B(n29793), .Z(n29794) );
  XOR U29618 ( .A(n29750), .B(n29603), .Z(n29751) );
  XOR U29619 ( .A(n29797), .B(n29798), .Z(n29603) );
  AND U29620 ( .A(n368), .B(n29799), .Z(n29797) );
  XOR U29621 ( .A(n29800), .B(n29798), .Z(n29799) );
  XNOR U29622 ( .A(n29801), .B(n29802), .Z(n29750) );
  NAND U29623 ( .A(n29803), .B(n29804), .Z(n29802) );
  XOR U29624 ( .A(n29805), .B(n29702), .Z(n29804) );
  XOR U29625 ( .A(n29778), .B(n29779), .Z(n29702) );
  XOR U29626 ( .A(n29806), .B(n29771), .Z(n29779) );
  XOR U29627 ( .A(n29807), .B(n29759), .Z(n29771) );
  XOR U29628 ( .A(n29808), .B(n29809), .Z(n29759) );
  ANDN U29629 ( .B(n29810), .A(n29811), .Z(n29808) );
  XOR U29630 ( .A(n29809), .B(n29812), .Z(n29810) );
  IV U29631 ( .A(n29757), .Z(n29807) );
  XOR U29632 ( .A(n29755), .B(n29813), .Z(n29757) );
  XOR U29633 ( .A(n29814), .B(n29815), .Z(n29813) );
  ANDN U29634 ( .B(n29816), .A(n29817), .Z(n29814) );
  XOR U29635 ( .A(n29818), .B(n29815), .Z(n29816) );
  IV U29636 ( .A(n29758), .Z(n29755) );
  XOR U29637 ( .A(n29819), .B(n29820), .Z(n29758) );
  ANDN U29638 ( .B(n29821), .A(n29822), .Z(n29819) );
  XOR U29639 ( .A(n29820), .B(n29823), .Z(n29821) );
  IV U29640 ( .A(n29770), .Z(n29806) );
  XOR U29641 ( .A(n29824), .B(n29825), .Z(n29770) );
  XNOR U29642 ( .A(n29765), .B(n29826), .Z(n29825) );
  IV U29643 ( .A(n29768), .Z(n29826) );
  XOR U29644 ( .A(n29827), .B(n29828), .Z(n29768) );
  ANDN U29645 ( .B(n29829), .A(n29830), .Z(n29827) );
  XOR U29646 ( .A(n29828), .B(n29831), .Z(n29829) );
  XNOR U29647 ( .A(n29832), .B(n29833), .Z(n29765) );
  ANDN U29648 ( .B(n29834), .A(n29835), .Z(n29832) );
  XOR U29649 ( .A(n29833), .B(n29836), .Z(n29834) );
  IV U29650 ( .A(n29764), .Z(n29824) );
  XOR U29651 ( .A(n29762), .B(n29837), .Z(n29764) );
  XOR U29652 ( .A(n29838), .B(n29839), .Z(n29837) );
  ANDN U29653 ( .B(n29840), .A(n29841), .Z(n29838) );
  XOR U29654 ( .A(n29842), .B(n29839), .Z(n29840) );
  IV U29655 ( .A(n29766), .Z(n29762) );
  XOR U29656 ( .A(n29843), .B(n29844), .Z(n29766) );
  ANDN U29657 ( .B(n29845), .A(n29846), .Z(n29843) );
  XOR U29658 ( .A(n29847), .B(n29844), .Z(n29845) );
  XOR U29659 ( .A(n29848), .B(n29849), .Z(n29778) );
  XOR U29660 ( .A(n29796), .B(n29850), .Z(n29849) );
  IV U29661 ( .A(n29776), .Z(n29850) );
  XOR U29662 ( .A(n29851), .B(n29852), .Z(n29776) );
  ANDN U29663 ( .B(n29853), .A(n29854), .Z(n29851) );
  XOR U29664 ( .A(n29852), .B(n29855), .Z(n29853) );
  XOR U29665 ( .A(n29856), .B(n29784), .Z(n29796) );
  XOR U29666 ( .A(n29857), .B(n29858), .Z(n29784) );
  ANDN U29667 ( .B(n29859), .A(n29860), .Z(n29857) );
  XOR U29668 ( .A(n29858), .B(n29861), .Z(n29859) );
  IV U29669 ( .A(n29783), .Z(n29856) );
  XOR U29670 ( .A(n29862), .B(n29863), .Z(n29783) );
  XOR U29671 ( .A(n29864), .B(n29865), .Z(n29863) );
  ANDN U29672 ( .B(n29866), .A(n29867), .Z(n29864) );
  XOR U29673 ( .A(n29868), .B(n29865), .Z(n29866) );
  IV U29674 ( .A(n29781), .Z(n29862) );
  XOR U29675 ( .A(n29869), .B(n29870), .Z(n29781) );
  ANDN U29676 ( .B(n29871), .A(n29872), .Z(n29869) );
  XOR U29677 ( .A(n29870), .B(n29873), .Z(n29871) );
  IV U29678 ( .A(n29795), .Z(n29848) );
  XOR U29679 ( .A(n29874), .B(n29875), .Z(n29795) );
  XNOR U29680 ( .A(n29790), .B(n29876), .Z(n29875) );
  IV U29681 ( .A(n29793), .Z(n29876) );
  XOR U29682 ( .A(n29877), .B(n29878), .Z(n29793) );
  ANDN U29683 ( .B(n29879), .A(n29880), .Z(n29877) );
  XOR U29684 ( .A(n29881), .B(n29878), .Z(n29879) );
  XNOR U29685 ( .A(n29882), .B(n29883), .Z(n29790) );
  ANDN U29686 ( .B(n29884), .A(n29885), .Z(n29882) );
  XOR U29687 ( .A(n29883), .B(n29886), .Z(n29884) );
  IV U29688 ( .A(n29789), .Z(n29874) );
  XOR U29689 ( .A(n29787), .B(n29887), .Z(n29789) );
  XOR U29690 ( .A(n29888), .B(n29889), .Z(n29887) );
  ANDN U29691 ( .B(n29890), .A(n29891), .Z(n29888) );
  XOR U29692 ( .A(n29892), .B(n29889), .Z(n29890) );
  IV U29693 ( .A(n29791), .Z(n29787) );
  XOR U29694 ( .A(n29893), .B(n29894), .Z(n29791) );
  ANDN U29695 ( .B(n29895), .A(n29896), .Z(n29893) );
  XOR U29696 ( .A(n29897), .B(n29894), .Z(n29895) );
  IV U29697 ( .A(n29801), .Z(n29805) );
  XOR U29698 ( .A(n29801), .B(n29704), .Z(n29803) );
  XOR U29699 ( .A(n29898), .B(n29899), .Z(n29704) );
  AND U29700 ( .A(n368), .B(n29900), .Z(n29898) );
  XOR U29701 ( .A(n29901), .B(n29899), .Z(n29900) );
  NANDN U29702 ( .A(n29706), .B(n29708), .Z(n29801) );
  XOR U29703 ( .A(n29902), .B(n29903), .Z(n29708) );
  AND U29704 ( .A(n368), .B(n29904), .Z(n29902) );
  XOR U29705 ( .A(n29903), .B(n29905), .Z(n29904) );
  XNOR U29706 ( .A(n29906), .B(n29907), .Z(n368) );
  AND U29707 ( .A(n29908), .B(n29909), .Z(n29906) );
  XOR U29708 ( .A(n29907), .B(n29719), .Z(n29909) );
  XNOR U29709 ( .A(n29910), .B(n29911), .Z(n29719) );
  ANDN U29710 ( .B(n29912), .A(n29913), .Z(n29910) );
  XOR U29711 ( .A(n29911), .B(n29914), .Z(n29912) );
  XNOR U29712 ( .A(n29907), .B(n29721), .Z(n29908) );
  XOR U29713 ( .A(n29915), .B(n29916), .Z(n29721) );
  AND U29714 ( .A(n372), .B(n29917), .Z(n29915) );
  XOR U29715 ( .A(n29918), .B(n29916), .Z(n29917) );
  XOR U29716 ( .A(n29919), .B(n29920), .Z(n29907) );
  AND U29717 ( .A(n29921), .B(n29922), .Z(n29919) );
  XOR U29718 ( .A(n29920), .B(n29746), .Z(n29922) );
  XOR U29719 ( .A(n29913), .B(n29914), .Z(n29746) );
  XNOR U29720 ( .A(n29923), .B(n29924), .Z(n29914) );
  ANDN U29721 ( .B(n29925), .A(n29926), .Z(n29923) );
  XOR U29722 ( .A(n29927), .B(n29928), .Z(n29925) );
  XOR U29723 ( .A(n29929), .B(n29930), .Z(n29913) );
  XNOR U29724 ( .A(n29931), .B(n29932), .Z(n29930) );
  ANDN U29725 ( .B(n29933), .A(n29934), .Z(n29931) );
  XNOR U29726 ( .A(n29935), .B(n29936), .Z(n29933) );
  IV U29727 ( .A(n29911), .Z(n29929) );
  XOR U29728 ( .A(n29937), .B(n29938), .Z(n29911) );
  ANDN U29729 ( .B(n29939), .A(n29940), .Z(n29937) );
  XOR U29730 ( .A(n29938), .B(n29941), .Z(n29939) );
  XNOR U29731 ( .A(n29920), .B(n29748), .Z(n29921) );
  XOR U29732 ( .A(n29942), .B(n29943), .Z(n29748) );
  AND U29733 ( .A(n372), .B(n29944), .Z(n29942) );
  XOR U29734 ( .A(n29945), .B(n29943), .Z(n29944) );
  XNOR U29735 ( .A(n29946), .B(n29947), .Z(n29920) );
  AND U29736 ( .A(n29948), .B(n29949), .Z(n29946) );
  XNOR U29737 ( .A(n29947), .B(n29798), .Z(n29949) );
  XOR U29738 ( .A(n29940), .B(n29941), .Z(n29798) );
  XOR U29739 ( .A(n29950), .B(n29928), .Z(n29941) );
  XNOR U29740 ( .A(n29951), .B(n29952), .Z(n29928) );
  ANDN U29741 ( .B(n29953), .A(n29954), .Z(n29951) );
  XOR U29742 ( .A(n29955), .B(n29956), .Z(n29953) );
  IV U29743 ( .A(n29926), .Z(n29950) );
  XOR U29744 ( .A(n29924), .B(n29957), .Z(n29926) );
  XNOR U29745 ( .A(n29958), .B(n29959), .Z(n29957) );
  ANDN U29746 ( .B(n29960), .A(n29961), .Z(n29958) );
  XNOR U29747 ( .A(n29962), .B(n29963), .Z(n29960) );
  IV U29748 ( .A(n29927), .Z(n29924) );
  XOR U29749 ( .A(n29964), .B(n29965), .Z(n29927) );
  ANDN U29750 ( .B(n29966), .A(n29967), .Z(n29964) );
  XOR U29751 ( .A(n29965), .B(n29968), .Z(n29966) );
  XOR U29752 ( .A(n29969), .B(n29970), .Z(n29940) );
  XNOR U29753 ( .A(n29935), .B(n29971), .Z(n29970) );
  IV U29754 ( .A(n29938), .Z(n29971) );
  XOR U29755 ( .A(n29972), .B(n29973), .Z(n29938) );
  ANDN U29756 ( .B(n29974), .A(n29975), .Z(n29972) );
  XOR U29757 ( .A(n29973), .B(n29976), .Z(n29974) );
  XNOR U29758 ( .A(n29977), .B(n29978), .Z(n29935) );
  ANDN U29759 ( .B(n29979), .A(n29980), .Z(n29977) );
  XOR U29760 ( .A(n29978), .B(n29981), .Z(n29979) );
  IV U29761 ( .A(n29934), .Z(n29969) );
  XOR U29762 ( .A(n29932), .B(n29982), .Z(n29934) );
  XNOR U29763 ( .A(n29983), .B(n29984), .Z(n29982) );
  ANDN U29764 ( .B(n29985), .A(n29986), .Z(n29983) );
  XNOR U29765 ( .A(n29987), .B(n29988), .Z(n29985) );
  IV U29766 ( .A(n29936), .Z(n29932) );
  XOR U29767 ( .A(n29989), .B(n29990), .Z(n29936) );
  ANDN U29768 ( .B(n29991), .A(n29992), .Z(n29989) );
  XOR U29769 ( .A(n29993), .B(n29990), .Z(n29991) );
  XOR U29770 ( .A(n29947), .B(n29800), .Z(n29948) );
  XOR U29771 ( .A(n29994), .B(n29995), .Z(n29800) );
  AND U29772 ( .A(n372), .B(n29996), .Z(n29994) );
  XOR U29773 ( .A(n29997), .B(n29995), .Z(n29996) );
  XNOR U29774 ( .A(n29998), .B(n29999), .Z(n29947) );
  NAND U29775 ( .A(n30000), .B(n30001), .Z(n29999) );
  XOR U29776 ( .A(n30002), .B(n29899), .Z(n30001) );
  XOR U29777 ( .A(n29975), .B(n29976), .Z(n29899) );
  XOR U29778 ( .A(n30003), .B(n29968), .Z(n29976) );
  XOR U29779 ( .A(n30004), .B(n29956), .Z(n29968) );
  XOR U29780 ( .A(n30005), .B(n30006), .Z(n29956) );
  ANDN U29781 ( .B(n30007), .A(n30008), .Z(n30005) );
  XOR U29782 ( .A(n30006), .B(n30009), .Z(n30007) );
  IV U29783 ( .A(n29954), .Z(n30004) );
  XOR U29784 ( .A(n29952), .B(n30010), .Z(n29954) );
  XOR U29785 ( .A(n30011), .B(n30012), .Z(n30010) );
  ANDN U29786 ( .B(n30013), .A(n30014), .Z(n30011) );
  XOR U29787 ( .A(n30015), .B(n30012), .Z(n30013) );
  IV U29788 ( .A(n29955), .Z(n29952) );
  XOR U29789 ( .A(n30016), .B(n30017), .Z(n29955) );
  ANDN U29790 ( .B(n30018), .A(n30019), .Z(n30016) );
  XOR U29791 ( .A(n30017), .B(n30020), .Z(n30018) );
  IV U29792 ( .A(n29967), .Z(n30003) );
  XOR U29793 ( .A(n30021), .B(n30022), .Z(n29967) );
  XNOR U29794 ( .A(n29962), .B(n30023), .Z(n30022) );
  IV U29795 ( .A(n29965), .Z(n30023) );
  XOR U29796 ( .A(n30024), .B(n30025), .Z(n29965) );
  ANDN U29797 ( .B(n30026), .A(n30027), .Z(n30024) );
  XOR U29798 ( .A(n30025), .B(n30028), .Z(n30026) );
  XNOR U29799 ( .A(n30029), .B(n30030), .Z(n29962) );
  ANDN U29800 ( .B(n30031), .A(n30032), .Z(n30029) );
  XOR U29801 ( .A(n30030), .B(n30033), .Z(n30031) );
  IV U29802 ( .A(n29961), .Z(n30021) );
  XOR U29803 ( .A(n29959), .B(n30034), .Z(n29961) );
  XOR U29804 ( .A(n30035), .B(n30036), .Z(n30034) );
  ANDN U29805 ( .B(n30037), .A(n30038), .Z(n30035) );
  XOR U29806 ( .A(n30039), .B(n30036), .Z(n30037) );
  IV U29807 ( .A(n29963), .Z(n29959) );
  XOR U29808 ( .A(n30040), .B(n30041), .Z(n29963) );
  ANDN U29809 ( .B(n30042), .A(n30043), .Z(n30040) );
  XOR U29810 ( .A(n30044), .B(n30041), .Z(n30042) );
  XOR U29811 ( .A(n30045), .B(n30046), .Z(n29975) );
  XOR U29812 ( .A(n29993), .B(n30047), .Z(n30046) );
  IV U29813 ( .A(n29973), .Z(n30047) );
  XOR U29814 ( .A(n30048), .B(n30049), .Z(n29973) );
  ANDN U29815 ( .B(n30050), .A(n30051), .Z(n30048) );
  XOR U29816 ( .A(n30049), .B(n30052), .Z(n30050) );
  XOR U29817 ( .A(n30053), .B(n29981), .Z(n29993) );
  XOR U29818 ( .A(n30054), .B(n30055), .Z(n29981) );
  ANDN U29819 ( .B(n30056), .A(n30057), .Z(n30054) );
  XOR U29820 ( .A(n30055), .B(n30058), .Z(n30056) );
  IV U29821 ( .A(n29980), .Z(n30053) );
  XOR U29822 ( .A(n30059), .B(n30060), .Z(n29980) );
  XOR U29823 ( .A(n30061), .B(n30062), .Z(n30060) );
  ANDN U29824 ( .B(n30063), .A(n30064), .Z(n30061) );
  XOR U29825 ( .A(n30065), .B(n30062), .Z(n30063) );
  IV U29826 ( .A(n29978), .Z(n30059) );
  XOR U29827 ( .A(n30066), .B(n30067), .Z(n29978) );
  ANDN U29828 ( .B(n30068), .A(n30069), .Z(n30066) );
  XOR U29829 ( .A(n30067), .B(n30070), .Z(n30068) );
  IV U29830 ( .A(n29992), .Z(n30045) );
  XOR U29831 ( .A(n30071), .B(n30072), .Z(n29992) );
  XNOR U29832 ( .A(n29987), .B(n30073), .Z(n30072) );
  IV U29833 ( .A(n29990), .Z(n30073) );
  XOR U29834 ( .A(n30074), .B(n30075), .Z(n29990) );
  ANDN U29835 ( .B(n30076), .A(n30077), .Z(n30074) );
  XOR U29836 ( .A(n30078), .B(n30075), .Z(n30076) );
  XNOR U29837 ( .A(n30079), .B(n30080), .Z(n29987) );
  ANDN U29838 ( .B(n30081), .A(n30082), .Z(n30079) );
  XOR U29839 ( .A(n30080), .B(n30083), .Z(n30081) );
  IV U29840 ( .A(n29986), .Z(n30071) );
  XOR U29841 ( .A(n29984), .B(n30084), .Z(n29986) );
  XOR U29842 ( .A(n30085), .B(n30086), .Z(n30084) );
  ANDN U29843 ( .B(n30087), .A(n30088), .Z(n30085) );
  XOR U29844 ( .A(n30089), .B(n30086), .Z(n30087) );
  IV U29845 ( .A(n29988), .Z(n29984) );
  XOR U29846 ( .A(n30090), .B(n30091), .Z(n29988) );
  ANDN U29847 ( .B(n30092), .A(n30093), .Z(n30090) );
  XOR U29848 ( .A(n30094), .B(n30091), .Z(n30092) );
  IV U29849 ( .A(n29998), .Z(n30002) );
  XOR U29850 ( .A(n29998), .B(n29901), .Z(n30000) );
  XOR U29851 ( .A(n30095), .B(n30096), .Z(n29901) );
  AND U29852 ( .A(n372), .B(n30097), .Z(n30095) );
  XOR U29853 ( .A(n30098), .B(n30096), .Z(n30097) );
  NANDN U29854 ( .A(n29903), .B(n29905), .Z(n29998) );
  XOR U29855 ( .A(n30099), .B(n30100), .Z(n29905) );
  AND U29856 ( .A(n372), .B(n30101), .Z(n30099) );
  XOR U29857 ( .A(n30100), .B(n30102), .Z(n30101) );
  XNOR U29858 ( .A(n30103), .B(n30104), .Z(n372) );
  AND U29859 ( .A(n30105), .B(n30106), .Z(n30103) );
  XOR U29860 ( .A(n30104), .B(n29916), .Z(n30106) );
  XNOR U29861 ( .A(n30107), .B(n30108), .Z(n29916) );
  ANDN U29862 ( .B(n30109), .A(n30110), .Z(n30107) );
  XOR U29863 ( .A(n30108), .B(n30111), .Z(n30109) );
  XNOR U29864 ( .A(n30104), .B(n29918), .Z(n30105) );
  XOR U29865 ( .A(n30112), .B(n30113), .Z(n29918) );
  AND U29866 ( .A(n376), .B(n30114), .Z(n30112) );
  XOR U29867 ( .A(n30115), .B(n30113), .Z(n30114) );
  XOR U29868 ( .A(n30116), .B(n30117), .Z(n30104) );
  AND U29869 ( .A(n30118), .B(n30119), .Z(n30116) );
  XOR U29870 ( .A(n30117), .B(n29943), .Z(n30119) );
  XOR U29871 ( .A(n30110), .B(n30111), .Z(n29943) );
  XNOR U29872 ( .A(n30120), .B(n30121), .Z(n30111) );
  ANDN U29873 ( .B(n30122), .A(n30123), .Z(n30120) );
  XOR U29874 ( .A(n30124), .B(n30125), .Z(n30122) );
  XOR U29875 ( .A(n30126), .B(n30127), .Z(n30110) );
  XNOR U29876 ( .A(n30128), .B(n30129), .Z(n30127) );
  ANDN U29877 ( .B(n30130), .A(n30131), .Z(n30128) );
  XNOR U29878 ( .A(n30132), .B(n30133), .Z(n30130) );
  IV U29879 ( .A(n30108), .Z(n30126) );
  XOR U29880 ( .A(n30134), .B(n30135), .Z(n30108) );
  ANDN U29881 ( .B(n30136), .A(n30137), .Z(n30134) );
  XOR U29882 ( .A(n30135), .B(n30138), .Z(n30136) );
  XNOR U29883 ( .A(n30117), .B(n29945), .Z(n30118) );
  XOR U29884 ( .A(n30139), .B(n30140), .Z(n29945) );
  AND U29885 ( .A(n376), .B(n30141), .Z(n30139) );
  XOR U29886 ( .A(n30142), .B(n30140), .Z(n30141) );
  XNOR U29887 ( .A(n30143), .B(n30144), .Z(n30117) );
  AND U29888 ( .A(n30145), .B(n30146), .Z(n30143) );
  XNOR U29889 ( .A(n30144), .B(n29995), .Z(n30146) );
  XOR U29890 ( .A(n30137), .B(n30138), .Z(n29995) );
  XOR U29891 ( .A(n30147), .B(n30125), .Z(n30138) );
  XNOR U29892 ( .A(n30148), .B(n30149), .Z(n30125) );
  ANDN U29893 ( .B(n30150), .A(n30151), .Z(n30148) );
  XOR U29894 ( .A(n30152), .B(n30153), .Z(n30150) );
  IV U29895 ( .A(n30123), .Z(n30147) );
  XOR U29896 ( .A(n30121), .B(n30154), .Z(n30123) );
  XNOR U29897 ( .A(n30155), .B(n30156), .Z(n30154) );
  ANDN U29898 ( .B(n30157), .A(n30158), .Z(n30155) );
  XNOR U29899 ( .A(n30159), .B(n30160), .Z(n30157) );
  IV U29900 ( .A(n30124), .Z(n30121) );
  XOR U29901 ( .A(n30161), .B(n30162), .Z(n30124) );
  ANDN U29902 ( .B(n30163), .A(n30164), .Z(n30161) );
  XOR U29903 ( .A(n30162), .B(n30165), .Z(n30163) );
  XOR U29904 ( .A(n30166), .B(n30167), .Z(n30137) );
  XNOR U29905 ( .A(n30132), .B(n30168), .Z(n30167) );
  IV U29906 ( .A(n30135), .Z(n30168) );
  XOR U29907 ( .A(n30169), .B(n30170), .Z(n30135) );
  ANDN U29908 ( .B(n30171), .A(n30172), .Z(n30169) );
  XOR U29909 ( .A(n30170), .B(n30173), .Z(n30171) );
  XNOR U29910 ( .A(n30174), .B(n30175), .Z(n30132) );
  ANDN U29911 ( .B(n30176), .A(n30177), .Z(n30174) );
  XOR U29912 ( .A(n30175), .B(n30178), .Z(n30176) );
  IV U29913 ( .A(n30131), .Z(n30166) );
  XOR U29914 ( .A(n30129), .B(n30179), .Z(n30131) );
  XNOR U29915 ( .A(n30180), .B(n30181), .Z(n30179) );
  ANDN U29916 ( .B(n30182), .A(n30183), .Z(n30180) );
  XNOR U29917 ( .A(n30184), .B(n30185), .Z(n30182) );
  IV U29918 ( .A(n30133), .Z(n30129) );
  XOR U29919 ( .A(n30186), .B(n30187), .Z(n30133) );
  ANDN U29920 ( .B(n30188), .A(n30189), .Z(n30186) );
  XOR U29921 ( .A(n30190), .B(n30187), .Z(n30188) );
  XOR U29922 ( .A(n30144), .B(n29997), .Z(n30145) );
  XOR U29923 ( .A(n30191), .B(n30192), .Z(n29997) );
  AND U29924 ( .A(n376), .B(n30193), .Z(n30191) );
  XOR U29925 ( .A(n30194), .B(n30192), .Z(n30193) );
  XNOR U29926 ( .A(n30195), .B(n30196), .Z(n30144) );
  NAND U29927 ( .A(n30197), .B(n30198), .Z(n30196) );
  XOR U29928 ( .A(n30199), .B(n30096), .Z(n30198) );
  XOR U29929 ( .A(n30172), .B(n30173), .Z(n30096) );
  XOR U29930 ( .A(n30200), .B(n30165), .Z(n30173) );
  XOR U29931 ( .A(n30201), .B(n30153), .Z(n30165) );
  XOR U29932 ( .A(n30202), .B(n30203), .Z(n30153) );
  ANDN U29933 ( .B(n30204), .A(n30205), .Z(n30202) );
  XOR U29934 ( .A(n30203), .B(n30206), .Z(n30204) );
  IV U29935 ( .A(n30151), .Z(n30201) );
  XOR U29936 ( .A(n30149), .B(n30207), .Z(n30151) );
  XOR U29937 ( .A(n30208), .B(n30209), .Z(n30207) );
  ANDN U29938 ( .B(n30210), .A(n30211), .Z(n30208) );
  XOR U29939 ( .A(n30212), .B(n30209), .Z(n30210) );
  IV U29940 ( .A(n30152), .Z(n30149) );
  XOR U29941 ( .A(n30213), .B(n30214), .Z(n30152) );
  ANDN U29942 ( .B(n30215), .A(n30216), .Z(n30213) );
  XOR U29943 ( .A(n30214), .B(n30217), .Z(n30215) );
  IV U29944 ( .A(n30164), .Z(n30200) );
  XOR U29945 ( .A(n30218), .B(n30219), .Z(n30164) );
  XNOR U29946 ( .A(n30159), .B(n30220), .Z(n30219) );
  IV U29947 ( .A(n30162), .Z(n30220) );
  XOR U29948 ( .A(n30221), .B(n30222), .Z(n30162) );
  ANDN U29949 ( .B(n30223), .A(n30224), .Z(n30221) );
  XOR U29950 ( .A(n30222), .B(n30225), .Z(n30223) );
  XNOR U29951 ( .A(n30226), .B(n30227), .Z(n30159) );
  ANDN U29952 ( .B(n30228), .A(n30229), .Z(n30226) );
  XOR U29953 ( .A(n30227), .B(n30230), .Z(n30228) );
  IV U29954 ( .A(n30158), .Z(n30218) );
  XOR U29955 ( .A(n30156), .B(n30231), .Z(n30158) );
  XOR U29956 ( .A(n30232), .B(n30233), .Z(n30231) );
  ANDN U29957 ( .B(n30234), .A(n30235), .Z(n30232) );
  XOR U29958 ( .A(n30236), .B(n30233), .Z(n30234) );
  IV U29959 ( .A(n30160), .Z(n30156) );
  XOR U29960 ( .A(n30237), .B(n30238), .Z(n30160) );
  ANDN U29961 ( .B(n30239), .A(n30240), .Z(n30237) );
  XOR U29962 ( .A(n30241), .B(n30238), .Z(n30239) );
  XOR U29963 ( .A(n30242), .B(n30243), .Z(n30172) );
  XOR U29964 ( .A(n30190), .B(n30244), .Z(n30243) );
  IV U29965 ( .A(n30170), .Z(n30244) );
  XOR U29966 ( .A(n30245), .B(n30246), .Z(n30170) );
  ANDN U29967 ( .B(n30247), .A(n30248), .Z(n30245) );
  XOR U29968 ( .A(n30246), .B(n30249), .Z(n30247) );
  XOR U29969 ( .A(n30250), .B(n30178), .Z(n30190) );
  XOR U29970 ( .A(n30251), .B(n30252), .Z(n30178) );
  ANDN U29971 ( .B(n30253), .A(n30254), .Z(n30251) );
  XOR U29972 ( .A(n30252), .B(n30255), .Z(n30253) );
  IV U29973 ( .A(n30177), .Z(n30250) );
  XOR U29974 ( .A(n30256), .B(n30257), .Z(n30177) );
  XOR U29975 ( .A(n30258), .B(n30259), .Z(n30257) );
  ANDN U29976 ( .B(n30260), .A(n30261), .Z(n30258) );
  XOR U29977 ( .A(n30262), .B(n30259), .Z(n30260) );
  IV U29978 ( .A(n30175), .Z(n30256) );
  XOR U29979 ( .A(n30263), .B(n30264), .Z(n30175) );
  ANDN U29980 ( .B(n30265), .A(n30266), .Z(n30263) );
  XOR U29981 ( .A(n30264), .B(n30267), .Z(n30265) );
  IV U29982 ( .A(n30189), .Z(n30242) );
  XOR U29983 ( .A(n30268), .B(n30269), .Z(n30189) );
  XNOR U29984 ( .A(n30184), .B(n30270), .Z(n30269) );
  IV U29985 ( .A(n30187), .Z(n30270) );
  XOR U29986 ( .A(n30271), .B(n30272), .Z(n30187) );
  ANDN U29987 ( .B(n30273), .A(n30274), .Z(n30271) );
  XOR U29988 ( .A(n30275), .B(n30272), .Z(n30273) );
  XNOR U29989 ( .A(n30276), .B(n30277), .Z(n30184) );
  ANDN U29990 ( .B(n30278), .A(n30279), .Z(n30276) );
  XOR U29991 ( .A(n30277), .B(n30280), .Z(n30278) );
  IV U29992 ( .A(n30183), .Z(n30268) );
  XOR U29993 ( .A(n30181), .B(n30281), .Z(n30183) );
  XOR U29994 ( .A(n30282), .B(n30283), .Z(n30281) );
  ANDN U29995 ( .B(n30284), .A(n30285), .Z(n30282) );
  XOR U29996 ( .A(n30286), .B(n30283), .Z(n30284) );
  IV U29997 ( .A(n30185), .Z(n30181) );
  XOR U29998 ( .A(n30287), .B(n30288), .Z(n30185) );
  ANDN U29999 ( .B(n30289), .A(n30290), .Z(n30287) );
  XOR U30000 ( .A(n30291), .B(n30288), .Z(n30289) );
  IV U30001 ( .A(n30195), .Z(n30199) );
  XOR U30002 ( .A(n30195), .B(n30098), .Z(n30197) );
  XOR U30003 ( .A(n30292), .B(n30293), .Z(n30098) );
  AND U30004 ( .A(n376), .B(n30294), .Z(n30292) );
  XOR U30005 ( .A(n30295), .B(n30293), .Z(n30294) );
  NANDN U30006 ( .A(n30100), .B(n30102), .Z(n30195) );
  XOR U30007 ( .A(n30296), .B(n30297), .Z(n30102) );
  AND U30008 ( .A(n376), .B(n30298), .Z(n30296) );
  XOR U30009 ( .A(n30297), .B(n30299), .Z(n30298) );
  XNOR U30010 ( .A(n30300), .B(n30301), .Z(n376) );
  AND U30011 ( .A(n30302), .B(n30303), .Z(n30300) );
  XOR U30012 ( .A(n30301), .B(n30113), .Z(n30303) );
  XNOR U30013 ( .A(n30304), .B(n30305), .Z(n30113) );
  ANDN U30014 ( .B(n30306), .A(n30307), .Z(n30304) );
  XOR U30015 ( .A(n30305), .B(n30308), .Z(n30306) );
  XNOR U30016 ( .A(n30301), .B(n30115), .Z(n30302) );
  XOR U30017 ( .A(n30309), .B(n30310), .Z(n30115) );
  AND U30018 ( .A(n380), .B(n30311), .Z(n30309) );
  XOR U30019 ( .A(n30312), .B(n30310), .Z(n30311) );
  XOR U30020 ( .A(n30313), .B(n30314), .Z(n30301) );
  AND U30021 ( .A(n30315), .B(n30316), .Z(n30313) );
  XOR U30022 ( .A(n30314), .B(n30140), .Z(n30316) );
  XOR U30023 ( .A(n30307), .B(n30308), .Z(n30140) );
  XNOR U30024 ( .A(n30317), .B(n30318), .Z(n30308) );
  ANDN U30025 ( .B(n30319), .A(n30320), .Z(n30317) );
  XOR U30026 ( .A(n30321), .B(n30322), .Z(n30319) );
  XOR U30027 ( .A(n30323), .B(n30324), .Z(n30307) );
  XNOR U30028 ( .A(n30325), .B(n30326), .Z(n30324) );
  ANDN U30029 ( .B(n30327), .A(n30328), .Z(n30325) );
  XNOR U30030 ( .A(n30329), .B(n30330), .Z(n30327) );
  IV U30031 ( .A(n30305), .Z(n30323) );
  XOR U30032 ( .A(n30331), .B(n30332), .Z(n30305) );
  ANDN U30033 ( .B(n30333), .A(n30334), .Z(n30331) );
  XOR U30034 ( .A(n30332), .B(n30335), .Z(n30333) );
  XNOR U30035 ( .A(n30314), .B(n30142), .Z(n30315) );
  XOR U30036 ( .A(n30336), .B(n30337), .Z(n30142) );
  AND U30037 ( .A(n380), .B(n30338), .Z(n30336) );
  XOR U30038 ( .A(n30339), .B(n30337), .Z(n30338) );
  XNOR U30039 ( .A(n30340), .B(n30341), .Z(n30314) );
  AND U30040 ( .A(n30342), .B(n30343), .Z(n30340) );
  XNOR U30041 ( .A(n30341), .B(n30192), .Z(n30343) );
  XOR U30042 ( .A(n30334), .B(n30335), .Z(n30192) );
  XOR U30043 ( .A(n30344), .B(n30322), .Z(n30335) );
  XNOR U30044 ( .A(n30345), .B(n30346), .Z(n30322) );
  ANDN U30045 ( .B(n30347), .A(n30348), .Z(n30345) );
  XOR U30046 ( .A(n30349), .B(n30350), .Z(n30347) );
  IV U30047 ( .A(n30320), .Z(n30344) );
  XOR U30048 ( .A(n30318), .B(n30351), .Z(n30320) );
  XNOR U30049 ( .A(n30352), .B(n30353), .Z(n30351) );
  ANDN U30050 ( .B(n30354), .A(n30355), .Z(n30352) );
  XNOR U30051 ( .A(n30356), .B(n30357), .Z(n30354) );
  IV U30052 ( .A(n30321), .Z(n30318) );
  XOR U30053 ( .A(n30358), .B(n30359), .Z(n30321) );
  ANDN U30054 ( .B(n30360), .A(n30361), .Z(n30358) );
  XOR U30055 ( .A(n30359), .B(n30362), .Z(n30360) );
  XOR U30056 ( .A(n30363), .B(n30364), .Z(n30334) );
  XNOR U30057 ( .A(n30329), .B(n30365), .Z(n30364) );
  IV U30058 ( .A(n30332), .Z(n30365) );
  XOR U30059 ( .A(n30366), .B(n30367), .Z(n30332) );
  ANDN U30060 ( .B(n30368), .A(n30369), .Z(n30366) );
  XOR U30061 ( .A(n30367), .B(n30370), .Z(n30368) );
  XNOR U30062 ( .A(n30371), .B(n30372), .Z(n30329) );
  ANDN U30063 ( .B(n30373), .A(n30374), .Z(n30371) );
  XOR U30064 ( .A(n30372), .B(n30375), .Z(n30373) );
  IV U30065 ( .A(n30328), .Z(n30363) );
  XOR U30066 ( .A(n30326), .B(n30376), .Z(n30328) );
  XNOR U30067 ( .A(n30377), .B(n30378), .Z(n30376) );
  ANDN U30068 ( .B(n30379), .A(n30380), .Z(n30377) );
  XNOR U30069 ( .A(n30381), .B(n30382), .Z(n30379) );
  IV U30070 ( .A(n30330), .Z(n30326) );
  XOR U30071 ( .A(n30383), .B(n30384), .Z(n30330) );
  ANDN U30072 ( .B(n30385), .A(n30386), .Z(n30383) );
  XOR U30073 ( .A(n30387), .B(n30384), .Z(n30385) );
  XOR U30074 ( .A(n30341), .B(n30194), .Z(n30342) );
  XOR U30075 ( .A(n30388), .B(n30389), .Z(n30194) );
  AND U30076 ( .A(n380), .B(n30390), .Z(n30388) );
  XOR U30077 ( .A(n30391), .B(n30389), .Z(n30390) );
  XNOR U30078 ( .A(n30392), .B(n30393), .Z(n30341) );
  NAND U30079 ( .A(n30394), .B(n30395), .Z(n30393) );
  XOR U30080 ( .A(n30396), .B(n30293), .Z(n30395) );
  XOR U30081 ( .A(n30369), .B(n30370), .Z(n30293) );
  XOR U30082 ( .A(n30397), .B(n30362), .Z(n30370) );
  XOR U30083 ( .A(n30398), .B(n30350), .Z(n30362) );
  XOR U30084 ( .A(n30399), .B(n30400), .Z(n30350) );
  ANDN U30085 ( .B(n30401), .A(n30402), .Z(n30399) );
  XOR U30086 ( .A(n30400), .B(n30403), .Z(n30401) );
  IV U30087 ( .A(n30348), .Z(n30398) );
  XOR U30088 ( .A(n30346), .B(n30404), .Z(n30348) );
  XOR U30089 ( .A(n30405), .B(n30406), .Z(n30404) );
  ANDN U30090 ( .B(n30407), .A(n30408), .Z(n30405) );
  XOR U30091 ( .A(n30409), .B(n30406), .Z(n30407) );
  IV U30092 ( .A(n30349), .Z(n30346) );
  XOR U30093 ( .A(n30410), .B(n30411), .Z(n30349) );
  ANDN U30094 ( .B(n30412), .A(n30413), .Z(n30410) );
  XOR U30095 ( .A(n30411), .B(n30414), .Z(n30412) );
  IV U30096 ( .A(n30361), .Z(n30397) );
  XOR U30097 ( .A(n30415), .B(n30416), .Z(n30361) );
  XNOR U30098 ( .A(n30356), .B(n30417), .Z(n30416) );
  IV U30099 ( .A(n30359), .Z(n30417) );
  XOR U30100 ( .A(n30418), .B(n30419), .Z(n30359) );
  ANDN U30101 ( .B(n30420), .A(n30421), .Z(n30418) );
  XOR U30102 ( .A(n30419), .B(n30422), .Z(n30420) );
  XNOR U30103 ( .A(n30423), .B(n30424), .Z(n30356) );
  ANDN U30104 ( .B(n30425), .A(n30426), .Z(n30423) );
  XOR U30105 ( .A(n30424), .B(n30427), .Z(n30425) );
  IV U30106 ( .A(n30355), .Z(n30415) );
  XOR U30107 ( .A(n30353), .B(n30428), .Z(n30355) );
  XOR U30108 ( .A(n30429), .B(n30430), .Z(n30428) );
  ANDN U30109 ( .B(n30431), .A(n30432), .Z(n30429) );
  XOR U30110 ( .A(n30433), .B(n30430), .Z(n30431) );
  IV U30111 ( .A(n30357), .Z(n30353) );
  XOR U30112 ( .A(n30434), .B(n30435), .Z(n30357) );
  ANDN U30113 ( .B(n30436), .A(n30437), .Z(n30434) );
  XOR U30114 ( .A(n30438), .B(n30435), .Z(n30436) );
  XOR U30115 ( .A(n30439), .B(n30440), .Z(n30369) );
  XOR U30116 ( .A(n30387), .B(n30441), .Z(n30440) );
  IV U30117 ( .A(n30367), .Z(n30441) );
  XOR U30118 ( .A(n30442), .B(n30443), .Z(n30367) );
  ANDN U30119 ( .B(n30444), .A(n30445), .Z(n30442) );
  XOR U30120 ( .A(n30443), .B(n30446), .Z(n30444) );
  XOR U30121 ( .A(n30447), .B(n30375), .Z(n30387) );
  XOR U30122 ( .A(n30448), .B(n30449), .Z(n30375) );
  ANDN U30123 ( .B(n30450), .A(n30451), .Z(n30448) );
  XOR U30124 ( .A(n30449), .B(n30452), .Z(n30450) );
  IV U30125 ( .A(n30374), .Z(n30447) );
  XOR U30126 ( .A(n30453), .B(n30454), .Z(n30374) );
  XOR U30127 ( .A(n30455), .B(n30456), .Z(n30454) );
  ANDN U30128 ( .B(n30457), .A(n30458), .Z(n30455) );
  XOR U30129 ( .A(n30459), .B(n30456), .Z(n30457) );
  IV U30130 ( .A(n30372), .Z(n30453) );
  XOR U30131 ( .A(n30460), .B(n30461), .Z(n30372) );
  ANDN U30132 ( .B(n30462), .A(n30463), .Z(n30460) );
  XOR U30133 ( .A(n30461), .B(n30464), .Z(n30462) );
  IV U30134 ( .A(n30386), .Z(n30439) );
  XOR U30135 ( .A(n30465), .B(n30466), .Z(n30386) );
  XNOR U30136 ( .A(n30381), .B(n30467), .Z(n30466) );
  IV U30137 ( .A(n30384), .Z(n30467) );
  XOR U30138 ( .A(n30468), .B(n30469), .Z(n30384) );
  ANDN U30139 ( .B(n30470), .A(n30471), .Z(n30468) );
  XOR U30140 ( .A(n30472), .B(n30469), .Z(n30470) );
  XNOR U30141 ( .A(n30473), .B(n30474), .Z(n30381) );
  ANDN U30142 ( .B(n30475), .A(n30476), .Z(n30473) );
  XOR U30143 ( .A(n30474), .B(n30477), .Z(n30475) );
  IV U30144 ( .A(n30380), .Z(n30465) );
  XOR U30145 ( .A(n30378), .B(n30478), .Z(n30380) );
  XOR U30146 ( .A(n30479), .B(n30480), .Z(n30478) );
  ANDN U30147 ( .B(n30481), .A(n30482), .Z(n30479) );
  XOR U30148 ( .A(n30483), .B(n30480), .Z(n30481) );
  IV U30149 ( .A(n30382), .Z(n30378) );
  XOR U30150 ( .A(n30484), .B(n30485), .Z(n30382) );
  ANDN U30151 ( .B(n30486), .A(n30487), .Z(n30484) );
  XOR U30152 ( .A(n30488), .B(n30485), .Z(n30486) );
  IV U30153 ( .A(n30392), .Z(n30396) );
  XOR U30154 ( .A(n30392), .B(n30295), .Z(n30394) );
  XOR U30155 ( .A(n30489), .B(n30490), .Z(n30295) );
  AND U30156 ( .A(n380), .B(n30491), .Z(n30489) );
  XOR U30157 ( .A(n30492), .B(n30490), .Z(n30491) );
  NANDN U30158 ( .A(n30297), .B(n30299), .Z(n30392) );
  XOR U30159 ( .A(n30493), .B(n30494), .Z(n30299) );
  AND U30160 ( .A(n380), .B(n30495), .Z(n30493) );
  XOR U30161 ( .A(n30494), .B(n30496), .Z(n30495) );
  XNOR U30162 ( .A(n30497), .B(n30498), .Z(n380) );
  AND U30163 ( .A(n30499), .B(n30500), .Z(n30497) );
  XOR U30164 ( .A(n30498), .B(n30310), .Z(n30500) );
  XNOR U30165 ( .A(n30501), .B(n30502), .Z(n30310) );
  ANDN U30166 ( .B(n30503), .A(n30504), .Z(n30501) );
  XOR U30167 ( .A(n30502), .B(n30505), .Z(n30503) );
  XNOR U30168 ( .A(n30498), .B(n30312), .Z(n30499) );
  XOR U30169 ( .A(n30506), .B(n30507), .Z(n30312) );
  AND U30170 ( .A(n384), .B(n30508), .Z(n30506) );
  XOR U30171 ( .A(n30509), .B(n30507), .Z(n30508) );
  XOR U30172 ( .A(n30510), .B(n30511), .Z(n30498) );
  AND U30173 ( .A(n30512), .B(n30513), .Z(n30510) );
  XOR U30174 ( .A(n30511), .B(n30337), .Z(n30513) );
  XOR U30175 ( .A(n30504), .B(n30505), .Z(n30337) );
  XNOR U30176 ( .A(n30514), .B(n30515), .Z(n30505) );
  ANDN U30177 ( .B(n30516), .A(n30517), .Z(n30514) );
  XOR U30178 ( .A(n30518), .B(n30519), .Z(n30516) );
  XOR U30179 ( .A(n30520), .B(n30521), .Z(n30504) );
  XNOR U30180 ( .A(n30522), .B(n30523), .Z(n30521) );
  ANDN U30181 ( .B(n30524), .A(n30525), .Z(n30522) );
  XNOR U30182 ( .A(n30526), .B(n30527), .Z(n30524) );
  IV U30183 ( .A(n30502), .Z(n30520) );
  XOR U30184 ( .A(n30528), .B(n30529), .Z(n30502) );
  ANDN U30185 ( .B(n30530), .A(n30531), .Z(n30528) );
  XOR U30186 ( .A(n30529), .B(n30532), .Z(n30530) );
  XNOR U30187 ( .A(n30511), .B(n30339), .Z(n30512) );
  XOR U30188 ( .A(n30533), .B(n30534), .Z(n30339) );
  AND U30189 ( .A(n384), .B(n30535), .Z(n30533) );
  XOR U30190 ( .A(n30536), .B(n30534), .Z(n30535) );
  XNOR U30191 ( .A(n30537), .B(n30538), .Z(n30511) );
  AND U30192 ( .A(n30539), .B(n30540), .Z(n30537) );
  XNOR U30193 ( .A(n30538), .B(n30389), .Z(n30540) );
  XOR U30194 ( .A(n30531), .B(n30532), .Z(n30389) );
  XOR U30195 ( .A(n30541), .B(n30519), .Z(n30532) );
  XNOR U30196 ( .A(n30542), .B(n30543), .Z(n30519) );
  ANDN U30197 ( .B(n30544), .A(n30545), .Z(n30542) );
  XOR U30198 ( .A(n30546), .B(n30547), .Z(n30544) );
  IV U30199 ( .A(n30517), .Z(n30541) );
  XOR U30200 ( .A(n30515), .B(n30548), .Z(n30517) );
  XNOR U30201 ( .A(n30549), .B(n30550), .Z(n30548) );
  ANDN U30202 ( .B(n30551), .A(n30552), .Z(n30549) );
  XNOR U30203 ( .A(n30553), .B(n30554), .Z(n30551) );
  IV U30204 ( .A(n30518), .Z(n30515) );
  XOR U30205 ( .A(n30555), .B(n30556), .Z(n30518) );
  ANDN U30206 ( .B(n30557), .A(n30558), .Z(n30555) );
  XOR U30207 ( .A(n30556), .B(n30559), .Z(n30557) );
  XOR U30208 ( .A(n30560), .B(n30561), .Z(n30531) );
  XNOR U30209 ( .A(n30526), .B(n30562), .Z(n30561) );
  IV U30210 ( .A(n30529), .Z(n30562) );
  XOR U30211 ( .A(n30563), .B(n30564), .Z(n30529) );
  ANDN U30212 ( .B(n30565), .A(n30566), .Z(n30563) );
  XOR U30213 ( .A(n30564), .B(n30567), .Z(n30565) );
  XNOR U30214 ( .A(n30568), .B(n30569), .Z(n30526) );
  ANDN U30215 ( .B(n30570), .A(n30571), .Z(n30568) );
  XOR U30216 ( .A(n30569), .B(n30572), .Z(n30570) );
  IV U30217 ( .A(n30525), .Z(n30560) );
  XOR U30218 ( .A(n30523), .B(n30573), .Z(n30525) );
  XNOR U30219 ( .A(n30574), .B(n30575), .Z(n30573) );
  ANDN U30220 ( .B(n30576), .A(n30577), .Z(n30574) );
  XNOR U30221 ( .A(n30578), .B(n30579), .Z(n30576) );
  IV U30222 ( .A(n30527), .Z(n30523) );
  XOR U30223 ( .A(n30580), .B(n30581), .Z(n30527) );
  ANDN U30224 ( .B(n30582), .A(n30583), .Z(n30580) );
  XOR U30225 ( .A(n30584), .B(n30581), .Z(n30582) );
  XOR U30226 ( .A(n30538), .B(n30391), .Z(n30539) );
  XOR U30227 ( .A(n30585), .B(n30586), .Z(n30391) );
  AND U30228 ( .A(n384), .B(n30587), .Z(n30585) );
  XOR U30229 ( .A(n30588), .B(n30586), .Z(n30587) );
  XNOR U30230 ( .A(n30589), .B(n30590), .Z(n30538) );
  NAND U30231 ( .A(n30591), .B(n30592), .Z(n30590) );
  XOR U30232 ( .A(n30593), .B(n30490), .Z(n30592) );
  XOR U30233 ( .A(n30566), .B(n30567), .Z(n30490) );
  XOR U30234 ( .A(n30594), .B(n30559), .Z(n30567) );
  XOR U30235 ( .A(n30595), .B(n30547), .Z(n30559) );
  XOR U30236 ( .A(n30596), .B(n30597), .Z(n30547) );
  ANDN U30237 ( .B(n30598), .A(n30599), .Z(n30596) );
  XOR U30238 ( .A(n30597), .B(n30600), .Z(n30598) );
  IV U30239 ( .A(n30545), .Z(n30595) );
  XOR U30240 ( .A(n30543), .B(n30601), .Z(n30545) );
  XOR U30241 ( .A(n30602), .B(n30603), .Z(n30601) );
  ANDN U30242 ( .B(n30604), .A(n30605), .Z(n30602) );
  XOR U30243 ( .A(n30606), .B(n30603), .Z(n30604) );
  IV U30244 ( .A(n30546), .Z(n30543) );
  XOR U30245 ( .A(n30607), .B(n30608), .Z(n30546) );
  ANDN U30246 ( .B(n30609), .A(n30610), .Z(n30607) );
  XOR U30247 ( .A(n30608), .B(n30611), .Z(n30609) );
  IV U30248 ( .A(n30558), .Z(n30594) );
  XOR U30249 ( .A(n30612), .B(n30613), .Z(n30558) );
  XNOR U30250 ( .A(n30553), .B(n30614), .Z(n30613) );
  IV U30251 ( .A(n30556), .Z(n30614) );
  XOR U30252 ( .A(n30615), .B(n30616), .Z(n30556) );
  ANDN U30253 ( .B(n30617), .A(n30618), .Z(n30615) );
  XOR U30254 ( .A(n30616), .B(n30619), .Z(n30617) );
  XNOR U30255 ( .A(n30620), .B(n30621), .Z(n30553) );
  ANDN U30256 ( .B(n30622), .A(n30623), .Z(n30620) );
  XOR U30257 ( .A(n30621), .B(n30624), .Z(n30622) );
  IV U30258 ( .A(n30552), .Z(n30612) );
  XOR U30259 ( .A(n30550), .B(n30625), .Z(n30552) );
  XOR U30260 ( .A(n30626), .B(n30627), .Z(n30625) );
  ANDN U30261 ( .B(n30628), .A(n30629), .Z(n30626) );
  XOR U30262 ( .A(n30630), .B(n30627), .Z(n30628) );
  IV U30263 ( .A(n30554), .Z(n30550) );
  XOR U30264 ( .A(n30631), .B(n30632), .Z(n30554) );
  ANDN U30265 ( .B(n30633), .A(n30634), .Z(n30631) );
  XOR U30266 ( .A(n30635), .B(n30632), .Z(n30633) );
  XOR U30267 ( .A(n30636), .B(n30637), .Z(n30566) );
  XOR U30268 ( .A(n30584), .B(n30638), .Z(n30637) );
  IV U30269 ( .A(n30564), .Z(n30638) );
  XOR U30270 ( .A(n30639), .B(n30640), .Z(n30564) );
  ANDN U30271 ( .B(n30641), .A(n30642), .Z(n30639) );
  XOR U30272 ( .A(n30640), .B(n30643), .Z(n30641) );
  XOR U30273 ( .A(n30644), .B(n30572), .Z(n30584) );
  XOR U30274 ( .A(n30645), .B(n30646), .Z(n30572) );
  ANDN U30275 ( .B(n30647), .A(n30648), .Z(n30645) );
  XOR U30276 ( .A(n30646), .B(n30649), .Z(n30647) );
  IV U30277 ( .A(n30571), .Z(n30644) );
  XOR U30278 ( .A(n30650), .B(n30651), .Z(n30571) );
  XOR U30279 ( .A(n30652), .B(n30653), .Z(n30651) );
  ANDN U30280 ( .B(n30654), .A(n30655), .Z(n30652) );
  XOR U30281 ( .A(n30656), .B(n30653), .Z(n30654) );
  IV U30282 ( .A(n30569), .Z(n30650) );
  XOR U30283 ( .A(n30657), .B(n30658), .Z(n30569) );
  ANDN U30284 ( .B(n30659), .A(n30660), .Z(n30657) );
  XOR U30285 ( .A(n30658), .B(n30661), .Z(n30659) );
  IV U30286 ( .A(n30583), .Z(n30636) );
  XOR U30287 ( .A(n30662), .B(n30663), .Z(n30583) );
  XNOR U30288 ( .A(n30578), .B(n30664), .Z(n30663) );
  IV U30289 ( .A(n30581), .Z(n30664) );
  XOR U30290 ( .A(n30665), .B(n30666), .Z(n30581) );
  ANDN U30291 ( .B(n30667), .A(n30668), .Z(n30665) );
  XOR U30292 ( .A(n30669), .B(n30666), .Z(n30667) );
  XNOR U30293 ( .A(n30670), .B(n30671), .Z(n30578) );
  ANDN U30294 ( .B(n30672), .A(n30673), .Z(n30670) );
  XOR U30295 ( .A(n30671), .B(n30674), .Z(n30672) );
  IV U30296 ( .A(n30577), .Z(n30662) );
  XOR U30297 ( .A(n30575), .B(n30675), .Z(n30577) );
  XOR U30298 ( .A(n30676), .B(n30677), .Z(n30675) );
  ANDN U30299 ( .B(n30678), .A(n30679), .Z(n30676) );
  XOR U30300 ( .A(n30680), .B(n30677), .Z(n30678) );
  IV U30301 ( .A(n30579), .Z(n30575) );
  XOR U30302 ( .A(n30681), .B(n30682), .Z(n30579) );
  ANDN U30303 ( .B(n30683), .A(n30684), .Z(n30681) );
  XOR U30304 ( .A(n30685), .B(n30682), .Z(n30683) );
  IV U30305 ( .A(n30589), .Z(n30593) );
  XOR U30306 ( .A(n30589), .B(n30492), .Z(n30591) );
  XOR U30307 ( .A(n30686), .B(n30687), .Z(n30492) );
  AND U30308 ( .A(n384), .B(n30688), .Z(n30686) );
  XOR U30309 ( .A(n30689), .B(n30687), .Z(n30688) );
  NANDN U30310 ( .A(n30494), .B(n30496), .Z(n30589) );
  XOR U30311 ( .A(n30690), .B(n30691), .Z(n30496) );
  AND U30312 ( .A(n384), .B(n30692), .Z(n30690) );
  XOR U30313 ( .A(n30691), .B(n30693), .Z(n30692) );
  XNOR U30314 ( .A(n30694), .B(n30695), .Z(n384) );
  AND U30315 ( .A(n30696), .B(n30697), .Z(n30694) );
  XOR U30316 ( .A(n30695), .B(n30507), .Z(n30697) );
  XNOR U30317 ( .A(n30698), .B(n30699), .Z(n30507) );
  ANDN U30318 ( .B(n30700), .A(n30701), .Z(n30698) );
  XOR U30319 ( .A(n30699), .B(n30702), .Z(n30700) );
  XNOR U30320 ( .A(n30695), .B(n30509), .Z(n30696) );
  XOR U30321 ( .A(n30703), .B(n30704), .Z(n30509) );
  AND U30322 ( .A(n388), .B(n30705), .Z(n30703) );
  XOR U30323 ( .A(n30706), .B(n30704), .Z(n30705) );
  XOR U30324 ( .A(n30707), .B(n30708), .Z(n30695) );
  AND U30325 ( .A(n30709), .B(n30710), .Z(n30707) );
  XOR U30326 ( .A(n30708), .B(n30534), .Z(n30710) );
  XOR U30327 ( .A(n30701), .B(n30702), .Z(n30534) );
  XNOR U30328 ( .A(n30711), .B(n30712), .Z(n30702) );
  ANDN U30329 ( .B(n30713), .A(n30714), .Z(n30711) );
  XOR U30330 ( .A(n30715), .B(n30716), .Z(n30713) );
  XOR U30331 ( .A(n30717), .B(n30718), .Z(n30701) );
  XNOR U30332 ( .A(n30719), .B(n30720), .Z(n30718) );
  ANDN U30333 ( .B(n30721), .A(n30722), .Z(n30719) );
  XNOR U30334 ( .A(n30723), .B(n30724), .Z(n30721) );
  IV U30335 ( .A(n30699), .Z(n30717) );
  XOR U30336 ( .A(n30725), .B(n30726), .Z(n30699) );
  ANDN U30337 ( .B(n30727), .A(n30728), .Z(n30725) );
  XOR U30338 ( .A(n30726), .B(n30729), .Z(n30727) );
  XNOR U30339 ( .A(n30708), .B(n30536), .Z(n30709) );
  XOR U30340 ( .A(n30730), .B(n30731), .Z(n30536) );
  AND U30341 ( .A(n388), .B(n30732), .Z(n30730) );
  XOR U30342 ( .A(n30733), .B(n30731), .Z(n30732) );
  XNOR U30343 ( .A(n30734), .B(n30735), .Z(n30708) );
  AND U30344 ( .A(n30736), .B(n30737), .Z(n30734) );
  XNOR U30345 ( .A(n30735), .B(n30586), .Z(n30737) );
  XOR U30346 ( .A(n30728), .B(n30729), .Z(n30586) );
  XOR U30347 ( .A(n30738), .B(n30716), .Z(n30729) );
  XNOR U30348 ( .A(n30739), .B(n30740), .Z(n30716) );
  ANDN U30349 ( .B(n30741), .A(n30742), .Z(n30739) );
  XOR U30350 ( .A(n30743), .B(n30744), .Z(n30741) );
  IV U30351 ( .A(n30714), .Z(n30738) );
  XOR U30352 ( .A(n30712), .B(n30745), .Z(n30714) );
  XNOR U30353 ( .A(n30746), .B(n30747), .Z(n30745) );
  ANDN U30354 ( .B(n30748), .A(n30749), .Z(n30746) );
  XNOR U30355 ( .A(n30750), .B(n30751), .Z(n30748) );
  IV U30356 ( .A(n30715), .Z(n30712) );
  XOR U30357 ( .A(n30752), .B(n30753), .Z(n30715) );
  ANDN U30358 ( .B(n30754), .A(n30755), .Z(n30752) );
  XOR U30359 ( .A(n30753), .B(n30756), .Z(n30754) );
  XOR U30360 ( .A(n30757), .B(n30758), .Z(n30728) );
  XNOR U30361 ( .A(n30723), .B(n30759), .Z(n30758) );
  IV U30362 ( .A(n30726), .Z(n30759) );
  XOR U30363 ( .A(n30760), .B(n30761), .Z(n30726) );
  ANDN U30364 ( .B(n30762), .A(n30763), .Z(n30760) );
  XOR U30365 ( .A(n30761), .B(n30764), .Z(n30762) );
  XNOR U30366 ( .A(n30765), .B(n30766), .Z(n30723) );
  ANDN U30367 ( .B(n30767), .A(n30768), .Z(n30765) );
  XOR U30368 ( .A(n30766), .B(n30769), .Z(n30767) );
  IV U30369 ( .A(n30722), .Z(n30757) );
  XOR U30370 ( .A(n30720), .B(n30770), .Z(n30722) );
  XNOR U30371 ( .A(n30771), .B(n30772), .Z(n30770) );
  ANDN U30372 ( .B(n30773), .A(n30774), .Z(n30771) );
  XNOR U30373 ( .A(n30775), .B(n30776), .Z(n30773) );
  IV U30374 ( .A(n30724), .Z(n30720) );
  XOR U30375 ( .A(n30777), .B(n30778), .Z(n30724) );
  ANDN U30376 ( .B(n30779), .A(n30780), .Z(n30777) );
  XOR U30377 ( .A(n30781), .B(n30778), .Z(n30779) );
  XOR U30378 ( .A(n30735), .B(n30588), .Z(n30736) );
  XOR U30379 ( .A(n30782), .B(n30783), .Z(n30588) );
  AND U30380 ( .A(n388), .B(n30784), .Z(n30782) );
  XOR U30381 ( .A(n30785), .B(n30783), .Z(n30784) );
  XNOR U30382 ( .A(n30786), .B(n30787), .Z(n30735) );
  NAND U30383 ( .A(n30788), .B(n30789), .Z(n30787) );
  XOR U30384 ( .A(n30790), .B(n30687), .Z(n30789) );
  XOR U30385 ( .A(n30763), .B(n30764), .Z(n30687) );
  XOR U30386 ( .A(n30791), .B(n30756), .Z(n30764) );
  XOR U30387 ( .A(n30792), .B(n30744), .Z(n30756) );
  XOR U30388 ( .A(n30793), .B(n30794), .Z(n30744) );
  ANDN U30389 ( .B(n30795), .A(n30796), .Z(n30793) );
  XOR U30390 ( .A(n30794), .B(n30797), .Z(n30795) );
  IV U30391 ( .A(n30742), .Z(n30792) );
  XOR U30392 ( .A(n30740), .B(n30798), .Z(n30742) );
  XOR U30393 ( .A(n30799), .B(n30800), .Z(n30798) );
  ANDN U30394 ( .B(n30801), .A(n30802), .Z(n30799) );
  XOR U30395 ( .A(n30803), .B(n30800), .Z(n30801) );
  IV U30396 ( .A(n30743), .Z(n30740) );
  XOR U30397 ( .A(n30804), .B(n30805), .Z(n30743) );
  ANDN U30398 ( .B(n30806), .A(n30807), .Z(n30804) );
  XOR U30399 ( .A(n30805), .B(n30808), .Z(n30806) );
  IV U30400 ( .A(n30755), .Z(n30791) );
  XOR U30401 ( .A(n30809), .B(n30810), .Z(n30755) );
  XNOR U30402 ( .A(n30750), .B(n30811), .Z(n30810) );
  IV U30403 ( .A(n30753), .Z(n30811) );
  XOR U30404 ( .A(n30812), .B(n30813), .Z(n30753) );
  ANDN U30405 ( .B(n30814), .A(n30815), .Z(n30812) );
  XOR U30406 ( .A(n30813), .B(n30816), .Z(n30814) );
  XNOR U30407 ( .A(n30817), .B(n30818), .Z(n30750) );
  ANDN U30408 ( .B(n30819), .A(n30820), .Z(n30817) );
  XOR U30409 ( .A(n30818), .B(n30821), .Z(n30819) );
  IV U30410 ( .A(n30749), .Z(n30809) );
  XOR U30411 ( .A(n30747), .B(n30822), .Z(n30749) );
  XOR U30412 ( .A(n30823), .B(n30824), .Z(n30822) );
  ANDN U30413 ( .B(n30825), .A(n30826), .Z(n30823) );
  XOR U30414 ( .A(n30827), .B(n30824), .Z(n30825) );
  IV U30415 ( .A(n30751), .Z(n30747) );
  XOR U30416 ( .A(n30828), .B(n30829), .Z(n30751) );
  ANDN U30417 ( .B(n30830), .A(n30831), .Z(n30828) );
  XOR U30418 ( .A(n30832), .B(n30829), .Z(n30830) );
  XOR U30419 ( .A(n30833), .B(n30834), .Z(n30763) );
  XOR U30420 ( .A(n30781), .B(n30835), .Z(n30834) );
  IV U30421 ( .A(n30761), .Z(n30835) );
  XOR U30422 ( .A(n30836), .B(n30837), .Z(n30761) );
  ANDN U30423 ( .B(n30838), .A(n30839), .Z(n30836) );
  XOR U30424 ( .A(n30837), .B(n30840), .Z(n30838) );
  XOR U30425 ( .A(n30841), .B(n30769), .Z(n30781) );
  XOR U30426 ( .A(n30842), .B(n30843), .Z(n30769) );
  ANDN U30427 ( .B(n30844), .A(n30845), .Z(n30842) );
  XOR U30428 ( .A(n30843), .B(n30846), .Z(n30844) );
  IV U30429 ( .A(n30768), .Z(n30841) );
  XOR U30430 ( .A(n30847), .B(n30848), .Z(n30768) );
  XOR U30431 ( .A(n30849), .B(n30850), .Z(n30848) );
  ANDN U30432 ( .B(n30851), .A(n30852), .Z(n30849) );
  XOR U30433 ( .A(n30853), .B(n30850), .Z(n30851) );
  IV U30434 ( .A(n30766), .Z(n30847) );
  XOR U30435 ( .A(n30854), .B(n30855), .Z(n30766) );
  ANDN U30436 ( .B(n30856), .A(n30857), .Z(n30854) );
  XOR U30437 ( .A(n30855), .B(n30858), .Z(n30856) );
  IV U30438 ( .A(n30780), .Z(n30833) );
  XOR U30439 ( .A(n30859), .B(n30860), .Z(n30780) );
  XNOR U30440 ( .A(n30775), .B(n30861), .Z(n30860) );
  IV U30441 ( .A(n30778), .Z(n30861) );
  XOR U30442 ( .A(n30862), .B(n30863), .Z(n30778) );
  ANDN U30443 ( .B(n30864), .A(n30865), .Z(n30862) );
  XOR U30444 ( .A(n30866), .B(n30863), .Z(n30864) );
  XNOR U30445 ( .A(n30867), .B(n30868), .Z(n30775) );
  ANDN U30446 ( .B(n30869), .A(n30870), .Z(n30867) );
  XOR U30447 ( .A(n30868), .B(n30871), .Z(n30869) );
  IV U30448 ( .A(n30774), .Z(n30859) );
  XOR U30449 ( .A(n30772), .B(n30872), .Z(n30774) );
  XOR U30450 ( .A(n30873), .B(n30874), .Z(n30872) );
  ANDN U30451 ( .B(n30875), .A(n30876), .Z(n30873) );
  XOR U30452 ( .A(n30877), .B(n30874), .Z(n30875) );
  IV U30453 ( .A(n30776), .Z(n30772) );
  XOR U30454 ( .A(n30878), .B(n30879), .Z(n30776) );
  ANDN U30455 ( .B(n30880), .A(n30881), .Z(n30878) );
  XOR U30456 ( .A(n30882), .B(n30879), .Z(n30880) );
  IV U30457 ( .A(n30786), .Z(n30790) );
  XOR U30458 ( .A(n30786), .B(n30689), .Z(n30788) );
  XOR U30459 ( .A(n30883), .B(n30884), .Z(n30689) );
  AND U30460 ( .A(n388), .B(n30885), .Z(n30883) );
  XOR U30461 ( .A(n30886), .B(n30884), .Z(n30885) );
  NANDN U30462 ( .A(n30691), .B(n30693), .Z(n30786) );
  XOR U30463 ( .A(n30887), .B(n30888), .Z(n30693) );
  AND U30464 ( .A(n388), .B(n30889), .Z(n30887) );
  XOR U30465 ( .A(n30888), .B(n30890), .Z(n30889) );
  XNOR U30466 ( .A(n30891), .B(n30892), .Z(n388) );
  AND U30467 ( .A(n30893), .B(n30894), .Z(n30891) );
  XOR U30468 ( .A(n30892), .B(n30704), .Z(n30894) );
  XNOR U30469 ( .A(n30895), .B(n30896), .Z(n30704) );
  ANDN U30470 ( .B(n30897), .A(n30898), .Z(n30895) );
  XOR U30471 ( .A(n30896), .B(n30899), .Z(n30897) );
  XNOR U30472 ( .A(n30892), .B(n30706), .Z(n30893) );
  XOR U30473 ( .A(n30900), .B(n30901), .Z(n30706) );
  AND U30474 ( .A(n392), .B(n30902), .Z(n30900) );
  XOR U30475 ( .A(n30903), .B(n30901), .Z(n30902) );
  XOR U30476 ( .A(n30904), .B(n30905), .Z(n30892) );
  AND U30477 ( .A(n30906), .B(n30907), .Z(n30904) );
  XOR U30478 ( .A(n30905), .B(n30731), .Z(n30907) );
  XOR U30479 ( .A(n30898), .B(n30899), .Z(n30731) );
  XNOR U30480 ( .A(n30908), .B(n30909), .Z(n30899) );
  ANDN U30481 ( .B(n30910), .A(n30911), .Z(n30908) );
  XOR U30482 ( .A(n30912), .B(n30913), .Z(n30910) );
  XOR U30483 ( .A(n30914), .B(n30915), .Z(n30898) );
  XNOR U30484 ( .A(n30916), .B(n30917), .Z(n30915) );
  ANDN U30485 ( .B(n30918), .A(n30919), .Z(n30916) );
  XNOR U30486 ( .A(n30920), .B(n30921), .Z(n30918) );
  IV U30487 ( .A(n30896), .Z(n30914) );
  XOR U30488 ( .A(n30922), .B(n30923), .Z(n30896) );
  ANDN U30489 ( .B(n30924), .A(n30925), .Z(n30922) );
  XOR U30490 ( .A(n30923), .B(n30926), .Z(n30924) );
  XNOR U30491 ( .A(n30905), .B(n30733), .Z(n30906) );
  XOR U30492 ( .A(n30927), .B(n30928), .Z(n30733) );
  AND U30493 ( .A(n392), .B(n30929), .Z(n30927) );
  XOR U30494 ( .A(n30930), .B(n30928), .Z(n30929) );
  XNOR U30495 ( .A(n30931), .B(n30932), .Z(n30905) );
  AND U30496 ( .A(n30933), .B(n30934), .Z(n30931) );
  XNOR U30497 ( .A(n30932), .B(n30783), .Z(n30934) );
  XOR U30498 ( .A(n30925), .B(n30926), .Z(n30783) );
  XOR U30499 ( .A(n30935), .B(n30913), .Z(n30926) );
  XNOR U30500 ( .A(n30936), .B(n30937), .Z(n30913) );
  ANDN U30501 ( .B(n30938), .A(n30939), .Z(n30936) );
  XOR U30502 ( .A(n30940), .B(n30941), .Z(n30938) );
  IV U30503 ( .A(n30911), .Z(n30935) );
  XOR U30504 ( .A(n30909), .B(n30942), .Z(n30911) );
  XNOR U30505 ( .A(n30943), .B(n30944), .Z(n30942) );
  ANDN U30506 ( .B(n30945), .A(n30946), .Z(n30943) );
  XNOR U30507 ( .A(n30947), .B(n30948), .Z(n30945) );
  IV U30508 ( .A(n30912), .Z(n30909) );
  XOR U30509 ( .A(n30949), .B(n30950), .Z(n30912) );
  ANDN U30510 ( .B(n30951), .A(n30952), .Z(n30949) );
  XOR U30511 ( .A(n30950), .B(n30953), .Z(n30951) );
  XOR U30512 ( .A(n30954), .B(n30955), .Z(n30925) );
  XNOR U30513 ( .A(n30920), .B(n30956), .Z(n30955) );
  IV U30514 ( .A(n30923), .Z(n30956) );
  XOR U30515 ( .A(n30957), .B(n30958), .Z(n30923) );
  ANDN U30516 ( .B(n30959), .A(n30960), .Z(n30957) );
  XOR U30517 ( .A(n30958), .B(n30961), .Z(n30959) );
  XNOR U30518 ( .A(n30962), .B(n30963), .Z(n30920) );
  ANDN U30519 ( .B(n30964), .A(n30965), .Z(n30962) );
  XOR U30520 ( .A(n30963), .B(n30966), .Z(n30964) );
  IV U30521 ( .A(n30919), .Z(n30954) );
  XOR U30522 ( .A(n30917), .B(n30967), .Z(n30919) );
  XNOR U30523 ( .A(n30968), .B(n30969), .Z(n30967) );
  ANDN U30524 ( .B(n30970), .A(n30971), .Z(n30968) );
  XNOR U30525 ( .A(n30972), .B(n30973), .Z(n30970) );
  IV U30526 ( .A(n30921), .Z(n30917) );
  XOR U30527 ( .A(n30974), .B(n30975), .Z(n30921) );
  ANDN U30528 ( .B(n30976), .A(n30977), .Z(n30974) );
  XOR U30529 ( .A(n30978), .B(n30975), .Z(n30976) );
  XOR U30530 ( .A(n30932), .B(n30785), .Z(n30933) );
  XOR U30531 ( .A(n30979), .B(n30980), .Z(n30785) );
  AND U30532 ( .A(n392), .B(n30981), .Z(n30979) );
  XOR U30533 ( .A(n30982), .B(n30980), .Z(n30981) );
  XNOR U30534 ( .A(n30983), .B(n30984), .Z(n30932) );
  NAND U30535 ( .A(n30985), .B(n30986), .Z(n30984) );
  XOR U30536 ( .A(n30987), .B(n30884), .Z(n30986) );
  XOR U30537 ( .A(n30960), .B(n30961), .Z(n30884) );
  XOR U30538 ( .A(n30988), .B(n30953), .Z(n30961) );
  XOR U30539 ( .A(n30989), .B(n30941), .Z(n30953) );
  XOR U30540 ( .A(n30990), .B(n30991), .Z(n30941) );
  ANDN U30541 ( .B(n30992), .A(n30993), .Z(n30990) );
  XOR U30542 ( .A(n30991), .B(n30994), .Z(n30992) );
  IV U30543 ( .A(n30939), .Z(n30989) );
  XOR U30544 ( .A(n30937), .B(n30995), .Z(n30939) );
  XOR U30545 ( .A(n30996), .B(n30997), .Z(n30995) );
  ANDN U30546 ( .B(n30998), .A(n30999), .Z(n30996) );
  XOR U30547 ( .A(n31000), .B(n30997), .Z(n30998) );
  IV U30548 ( .A(n30940), .Z(n30937) );
  XOR U30549 ( .A(n31001), .B(n31002), .Z(n30940) );
  ANDN U30550 ( .B(n31003), .A(n31004), .Z(n31001) );
  XOR U30551 ( .A(n31002), .B(n31005), .Z(n31003) );
  IV U30552 ( .A(n30952), .Z(n30988) );
  XOR U30553 ( .A(n31006), .B(n31007), .Z(n30952) );
  XNOR U30554 ( .A(n30947), .B(n31008), .Z(n31007) );
  IV U30555 ( .A(n30950), .Z(n31008) );
  XOR U30556 ( .A(n31009), .B(n31010), .Z(n30950) );
  ANDN U30557 ( .B(n31011), .A(n31012), .Z(n31009) );
  XOR U30558 ( .A(n31010), .B(n31013), .Z(n31011) );
  XNOR U30559 ( .A(n31014), .B(n31015), .Z(n30947) );
  ANDN U30560 ( .B(n31016), .A(n31017), .Z(n31014) );
  XOR U30561 ( .A(n31015), .B(n31018), .Z(n31016) );
  IV U30562 ( .A(n30946), .Z(n31006) );
  XOR U30563 ( .A(n30944), .B(n31019), .Z(n30946) );
  XOR U30564 ( .A(n31020), .B(n31021), .Z(n31019) );
  ANDN U30565 ( .B(n31022), .A(n31023), .Z(n31020) );
  XOR U30566 ( .A(n31024), .B(n31021), .Z(n31022) );
  IV U30567 ( .A(n30948), .Z(n30944) );
  XOR U30568 ( .A(n31025), .B(n31026), .Z(n30948) );
  ANDN U30569 ( .B(n31027), .A(n31028), .Z(n31025) );
  XOR U30570 ( .A(n31029), .B(n31026), .Z(n31027) );
  XOR U30571 ( .A(n31030), .B(n31031), .Z(n30960) );
  XOR U30572 ( .A(n30978), .B(n31032), .Z(n31031) );
  IV U30573 ( .A(n30958), .Z(n31032) );
  XOR U30574 ( .A(n31033), .B(n31034), .Z(n30958) );
  ANDN U30575 ( .B(n31035), .A(n31036), .Z(n31033) );
  XOR U30576 ( .A(n31034), .B(n31037), .Z(n31035) );
  XOR U30577 ( .A(n31038), .B(n30966), .Z(n30978) );
  XOR U30578 ( .A(n31039), .B(n31040), .Z(n30966) );
  ANDN U30579 ( .B(n31041), .A(n31042), .Z(n31039) );
  XOR U30580 ( .A(n31040), .B(n31043), .Z(n31041) );
  IV U30581 ( .A(n30965), .Z(n31038) );
  XOR U30582 ( .A(n31044), .B(n31045), .Z(n30965) );
  XOR U30583 ( .A(n31046), .B(n31047), .Z(n31045) );
  ANDN U30584 ( .B(n31048), .A(n31049), .Z(n31046) );
  XOR U30585 ( .A(n31050), .B(n31047), .Z(n31048) );
  IV U30586 ( .A(n30963), .Z(n31044) );
  XOR U30587 ( .A(n31051), .B(n31052), .Z(n30963) );
  ANDN U30588 ( .B(n31053), .A(n31054), .Z(n31051) );
  XOR U30589 ( .A(n31052), .B(n31055), .Z(n31053) );
  IV U30590 ( .A(n30977), .Z(n31030) );
  XOR U30591 ( .A(n31056), .B(n31057), .Z(n30977) );
  XNOR U30592 ( .A(n30972), .B(n31058), .Z(n31057) );
  IV U30593 ( .A(n30975), .Z(n31058) );
  XOR U30594 ( .A(n31059), .B(n31060), .Z(n30975) );
  ANDN U30595 ( .B(n31061), .A(n31062), .Z(n31059) );
  XOR U30596 ( .A(n31063), .B(n31060), .Z(n31061) );
  XNOR U30597 ( .A(n31064), .B(n31065), .Z(n30972) );
  ANDN U30598 ( .B(n31066), .A(n31067), .Z(n31064) );
  XOR U30599 ( .A(n31065), .B(n31068), .Z(n31066) );
  IV U30600 ( .A(n30971), .Z(n31056) );
  XOR U30601 ( .A(n30969), .B(n31069), .Z(n30971) );
  XOR U30602 ( .A(n31070), .B(n31071), .Z(n31069) );
  ANDN U30603 ( .B(n31072), .A(n31073), .Z(n31070) );
  XOR U30604 ( .A(n31074), .B(n31071), .Z(n31072) );
  IV U30605 ( .A(n30973), .Z(n30969) );
  XOR U30606 ( .A(n31075), .B(n31076), .Z(n30973) );
  ANDN U30607 ( .B(n31077), .A(n31078), .Z(n31075) );
  XOR U30608 ( .A(n31079), .B(n31076), .Z(n31077) );
  IV U30609 ( .A(n30983), .Z(n30987) );
  XOR U30610 ( .A(n30983), .B(n30886), .Z(n30985) );
  XOR U30611 ( .A(n31080), .B(n31081), .Z(n30886) );
  AND U30612 ( .A(n392), .B(n31082), .Z(n31080) );
  XOR U30613 ( .A(n31083), .B(n31081), .Z(n31082) );
  NANDN U30614 ( .A(n30888), .B(n30890), .Z(n30983) );
  XOR U30615 ( .A(n31084), .B(n31085), .Z(n30890) );
  AND U30616 ( .A(n392), .B(n31086), .Z(n31084) );
  XOR U30617 ( .A(n31085), .B(n31087), .Z(n31086) );
  XNOR U30618 ( .A(n31088), .B(n31089), .Z(n392) );
  AND U30619 ( .A(n31090), .B(n31091), .Z(n31088) );
  XOR U30620 ( .A(n31089), .B(n30901), .Z(n31091) );
  XNOR U30621 ( .A(n31092), .B(n31093), .Z(n30901) );
  ANDN U30622 ( .B(n31094), .A(n31095), .Z(n31092) );
  XOR U30623 ( .A(n31093), .B(n31096), .Z(n31094) );
  XNOR U30624 ( .A(n31089), .B(n30903), .Z(n31090) );
  XOR U30625 ( .A(n31097), .B(n31098), .Z(n30903) );
  AND U30626 ( .A(n396), .B(n31099), .Z(n31097) );
  XOR U30627 ( .A(n31100), .B(n31098), .Z(n31099) );
  XOR U30628 ( .A(n31101), .B(n31102), .Z(n31089) );
  AND U30629 ( .A(n31103), .B(n31104), .Z(n31101) );
  XOR U30630 ( .A(n31102), .B(n30928), .Z(n31104) );
  XOR U30631 ( .A(n31095), .B(n31096), .Z(n30928) );
  XNOR U30632 ( .A(n31105), .B(n31106), .Z(n31096) );
  ANDN U30633 ( .B(n31107), .A(n31108), .Z(n31105) );
  XOR U30634 ( .A(n31109), .B(n31110), .Z(n31107) );
  XOR U30635 ( .A(n31111), .B(n31112), .Z(n31095) );
  XNOR U30636 ( .A(n31113), .B(n31114), .Z(n31112) );
  ANDN U30637 ( .B(n31115), .A(n31116), .Z(n31113) );
  XNOR U30638 ( .A(n31117), .B(n31118), .Z(n31115) );
  IV U30639 ( .A(n31093), .Z(n31111) );
  XOR U30640 ( .A(n31119), .B(n31120), .Z(n31093) );
  ANDN U30641 ( .B(n31121), .A(n31122), .Z(n31119) );
  XOR U30642 ( .A(n31120), .B(n31123), .Z(n31121) );
  XNOR U30643 ( .A(n31102), .B(n30930), .Z(n31103) );
  XOR U30644 ( .A(n31124), .B(n31125), .Z(n30930) );
  AND U30645 ( .A(n396), .B(n31126), .Z(n31124) );
  XOR U30646 ( .A(n31127), .B(n31125), .Z(n31126) );
  XNOR U30647 ( .A(n31128), .B(n31129), .Z(n31102) );
  AND U30648 ( .A(n31130), .B(n31131), .Z(n31128) );
  XNOR U30649 ( .A(n31129), .B(n30980), .Z(n31131) );
  XOR U30650 ( .A(n31122), .B(n31123), .Z(n30980) );
  XOR U30651 ( .A(n31132), .B(n31110), .Z(n31123) );
  XNOR U30652 ( .A(n31133), .B(n31134), .Z(n31110) );
  ANDN U30653 ( .B(n31135), .A(n31136), .Z(n31133) );
  XOR U30654 ( .A(n31137), .B(n31138), .Z(n31135) );
  IV U30655 ( .A(n31108), .Z(n31132) );
  XOR U30656 ( .A(n31106), .B(n31139), .Z(n31108) );
  XNOR U30657 ( .A(n31140), .B(n31141), .Z(n31139) );
  ANDN U30658 ( .B(n31142), .A(n31143), .Z(n31140) );
  XNOR U30659 ( .A(n31144), .B(n31145), .Z(n31142) );
  IV U30660 ( .A(n31109), .Z(n31106) );
  XOR U30661 ( .A(n31146), .B(n31147), .Z(n31109) );
  ANDN U30662 ( .B(n31148), .A(n31149), .Z(n31146) );
  XOR U30663 ( .A(n31147), .B(n31150), .Z(n31148) );
  XOR U30664 ( .A(n31151), .B(n31152), .Z(n31122) );
  XNOR U30665 ( .A(n31117), .B(n31153), .Z(n31152) );
  IV U30666 ( .A(n31120), .Z(n31153) );
  XOR U30667 ( .A(n31154), .B(n31155), .Z(n31120) );
  ANDN U30668 ( .B(n31156), .A(n31157), .Z(n31154) );
  XOR U30669 ( .A(n31155), .B(n31158), .Z(n31156) );
  XNOR U30670 ( .A(n31159), .B(n31160), .Z(n31117) );
  ANDN U30671 ( .B(n31161), .A(n31162), .Z(n31159) );
  XOR U30672 ( .A(n31160), .B(n31163), .Z(n31161) );
  IV U30673 ( .A(n31116), .Z(n31151) );
  XOR U30674 ( .A(n31114), .B(n31164), .Z(n31116) );
  XNOR U30675 ( .A(n31165), .B(n31166), .Z(n31164) );
  ANDN U30676 ( .B(n31167), .A(n31168), .Z(n31165) );
  XNOR U30677 ( .A(n31169), .B(n31170), .Z(n31167) );
  IV U30678 ( .A(n31118), .Z(n31114) );
  XOR U30679 ( .A(n31171), .B(n31172), .Z(n31118) );
  ANDN U30680 ( .B(n31173), .A(n31174), .Z(n31171) );
  XOR U30681 ( .A(n31175), .B(n31172), .Z(n31173) );
  XOR U30682 ( .A(n31129), .B(n30982), .Z(n31130) );
  XOR U30683 ( .A(n31176), .B(n31177), .Z(n30982) );
  AND U30684 ( .A(n396), .B(n31178), .Z(n31176) );
  XOR U30685 ( .A(n31179), .B(n31177), .Z(n31178) );
  XNOR U30686 ( .A(n31180), .B(n31181), .Z(n31129) );
  NAND U30687 ( .A(n31182), .B(n31183), .Z(n31181) );
  XOR U30688 ( .A(n31184), .B(n31081), .Z(n31183) );
  XOR U30689 ( .A(n31157), .B(n31158), .Z(n31081) );
  XOR U30690 ( .A(n31185), .B(n31150), .Z(n31158) );
  XOR U30691 ( .A(n31186), .B(n31138), .Z(n31150) );
  XOR U30692 ( .A(n31187), .B(n31188), .Z(n31138) );
  ANDN U30693 ( .B(n31189), .A(n31190), .Z(n31187) );
  XOR U30694 ( .A(n31188), .B(n31191), .Z(n31189) );
  IV U30695 ( .A(n31136), .Z(n31186) );
  XOR U30696 ( .A(n31134), .B(n31192), .Z(n31136) );
  XOR U30697 ( .A(n31193), .B(n31194), .Z(n31192) );
  ANDN U30698 ( .B(n31195), .A(n31196), .Z(n31193) );
  XOR U30699 ( .A(n31197), .B(n31194), .Z(n31195) );
  IV U30700 ( .A(n31137), .Z(n31134) );
  XOR U30701 ( .A(n31198), .B(n31199), .Z(n31137) );
  ANDN U30702 ( .B(n31200), .A(n31201), .Z(n31198) );
  XOR U30703 ( .A(n31199), .B(n31202), .Z(n31200) );
  IV U30704 ( .A(n31149), .Z(n31185) );
  XOR U30705 ( .A(n31203), .B(n31204), .Z(n31149) );
  XNOR U30706 ( .A(n31144), .B(n31205), .Z(n31204) );
  IV U30707 ( .A(n31147), .Z(n31205) );
  XOR U30708 ( .A(n31206), .B(n31207), .Z(n31147) );
  ANDN U30709 ( .B(n31208), .A(n31209), .Z(n31206) );
  XOR U30710 ( .A(n31207), .B(n31210), .Z(n31208) );
  XNOR U30711 ( .A(n31211), .B(n31212), .Z(n31144) );
  ANDN U30712 ( .B(n31213), .A(n31214), .Z(n31211) );
  XOR U30713 ( .A(n31212), .B(n31215), .Z(n31213) );
  IV U30714 ( .A(n31143), .Z(n31203) );
  XOR U30715 ( .A(n31141), .B(n31216), .Z(n31143) );
  XOR U30716 ( .A(n31217), .B(n31218), .Z(n31216) );
  ANDN U30717 ( .B(n31219), .A(n31220), .Z(n31217) );
  XOR U30718 ( .A(n31221), .B(n31218), .Z(n31219) );
  IV U30719 ( .A(n31145), .Z(n31141) );
  XOR U30720 ( .A(n31222), .B(n31223), .Z(n31145) );
  ANDN U30721 ( .B(n31224), .A(n31225), .Z(n31222) );
  XOR U30722 ( .A(n31226), .B(n31223), .Z(n31224) );
  XOR U30723 ( .A(n31227), .B(n31228), .Z(n31157) );
  XOR U30724 ( .A(n31175), .B(n31229), .Z(n31228) );
  IV U30725 ( .A(n31155), .Z(n31229) );
  XOR U30726 ( .A(n31230), .B(n31231), .Z(n31155) );
  ANDN U30727 ( .B(n31232), .A(n31233), .Z(n31230) );
  XOR U30728 ( .A(n31231), .B(n31234), .Z(n31232) );
  XOR U30729 ( .A(n31235), .B(n31163), .Z(n31175) );
  XOR U30730 ( .A(n31236), .B(n31237), .Z(n31163) );
  ANDN U30731 ( .B(n31238), .A(n31239), .Z(n31236) );
  XOR U30732 ( .A(n31237), .B(n31240), .Z(n31238) );
  IV U30733 ( .A(n31162), .Z(n31235) );
  XOR U30734 ( .A(n31241), .B(n31242), .Z(n31162) );
  XOR U30735 ( .A(n31243), .B(n31244), .Z(n31242) );
  ANDN U30736 ( .B(n31245), .A(n31246), .Z(n31243) );
  XOR U30737 ( .A(n31247), .B(n31244), .Z(n31245) );
  IV U30738 ( .A(n31160), .Z(n31241) );
  XOR U30739 ( .A(n31248), .B(n31249), .Z(n31160) );
  ANDN U30740 ( .B(n31250), .A(n31251), .Z(n31248) );
  XOR U30741 ( .A(n31249), .B(n31252), .Z(n31250) );
  IV U30742 ( .A(n31174), .Z(n31227) );
  XOR U30743 ( .A(n31253), .B(n31254), .Z(n31174) );
  XNOR U30744 ( .A(n31169), .B(n31255), .Z(n31254) );
  IV U30745 ( .A(n31172), .Z(n31255) );
  XOR U30746 ( .A(n31256), .B(n31257), .Z(n31172) );
  ANDN U30747 ( .B(n31258), .A(n31259), .Z(n31256) );
  XOR U30748 ( .A(n31260), .B(n31257), .Z(n31258) );
  XNOR U30749 ( .A(n31261), .B(n31262), .Z(n31169) );
  ANDN U30750 ( .B(n31263), .A(n31264), .Z(n31261) );
  XOR U30751 ( .A(n31262), .B(n31265), .Z(n31263) );
  IV U30752 ( .A(n31168), .Z(n31253) );
  XOR U30753 ( .A(n31166), .B(n31266), .Z(n31168) );
  XOR U30754 ( .A(n31267), .B(n31268), .Z(n31266) );
  ANDN U30755 ( .B(n31269), .A(n31270), .Z(n31267) );
  XOR U30756 ( .A(n31271), .B(n31268), .Z(n31269) );
  IV U30757 ( .A(n31170), .Z(n31166) );
  XOR U30758 ( .A(n31272), .B(n31273), .Z(n31170) );
  ANDN U30759 ( .B(n31274), .A(n31275), .Z(n31272) );
  XOR U30760 ( .A(n31276), .B(n31273), .Z(n31274) );
  IV U30761 ( .A(n31180), .Z(n31184) );
  XOR U30762 ( .A(n31180), .B(n31083), .Z(n31182) );
  XOR U30763 ( .A(n31277), .B(n31278), .Z(n31083) );
  AND U30764 ( .A(n396), .B(n31279), .Z(n31277) );
  XOR U30765 ( .A(n31280), .B(n31278), .Z(n31279) );
  NANDN U30766 ( .A(n31085), .B(n31087), .Z(n31180) );
  XOR U30767 ( .A(n31281), .B(n31282), .Z(n31087) );
  AND U30768 ( .A(n396), .B(n31283), .Z(n31281) );
  XOR U30769 ( .A(n31282), .B(n31284), .Z(n31283) );
  XNOR U30770 ( .A(n31285), .B(n31286), .Z(n396) );
  AND U30771 ( .A(n31287), .B(n31288), .Z(n31285) );
  XOR U30772 ( .A(n31286), .B(n31098), .Z(n31288) );
  XNOR U30773 ( .A(n31289), .B(n31290), .Z(n31098) );
  ANDN U30774 ( .B(n31291), .A(n31292), .Z(n31289) );
  XOR U30775 ( .A(n31290), .B(n31293), .Z(n31291) );
  XNOR U30776 ( .A(n31286), .B(n31100), .Z(n31287) );
  XOR U30777 ( .A(n31294), .B(n31295), .Z(n31100) );
  AND U30778 ( .A(n400), .B(n31296), .Z(n31294) );
  XOR U30779 ( .A(n31297), .B(n31295), .Z(n31296) );
  XOR U30780 ( .A(n31298), .B(n31299), .Z(n31286) );
  AND U30781 ( .A(n31300), .B(n31301), .Z(n31298) );
  XOR U30782 ( .A(n31299), .B(n31125), .Z(n31301) );
  XOR U30783 ( .A(n31292), .B(n31293), .Z(n31125) );
  XNOR U30784 ( .A(n31302), .B(n31303), .Z(n31293) );
  ANDN U30785 ( .B(n31304), .A(n31305), .Z(n31302) );
  XOR U30786 ( .A(n31306), .B(n31307), .Z(n31304) );
  XOR U30787 ( .A(n31308), .B(n31309), .Z(n31292) );
  XNOR U30788 ( .A(n31310), .B(n31311), .Z(n31309) );
  ANDN U30789 ( .B(n31312), .A(n31313), .Z(n31310) );
  XNOR U30790 ( .A(n31314), .B(n31315), .Z(n31312) );
  IV U30791 ( .A(n31290), .Z(n31308) );
  XOR U30792 ( .A(n31316), .B(n31317), .Z(n31290) );
  ANDN U30793 ( .B(n31318), .A(n31319), .Z(n31316) );
  XOR U30794 ( .A(n31317), .B(n31320), .Z(n31318) );
  XNOR U30795 ( .A(n31299), .B(n31127), .Z(n31300) );
  XOR U30796 ( .A(n31321), .B(n31322), .Z(n31127) );
  AND U30797 ( .A(n400), .B(n31323), .Z(n31321) );
  XOR U30798 ( .A(n31324), .B(n31322), .Z(n31323) );
  XNOR U30799 ( .A(n31325), .B(n31326), .Z(n31299) );
  AND U30800 ( .A(n31327), .B(n31328), .Z(n31325) );
  XNOR U30801 ( .A(n31326), .B(n31177), .Z(n31328) );
  XOR U30802 ( .A(n31319), .B(n31320), .Z(n31177) );
  XOR U30803 ( .A(n31329), .B(n31307), .Z(n31320) );
  XNOR U30804 ( .A(n31330), .B(n31331), .Z(n31307) );
  ANDN U30805 ( .B(n31332), .A(n31333), .Z(n31330) );
  XOR U30806 ( .A(n31334), .B(n31335), .Z(n31332) );
  IV U30807 ( .A(n31305), .Z(n31329) );
  XOR U30808 ( .A(n31303), .B(n31336), .Z(n31305) );
  XNOR U30809 ( .A(n31337), .B(n31338), .Z(n31336) );
  ANDN U30810 ( .B(n31339), .A(n31340), .Z(n31337) );
  XNOR U30811 ( .A(n31341), .B(n31342), .Z(n31339) );
  IV U30812 ( .A(n31306), .Z(n31303) );
  XOR U30813 ( .A(n31343), .B(n31344), .Z(n31306) );
  ANDN U30814 ( .B(n31345), .A(n31346), .Z(n31343) );
  XOR U30815 ( .A(n31344), .B(n31347), .Z(n31345) );
  XOR U30816 ( .A(n31348), .B(n31349), .Z(n31319) );
  XNOR U30817 ( .A(n31314), .B(n31350), .Z(n31349) );
  IV U30818 ( .A(n31317), .Z(n31350) );
  XOR U30819 ( .A(n31351), .B(n31352), .Z(n31317) );
  ANDN U30820 ( .B(n31353), .A(n31354), .Z(n31351) );
  XOR U30821 ( .A(n31352), .B(n31355), .Z(n31353) );
  XNOR U30822 ( .A(n31356), .B(n31357), .Z(n31314) );
  ANDN U30823 ( .B(n31358), .A(n31359), .Z(n31356) );
  XOR U30824 ( .A(n31357), .B(n31360), .Z(n31358) );
  IV U30825 ( .A(n31313), .Z(n31348) );
  XOR U30826 ( .A(n31311), .B(n31361), .Z(n31313) );
  XNOR U30827 ( .A(n31362), .B(n31363), .Z(n31361) );
  ANDN U30828 ( .B(n31364), .A(n31365), .Z(n31362) );
  XNOR U30829 ( .A(n31366), .B(n31367), .Z(n31364) );
  IV U30830 ( .A(n31315), .Z(n31311) );
  XOR U30831 ( .A(n31368), .B(n31369), .Z(n31315) );
  ANDN U30832 ( .B(n31370), .A(n31371), .Z(n31368) );
  XOR U30833 ( .A(n31372), .B(n31369), .Z(n31370) );
  XOR U30834 ( .A(n31326), .B(n31179), .Z(n31327) );
  XOR U30835 ( .A(n31373), .B(n31374), .Z(n31179) );
  AND U30836 ( .A(n400), .B(n31375), .Z(n31373) );
  XOR U30837 ( .A(n31376), .B(n31374), .Z(n31375) );
  XNOR U30838 ( .A(n31377), .B(n31378), .Z(n31326) );
  NAND U30839 ( .A(n31379), .B(n31380), .Z(n31378) );
  XOR U30840 ( .A(n31381), .B(n31278), .Z(n31380) );
  XOR U30841 ( .A(n31354), .B(n31355), .Z(n31278) );
  XOR U30842 ( .A(n31382), .B(n31347), .Z(n31355) );
  XOR U30843 ( .A(n31383), .B(n31335), .Z(n31347) );
  XOR U30844 ( .A(n31384), .B(n31385), .Z(n31335) );
  ANDN U30845 ( .B(n31386), .A(n31387), .Z(n31384) );
  XOR U30846 ( .A(n31385), .B(n31388), .Z(n31386) );
  IV U30847 ( .A(n31333), .Z(n31383) );
  XOR U30848 ( .A(n31331), .B(n31389), .Z(n31333) );
  XOR U30849 ( .A(n31390), .B(n31391), .Z(n31389) );
  ANDN U30850 ( .B(n31392), .A(n31393), .Z(n31390) );
  XOR U30851 ( .A(n31394), .B(n31391), .Z(n31392) );
  IV U30852 ( .A(n31334), .Z(n31331) );
  XOR U30853 ( .A(n31395), .B(n31396), .Z(n31334) );
  ANDN U30854 ( .B(n31397), .A(n31398), .Z(n31395) );
  XOR U30855 ( .A(n31396), .B(n31399), .Z(n31397) );
  IV U30856 ( .A(n31346), .Z(n31382) );
  XOR U30857 ( .A(n31400), .B(n31401), .Z(n31346) );
  XNOR U30858 ( .A(n31341), .B(n31402), .Z(n31401) );
  IV U30859 ( .A(n31344), .Z(n31402) );
  XOR U30860 ( .A(n31403), .B(n31404), .Z(n31344) );
  ANDN U30861 ( .B(n31405), .A(n31406), .Z(n31403) );
  XOR U30862 ( .A(n31404), .B(n31407), .Z(n31405) );
  XNOR U30863 ( .A(n31408), .B(n31409), .Z(n31341) );
  ANDN U30864 ( .B(n31410), .A(n31411), .Z(n31408) );
  XOR U30865 ( .A(n31409), .B(n31412), .Z(n31410) );
  IV U30866 ( .A(n31340), .Z(n31400) );
  XOR U30867 ( .A(n31338), .B(n31413), .Z(n31340) );
  XOR U30868 ( .A(n31414), .B(n31415), .Z(n31413) );
  ANDN U30869 ( .B(n31416), .A(n31417), .Z(n31414) );
  XOR U30870 ( .A(n31418), .B(n31415), .Z(n31416) );
  IV U30871 ( .A(n31342), .Z(n31338) );
  XOR U30872 ( .A(n31419), .B(n31420), .Z(n31342) );
  ANDN U30873 ( .B(n31421), .A(n31422), .Z(n31419) );
  XOR U30874 ( .A(n31423), .B(n31420), .Z(n31421) );
  XOR U30875 ( .A(n31424), .B(n31425), .Z(n31354) );
  XOR U30876 ( .A(n31372), .B(n31426), .Z(n31425) );
  IV U30877 ( .A(n31352), .Z(n31426) );
  XOR U30878 ( .A(n31427), .B(n31428), .Z(n31352) );
  ANDN U30879 ( .B(n31429), .A(n31430), .Z(n31427) );
  XOR U30880 ( .A(n31428), .B(n31431), .Z(n31429) );
  XOR U30881 ( .A(n31432), .B(n31360), .Z(n31372) );
  XOR U30882 ( .A(n31433), .B(n31434), .Z(n31360) );
  ANDN U30883 ( .B(n31435), .A(n31436), .Z(n31433) );
  XOR U30884 ( .A(n31434), .B(n31437), .Z(n31435) );
  IV U30885 ( .A(n31359), .Z(n31432) );
  XOR U30886 ( .A(n31438), .B(n31439), .Z(n31359) );
  XOR U30887 ( .A(n31440), .B(n31441), .Z(n31439) );
  ANDN U30888 ( .B(n31442), .A(n31443), .Z(n31440) );
  XOR U30889 ( .A(n31444), .B(n31441), .Z(n31442) );
  IV U30890 ( .A(n31357), .Z(n31438) );
  XOR U30891 ( .A(n31445), .B(n31446), .Z(n31357) );
  ANDN U30892 ( .B(n31447), .A(n31448), .Z(n31445) );
  XOR U30893 ( .A(n31446), .B(n31449), .Z(n31447) );
  IV U30894 ( .A(n31371), .Z(n31424) );
  XOR U30895 ( .A(n31450), .B(n31451), .Z(n31371) );
  XNOR U30896 ( .A(n31366), .B(n31452), .Z(n31451) );
  IV U30897 ( .A(n31369), .Z(n31452) );
  XOR U30898 ( .A(n31453), .B(n31454), .Z(n31369) );
  ANDN U30899 ( .B(n31455), .A(n31456), .Z(n31453) );
  XOR U30900 ( .A(n31457), .B(n31454), .Z(n31455) );
  XNOR U30901 ( .A(n31458), .B(n31459), .Z(n31366) );
  ANDN U30902 ( .B(n31460), .A(n31461), .Z(n31458) );
  XOR U30903 ( .A(n31459), .B(n31462), .Z(n31460) );
  IV U30904 ( .A(n31365), .Z(n31450) );
  XOR U30905 ( .A(n31363), .B(n31463), .Z(n31365) );
  XOR U30906 ( .A(n31464), .B(n31465), .Z(n31463) );
  ANDN U30907 ( .B(n31466), .A(n31467), .Z(n31464) );
  XOR U30908 ( .A(n31468), .B(n31465), .Z(n31466) );
  IV U30909 ( .A(n31367), .Z(n31363) );
  XOR U30910 ( .A(n31469), .B(n31470), .Z(n31367) );
  ANDN U30911 ( .B(n31471), .A(n31472), .Z(n31469) );
  XOR U30912 ( .A(n31473), .B(n31470), .Z(n31471) );
  IV U30913 ( .A(n31377), .Z(n31381) );
  XOR U30914 ( .A(n31377), .B(n31280), .Z(n31379) );
  XOR U30915 ( .A(n31474), .B(n31475), .Z(n31280) );
  AND U30916 ( .A(n400), .B(n31476), .Z(n31474) );
  XOR U30917 ( .A(n31477), .B(n31475), .Z(n31476) );
  NANDN U30918 ( .A(n31282), .B(n31284), .Z(n31377) );
  XOR U30919 ( .A(n31478), .B(n31479), .Z(n31284) );
  AND U30920 ( .A(n400), .B(n31480), .Z(n31478) );
  XOR U30921 ( .A(n31479), .B(n31481), .Z(n31480) );
  XNOR U30922 ( .A(n31482), .B(n31483), .Z(n400) );
  AND U30923 ( .A(n31484), .B(n31485), .Z(n31482) );
  XOR U30924 ( .A(n31483), .B(n31295), .Z(n31485) );
  XNOR U30925 ( .A(n31486), .B(n31487), .Z(n31295) );
  ANDN U30926 ( .B(n31488), .A(n31489), .Z(n31486) );
  XOR U30927 ( .A(n31487), .B(n31490), .Z(n31488) );
  XNOR U30928 ( .A(n31483), .B(n31297), .Z(n31484) );
  XOR U30929 ( .A(n31491), .B(n31492), .Z(n31297) );
  AND U30930 ( .A(n404), .B(n31493), .Z(n31491) );
  XOR U30931 ( .A(n31494), .B(n31492), .Z(n31493) );
  XOR U30932 ( .A(n31495), .B(n31496), .Z(n31483) );
  AND U30933 ( .A(n31497), .B(n31498), .Z(n31495) );
  XOR U30934 ( .A(n31496), .B(n31322), .Z(n31498) );
  XOR U30935 ( .A(n31489), .B(n31490), .Z(n31322) );
  XNOR U30936 ( .A(n31499), .B(n31500), .Z(n31490) );
  ANDN U30937 ( .B(n31501), .A(n31502), .Z(n31499) );
  XOR U30938 ( .A(n31503), .B(n31504), .Z(n31501) );
  XOR U30939 ( .A(n31505), .B(n31506), .Z(n31489) );
  XNOR U30940 ( .A(n31507), .B(n31508), .Z(n31506) );
  ANDN U30941 ( .B(n31509), .A(n31510), .Z(n31507) );
  XNOR U30942 ( .A(n31511), .B(n31512), .Z(n31509) );
  IV U30943 ( .A(n31487), .Z(n31505) );
  XOR U30944 ( .A(n31513), .B(n31514), .Z(n31487) );
  ANDN U30945 ( .B(n31515), .A(n31516), .Z(n31513) );
  XOR U30946 ( .A(n31514), .B(n31517), .Z(n31515) );
  XNOR U30947 ( .A(n31496), .B(n31324), .Z(n31497) );
  XOR U30948 ( .A(n31518), .B(n31519), .Z(n31324) );
  AND U30949 ( .A(n404), .B(n31520), .Z(n31518) );
  XOR U30950 ( .A(n31521), .B(n31519), .Z(n31520) );
  XNOR U30951 ( .A(n31522), .B(n31523), .Z(n31496) );
  AND U30952 ( .A(n31524), .B(n31525), .Z(n31522) );
  XNOR U30953 ( .A(n31523), .B(n31374), .Z(n31525) );
  XOR U30954 ( .A(n31516), .B(n31517), .Z(n31374) );
  XOR U30955 ( .A(n31526), .B(n31504), .Z(n31517) );
  XNOR U30956 ( .A(n31527), .B(n31528), .Z(n31504) );
  ANDN U30957 ( .B(n31529), .A(n31530), .Z(n31527) );
  XOR U30958 ( .A(n31531), .B(n31532), .Z(n31529) );
  IV U30959 ( .A(n31502), .Z(n31526) );
  XOR U30960 ( .A(n31500), .B(n31533), .Z(n31502) );
  XNOR U30961 ( .A(n31534), .B(n31535), .Z(n31533) );
  ANDN U30962 ( .B(n31536), .A(n31537), .Z(n31534) );
  XNOR U30963 ( .A(n31538), .B(n31539), .Z(n31536) );
  IV U30964 ( .A(n31503), .Z(n31500) );
  XOR U30965 ( .A(n31540), .B(n31541), .Z(n31503) );
  ANDN U30966 ( .B(n31542), .A(n31543), .Z(n31540) );
  XOR U30967 ( .A(n31541), .B(n31544), .Z(n31542) );
  XOR U30968 ( .A(n31545), .B(n31546), .Z(n31516) );
  XNOR U30969 ( .A(n31511), .B(n31547), .Z(n31546) );
  IV U30970 ( .A(n31514), .Z(n31547) );
  XOR U30971 ( .A(n31548), .B(n31549), .Z(n31514) );
  ANDN U30972 ( .B(n31550), .A(n31551), .Z(n31548) );
  XOR U30973 ( .A(n31549), .B(n31552), .Z(n31550) );
  XNOR U30974 ( .A(n31553), .B(n31554), .Z(n31511) );
  ANDN U30975 ( .B(n31555), .A(n31556), .Z(n31553) );
  XOR U30976 ( .A(n31554), .B(n31557), .Z(n31555) );
  IV U30977 ( .A(n31510), .Z(n31545) );
  XOR U30978 ( .A(n31508), .B(n31558), .Z(n31510) );
  XNOR U30979 ( .A(n31559), .B(n31560), .Z(n31558) );
  ANDN U30980 ( .B(n31561), .A(n31562), .Z(n31559) );
  XNOR U30981 ( .A(n31563), .B(n31564), .Z(n31561) );
  IV U30982 ( .A(n31512), .Z(n31508) );
  XOR U30983 ( .A(n31565), .B(n31566), .Z(n31512) );
  ANDN U30984 ( .B(n31567), .A(n31568), .Z(n31565) );
  XOR U30985 ( .A(n31569), .B(n31566), .Z(n31567) );
  XOR U30986 ( .A(n31523), .B(n31376), .Z(n31524) );
  XOR U30987 ( .A(n31570), .B(n31571), .Z(n31376) );
  AND U30988 ( .A(n404), .B(n31572), .Z(n31570) );
  XOR U30989 ( .A(n31573), .B(n31571), .Z(n31572) );
  XNOR U30990 ( .A(n31574), .B(n31575), .Z(n31523) );
  NAND U30991 ( .A(n31576), .B(n31577), .Z(n31575) );
  XOR U30992 ( .A(n31578), .B(n31475), .Z(n31577) );
  XOR U30993 ( .A(n31551), .B(n31552), .Z(n31475) );
  XOR U30994 ( .A(n31579), .B(n31544), .Z(n31552) );
  XOR U30995 ( .A(n31580), .B(n31532), .Z(n31544) );
  XOR U30996 ( .A(n31581), .B(n31582), .Z(n31532) );
  ANDN U30997 ( .B(n31583), .A(n31584), .Z(n31581) );
  XOR U30998 ( .A(n31582), .B(n31585), .Z(n31583) );
  IV U30999 ( .A(n31530), .Z(n31580) );
  XOR U31000 ( .A(n31528), .B(n31586), .Z(n31530) );
  XOR U31001 ( .A(n31587), .B(n31588), .Z(n31586) );
  ANDN U31002 ( .B(n31589), .A(n31590), .Z(n31587) );
  XOR U31003 ( .A(n31591), .B(n31588), .Z(n31589) );
  IV U31004 ( .A(n31531), .Z(n31528) );
  XOR U31005 ( .A(n31592), .B(n31593), .Z(n31531) );
  ANDN U31006 ( .B(n31594), .A(n31595), .Z(n31592) );
  XOR U31007 ( .A(n31593), .B(n31596), .Z(n31594) );
  IV U31008 ( .A(n31543), .Z(n31579) );
  XOR U31009 ( .A(n31597), .B(n31598), .Z(n31543) );
  XNOR U31010 ( .A(n31538), .B(n31599), .Z(n31598) );
  IV U31011 ( .A(n31541), .Z(n31599) );
  XOR U31012 ( .A(n31600), .B(n31601), .Z(n31541) );
  ANDN U31013 ( .B(n31602), .A(n31603), .Z(n31600) );
  XOR U31014 ( .A(n31601), .B(n31604), .Z(n31602) );
  XNOR U31015 ( .A(n31605), .B(n31606), .Z(n31538) );
  ANDN U31016 ( .B(n31607), .A(n31608), .Z(n31605) );
  XOR U31017 ( .A(n31606), .B(n31609), .Z(n31607) );
  IV U31018 ( .A(n31537), .Z(n31597) );
  XOR U31019 ( .A(n31535), .B(n31610), .Z(n31537) );
  XOR U31020 ( .A(n31611), .B(n31612), .Z(n31610) );
  ANDN U31021 ( .B(n31613), .A(n31614), .Z(n31611) );
  XOR U31022 ( .A(n31615), .B(n31612), .Z(n31613) );
  IV U31023 ( .A(n31539), .Z(n31535) );
  XOR U31024 ( .A(n31616), .B(n31617), .Z(n31539) );
  ANDN U31025 ( .B(n31618), .A(n31619), .Z(n31616) );
  XOR U31026 ( .A(n31620), .B(n31617), .Z(n31618) );
  XOR U31027 ( .A(n31621), .B(n31622), .Z(n31551) );
  XOR U31028 ( .A(n31569), .B(n31623), .Z(n31622) );
  IV U31029 ( .A(n31549), .Z(n31623) );
  XOR U31030 ( .A(n31624), .B(n31625), .Z(n31549) );
  ANDN U31031 ( .B(n31626), .A(n31627), .Z(n31624) );
  XOR U31032 ( .A(n31625), .B(n31628), .Z(n31626) );
  XOR U31033 ( .A(n31629), .B(n31557), .Z(n31569) );
  XOR U31034 ( .A(n31630), .B(n31631), .Z(n31557) );
  ANDN U31035 ( .B(n31632), .A(n31633), .Z(n31630) );
  XOR U31036 ( .A(n31631), .B(n31634), .Z(n31632) );
  IV U31037 ( .A(n31556), .Z(n31629) );
  XOR U31038 ( .A(n31635), .B(n31636), .Z(n31556) );
  XOR U31039 ( .A(n31637), .B(n31638), .Z(n31636) );
  ANDN U31040 ( .B(n31639), .A(n31640), .Z(n31637) );
  XOR U31041 ( .A(n31641), .B(n31638), .Z(n31639) );
  IV U31042 ( .A(n31554), .Z(n31635) );
  XOR U31043 ( .A(n31642), .B(n31643), .Z(n31554) );
  ANDN U31044 ( .B(n31644), .A(n31645), .Z(n31642) );
  XOR U31045 ( .A(n31643), .B(n31646), .Z(n31644) );
  IV U31046 ( .A(n31568), .Z(n31621) );
  XOR U31047 ( .A(n31647), .B(n31648), .Z(n31568) );
  XNOR U31048 ( .A(n31563), .B(n31649), .Z(n31648) );
  IV U31049 ( .A(n31566), .Z(n31649) );
  XOR U31050 ( .A(n31650), .B(n31651), .Z(n31566) );
  ANDN U31051 ( .B(n31652), .A(n31653), .Z(n31650) );
  XOR U31052 ( .A(n31654), .B(n31651), .Z(n31652) );
  XNOR U31053 ( .A(n31655), .B(n31656), .Z(n31563) );
  ANDN U31054 ( .B(n31657), .A(n31658), .Z(n31655) );
  XOR U31055 ( .A(n31656), .B(n31659), .Z(n31657) );
  IV U31056 ( .A(n31562), .Z(n31647) );
  XOR U31057 ( .A(n31560), .B(n31660), .Z(n31562) );
  XOR U31058 ( .A(n31661), .B(n31662), .Z(n31660) );
  ANDN U31059 ( .B(n31663), .A(n31664), .Z(n31661) );
  XOR U31060 ( .A(n31665), .B(n31662), .Z(n31663) );
  IV U31061 ( .A(n31564), .Z(n31560) );
  XOR U31062 ( .A(n31666), .B(n31667), .Z(n31564) );
  ANDN U31063 ( .B(n31668), .A(n31669), .Z(n31666) );
  XOR U31064 ( .A(n31670), .B(n31667), .Z(n31668) );
  IV U31065 ( .A(n31574), .Z(n31578) );
  XOR U31066 ( .A(n31574), .B(n31477), .Z(n31576) );
  XOR U31067 ( .A(n31671), .B(n31672), .Z(n31477) );
  AND U31068 ( .A(n404), .B(n31673), .Z(n31671) );
  XOR U31069 ( .A(n31674), .B(n31672), .Z(n31673) );
  NANDN U31070 ( .A(n31479), .B(n31481), .Z(n31574) );
  XOR U31071 ( .A(n31675), .B(n31676), .Z(n31481) );
  AND U31072 ( .A(n404), .B(n31677), .Z(n31675) );
  XOR U31073 ( .A(n31676), .B(n31678), .Z(n31677) );
  XNOR U31074 ( .A(n31679), .B(n31680), .Z(n404) );
  AND U31075 ( .A(n31681), .B(n31682), .Z(n31679) );
  XOR U31076 ( .A(n31680), .B(n31492), .Z(n31682) );
  XNOR U31077 ( .A(n31683), .B(n31684), .Z(n31492) );
  ANDN U31078 ( .B(n31685), .A(n31686), .Z(n31683) );
  XOR U31079 ( .A(n31684), .B(n31687), .Z(n31685) );
  XNOR U31080 ( .A(n31680), .B(n31494), .Z(n31681) );
  XOR U31081 ( .A(n31688), .B(n31689), .Z(n31494) );
  AND U31082 ( .A(n408), .B(n31690), .Z(n31688) );
  XOR U31083 ( .A(n31691), .B(n31689), .Z(n31690) );
  XOR U31084 ( .A(n31692), .B(n31693), .Z(n31680) );
  AND U31085 ( .A(n31694), .B(n31695), .Z(n31692) );
  XOR U31086 ( .A(n31693), .B(n31519), .Z(n31695) );
  XOR U31087 ( .A(n31686), .B(n31687), .Z(n31519) );
  XNOR U31088 ( .A(n31696), .B(n31697), .Z(n31687) );
  ANDN U31089 ( .B(n31698), .A(n31699), .Z(n31696) );
  XOR U31090 ( .A(n31700), .B(n31701), .Z(n31698) );
  XOR U31091 ( .A(n31702), .B(n31703), .Z(n31686) );
  XNOR U31092 ( .A(n31704), .B(n31705), .Z(n31703) );
  ANDN U31093 ( .B(n31706), .A(n31707), .Z(n31704) );
  XNOR U31094 ( .A(n31708), .B(n31709), .Z(n31706) );
  IV U31095 ( .A(n31684), .Z(n31702) );
  XOR U31096 ( .A(n31710), .B(n31711), .Z(n31684) );
  ANDN U31097 ( .B(n31712), .A(n31713), .Z(n31710) );
  XOR U31098 ( .A(n31711), .B(n31714), .Z(n31712) );
  XNOR U31099 ( .A(n31693), .B(n31521), .Z(n31694) );
  XOR U31100 ( .A(n31715), .B(n31716), .Z(n31521) );
  AND U31101 ( .A(n408), .B(n31717), .Z(n31715) );
  XOR U31102 ( .A(n31718), .B(n31716), .Z(n31717) );
  XNOR U31103 ( .A(n31719), .B(n31720), .Z(n31693) );
  AND U31104 ( .A(n31721), .B(n31722), .Z(n31719) );
  XNOR U31105 ( .A(n31720), .B(n31571), .Z(n31722) );
  XOR U31106 ( .A(n31713), .B(n31714), .Z(n31571) );
  XOR U31107 ( .A(n31723), .B(n31701), .Z(n31714) );
  XNOR U31108 ( .A(n31724), .B(n31725), .Z(n31701) );
  ANDN U31109 ( .B(n31726), .A(n31727), .Z(n31724) );
  XOR U31110 ( .A(n31728), .B(n31729), .Z(n31726) );
  IV U31111 ( .A(n31699), .Z(n31723) );
  XOR U31112 ( .A(n31697), .B(n31730), .Z(n31699) );
  XNOR U31113 ( .A(n31731), .B(n31732), .Z(n31730) );
  ANDN U31114 ( .B(n31733), .A(n31734), .Z(n31731) );
  XNOR U31115 ( .A(n31735), .B(n31736), .Z(n31733) );
  IV U31116 ( .A(n31700), .Z(n31697) );
  XOR U31117 ( .A(n31737), .B(n31738), .Z(n31700) );
  ANDN U31118 ( .B(n31739), .A(n31740), .Z(n31737) );
  XOR U31119 ( .A(n31738), .B(n31741), .Z(n31739) );
  XOR U31120 ( .A(n31742), .B(n31743), .Z(n31713) );
  XNOR U31121 ( .A(n31708), .B(n31744), .Z(n31743) );
  IV U31122 ( .A(n31711), .Z(n31744) );
  XOR U31123 ( .A(n31745), .B(n31746), .Z(n31711) );
  ANDN U31124 ( .B(n31747), .A(n31748), .Z(n31745) );
  XOR U31125 ( .A(n31746), .B(n31749), .Z(n31747) );
  XNOR U31126 ( .A(n31750), .B(n31751), .Z(n31708) );
  ANDN U31127 ( .B(n31752), .A(n31753), .Z(n31750) );
  XOR U31128 ( .A(n31751), .B(n31754), .Z(n31752) );
  IV U31129 ( .A(n31707), .Z(n31742) );
  XOR U31130 ( .A(n31705), .B(n31755), .Z(n31707) );
  XNOR U31131 ( .A(n31756), .B(n31757), .Z(n31755) );
  ANDN U31132 ( .B(n31758), .A(n31759), .Z(n31756) );
  XNOR U31133 ( .A(n31760), .B(n31761), .Z(n31758) );
  IV U31134 ( .A(n31709), .Z(n31705) );
  XOR U31135 ( .A(n31762), .B(n31763), .Z(n31709) );
  ANDN U31136 ( .B(n31764), .A(n31765), .Z(n31762) );
  XOR U31137 ( .A(n31766), .B(n31763), .Z(n31764) );
  XOR U31138 ( .A(n31720), .B(n31573), .Z(n31721) );
  XOR U31139 ( .A(n31767), .B(n31768), .Z(n31573) );
  AND U31140 ( .A(n408), .B(n31769), .Z(n31767) );
  XOR U31141 ( .A(n31770), .B(n31768), .Z(n31769) );
  XNOR U31142 ( .A(n31771), .B(n31772), .Z(n31720) );
  NAND U31143 ( .A(n31773), .B(n31774), .Z(n31772) );
  XOR U31144 ( .A(n31775), .B(n31672), .Z(n31774) );
  XOR U31145 ( .A(n31748), .B(n31749), .Z(n31672) );
  XOR U31146 ( .A(n31776), .B(n31741), .Z(n31749) );
  XOR U31147 ( .A(n31777), .B(n31729), .Z(n31741) );
  XOR U31148 ( .A(n31778), .B(n31779), .Z(n31729) );
  ANDN U31149 ( .B(n31780), .A(n31781), .Z(n31778) );
  XOR U31150 ( .A(n31779), .B(n31782), .Z(n31780) );
  IV U31151 ( .A(n31727), .Z(n31777) );
  XOR U31152 ( .A(n31725), .B(n31783), .Z(n31727) );
  XOR U31153 ( .A(n31784), .B(n31785), .Z(n31783) );
  ANDN U31154 ( .B(n31786), .A(n31787), .Z(n31784) );
  XOR U31155 ( .A(n31788), .B(n31785), .Z(n31786) );
  IV U31156 ( .A(n31728), .Z(n31725) );
  XOR U31157 ( .A(n31789), .B(n31790), .Z(n31728) );
  ANDN U31158 ( .B(n31791), .A(n31792), .Z(n31789) );
  XOR U31159 ( .A(n31790), .B(n31793), .Z(n31791) );
  IV U31160 ( .A(n31740), .Z(n31776) );
  XOR U31161 ( .A(n31794), .B(n31795), .Z(n31740) );
  XNOR U31162 ( .A(n31735), .B(n31796), .Z(n31795) );
  IV U31163 ( .A(n31738), .Z(n31796) );
  XOR U31164 ( .A(n31797), .B(n31798), .Z(n31738) );
  ANDN U31165 ( .B(n31799), .A(n31800), .Z(n31797) );
  XOR U31166 ( .A(n31798), .B(n31801), .Z(n31799) );
  XNOR U31167 ( .A(n31802), .B(n31803), .Z(n31735) );
  ANDN U31168 ( .B(n31804), .A(n31805), .Z(n31802) );
  XOR U31169 ( .A(n31803), .B(n31806), .Z(n31804) );
  IV U31170 ( .A(n31734), .Z(n31794) );
  XOR U31171 ( .A(n31732), .B(n31807), .Z(n31734) );
  XOR U31172 ( .A(n31808), .B(n31809), .Z(n31807) );
  ANDN U31173 ( .B(n31810), .A(n31811), .Z(n31808) );
  XOR U31174 ( .A(n31812), .B(n31809), .Z(n31810) );
  IV U31175 ( .A(n31736), .Z(n31732) );
  XOR U31176 ( .A(n31813), .B(n31814), .Z(n31736) );
  ANDN U31177 ( .B(n31815), .A(n31816), .Z(n31813) );
  XOR U31178 ( .A(n31817), .B(n31814), .Z(n31815) );
  XOR U31179 ( .A(n31818), .B(n31819), .Z(n31748) );
  XOR U31180 ( .A(n31766), .B(n31820), .Z(n31819) );
  IV U31181 ( .A(n31746), .Z(n31820) );
  XOR U31182 ( .A(n31821), .B(n31822), .Z(n31746) );
  ANDN U31183 ( .B(n31823), .A(n31824), .Z(n31821) );
  XOR U31184 ( .A(n31822), .B(n31825), .Z(n31823) );
  XOR U31185 ( .A(n31826), .B(n31754), .Z(n31766) );
  XOR U31186 ( .A(n31827), .B(n31828), .Z(n31754) );
  ANDN U31187 ( .B(n31829), .A(n31830), .Z(n31827) );
  XOR U31188 ( .A(n31828), .B(n31831), .Z(n31829) );
  IV U31189 ( .A(n31753), .Z(n31826) );
  XOR U31190 ( .A(n31832), .B(n31833), .Z(n31753) );
  XOR U31191 ( .A(n31834), .B(n31835), .Z(n31833) );
  ANDN U31192 ( .B(n31836), .A(n31837), .Z(n31834) );
  XOR U31193 ( .A(n31838), .B(n31835), .Z(n31836) );
  IV U31194 ( .A(n31751), .Z(n31832) );
  XOR U31195 ( .A(n31839), .B(n31840), .Z(n31751) );
  ANDN U31196 ( .B(n31841), .A(n31842), .Z(n31839) );
  XOR U31197 ( .A(n31840), .B(n31843), .Z(n31841) );
  IV U31198 ( .A(n31765), .Z(n31818) );
  XOR U31199 ( .A(n31844), .B(n31845), .Z(n31765) );
  XNOR U31200 ( .A(n31760), .B(n31846), .Z(n31845) );
  IV U31201 ( .A(n31763), .Z(n31846) );
  XOR U31202 ( .A(n31847), .B(n31848), .Z(n31763) );
  ANDN U31203 ( .B(n31849), .A(n31850), .Z(n31847) );
  XOR U31204 ( .A(n31851), .B(n31848), .Z(n31849) );
  XNOR U31205 ( .A(n31852), .B(n31853), .Z(n31760) );
  ANDN U31206 ( .B(n31854), .A(n31855), .Z(n31852) );
  XOR U31207 ( .A(n31853), .B(n31856), .Z(n31854) );
  IV U31208 ( .A(n31759), .Z(n31844) );
  XOR U31209 ( .A(n31757), .B(n31857), .Z(n31759) );
  XOR U31210 ( .A(n31858), .B(n31859), .Z(n31857) );
  ANDN U31211 ( .B(n31860), .A(n31861), .Z(n31858) );
  XOR U31212 ( .A(n31862), .B(n31859), .Z(n31860) );
  IV U31213 ( .A(n31761), .Z(n31757) );
  XOR U31214 ( .A(n31863), .B(n31864), .Z(n31761) );
  ANDN U31215 ( .B(n31865), .A(n31866), .Z(n31863) );
  XOR U31216 ( .A(n31867), .B(n31864), .Z(n31865) );
  IV U31217 ( .A(n31771), .Z(n31775) );
  XOR U31218 ( .A(n31771), .B(n31674), .Z(n31773) );
  XOR U31219 ( .A(n31868), .B(n31869), .Z(n31674) );
  AND U31220 ( .A(n408), .B(n31870), .Z(n31868) );
  XOR U31221 ( .A(n31871), .B(n31869), .Z(n31870) );
  NANDN U31222 ( .A(n31676), .B(n31678), .Z(n31771) );
  XOR U31223 ( .A(n31872), .B(n31873), .Z(n31678) );
  AND U31224 ( .A(n408), .B(n31874), .Z(n31872) );
  XOR U31225 ( .A(n31873), .B(n31875), .Z(n31874) );
  XNOR U31226 ( .A(n31876), .B(n31877), .Z(n408) );
  AND U31227 ( .A(n31878), .B(n31879), .Z(n31876) );
  XOR U31228 ( .A(n31877), .B(n31689), .Z(n31879) );
  XNOR U31229 ( .A(n31880), .B(n31881), .Z(n31689) );
  ANDN U31230 ( .B(n31882), .A(n31883), .Z(n31880) );
  XOR U31231 ( .A(n31881), .B(n31884), .Z(n31882) );
  XNOR U31232 ( .A(n31877), .B(n31691), .Z(n31878) );
  XOR U31233 ( .A(n31885), .B(n31886), .Z(n31691) );
  AND U31234 ( .A(n412), .B(n31887), .Z(n31885) );
  XOR U31235 ( .A(n31888), .B(n31886), .Z(n31887) );
  XOR U31236 ( .A(n31889), .B(n31890), .Z(n31877) );
  AND U31237 ( .A(n31891), .B(n31892), .Z(n31889) );
  XOR U31238 ( .A(n31890), .B(n31716), .Z(n31892) );
  XOR U31239 ( .A(n31883), .B(n31884), .Z(n31716) );
  XNOR U31240 ( .A(n31893), .B(n31894), .Z(n31884) );
  ANDN U31241 ( .B(n31895), .A(n31896), .Z(n31893) );
  XOR U31242 ( .A(n31897), .B(n31898), .Z(n31895) );
  XOR U31243 ( .A(n31899), .B(n31900), .Z(n31883) );
  XNOR U31244 ( .A(n31901), .B(n31902), .Z(n31900) );
  ANDN U31245 ( .B(n31903), .A(n31904), .Z(n31901) );
  XNOR U31246 ( .A(n31905), .B(n31906), .Z(n31903) );
  IV U31247 ( .A(n31881), .Z(n31899) );
  XOR U31248 ( .A(n31907), .B(n31908), .Z(n31881) );
  ANDN U31249 ( .B(n31909), .A(n31910), .Z(n31907) );
  XOR U31250 ( .A(n31908), .B(n31911), .Z(n31909) );
  XNOR U31251 ( .A(n31890), .B(n31718), .Z(n31891) );
  XOR U31252 ( .A(n31912), .B(n31913), .Z(n31718) );
  AND U31253 ( .A(n412), .B(n31914), .Z(n31912) );
  XOR U31254 ( .A(n31915), .B(n31913), .Z(n31914) );
  XNOR U31255 ( .A(n31916), .B(n31917), .Z(n31890) );
  AND U31256 ( .A(n31918), .B(n31919), .Z(n31916) );
  XNOR U31257 ( .A(n31917), .B(n31768), .Z(n31919) );
  XOR U31258 ( .A(n31910), .B(n31911), .Z(n31768) );
  XOR U31259 ( .A(n31920), .B(n31898), .Z(n31911) );
  XNOR U31260 ( .A(n31921), .B(n31922), .Z(n31898) );
  ANDN U31261 ( .B(n31923), .A(n31924), .Z(n31921) );
  XOR U31262 ( .A(n31925), .B(n31926), .Z(n31923) );
  IV U31263 ( .A(n31896), .Z(n31920) );
  XOR U31264 ( .A(n31894), .B(n31927), .Z(n31896) );
  XNOR U31265 ( .A(n31928), .B(n31929), .Z(n31927) );
  ANDN U31266 ( .B(n31930), .A(n31931), .Z(n31928) );
  XNOR U31267 ( .A(n31932), .B(n31933), .Z(n31930) );
  IV U31268 ( .A(n31897), .Z(n31894) );
  XOR U31269 ( .A(n31934), .B(n31935), .Z(n31897) );
  ANDN U31270 ( .B(n31936), .A(n31937), .Z(n31934) );
  XOR U31271 ( .A(n31935), .B(n31938), .Z(n31936) );
  XOR U31272 ( .A(n31939), .B(n31940), .Z(n31910) );
  XNOR U31273 ( .A(n31905), .B(n31941), .Z(n31940) );
  IV U31274 ( .A(n31908), .Z(n31941) );
  XOR U31275 ( .A(n31942), .B(n31943), .Z(n31908) );
  ANDN U31276 ( .B(n31944), .A(n31945), .Z(n31942) );
  XOR U31277 ( .A(n31943), .B(n31946), .Z(n31944) );
  XNOR U31278 ( .A(n31947), .B(n31948), .Z(n31905) );
  ANDN U31279 ( .B(n31949), .A(n31950), .Z(n31947) );
  XOR U31280 ( .A(n31948), .B(n31951), .Z(n31949) );
  IV U31281 ( .A(n31904), .Z(n31939) );
  XOR U31282 ( .A(n31902), .B(n31952), .Z(n31904) );
  XNOR U31283 ( .A(n31953), .B(n31954), .Z(n31952) );
  ANDN U31284 ( .B(n31955), .A(n31956), .Z(n31953) );
  XNOR U31285 ( .A(n31957), .B(n31958), .Z(n31955) );
  IV U31286 ( .A(n31906), .Z(n31902) );
  XOR U31287 ( .A(n31959), .B(n31960), .Z(n31906) );
  ANDN U31288 ( .B(n31961), .A(n31962), .Z(n31959) );
  XOR U31289 ( .A(n31963), .B(n31960), .Z(n31961) );
  XOR U31290 ( .A(n31917), .B(n31770), .Z(n31918) );
  XOR U31291 ( .A(n31964), .B(n31965), .Z(n31770) );
  AND U31292 ( .A(n412), .B(n31966), .Z(n31964) );
  XOR U31293 ( .A(n31967), .B(n31965), .Z(n31966) );
  XNOR U31294 ( .A(n31968), .B(n31969), .Z(n31917) );
  NAND U31295 ( .A(n31970), .B(n31971), .Z(n31969) );
  XOR U31296 ( .A(n31972), .B(n31869), .Z(n31971) );
  XOR U31297 ( .A(n31945), .B(n31946), .Z(n31869) );
  XOR U31298 ( .A(n31973), .B(n31938), .Z(n31946) );
  XOR U31299 ( .A(n31974), .B(n31926), .Z(n31938) );
  XOR U31300 ( .A(n31975), .B(n31976), .Z(n31926) );
  ANDN U31301 ( .B(n31977), .A(n31978), .Z(n31975) );
  XOR U31302 ( .A(n31976), .B(n31979), .Z(n31977) );
  IV U31303 ( .A(n31924), .Z(n31974) );
  XOR U31304 ( .A(n31922), .B(n31980), .Z(n31924) );
  XOR U31305 ( .A(n31981), .B(n31982), .Z(n31980) );
  ANDN U31306 ( .B(n31983), .A(n31984), .Z(n31981) );
  XOR U31307 ( .A(n31985), .B(n31982), .Z(n31983) );
  IV U31308 ( .A(n31925), .Z(n31922) );
  XOR U31309 ( .A(n31986), .B(n31987), .Z(n31925) );
  ANDN U31310 ( .B(n31988), .A(n31989), .Z(n31986) );
  XOR U31311 ( .A(n31987), .B(n31990), .Z(n31988) );
  IV U31312 ( .A(n31937), .Z(n31973) );
  XOR U31313 ( .A(n31991), .B(n31992), .Z(n31937) );
  XNOR U31314 ( .A(n31932), .B(n31993), .Z(n31992) );
  IV U31315 ( .A(n31935), .Z(n31993) );
  XOR U31316 ( .A(n31994), .B(n31995), .Z(n31935) );
  ANDN U31317 ( .B(n31996), .A(n31997), .Z(n31994) );
  XOR U31318 ( .A(n31995), .B(n31998), .Z(n31996) );
  XNOR U31319 ( .A(n31999), .B(n32000), .Z(n31932) );
  ANDN U31320 ( .B(n32001), .A(n32002), .Z(n31999) );
  XOR U31321 ( .A(n32000), .B(n32003), .Z(n32001) );
  IV U31322 ( .A(n31931), .Z(n31991) );
  XOR U31323 ( .A(n31929), .B(n32004), .Z(n31931) );
  XOR U31324 ( .A(n32005), .B(n32006), .Z(n32004) );
  ANDN U31325 ( .B(n32007), .A(n32008), .Z(n32005) );
  XOR U31326 ( .A(n32009), .B(n32006), .Z(n32007) );
  IV U31327 ( .A(n31933), .Z(n31929) );
  XOR U31328 ( .A(n32010), .B(n32011), .Z(n31933) );
  ANDN U31329 ( .B(n32012), .A(n32013), .Z(n32010) );
  XOR U31330 ( .A(n32014), .B(n32011), .Z(n32012) );
  XOR U31331 ( .A(n32015), .B(n32016), .Z(n31945) );
  XOR U31332 ( .A(n31963), .B(n32017), .Z(n32016) );
  IV U31333 ( .A(n31943), .Z(n32017) );
  XOR U31334 ( .A(n32018), .B(n32019), .Z(n31943) );
  ANDN U31335 ( .B(n32020), .A(n32021), .Z(n32018) );
  XOR U31336 ( .A(n32019), .B(n32022), .Z(n32020) );
  XOR U31337 ( .A(n32023), .B(n31951), .Z(n31963) );
  XOR U31338 ( .A(n32024), .B(n32025), .Z(n31951) );
  ANDN U31339 ( .B(n32026), .A(n32027), .Z(n32024) );
  XOR U31340 ( .A(n32025), .B(n32028), .Z(n32026) );
  IV U31341 ( .A(n31950), .Z(n32023) );
  XOR U31342 ( .A(n32029), .B(n32030), .Z(n31950) );
  XOR U31343 ( .A(n32031), .B(n32032), .Z(n32030) );
  ANDN U31344 ( .B(n32033), .A(n32034), .Z(n32031) );
  XOR U31345 ( .A(n32035), .B(n32032), .Z(n32033) );
  IV U31346 ( .A(n31948), .Z(n32029) );
  XOR U31347 ( .A(n32036), .B(n32037), .Z(n31948) );
  ANDN U31348 ( .B(n32038), .A(n32039), .Z(n32036) );
  XOR U31349 ( .A(n32037), .B(n32040), .Z(n32038) );
  IV U31350 ( .A(n31962), .Z(n32015) );
  XOR U31351 ( .A(n32041), .B(n32042), .Z(n31962) );
  XNOR U31352 ( .A(n31957), .B(n32043), .Z(n32042) );
  IV U31353 ( .A(n31960), .Z(n32043) );
  XOR U31354 ( .A(n32044), .B(n32045), .Z(n31960) );
  ANDN U31355 ( .B(n32046), .A(n32047), .Z(n32044) );
  XOR U31356 ( .A(n32048), .B(n32045), .Z(n32046) );
  XNOR U31357 ( .A(n32049), .B(n32050), .Z(n31957) );
  ANDN U31358 ( .B(n32051), .A(n32052), .Z(n32049) );
  XOR U31359 ( .A(n32050), .B(n32053), .Z(n32051) );
  IV U31360 ( .A(n31956), .Z(n32041) );
  XOR U31361 ( .A(n31954), .B(n32054), .Z(n31956) );
  XOR U31362 ( .A(n32055), .B(n32056), .Z(n32054) );
  ANDN U31363 ( .B(n32057), .A(n32058), .Z(n32055) );
  XOR U31364 ( .A(n32059), .B(n32056), .Z(n32057) );
  IV U31365 ( .A(n31958), .Z(n31954) );
  XOR U31366 ( .A(n32060), .B(n32061), .Z(n31958) );
  ANDN U31367 ( .B(n32062), .A(n32063), .Z(n32060) );
  XOR U31368 ( .A(n32064), .B(n32061), .Z(n32062) );
  IV U31369 ( .A(n31968), .Z(n31972) );
  XOR U31370 ( .A(n31968), .B(n31871), .Z(n31970) );
  XOR U31371 ( .A(n32065), .B(n32066), .Z(n31871) );
  AND U31372 ( .A(n412), .B(n32067), .Z(n32065) );
  XOR U31373 ( .A(n32068), .B(n32066), .Z(n32067) );
  NANDN U31374 ( .A(n31873), .B(n31875), .Z(n31968) );
  XOR U31375 ( .A(n32069), .B(n32070), .Z(n31875) );
  AND U31376 ( .A(n412), .B(n32071), .Z(n32069) );
  XOR U31377 ( .A(n32070), .B(n32072), .Z(n32071) );
  XNOR U31378 ( .A(n32073), .B(n32074), .Z(n412) );
  AND U31379 ( .A(n32075), .B(n32076), .Z(n32073) );
  XOR U31380 ( .A(n32074), .B(n31886), .Z(n32076) );
  XNOR U31381 ( .A(n32077), .B(n32078), .Z(n31886) );
  ANDN U31382 ( .B(n32079), .A(n32080), .Z(n32077) );
  XOR U31383 ( .A(n32078), .B(n32081), .Z(n32079) );
  XNOR U31384 ( .A(n32074), .B(n31888), .Z(n32075) );
  XOR U31385 ( .A(n32082), .B(n32083), .Z(n31888) );
  AND U31386 ( .A(n416), .B(n32084), .Z(n32082) );
  XOR U31387 ( .A(n32085), .B(n32083), .Z(n32084) );
  XOR U31388 ( .A(n32086), .B(n32087), .Z(n32074) );
  AND U31389 ( .A(n32088), .B(n32089), .Z(n32086) );
  XOR U31390 ( .A(n32087), .B(n31913), .Z(n32089) );
  XOR U31391 ( .A(n32080), .B(n32081), .Z(n31913) );
  XNOR U31392 ( .A(n32090), .B(n32091), .Z(n32081) );
  ANDN U31393 ( .B(n32092), .A(n32093), .Z(n32090) );
  XOR U31394 ( .A(n32094), .B(n32095), .Z(n32092) );
  XOR U31395 ( .A(n32096), .B(n32097), .Z(n32080) );
  XNOR U31396 ( .A(n32098), .B(n32099), .Z(n32097) );
  ANDN U31397 ( .B(n32100), .A(n32101), .Z(n32098) );
  XNOR U31398 ( .A(n32102), .B(n32103), .Z(n32100) );
  IV U31399 ( .A(n32078), .Z(n32096) );
  XOR U31400 ( .A(n32104), .B(n32105), .Z(n32078) );
  ANDN U31401 ( .B(n32106), .A(n32107), .Z(n32104) );
  XOR U31402 ( .A(n32105), .B(n32108), .Z(n32106) );
  XNOR U31403 ( .A(n32087), .B(n31915), .Z(n32088) );
  XOR U31404 ( .A(n32109), .B(n32110), .Z(n31915) );
  AND U31405 ( .A(n416), .B(n32111), .Z(n32109) );
  XOR U31406 ( .A(n32112), .B(n32110), .Z(n32111) );
  XNOR U31407 ( .A(n32113), .B(n32114), .Z(n32087) );
  AND U31408 ( .A(n32115), .B(n32116), .Z(n32113) );
  XNOR U31409 ( .A(n32114), .B(n31965), .Z(n32116) );
  XOR U31410 ( .A(n32107), .B(n32108), .Z(n31965) );
  XOR U31411 ( .A(n32117), .B(n32095), .Z(n32108) );
  XNOR U31412 ( .A(n32118), .B(n32119), .Z(n32095) );
  ANDN U31413 ( .B(n32120), .A(n32121), .Z(n32118) );
  XOR U31414 ( .A(n32122), .B(n32123), .Z(n32120) );
  IV U31415 ( .A(n32093), .Z(n32117) );
  XOR U31416 ( .A(n32091), .B(n32124), .Z(n32093) );
  XNOR U31417 ( .A(n32125), .B(n32126), .Z(n32124) );
  ANDN U31418 ( .B(n32127), .A(n32128), .Z(n32125) );
  XNOR U31419 ( .A(n32129), .B(n32130), .Z(n32127) );
  IV U31420 ( .A(n32094), .Z(n32091) );
  XOR U31421 ( .A(n32131), .B(n32132), .Z(n32094) );
  ANDN U31422 ( .B(n32133), .A(n32134), .Z(n32131) );
  XOR U31423 ( .A(n32132), .B(n32135), .Z(n32133) );
  XOR U31424 ( .A(n32136), .B(n32137), .Z(n32107) );
  XNOR U31425 ( .A(n32102), .B(n32138), .Z(n32137) );
  IV U31426 ( .A(n32105), .Z(n32138) );
  XOR U31427 ( .A(n32139), .B(n32140), .Z(n32105) );
  ANDN U31428 ( .B(n32141), .A(n32142), .Z(n32139) );
  XOR U31429 ( .A(n32140), .B(n32143), .Z(n32141) );
  XNOR U31430 ( .A(n32144), .B(n32145), .Z(n32102) );
  ANDN U31431 ( .B(n32146), .A(n32147), .Z(n32144) );
  XOR U31432 ( .A(n32145), .B(n32148), .Z(n32146) );
  IV U31433 ( .A(n32101), .Z(n32136) );
  XOR U31434 ( .A(n32099), .B(n32149), .Z(n32101) );
  XNOR U31435 ( .A(n32150), .B(n32151), .Z(n32149) );
  ANDN U31436 ( .B(n32152), .A(n32153), .Z(n32150) );
  XNOR U31437 ( .A(n32154), .B(n32155), .Z(n32152) );
  IV U31438 ( .A(n32103), .Z(n32099) );
  XOR U31439 ( .A(n32156), .B(n32157), .Z(n32103) );
  ANDN U31440 ( .B(n32158), .A(n32159), .Z(n32156) );
  XOR U31441 ( .A(n32160), .B(n32157), .Z(n32158) );
  XOR U31442 ( .A(n32114), .B(n31967), .Z(n32115) );
  XOR U31443 ( .A(n32161), .B(n32162), .Z(n31967) );
  AND U31444 ( .A(n416), .B(n32163), .Z(n32161) );
  XOR U31445 ( .A(n32164), .B(n32162), .Z(n32163) );
  XNOR U31446 ( .A(n32165), .B(n32166), .Z(n32114) );
  NAND U31447 ( .A(n32167), .B(n32168), .Z(n32166) );
  XOR U31448 ( .A(n32169), .B(n32066), .Z(n32168) );
  XOR U31449 ( .A(n32142), .B(n32143), .Z(n32066) );
  XOR U31450 ( .A(n32170), .B(n32135), .Z(n32143) );
  XOR U31451 ( .A(n32171), .B(n32123), .Z(n32135) );
  XOR U31452 ( .A(n32172), .B(n32173), .Z(n32123) );
  ANDN U31453 ( .B(n32174), .A(n32175), .Z(n32172) );
  XOR U31454 ( .A(n32173), .B(n32176), .Z(n32174) );
  IV U31455 ( .A(n32121), .Z(n32171) );
  XOR U31456 ( .A(n32119), .B(n32177), .Z(n32121) );
  XOR U31457 ( .A(n32178), .B(n32179), .Z(n32177) );
  ANDN U31458 ( .B(n32180), .A(n32181), .Z(n32178) );
  XOR U31459 ( .A(n32182), .B(n32179), .Z(n32180) );
  IV U31460 ( .A(n32122), .Z(n32119) );
  XOR U31461 ( .A(n32183), .B(n32184), .Z(n32122) );
  ANDN U31462 ( .B(n32185), .A(n32186), .Z(n32183) );
  XOR U31463 ( .A(n32184), .B(n32187), .Z(n32185) );
  IV U31464 ( .A(n32134), .Z(n32170) );
  XOR U31465 ( .A(n32188), .B(n32189), .Z(n32134) );
  XNOR U31466 ( .A(n32129), .B(n32190), .Z(n32189) );
  IV U31467 ( .A(n32132), .Z(n32190) );
  XOR U31468 ( .A(n32191), .B(n32192), .Z(n32132) );
  ANDN U31469 ( .B(n32193), .A(n32194), .Z(n32191) );
  XOR U31470 ( .A(n32192), .B(n32195), .Z(n32193) );
  XNOR U31471 ( .A(n32196), .B(n32197), .Z(n32129) );
  ANDN U31472 ( .B(n32198), .A(n32199), .Z(n32196) );
  XOR U31473 ( .A(n32197), .B(n32200), .Z(n32198) );
  IV U31474 ( .A(n32128), .Z(n32188) );
  XOR U31475 ( .A(n32126), .B(n32201), .Z(n32128) );
  XOR U31476 ( .A(n32202), .B(n32203), .Z(n32201) );
  ANDN U31477 ( .B(n32204), .A(n32205), .Z(n32202) );
  XOR U31478 ( .A(n32206), .B(n32203), .Z(n32204) );
  IV U31479 ( .A(n32130), .Z(n32126) );
  XOR U31480 ( .A(n32207), .B(n32208), .Z(n32130) );
  ANDN U31481 ( .B(n32209), .A(n32210), .Z(n32207) );
  XOR U31482 ( .A(n32211), .B(n32208), .Z(n32209) );
  XOR U31483 ( .A(n32212), .B(n32213), .Z(n32142) );
  XOR U31484 ( .A(n32160), .B(n32214), .Z(n32213) );
  IV U31485 ( .A(n32140), .Z(n32214) );
  XOR U31486 ( .A(n32215), .B(n32216), .Z(n32140) );
  ANDN U31487 ( .B(n32217), .A(n32218), .Z(n32215) );
  XOR U31488 ( .A(n32216), .B(n32219), .Z(n32217) );
  XOR U31489 ( .A(n32220), .B(n32148), .Z(n32160) );
  XOR U31490 ( .A(n32221), .B(n32222), .Z(n32148) );
  ANDN U31491 ( .B(n32223), .A(n32224), .Z(n32221) );
  XOR U31492 ( .A(n32222), .B(n32225), .Z(n32223) );
  IV U31493 ( .A(n32147), .Z(n32220) );
  XOR U31494 ( .A(n32226), .B(n32227), .Z(n32147) );
  XOR U31495 ( .A(n32228), .B(n32229), .Z(n32227) );
  ANDN U31496 ( .B(n32230), .A(n32231), .Z(n32228) );
  XOR U31497 ( .A(n32232), .B(n32229), .Z(n32230) );
  IV U31498 ( .A(n32145), .Z(n32226) );
  XOR U31499 ( .A(n32233), .B(n32234), .Z(n32145) );
  ANDN U31500 ( .B(n32235), .A(n32236), .Z(n32233) );
  XOR U31501 ( .A(n32234), .B(n32237), .Z(n32235) );
  IV U31502 ( .A(n32159), .Z(n32212) );
  XOR U31503 ( .A(n32238), .B(n32239), .Z(n32159) );
  XNOR U31504 ( .A(n32154), .B(n32240), .Z(n32239) );
  IV U31505 ( .A(n32157), .Z(n32240) );
  XOR U31506 ( .A(n32241), .B(n32242), .Z(n32157) );
  ANDN U31507 ( .B(n32243), .A(n32244), .Z(n32241) );
  XOR U31508 ( .A(n32245), .B(n32242), .Z(n32243) );
  XNOR U31509 ( .A(n32246), .B(n32247), .Z(n32154) );
  ANDN U31510 ( .B(n32248), .A(n32249), .Z(n32246) );
  XOR U31511 ( .A(n32247), .B(n32250), .Z(n32248) );
  IV U31512 ( .A(n32153), .Z(n32238) );
  XOR U31513 ( .A(n32151), .B(n32251), .Z(n32153) );
  XOR U31514 ( .A(n32252), .B(n32253), .Z(n32251) );
  ANDN U31515 ( .B(n32254), .A(n32255), .Z(n32252) );
  XOR U31516 ( .A(n32256), .B(n32253), .Z(n32254) );
  IV U31517 ( .A(n32155), .Z(n32151) );
  XOR U31518 ( .A(n32257), .B(n32258), .Z(n32155) );
  ANDN U31519 ( .B(n32259), .A(n32260), .Z(n32257) );
  XOR U31520 ( .A(n32261), .B(n32258), .Z(n32259) );
  IV U31521 ( .A(n32165), .Z(n32169) );
  XOR U31522 ( .A(n32165), .B(n32068), .Z(n32167) );
  XOR U31523 ( .A(n32262), .B(n32263), .Z(n32068) );
  AND U31524 ( .A(n416), .B(n32264), .Z(n32262) );
  XOR U31525 ( .A(n32265), .B(n32263), .Z(n32264) );
  NANDN U31526 ( .A(n32070), .B(n32072), .Z(n32165) );
  XOR U31527 ( .A(n32266), .B(n32267), .Z(n32072) );
  AND U31528 ( .A(n416), .B(n32268), .Z(n32266) );
  XOR U31529 ( .A(n32267), .B(n32269), .Z(n32268) );
  XNOR U31530 ( .A(n32270), .B(n32271), .Z(n416) );
  AND U31531 ( .A(n32272), .B(n32273), .Z(n32270) );
  XOR U31532 ( .A(n32271), .B(n32083), .Z(n32273) );
  XNOR U31533 ( .A(n32274), .B(n32275), .Z(n32083) );
  ANDN U31534 ( .B(n32276), .A(n32277), .Z(n32274) );
  XOR U31535 ( .A(n32275), .B(n32278), .Z(n32276) );
  XNOR U31536 ( .A(n32271), .B(n32085), .Z(n32272) );
  XOR U31537 ( .A(n32279), .B(n32280), .Z(n32085) );
  AND U31538 ( .A(n420), .B(n32281), .Z(n32279) );
  XOR U31539 ( .A(n32282), .B(n32280), .Z(n32281) );
  XOR U31540 ( .A(n32283), .B(n32284), .Z(n32271) );
  AND U31541 ( .A(n32285), .B(n32286), .Z(n32283) );
  XOR U31542 ( .A(n32284), .B(n32110), .Z(n32286) );
  XOR U31543 ( .A(n32277), .B(n32278), .Z(n32110) );
  XNOR U31544 ( .A(n32287), .B(n32288), .Z(n32278) );
  ANDN U31545 ( .B(n32289), .A(n32290), .Z(n32287) );
  XOR U31546 ( .A(n32291), .B(n32292), .Z(n32289) );
  XOR U31547 ( .A(n32293), .B(n32294), .Z(n32277) );
  XNOR U31548 ( .A(n32295), .B(n32296), .Z(n32294) );
  ANDN U31549 ( .B(n32297), .A(n32298), .Z(n32295) );
  XNOR U31550 ( .A(n32299), .B(n32300), .Z(n32297) );
  IV U31551 ( .A(n32275), .Z(n32293) );
  XOR U31552 ( .A(n32301), .B(n32302), .Z(n32275) );
  ANDN U31553 ( .B(n32303), .A(n32304), .Z(n32301) );
  XOR U31554 ( .A(n32302), .B(n32305), .Z(n32303) );
  XNOR U31555 ( .A(n32284), .B(n32112), .Z(n32285) );
  XOR U31556 ( .A(n32306), .B(n32307), .Z(n32112) );
  AND U31557 ( .A(n420), .B(n32308), .Z(n32306) );
  XOR U31558 ( .A(n32309), .B(n32307), .Z(n32308) );
  XNOR U31559 ( .A(n32310), .B(n32311), .Z(n32284) );
  AND U31560 ( .A(n32312), .B(n32313), .Z(n32310) );
  XNOR U31561 ( .A(n32311), .B(n32162), .Z(n32313) );
  XOR U31562 ( .A(n32304), .B(n32305), .Z(n32162) );
  XOR U31563 ( .A(n32314), .B(n32292), .Z(n32305) );
  XNOR U31564 ( .A(n32315), .B(n32316), .Z(n32292) );
  ANDN U31565 ( .B(n32317), .A(n32318), .Z(n32315) );
  XOR U31566 ( .A(n32319), .B(n32320), .Z(n32317) );
  IV U31567 ( .A(n32290), .Z(n32314) );
  XOR U31568 ( .A(n32288), .B(n32321), .Z(n32290) );
  XNOR U31569 ( .A(n32322), .B(n32323), .Z(n32321) );
  ANDN U31570 ( .B(n32324), .A(n32325), .Z(n32322) );
  XNOR U31571 ( .A(n32326), .B(n32327), .Z(n32324) );
  IV U31572 ( .A(n32291), .Z(n32288) );
  XOR U31573 ( .A(n32328), .B(n32329), .Z(n32291) );
  ANDN U31574 ( .B(n32330), .A(n32331), .Z(n32328) );
  XOR U31575 ( .A(n32329), .B(n32332), .Z(n32330) );
  XOR U31576 ( .A(n32333), .B(n32334), .Z(n32304) );
  XNOR U31577 ( .A(n32299), .B(n32335), .Z(n32334) );
  IV U31578 ( .A(n32302), .Z(n32335) );
  XOR U31579 ( .A(n32336), .B(n32337), .Z(n32302) );
  ANDN U31580 ( .B(n32338), .A(n32339), .Z(n32336) );
  XOR U31581 ( .A(n32337), .B(n32340), .Z(n32338) );
  XNOR U31582 ( .A(n32341), .B(n32342), .Z(n32299) );
  ANDN U31583 ( .B(n32343), .A(n32344), .Z(n32341) );
  XOR U31584 ( .A(n32342), .B(n32345), .Z(n32343) );
  IV U31585 ( .A(n32298), .Z(n32333) );
  XOR U31586 ( .A(n32296), .B(n32346), .Z(n32298) );
  XNOR U31587 ( .A(n32347), .B(n32348), .Z(n32346) );
  ANDN U31588 ( .B(n32349), .A(n32350), .Z(n32347) );
  XNOR U31589 ( .A(n32351), .B(n32352), .Z(n32349) );
  IV U31590 ( .A(n32300), .Z(n32296) );
  XOR U31591 ( .A(n32353), .B(n32354), .Z(n32300) );
  ANDN U31592 ( .B(n32355), .A(n32356), .Z(n32353) );
  XOR U31593 ( .A(n32357), .B(n32354), .Z(n32355) );
  XOR U31594 ( .A(n32311), .B(n32164), .Z(n32312) );
  XOR U31595 ( .A(n32358), .B(n32359), .Z(n32164) );
  AND U31596 ( .A(n420), .B(n32360), .Z(n32358) );
  XOR U31597 ( .A(n32361), .B(n32359), .Z(n32360) );
  XNOR U31598 ( .A(n32362), .B(n32363), .Z(n32311) );
  NAND U31599 ( .A(n32364), .B(n32365), .Z(n32363) );
  XOR U31600 ( .A(n32366), .B(n32263), .Z(n32365) );
  XOR U31601 ( .A(n32339), .B(n32340), .Z(n32263) );
  XOR U31602 ( .A(n32367), .B(n32332), .Z(n32340) );
  XOR U31603 ( .A(n32368), .B(n32320), .Z(n32332) );
  XOR U31604 ( .A(n32369), .B(n32370), .Z(n32320) );
  ANDN U31605 ( .B(n32371), .A(n32372), .Z(n32369) );
  XOR U31606 ( .A(n32370), .B(n32373), .Z(n32371) );
  IV U31607 ( .A(n32318), .Z(n32368) );
  XOR U31608 ( .A(n32316), .B(n32374), .Z(n32318) );
  XOR U31609 ( .A(n32375), .B(n32376), .Z(n32374) );
  ANDN U31610 ( .B(n32377), .A(n32378), .Z(n32375) );
  XOR U31611 ( .A(n32379), .B(n32376), .Z(n32377) );
  IV U31612 ( .A(n32319), .Z(n32316) );
  XOR U31613 ( .A(n32380), .B(n32381), .Z(n32319) );
  ANDN U31614 ( .B(n32382), .A(n32383), .Z(n32380) );
  XOR U31615 ( .A(n32381), .B(n32384), .Z(n32382) );
  IV U31616 ( .A(n32331), .Z(n32367) );
  XOR U31617 ( .A(n32385), .B(n32386), .Z(n32331) );
  XNOR U31618 ( .A(n32326), .B(n32387), .Z(n32386) );
  IV U31619 ( .A(n32329), .Z(n32387) );
  XOR U31620 ( .A(n32388), .B(n32389), .Z(n32329) );
  ANDN U31621 ( .B(n32390), .A(n32391), .Z(n32388) );
  XOR U31622 ( .A(n32389), .B(n32392), .Z(n32390) );
  XNOR U31623 ( .A(n32393), .B(n32394), .Z(n32326) );
  ANDN U31624 ( .B(n32395), .A(n32396), .Z(n32393) );
  XOR U31625 ( .A(n32394), .B(n32397), .Z(n32395) );
  IV U31626 ( .A(n32325), .Z(n32385) );
  XOR U31627 ( .A(n32323), .B(n32398), .Z(n32325) );
  XOR U31628 ( .A(n32399), .B(n32400), .Z(n32398) );
  ANDN U31629 ( .B(n32401), .A(n32402), .Z(n32399) );
  XOR U31630 ( .A(n32403), .B(n32400), .Z(n32401) );
  IV U31631 ( .A(n32327), .Z(n32323) );
  XOR U31632 ( .A(n32404), .B(n32405), .Z(n32327) );
  ANDN U31633 ( .B(n32406), .A(n32407), .Z(n32404) );
  XOR U31634 ( .A(n32408), .B(n32405), .Z(n32406) );
  XOR U31635 ( .A(n32409), .B(n32410), .Z(n32339) );
  XOR U31636 ( .A(n32357), .B(n32411), .Z(n32410) );
  IV U31637 ( .A(n32337), .Z(n32411) );
  XOR U31638 ( .A(n32412), .B(n32413), .Z(n32337) );
  ANDN U31639 ( .B(n32414), .A(n32415), .Z(n32412) );
  XOR U31640 ( .A(n32413), .B(n32416), .Z(n32414) );
  XOR U31641 ( .A(n32417), .B(n32345), .Z(n32357) );
  XOR U31642 ( .A(n32418), .B(n32419), .Z(n32345) );
  ANDN U31643 ( .B(n32420), .A(n32421), .Z(n32418) );
  XOR U31644 ( .A(n32419), .B(n32422), .Z(n32420) );
  IV U31645 ( .A(n32344), .Z(n32417) );
  XOR U31646 ( .A(n32423), .B(n32424), .Z(n32344) );
  XOR U31647 ( .A(n32425), .B(n32426), .Z(n32424) );
  ANDN U31648 ( .B(n32427), .A(n32428), .Z(n32425) );
  XOR U31649 ( .A(n32429), .B(n32426), .Z(n32427) );
  IV U31650 ( .A(n32342), .Z(n32423) );
  XOR U31651 ( .A(n32430), .B(n32431), .Z(n32342) );
  ANDN U31652 ( .B(n32432), .A(n32433), .Z(n32430) );
  XOR U31653 ( .A(n32431), .B(n32434), .Z(n32432) );
  IV U31654 ( .A(n32356), .Z(n32409) );
  XOR U31655 ( .A(n32435), .B(n32436), .Z(n32356) );
  XNOR U31656 ( .A(n32351), .B(n32437), .Z(n32436) );
  IV U31657 ( .A(n32354), .Z(n32437) );
  XOR U31658 ( .A(n32438), .B(n32439), .Z(n32354) );
  ANDN U31659 ( .B(n32440), .A(n32441), .Z(n32438) );
  XOR U31660 ( .A(n32442), .B(n32439), .Z(n32440) );
  XNOR U31661 ( .A(n32443), .B(n32444), .Z(n32351) );
  ANDN U31662 ( .B(n32445), .A(n32446), .Z(n32443) );
  XOR U31663 ( .A(n32444), .B(n32447), .Z(n32445) );
  IV U31664 ( .A(n32350), .Z(n32435) );
  XOR U31665 ( .A(n32348), .B(n32448), .Z(n32350) );
  XOR U31666 ( .A(n32449), .B(n32450), .Z(n32448) );
  ANDN U31667 ( .B(n32451), .A(n32452), .Z(n32449) );
  XOR U31668 ( .A(n32453), .B(n32450), .Z(n32451) );
  IV U31669 ( .A(n32352), .Z(n32348) );
  XOR U31670 ( .A(n32454), .B(n32455), .Z(n32352) );
  ANDN U31671 ( .B(n32456), .A(n32457), .Z(n32454) );
  XOR U31672 ( .A(n32458), .B(n32455), .Z(n32456) );
  IV U31673 ( .A(n32362), .Z(n32366) );
  XOR U31674 ( .A(n32362), .B(n32265), .Z(n32364) );
  XOR U31675 ( .A(n32459), .B(n32460), .Z(n32265) );
  AND U31676 ( .A(n420), .B(n32461), .Z(n32459) );
  XOR U31677 ( .A(n32462), .B(n32460), .Z(n32461) );
  NANDN U31678 ( .A(n32267), .B(n32269), .Z(n32362) );
  XOR U31679 ( .A(n32463), .B(n32464), .Z(n32269) );
  AND U31680 ( .A(n420), .B(n32465), .Z(n32463) );
  XOR U31681 ( .A(n32464), .B(n32466), .Z(n32465) );
  XNOR U31682 ( .A(n32467), .B(n32468), .Z(n420) );
  AND U31683 ( .A(n32469), .B(n32470), .Z(n32467) );
  XOR U31684 ( .A(n32468), .B(n32280), .Z(n32470) );
  XNOR U31685 ( .A(n32471), .B(n32472), .Z(n32280) );
  ANDN U31686 ( .B(n32473), .A(n32474), .Z(n32471) );
  XOR U31687 ( .A(n32472), .B(n32475), .Z(n32473) );
  XNOR U31688 ( .A(n32468), .B(n32282), .Z(n32469) );
  XOR U31689 ( .A(n32476), .B(n32477), .Z(n32282) );
  AND U31690 ( .A(n424), .B(n32478), .Z(n32476) );
  XOR U31691 ( .A(n32479), .B(n32477), .Z(n32478) );
  XOR U31692 ( .A(n32480), .B(n32481), .Z(n32468) );
  AND U31693 ( .A(n32482), .B(n32483), .Z(n32480) );
  XOR U31694 ( .A(n32481), .B(n32307), .Z(n32483) );
  XOR U31695 ( .A(n32474), .B(n32475), .Z(n32307) );
  XNOR U31696 ( .A(n32484), .B(n32485), .Z(n32475) );
  ANDN U31697 ( .B(n32486), .A(n32487), .Z(n32484) );
  XOR U31698 ( .A(n32488), .B(n32489), .Z(n32486) );
  XOR U31699 ( .A(n32490), .B(n32491), .Z(n32474) );
  XNOR U31700 ( .A(n32492), .B(n32493), .Z(n32491) );
  ANDN U31701 ( .B(n32494), .A(n32495), .Z(n32492) );
  XNOR U31702 ( .A(n32496), .B(n32497), .Z(n32494) );
  IV U31703 ( .A(n32472), .Z(n32490) );
  XOR U31704 ( .A(n32498), .B(n32499), .Z(n32472) );
  ANDN U31705 ( .B(n32500), .A(n32501), .Z(n32498) );
  XOR U31706 ( .A(n32499), .B(n32502), .Z(n32500) );
  XNOR U31707 ( .A(n32481), .B(n32309), .Z(n32482) );
  XOR U31708 ( .A(n32503), .B(n32504), .Z(n32309) );
  AND U31709 ( .A(n424), .B(n32505), .Z(n32503) );
  XOR U31710 ( .A(n32506), .B(n32504), .Z(n32505) );
  XNOR U31711 ( .A(n32507), .B(n32508), .Z(n32481) );
  AND U31712 ( .A(n32509), .B(n32510), .Z(n32507) );
  XNOR U31713 ( .A(n32508), .B(n32359), .Z(n32510) );
  XOR U31714 ( .A(n32501), .B(n32502), .Z(n32359) );
  XOR U31715 ( .A(n32511), .B(n32489), .Z(n32502) );
  XNOR U31716 ( .A(n32512), .B(n32513), .Z(n32489) );
  ANDN U31717 ( .B(n32514), .A(n32515), .Z(n32512) );
  XOR U31718 ( .A(n32516), .B(n32517), .Z(n32514) );
  IV U31719 ( .A(n32487), .Z(n32511) );
  XOR U31720 ( .A(n32485), .B(n32518), .Z(n32487) );
  XNOR U31721 ( .A(n32519), .B(n32520), .Z(n32518) );
  ANDN U31722 ( .B(n32521), .A(n32522), .Z(n32519) );
  XNOR U31723 ( .A(n32523), .B(n32524), .Z(n32521) );
  IV U31724 ( .A(n32488), .Z(n32485) );
  XOR U31725 ( .A(n32525), .B(n32526), .Z(n32488) );
  ANDN U31726 ( .B(n32527), .A(n32528), .Z(n32525) );
  XOR U31727 ( .A(n32526), .B(n32529), .Z(n32527) );
  XOR U31728 ( .A(n32530), .B(n32531), .Z(n32501) );
  XNOR U31729 ( .A(n32496), .B(n32532), .Z(n32531) );
  IV U31730 ( .A(n32499), .Z(n32532) );
  XOR U31731 ( .A(n32533), .B(n32534), .Z(n32499) );
  ANDN U31732 ( .B(n32535), .A(n32536), .Z(n32533) );
  XOR U31733 ( .A(n32534), .B(n32537), .Z(n32535) );
  XNOR U31734 ( .A(n32538), .B(n32539), .Z(n32496) );
  ANDN U31735 ( .B(n32540), .A(n32541), .Z(n32538) );
  XOR U31736 ( .A(n32539), .B(n32542), .Z(n32540) );
  IV U31737 ( .A(n32495), .Z(n32530) );
  XOR U31738 ( .A(n32493), .B(n32543), .Z(n32495) );
  XNOR U31739 ( .A(n32544), .B(n32545), .Z(n32543) );
  ANDN U31740 ( .B(n32546), .A(n32547), .Z(n32544) );
  XNOR U31741 ( .A(n32548), .B(n32549), .Z(n32546) );
  IV U31742 ( .A(n32497), .Z(n32493) );
  XOR U31743 ( .A(n32550), .B(n32551), .Z(n32497) );
  ANDN U31744 ( .B(n32552), .A(n32553), .Z(n32550) );
  XOR U31745 ( .A(n32554), .B(n32551), .Z(n32552) );
  XOR U31746 ( .A(n32508), .B(n32361), .Z(n32509) );
  XOR U31747 ( .A(n32555), .B(n32556), .Z(n32361) );
  AND U31748 ( .A(n424), .B(n32557), .Z(n32555) );
  XOR U31749 ( .A(n32558), .B(n32556), .Z(n32557) );
  XNOR U31750 ( .A(n32559), .B(n32560), .Z(n32508) );
  NAND U31751 ( .A(n32561), .B(n32562), .Z(n32560) );
  XOR U31752 ( .A(n32563), .B(n32460), .Z(n32562) );
  XOR U31753 ( .A(n32536), .B(n32537), .Z(n32460) );
  XOR U31754 ( .A(n32564), .B(n32529), .Z(n32537) );
  XOR U31755 ( .A(n32565), .B(n32517), .Z(n32529) );
  XOR U31756 ( .A(n32566), .B(n32567), .Z(n32517) );
  ANDN U31757 ( .B(n32568), .A(n32569), .Z(n32566) );
  XOR U31758 ( .A(n32567), .B(n32570), .Z(n32568) );
  IV U31759 ( .A(n32515), .Z(n32565) );
  XOR U31760 ( .A(n32513), .B(n32571), .Z(n32515) );
  XOR U31761 ( .A(n32572), .B(n32573), .Z(n32571) );
  ANDN U31762 ( .B(n32574), .A(n32575), .Z(n32572) );
  XOR U31763 ( .A(n32576), .B(n32573), .Z(n32574) );
  IV U31764 ( .A(n32516), .Z(n32513) );
  XOR U31765 ( .A(n32577), .B(n32578), .Z(n32516) );
  ANDN U31766 ( .B(n32579), .A(n32580), .Z(n32577) );
  XOR U31767 ( .A(n32578), .B(n32581), .Z(n32579) );
  IV U31768 ( .A(n32528), .Z(n32564) );
  XOR U31769 ( .A(n32582), .B(n32583), .Z(n32528) );
  XNOR U31770 ( .A(n32523), .B(n32584), .Z(n32583) );
  IV U31771 ( .A(n32526), .Z(n32584) );
  XOR U31772 ( .A(n32585), .B(n32586), .Z(n32526) );
  ANDN U31773 ( .B(n32587), .A(n32588), .Z(n32585) );
  XOR U31774 ( .A(n32586), .B(n32589), .Z(n32587) );
  XNOR U31775 ( .A(n32590), .B(n32591), .Z(n32523) );
  ANDN U31776 ( .B(n32592), .A(n32593), .Z(n32590) );
  XOR U31777 ( .A(n32591), .B(n32594), .Z(n32592) );
  IV U31778 ( .A(n32522), .Z(n32582) );
  XOR U31779 ( .A(n32520), .B(n32595), .Z(n32522) );
  XOR U31780 ( .A(n32596), .B(n32597), .Z(n32595) );
  ANDN U31781 ( .B(n32598), .A(n32599), .Z(n32596) );
  XOR U31782 ( .A(n32600), .B(n32597), .Z(n32598) );
  IV U31783 ( .A(n32524), .Z(n32520) );
  XOR U31784 ( .A(n32601), .B(n32602), .Z(n32524) );
  ANDN U31785 ( .B(n32603), .A(n32604), .Z(n32601) );
  XOR U31786 ( .A(n32605), .B(n32602), .Z(n32603) );
  XOR U31787 ( .A(n32606), .B(n32607), .Z(n32536) );
  XOR U31788 ( .A(n32554), .B(n32608), .Z(n32607) );
  IV U31789 ( .A(n32534), .Z(n32608) );
  XOR U31790 ( .A(n32609), .B(n32610), .Z(n32534) );
  ANDN U31791 ( .B(n32611), .A(n32612), .Z(n32609) );
  XOR U31792 ( .A(n32610), .B(n32613), .Z(n32611) );
  XOR U31793 ( .A(n32614), .B(n32542), .Z(n32554) );
  XOR U31794 ( .A(n32615), .B(n32616), .Z(n32542) );
  ANDN U31795 ( .B(n32617), .A(n32618), .Z(n32615) );
  XOR U31796 ( .A(n32616), .B(n32619), .Z(n32617) );
  IV U31797 ( .A(n32541), .Z(n32614) );
  XOR U31798 ( .A(n32620), .B(n32621), .Z(n32541) );
  XOR U31799 ( .A(n32622), .B(n32623), .Z(n32621) );
  ANDN U31800 ( .B(n32624), .A(n32625), .Z(n32622) );
  XOR U31801 ( .A(n32626), .B(n32623), .Z(n32624) );
  IV U31802 ( .A(n32539), .Z(n32620) );
  XOR U31803 ( .A(n32627), .B(n32628), .Z(n32539) );
  ANDN U31804 ( .B(n32629), .A(n32630), .Z(n32627) );
  XOR U31805 ( .A(n32628), .B(n32631), .Z(n32629) );
  IV U31806 ( .A(n32553), .Z(n32606) );
  XOR U31807 ( .A(n32632), .B(n32633), .Z(n32553) );
  XNOR U31808 ( .A(n32548), .B(n32634), .Z(n32633) );
  IV U31809 ( .A(n32551), .Z(n32634) );
  XOR U31810 ( .A(n32635), .B(n32636), .Z(n32551) );
  ANDN U31811 ( .B(n32637), .A(n32638), .Z(n32635) );
  XOR U31812 ( .A(n32639), .B(n32636), .Z(n32637) );
  XNOR U31813 ( .A(n32640), .B(n32641), .Z(n32548) );
  ANDN U31814 ( .B(n32642), .A(n32643), .Z(n32640) );
  XOR U31815 ( .A(n32641), .B(n32644), .Z(n32642) );
  IV U31816 ( .A(n32547), .Z(n32632) );
  XOR U31817 ( .A(n32545), .B(n32645), .Z(n32547) );
  XOR U31818 ( .A(n32646), .B(n32647), .Z(n32645) );
  ANDN U31819 ( .B(n32648), .A(n32649), .Z(n32646) );
  XOR U31820 ( .A(n32650), .B(n32647), .Z(n32648) );
  IV U31821 ( .A(n32549), .Z(n32545) );
  XOR U31822 ( .A(n32651), .B(n32652), .Z(n32549) );
  ANDN U31823 ( .B(n32653), .A(n32654), .Z(n32651) );
  XOR U31824 ( .A(n32655), .B(n32652), .Z(n32653) );
  IV U31825 ( .A(n32559), .Z(n32563) );
  XOR U31826 ( .A(n32559), .B(n32462), .Z(n32561) );
  XOR U31827 ( .A(n32656), .B(n32657), .Z(n32462) );
  AND U31828 ( .A(n424), .B(n32658), .Z(n32656) );
  XOR U31829 ( .A(n32659), .B(n32657), .Z(n32658) );
  NANDN U31830 ( .A(n32464), .B(n32466), .Z(n32559) );
  XOR U31831 ( .A(n32660), .B(n32661), .Z(n32466) );
  AND U31832 ( .A(n424), .B(n32662), .Z(n32660) );
  XOR U31833 ( .A(n32661), .B(n32663), .Z(n32662) );
  XNOR U31834 ( .A(n32664), .B(n32665), .Z(n424) );
  AND U31835 ( .A(n32666), .B(n32667), .Z(n32664) );
  XOR U31836 ( .A(n32665), .B(n32477), .Z(n32667) );
  XNOR U31837 ( .A(n32668), .B(n32669), .Z(n32477) );
  ANDN U31838 ( .B(n32670), .A(n32671), .Z(n32668) );
  XOR U31839 ( .A(n32669), .B(n32672), .Z(n32670) );
  XNOR U31840 ( .A(n32665), .B(n32479), .Z(n32666) );
  XOR U31841 ( .A(n32673), .B(n32674), .Z(n32479) );
  AND U31842 ( .A(n428), .B(n32675), .Z(n32673) );
  XOR U31843 ( .A(n32676), .B(n32674), .Z(n32675) );
  XOR U31844 ( .A(n32677), .B(n32678), .Z(n32665) );
  AND U31845 ( .A(n32679), .B(n32680), .Z(n32677) );
  XOR U31846 ( .A(n32678), .B(n32504), .Z(n32680) );
  XOR U31847 ( .A(n32671), .B(n32672), .Z(n32504) );
  XNOR U31848 ( .A(n32681), .B(n32682), .Z(n32672) );
  ANDN U31849 ( .B(n32683), .A(n32684), .Z(n32681) );
  XOR U31850 ( .A(n32685), .B(n32686), .Z(n32683) );
  XOR U31851 ( .A(n32687), .B(n32688), .Z(n32671) );
  XNOR U31852 ( .A(n32689), .B(n32690), .Z(n32688) );
  ANDN U31853 ( .B(n32691), .A(n32692), .Z(n32689) );
  XNOR U31854 ( .A(n32693), .B(n32694), .Z(n32691) );
  IV U31855 ( .A(n32669), .Z(n32687) );
  XOR U31856 ( .A(n32695), .B(n32696), .Z(n32669) );
  ANDN U31857 ( .B(n32697), .A(n32698), .Z(n32695) );
  XOR U31858 ( .A(n32696), .B(n32699), .Z(n32697) );
  XNOR U31859 ( .A(n32678), .B(n32506), .Z(n32679) );
  XOR U31860 ( .A(n32700), .B(n32701), .Z(n32506) );
  AND U31861 ( .A(n428), .B(n32702), .Z(n32700) );
  XOR U31862 ( .A(n32703), .B(n32701), .Z(n32702) );
  XNOR U31863 ( .A(n32704), .B(n32705), .Z(n32678) );
  AND U31864 ( .A(n32706), .B(n32707), .Z(n32704) );
  XNOR U31865 ( .A(n32705), .B(n32556), .Z(n32707) );
  XOR U31866 ( .A(n32698), .B(n32699), .Z(n32556) );
  XOR U31867 ( .A(n32708), .B(n32686), .Z(n32699) );
  XNOR U31868 ( .A(n32709), .B(n32710), .Z(n32686) );
  ANDN U31869 ( .B(n32711), .A(n32712), .Z(n32709) );
  XOR U31870 ( .A(n32713), .B(n32714), .Z(n32711) );
  IV U31871 ( .A(n32684), .Z(n32708) );
  XOR U31872 ( .A(n32682), .B(n32715), .Z(n32684) );
  XNOR U31873 ( .A(n32716), .B(n32717), .Z(n32715) );
  ANDN U31874 ( .B(n32718), .A(n32719), .Z(n32716) );
  XNOR U31875 ( .A(n32720), .B(n32721), .Z(n32718) );
  IV U31876 ( .A(n32685), .Z(n32682) );
  XOR U31877 ( .A(n32722), .B(n32723), .Z(n32685) );
  ANDN U31878 ( .B(n32724), .A(n32725), .Z(n32722) );
  XOR U31879 ( .A(n32723), .B(n32726), .Z(n32724) );
  XOR U31880 ( .A(n32727), .B(n32728), .Z(n32698) );
  XNOR U31881 ( .A(n32693), .B(n32729), .Z(n32728) );
  IV U31882 ( .A(n32696), .Z(n32729) );
  XOR U31883 ( .A(n32730), .B(n32731), .Z(n32696) );
  ANDN U31884 ( .B(n32732), .A(n32733), .Z(n32730) );
  XOR U31885 ( .A(n32731), .B(n32734), .Z(n32732) );
  XNOR U31886 ( .A(n32735), .B(n32736), .Z(n32693) );
  ANDN U31887 ( .B(n32737), .A(n32738), .Z(n32735) );
  XOR U31888 ( .A(n32736), .B(n32739), .Z(n32737) );
  IV U31889 ( .A(n32692), .Z(n32727) );
  XOR U31890 ( .A(n32690), .B(n32740), .Z(n32692) );
  XNOR U31891 ( .A(n32741), .B(n32742), .Z(n32740) );
  ANDN U31892 ( .B(n32743), .A(n32744), .Z(n32741) );
  XNOR U31893 ( .A(n32745), .B(n32746), .Z(n32743) );
  IV U31894 ( .A(n32694), .Z(n32690) );
  XOR U31895 ( .A(n32747), .B(n32748), .Z(n32694) );
  ANDN U31896 ( .B(n32749), .A(n32750), .Z(n32747) );
  XOR U31897 ( .A(n32751), .B(n32748), .Z(n32749) );
  XOR U31898 ( .A(n32705), .B(n32558), .Z(n32706) );
  XOR U31899 ( .A(n32752), .B(n32753), .Z(n32558) );
  AND U31900 ( .A(n428), .B(n32754), .Z(n32752) );
  XOR U31901 ( .A(n32755), .B(n32753), .Z(n32754) );
  XNOR U31902 ( .A(n32756), .B(n32757), .Z(n32705) );
  NAND U31903 ( .A(n32758), .B(n32759), .Z(n32757) );
  XOR U31904 ( .A(n32760), .B(n32657), .Z(n32759) );
  XOR U31905 ( .A(n32733), .B(n32734), .Z(n32657) );
  XOR U31906 ( .A(n32761), .B(n32726), .Z(n32734) );
  XOR U31907 ( .A(n32762), .B(n32714), .Z(n32726) );
  XOR U31908 ( .A(n32763), .B(n32764), .Z(n32714) );
  ANDN U31909 ( .B(n32765), .A(n32766), .Z(n32763) );
  XOR U31910 ( .A(n32764), .B(n32767), .Z(n32765) );
  IV U31911 ( .A(n32712), .Z(n32762) );
  XOR U31912 ( .A(n32710), .B(n32768), .Z(n32712) );
  XOR U31913 ( .A(n32769), .B(n32770), .Z(n32768) );
  ANDN U31914 ( .B(n32771), .A(n32772), .Z(n32769) );
  XOR U31915 ( .A(n32773), .B(n32770), .Z(n32771) );
  IV U31916 ( .A(n32713), .Z(n32710) );
  XOR U31917 ( .A(n32774), .B(n32775), .Z(n32713) );
  ANDN U31918 ( .B(n32776), .A(n32777), .Z(n32774) );
  XOR U31919 ( .A(n32775), .B(n32778), .Z(n32776) );
  IV U31920 ( .A(n32725), .Z(n32761) );
  XOR U31921 ( .A(n32779), .B(n32780), .Z(n32725) );
  XNOR U31922 ( .A(n32720), .B(n32781), .Z(n32780) );
  IV U31923 ( .A(n32723), .Z(n32781) );
  XOR U31924 ( .A(n32782), .B(n32783), .Z(n32723) );
  ANDN U31925 ( .B(n32784), .A(n32785), .Z(n32782) );
  XOR U31926 ( .A(n32783), .B(n32786), .Z(n32784) );
  XNOR U31927 ( .A(n32787), .B(n32788), .Z(n32720) );
  ANDN U31928 ( .B(n32789), .A(n32790), .Z(n32787) );
  XOR U31929 ( .A(n32788), .B(n32791), .Z(n32789) );
  IV U31930 ( .A(n32719), .Z(n32779) );
  XOR U31931 ( .A(n32717), .B(n32792), .Z(n32719) );
  XOR U31932 ( .A(n32793), .B(n32794), .Z(n32792) );
  ANDN U31933 ( .B(n32795), .A(n32796), .Z(n32793) );
  XOR U31934 ( .A(n32797), .B(n32794), .Z(n32795) );
  IV U31935 ( .A(n32721), .Z(n32717) );
  XOR U31936 ( .A(n32798), .B(n32799), .Z(n32721) );
  ANDN U31937 ( .B(n32800), .A(n32801), .Z(n32798) );
  XOR U31938 ( .A(n32802), .B(n32799), .Z(n32800) );
  XOR U31939 ( .A(n32803), .B(n32804), .Z(n32733) );
  XOR U31940 ( .A(n32751), .B(n32805), .Z(n32804) );
  IV U31941 ( .A(n32731), .Z(n32805) );
  XOR U31942 ( .A(n32806), .B(n32807), .Z(n32731) );
  ANDN U31943 ( .B(n32808), .A(n32809), .Z(n32806) );
  XOR U31944 ( .A(n32807), .B(n32810), .Z(n32808) );
  XOR U31945 ( .A(n32811), .B(n32739), .Z(n32751) );
  XOR U31946 ( .A(n32812), .B(n32813), .Z(n32739) );
  ANDN U31947 ( .B(n32814), .A(n32815), .Z(n32812) );
  XOR U31948 ( .A(n32813), .B(n32816), .Z(n32814) );
  IV U31949 ( .A(n32738), .Z(n32811) );
  XOR U31950 ( .A(n32817), .B(n32818), .Z(n32738) );
  XOR U31951 ( .A(n32819), .B(n32820), .Z(n32818) );
  ANDN U31952 ( .B(n32821), .A(n32822), .Z(n32819) );
  XOR U31953 ( .A(n32823), .B(n32820), .Z(n32821) );
  IV U31954 ( .A(n32736), .Z(n32817) );
  XOR U31955 ( .A(n32824), .B(n32825), .Z(n32736) );
  ANDN U31956 ( .B(n32826), .A(n32827), .Z(n32824) );
  XOR U31957 ( .A(n32825), .B(n32828), .Z(n32826) );
  IV U31958 ( .A(n32750), .Z(n32803) );
  XOR U31959 ( .A(n32829), .B(n32830), .Z(n32750) );
  XNOR U31960 ( .A(n32745), .B(n32831), .Z(n32830) );
  IV U31961 ( .A(n32748), .Z(n32831) );
  XOR U31962 ( .A(n32832), .B(n32833), .Z(n32748) );
  ANDN U31963 ( .B(n32834), .A(n32835), .Z(n32832) );
  XOR U31964 ( .A(n32836), .B(n32833), .Z(n32834) );
  XNOR U31965 ( .A(n32837), .B(n32838), .Z(n32745) );
  ANDN U31966 ( .B(n32839), .A(n32840), .Z(n32837) );
  XOR U31967 ( .A(n32838), .B(n32841), .Z(n32839) );
  IV U31968 ( .A(n32744), .Z(n32829) );
  XOR U31969 ( .A(n32742), .B(n32842), .Z(n32744) );
  XOR U31970 ( .A(n32843), .B(n32844), .Z(n32842) );
  ANDN U31971 ( .B(n32845), .A(n32846), .Z(n32843) );
  XOR U31972 ( .A(n32847), .B(n32844), .Z(n32845) );
  IV U31973 ( .A(n32746), .Z(n32742) );
  XOR U31974 ( .A(n32848), .B(n32849), .Z(n32746) );
  ANDN U31975 ( .B(n32850), .A(n32851), .Z(n32848) );
  XOR U31976 ( .A(n32852), .B(n32849), .Z(n32850) );
  IV U31977 ( .A(n32756), .Z(n32760) );
  XOR U31978 ( .A(n32756), .B(n32659), .Z(n32758) );
  XOR U31979 ( .A(n32853), .B(n32854), .Z(n32659) );
  AND U31980 ( .A(n428), .B(n32855), .Z(n32853) );
  XOR U31981 ( .A(n32856), .B(n32854), .Z(n32855) );
  NANDN U31982 ( .A(n32661), .B(n32663), .Z(n32756) );
  XOR U31983 ( .A(n32857), .B(n32858), .Z(n32663) );
  AND U31984 ( .A(n428), .B(n32859), .Z(n32857) );
  XOR U31985 ( .A(n32858), .B(n32860), .Z(n32859) );
  XNOR U31986 ( .A(n32861), .B(n32862), .Z(n428) );
  AND U31987 ( .A(n32863), .B(n32864), .Z(n32861) );
  XOR U31988 ( .A(n32862), .B(n32674), .Z(n32864) );
  XNOR U31989 ( .A(n32865), .B(n32866), .Z(n32674) );
  ANDN U31990 ( .B(n32867), .A(n32868), .Z(n32865) );
  XOR U31991 ( .A(n32866), .B(n32869), .Z(n32867) );
  XNOR U31992 ( .A(n32862), .B(n32676), .Z(n32863) );
  XOR U31993 ( .A(n32870), .B(n32871), .Z(n32676) );
  AND U31994 ( .A(n432), .B(n32872), .Z(n32870) );
  XOR U31995 ( .A(n32873), .B(n32871), .Z(n32872) );
  XOR U31996 ( .A(n32874), .B(n32875), .Z(n32862) );
  AND U31997 ( .A(n32876), .B(n32877), .Z(n32874) );
  XOR U31998 ( .A(n32875), .B(n32701), .Z(n32877) );
  XOR U31999 ( .A(n32868), .B(n32869), .Z(n32701) );
  XNOR U32000 ( .A(n32878), .B(n32879), .Z(n32869) );
  ANDN U32001 ( .B(n32880), .A(n32881), .Z(n32878) );
  XOR U32002 ( .A(n32882), .B(n32883), .Z(n32880) );
  XOR U32003 ( .A(n32884), .B(n32885), .Z(n32868) );
  XNOR U32004 ( .A(n32886), .B(n32887), .Z(n32885) );
  ANDN U32005 ( .B(n32888), .A(n32889), .Z(n32886) );
  XNOR U32006 ( .A(n32890), .B(n32891), .Z(n32888) );
  IV U32007 ( .A(n32866), .Z(n32884) );
  XOR U32008 ( .A(n32892), .B(n32893), .Z(n32866) );
  ANDN U32009 ( .B(n32894), .A(n32895), .Z(n32892) );
  XOR U32010 ( .A(n32893), .B(n32896), .Z(n32894) );
  XNOR U32011 ( .A(n32875), .B(n32703), .Z(n32876) );
  XOR U32012 ( .A(n32897), .B(n32898), .Z(n32703) );
  AND U32013 ( .A(n432), .B(n32899), .Z(n32897) );
  XOR U32014 ( .A(n32900), .B(n32898), .Z(n32899) );
  XNOR U32015 ( .A(n32901), .B(n32902), .Z(n32875) );
  AND U32016 ( .A(n32903), .B(n32904), .Z(n32901) );
  XNOR U32017 ( .A(n32902), .B(n32753), .Z(n32904) );
  XOR U32018 ( .A(n32895), .B(n32896), .Z(n32753) );
  XOR U32019 ( .A(n32905), .B(n32883), .Z(n32896) );
  XNOR U32020 ( .A(n32906), .B(n32907), .Z(n32883) );
  ANDN U32021 ( .B(n32908), .A(n32909), .Z(n32906) );
  XOR U32022 ( .A(n32910), .B(n32911), .Z(n32908) );
  IV U32023 ( .A(n32881), .Z(n32905) );
  XOR U32024 ( .A(n32879), .B(n32912), .Z(n32881) );
  XNOR U32025 ( .A(n32913), .B(n32914), .Z(n32912) );
  ANDN U32026 ( .B(n32915), .A(n32916), .Z(n32913) );
  XNOR U32027 ( .A(n32917), .B(n32918), .Z(n32915) );
  IV U32028 ( .A(n32882), .Z(n32879) );
  XOR U32029 ( .A(n32919), .B(n32920), .Z(n32882) );
  ANDN U32030 ( .B(n32921), .A(n32922), .Z(n32919) );
  XOR U32031 ( .A(n32920), .B(n32923), .Z(n32921) );
  XOR U32032 ( .A(n32924), .B(n32925), .Z(n32895) );
  XNOR U32033 ( .A(n32890), .B(n32926), .Z(n32925) );
  IV U32034 ( .A(n32893), .Z(n32926) );
  XOR U32035 ( .A(n32927), .B(n32928), .Z(n32893) );
  ANDN U32036 ( .B(n32929), .A(n32930), .Z(n32927) );
  XOR U32037 ( .A(n32928), .B(n32931), .Z(n32929) );
  XNOR U32038 ( .A(n32932), .B(n32933), .Z(n32890) );
  ANDN U32039 ( .B(n32934), .A(n32935), .Z(n32932) );
  XOR U32040 ( .A(n32933), .B(n32936), .Z(n32934) );
  IV U32041 ( .A(n32889), .Z(n32924) );
  XOR U32042 ( .A(n32887), .B(n32937), .Z(n32889) );
  XNOR U32043 ( .A(n32938), .B(n32939), .Z(n32937) );
  ANDN U32044 ( .B(n32940), .A(n32941), .Z(n32938) );
  XNOR U32045 ( .A(n32942), .B(n32943), .Z(n32940) );
  IV U32046 ( .A(n32891), .Z(n32887) );
  XOR U32047 ( .A(n32944), .B(n32945), .Z(n32891) );
  ANDN U32048 ( .B(n32946), .A(n32947), .Z(n32944) );
  XOR U32049 ( .A(n32948), .B(n32945), .Z(n32946) );
  XOR U32050 ( .A(n32902), .B(n32755), .Z(n32903) );
  XOR U32051 ( .A(n32949), .B(n32950), .Z(n32755) );
  AND U32052 ( .A(n432), .B(n32951), .Z(n32949) );
  XOR U32053 ( .A(n32952), .B(n32950), .Z(n32951) );
  XNOR U32054 ( .A(n32953), .B(n32954), .Z(n32902) );
  NAND U32055 ( .A(n32955), .B(n32956), .Z(n32954) );
  XOR U32056 ( .A(n32957), .B(n32854), .Z(n32956) );
  XOR U32057 ( .A(n32930), .B(n32931), .Z(n32854) );
  XOR U32058 ( .A(n32958), .B(n32923), .Z(n32931) );
  XOR U32059 ( .A(n32959), .B(n32911), .Z(n32923) );
  XOR U32060 ( .A(n32960), .B(n32961), .Z(n32911) );
  ANDN U32061 ( .B(n32962), .A(n32963), .Z(n32960) );
  XOR U32062 ( .A(n32961), .B(n32964), .Z(n32962) );
  IV U32063 ( .A(n32909), .Z(n32959) );
  XOR U32064 ( .A(n32907), .B(n32965), .Z(n32909) );
  XOR U32065 ( .A(n32966), .B(n32967), .Z(n32965) );
  ANDN U32066 ( .B(n32968), .A(n32969), .Z(n32966) );
  XOR U32067 ( .A(n32970), .B(n32967), .Z(n32968) );
  IV U32068 ( .A(n32910), .Z(n32907) );
  XOR U32069 ( .A(n32971), .B(n32972), .Z(n32910) );
  ANDN U32070 ( .B(n32973), .A(n32974), .Z(n32971) );
  XOR U32071 ( .A(n32972), .B(n32975), .Z(n32973) );
  IV U32072 ( .A(n32922), .Z(n32958) );
  XOR U32073 ( .A(n32976), .B(n32977), .Z(n32922) );
  XNOR U32074 ( .A(n32917), .B(n32978), .Z(n32977) );
  IV U32075 ( .A(n32920), .Z(n32978) );
  XOR U32076 ( .A(n32979), .B(n32980), .Z(n32920) );
  ANDN U32077 ( .B(n32981), .A(n32982), .Z(n32979) );
  XOR U32078 ( .A(n32980), .B(n32983), .Z(n32981) );
  XNOR U32079 ( .A(n32984), .B(n32985), .Z(n32917) );
  ANDN U32080 ( .B(n32986), .A(n32987), .Z(n32984) );
  XOR U32081 ( .A(n32985), .B(n32988), .Z(n32986) );
  IV U32082 ( .A(n32916), .Z(n32976) );
  XOR U32083 ( .A(n32914), .B(n32989), .Z(n32916) );
  XOR U32084 ( .A(n32990), .B(n32991), .Z(n32989) );
  ANDN U32085 ( .B(n32992), .A(n32993), .Z(n32990) );
  XOR U32086 ( .A(n32994), .B(n32991), .Z(n32992) );
  IV U32087 ( .A(n32918), .Z(n32914) );
  XOR U32088 ( .A(n32995), .B(n32996), .Z(n32918) );
  ANDN U32089 ( .B(n32997), .A(n32998), .Z(n32995) );
  XOR U32090 ( .A(n32999), .B(n32996), .Z(n32997) );
  XOR U32091 ( .A(n33000), .B(n33001), .Z(n32930) );
  XOR U32092 ( .A(n32948), .B(n33002), .Z(n33001) );
  IV U32093 ( .A(n32928), .Z(n33002) );
  XOR U32094 ( .A(n33003), .B(n33004), .Z(n32928) );
  ANDN U32095 ( .B(n33005), .A(n33006), .Z(n33003) );
  XOR U32096 ( .A(n33004), .B(n33007), .Z(n33005) );
  XOR U32097 ( .A(n33008), .B(n32936), .Z(n32948) );
  XOR U32098 ( .A(n33009), .B(n33010), .Z(n32936) );
  ANDN U32099 ( .B(n33011), .A(n33012), .Z(n33009) );
  XOR U32100 ( .A(n33010), .B(n33013), .Z(n33011) );
  IV U32101 ( .A(n32935), .Z(n33008) );
  XOR U32102 ( .A(n33014), .B(n33015), .Z(n32935) );
  XOR U32103 ( .A(n33016), .B(n33017), .Z(n33015) );
  ANDN U32104 ( .B(n33018), .A(n33019), .Z(n33016) );
  XOR U32105 ( .A(n33020), .B(n33017), .Z(n33018) );
  IV U32106 ( .A(n32933), .Z(n33014) );
  XOR U32107 ( .A(n33021), .B(n33022), .Z(n32933) );
  ANDN U32108 ( .B(n33023), .A(n33024), .Z(n33021) );
  XOR U32109 ( .A(n33022), .B(n33025), .Z(n33023) );
  IV U32110 ( .A(n32947), .Z(n33000) );
  XOR U32111 ( .A(n33026), .B(n33027), .Z(n32947) );
  XNOR U32112 ( .A(n32942), .B(n33028), .Z(n33027) );
  IV U32113 ( .A(n32945), .Z(n33028) );
  XOR U32114 ( .A(n33029), .B(n33030), .Z(n32945) );
  ANDN U32115 ( .B(n33031), .A(n33032), .Z(n33029) );
  XOR U32116 ( .A(n33033), .B(n33030), .Z(n33031) );
  XNOR U32117 ( .A(n33034), .B(n33035), .Z(n32942) );
  ANDN U32118 ( .B(n33036), .A(n33037), .Z(n33034) );
  XOR U32119 ( .A(n33035), .B(n33038), .Z(n33036) );
  IV U32120 ( .A(n32941), .Z(n33026) );
  XOR U32121 ( .A(n32939), .B(n33039), .Z(n32941) );
  XOR U32122 ( .A(n33040), .B(n33041), .Z(n33039) );
  ANDN U32123 ( .B(n33042), .A(n33043), .Z(n33040) );
  XOR U32124 ( .A(n33044), .B(n33041), .Z(n33042) );
  IV U32125 ( .A(n32943), .Z(n32939) );
  XOR U32126 ( .A(n33045), .B(n33046), .Z(n32943) );
  ANDN U32127 ( .B(n33047), .A(n33048), .Z(n33045) );
  XOR U32128 ( .A(n33049), .B(n33046), .Z(n33047) );
  IV U32129 ( .A(n32953), .Z(n32957) );
  XOR U32130 ( .A(n32953), .B(n32856), .Z(n32955) );
  XOR U32131 ( .A(n33050), .B(n33051), .Z(n32856) );
  AND U32132 ( .A(n432), .B(n33052), .Z(n33050) );
  XOR U32133 ( .A(n33053), .B(n33051), .Z(n33052) );
  NANDN U32134 ( .A(n32858), .B(n32860), .Z(n32953) );
  XOR U32135 ( .A(n33054), .B(n33055), .Z(n32860) );
  AND U32136 ( .A(n432), .B(n33056), .Z(n33054) );
  XOR U32137 ( .A(n33055), .B(n33057), .Z(n33056) );
  XNOR U32138 ( .A(n33058), .B(n33059), .Z(n432) );
  AND U32139 ( .A(n33060), .B(n33061), .Z(n33058) );
  XOR U32140 ( .A(n33059), .B(n32871), .Z(n33061) );
  XNOR U32141 ( .A(n33062), .B(n33063), .Z(n32871) );
  ANDN U32142 ( .B(n33064), .A(n33065), .Z(n33062) );
  XOR U32143 ( .A(n33063), .B(n33066), .Z(n33064) );
  XNOR U32144 ( .A(n33059), .B(n32873), .Z(n33060) );
  XOR U32145 ( .A(n33067), .B(n33068), .Z(n32873) );
  AND U32146 ( .A(n436), .B(n33069), .Z(n33067) );
  XOR U32147 ( .A(n33070), .B(n33068), .Z(n33069) );
  XOR U32148 ( .A(n33071), .B(n33072), .Z(n33059) );
  AND U32149 ( .A(n33073), .B(n33074), .Z(n33071) );
  XOR U32150 ( .A(n33072), .B(n32898), .Z(n33074) );
  XOR U32151 ( .A(n33065), .B(n33066), .Z(n32898) );
  XNOR U32152 ( .A(n33075), .B(n33076), .Z(n33066) );
  ANDN U32153 ( .B(n33077), .A(n33078), .Z(n33075) );
  XOR U32154 ( .A(n33079), .B(n33080), .Z(n33077) );
  XOR U32155 ( .A(n33081), .B(n33082), .Z(n33065) );
  XNOR U32156 ( .A(n33083), .B(n33084), .Z(n33082) );
  ANDN U32157 ( .B(n33085), .A(n33086), .Z(n33083) );
  XNOR U32158 ( .A(n33087), .B(n33088), .Z(n33085) );
  IV U32159 ( .A(n33063), .Z(n33081) );
  XOR U32160 ( .A(n33089), .B(n33090), .Z(n33063) );
  ANDN U32161 ( .B(n33091), .A(n33092), .Z(n33089) );
  XOR U32162 ( .A(n33090), .B(n33093), .Z(n33091) );
  XNOR U32163 ( .A(n33072), .B(n32900), .Z(n33073) );
  XOR U32164 ( .A(n33094), .B(n33095), .Z(n32900) );
  AND U32165 ( .A(n436), .B(n33096), .Z(n33094) );
  XOR U32166 ( .A(n33097), .B(n33095), .Z(n33096) );
  XNOR U32167 ( .A(n33098), .B(n33099), .Z(n33072) );
  AND U32168 ( .A(n33100), .B(n33101), .Z(n33098) );
  XNOR U32169 ( .A(n33099), .B(n32950), .Z(n33101) );
  XOR U32170 ( .A(n33092), .B(n33093), .Z(n32950) );
  XOR U32171 ( .A(n33102), .B(n33080), .Z(n33093) );
  XNOR U32172 ( .A(n33103), .B(n33104), .Z(n33080) );
  ANDN U32173 ( .B(n33105), .A(n33106), .Z(n33103) );
  XOR U32174 ( .A(n33107), .B(n33108), .Z(n33105) );
  IV U32175 ( .A(n33078), .Z(n33102) );
  XOR U32176 ( .A(n33076), .B(n33109), .Z(n33078) );
  XNOR U32177 ( .A(n33110), .B(n33111), .Z(n33109) );
  ANDN U32178 ( .B(n33112), .A(n33113), .Z(n33110) );
  XNOR U32179 ( .A(n33114), .B(n33115), .Z(n33112) );
  IV U32180 ( .A(n33079), .Z(n33076) );
  XOR U32181 ( .A(n33116), .B(n33117), .Z(n33079) );
  ANDN U32182 ( .B(n33118), .A(n33119), .Z(n33116) );
  XOR U32183 ( .A(n33117), .B(n33120), .Z(n33118) );
  XOR U32184 ( .A(n33121), .B(n33122), .Z(n33092) );
  XNOR U32185 ( .A(n33087), .B(n33123), .Z(n33122) );
  IV U32186 ( .A(n33090), .Z(n33123) );
  XOR U32187 ( .A(n33124), .B(n33125), .Z(n33090) );
  ANDN U32188 ( .B(n33126), .A(n33127), .Z(n33124) );
  XOR U32189 ( .A(n33125), .B(n33128), .Z(n33126) );
  XNOR U32190 ( .A(n33129), .B(n33130), .Z(n33087) );
  ANDN U32191 ( .B(n33131), .A(n33132), .Z(n33129) );
  XOR U32192 ( .A(n33130), .B(n33133), .Z(n33131) );
  IV U32193 ( .A(n33086), .Z(n33121) );
  XOR U32194 ( .A(n33084), .B(n33134), .Z(n33086) );
  XNOR U32195 ( .A(n33135), .B(n33136), .Z(n33134) );
  ANDN U32196 ( .B(n33137), .A(n33138), .Z(n33135) );
  XNOR U32197 ( .A(n33139), .B(n33140), .Z(n33137) );
  IV U32198 ( .A(n33088), .Z(n33084) );
  XOR U32199 ( .A(n33141), .B(n33142), .Z(n33088) );
  ANDN U32200 ( .B(n33143), .A(n33144), .Z(n33141) );
  XOR U32201 ( .A(n33145), .B(n33142), .Z(n33143) );
  XOR U32202 ( .A(n33099), .B(n32952), .Z(n33100) );
  XOR U32203 ( .A(n33146), .B(n33147), .Z(n32952) );
  AND U32204 ( .A(n436), .B(n33148), .Z(n33146) );
  XOR U32205 ( .A(n33149), .B(n33147), .Z(n33148) );
  XNOR U32206 ( .A(n33150), .B(n33151), .Z(n33099) );
  NAND U32207 ( .A(n33152), .B(n33153), .Z(n33151) );
  XOR U32208 ( .A(n33154), .B(n33051), .Z(n33153) );
  XOR U32209 ( .A(n33127), .B(n33128), .Z(n33051) );
  XOR U32210 ( .A(n33155), .B(n33120), .Z(n33128) );
  XOR U32211 ( .A(n33156), .B(n33108), .Z(n33120) );
  XOR U32212 ( .A(n33157), .B(n33158), .Z(n33108) );
  ANDN U32213 ( .B(n33159), .A(n33160), .Z(n33157) );
  XOR U32214 ( .A(n33158), .B(n33161), .Z(n33159) );
  IV U32215 ( .A(n33106), .Z(n33156) );
  XOR U32216 ( .A(n33104), .B(n33162), .Z(n33106) );
  XOR U32217 ( .A(n33163), .B(n33164), .Z(n33162) );
  ANDN U32218 ( .B(n33165), .A(n33166), .Z(n33163) );
  XOR U32219 ( .A(n33167), .B(n33164), .Z(n33165) );
  IV U32220 ( .A(n33107), .Z(n33104) );
  XOR U32221 ( .A(n33168), .B(n33169), .Z(n33107) );
  ANDN U32222 ( .B(n33170), .A(n33171), .Z(n33168) );
  XOR U32223 ( .A(n33169), .B(n33172), .Z(n33170) );
  IV U32224 ( .A(n33119), .Z(n33155) );
  XOR U32225 ( .A(n33173), .B(n33174), .Z(n33119) );
  XNOR U32226 ( .A(n33114), .B(n33175), .Z(n33174) );
  IV U32227 ( .A(n33117), .Z(n33175) );
  XOR U32228 ( .A(n33176), .B(n33177), .Z(n33117) );
  ANDN U32229 ( .B(n33178), .A(n33179), .Z(n33176) );
  XOR U32230 ( .A(n33177), .B(n33180), .Z(n33178) );
  XNOR U32231 ( .A(n33181), .B(n33182), .Z(n33114) );
  ANDN U32232 ( .B(n33183), .A(n33184), .Z(n33181) );
  XOR U32233 ( .A(n33182), .B(n33185), .Z(n33183) );
  IV U32234 ( .A(n33113), .Z(n33173) );
  XOR U32235 ( .A(n33111), .B(n33186), .Z(n33113) );
  XOR U32236 ( .A(n33187), .B(n33188), .Z(n33186) );
  ANDN U32237 ( .B(n33189), .A(n33190), .Z(n33187) );
  XOR U32238 ( .A(n33191), .B(n33188), .Z(n33189) );
  IV U32239 ( .A(n33115), .Z(n33111) );
  XOR U32240 ( .A(n33192), .B(n33193), .Z(n33115) );
  ANDN U32241 ( .B(n33194), .A(n33195), .Z(n33192) );
  XOR U32242 ( .A(n33196), .B(n33193), .Z(n33194) );
  XOR U32243 ( .A(n33197), .B(n33198), .Z(n33127) );
  XOR U32244 ( .A(n33145), .B(n33199), .Z(n33198) );
  IV U32245 ( .A(n33125), .Z(n33199) );
  XOR U32246 ( .A(n33200), .B(n33201), .Z(n33125) );
  ANDN U32247 ( .B(n33202), .A(n33203), .Z(n33200) );
  XOR U32248 ( .A(n33201), .B(n33204), .Z(n33202) );
  XOR U32249 ( .A(n33205), .B(n33133), .Z(n33145) );
  XOR U32250 ( .A(n33206), .B(n33207), .Z(n33133) );
  ANDN U32251 ( .B(n33208), .A(n33209), .Z(n33206) );
  XOR U32252 ( .A(n33207), .B(n33210), .Z(n33208) );
  IV U32253 ( .A(n33132), .Z(n33205) );
  XOR U32254 ( .A(n33211), .B(n33212), .Z(n33132) );
  XOR U32255 ( .A(n33213), .B(n33214), .Z(n33212) );
  ANDN U32256 ( .B(n33215), .A(n33216), .Z(n33213) );
  XOR U32257 ( .A(n33217), .B(n33214), .Z(n33215) );
  IV U32258 ( .A(n33130), .Z(n33211) );
  XOR U32259 ( .A(n33218), .B(n33219), .Z(n33130) );
  ANDN U32260 ( .B(n33220), .A(n33221), .Z(n33218) );
  XOR U32261 ( .A(n33219), .B(n33222), .Z(n33220) );
  IV U32262 ( .A(n33144), .Z(n33197) );
  XOR U32263 ( .A(n33223), .B(n33224), .Z(n33144) );
  XNOR U32264 ( .A(n33139), .B(n33225), .Z(n33224) );
  IV U32265 ( .A(n33142), .Z(n33225) );
  XOR U32266 ( .A(n33226), .B(n33227), .Z(n33142) );
  ANDN U32267 ( .B(n33228), .A(n33229), .Z(n33226) );
  XOR U32268 ( .A(n33230), .B(n33227), .Z(n33228) );
  XNOR U32269 ( .A(n33231), .B(n33232), .Z(n33139) );
  ANDN U32270 ( .B(n33233), .A(n33234), .Z(n33231) );
  XOR U32271 ( .A(n33232), .B(n33235), .Z(n33233) );
  IV U32272 ( .A(n33138), .Z(n33223) );
  XOR U32273 ( .A(n33136), .B(n33236), .Z(n33138) );
  XOR U32274 ( .A(n33237), .B(n33238), .Z(n33236) );
  ANDN U32275 ( .B(n33239), .A(n33240), .Z(n33237) );
  XOR U32276 ( .A(n33241), .B(n33238), .Z(n33239) );
  IV U32277 ( .A(n33140), .Z(n33136) );
  XOR U32278 ( .A(n33242), .B(n33243), .Z(n33140) );
  ANDN U32279 ( .B(n33244), .A(n33245), .Z(n33242) );
  XOR U32280 ( .A(n33246), .B(n33243), .Z(n33244) );
  IV U32281 ( .A(n33150), .Z(n33154) );
  XOR U32282 ( .A(n33150), .B(n33053), .Z(n33152) );
  XOR U32283 ( .A(n33247), .B(n33248), .Z(n33053) );
  AND U32284 ( .A(n436), .B(n33249), .Z(n33247) );
  XOR U32285 ( .A(n33250), .B(n33248), .Z(n33249) );
  NANDN U32286 ( .A(n33055), .B(n33057), .Z(n33150) );
  XOR U32287 ( .A(n33251), .B(n33252), .Z(n33057) );
  AND U32288 ( .A(n436), .B(n33253), .Z(n33251) );
  XOR U32289 ( .A(n33252), .B(n33254), .Z(n33253) );
  XNOR U32290 ( .A(n33255), .B(n33256), .Z(n436) );
  AND U32291 ( .A(n33257), .B(n33258), .Z(n33255) );
  XOR U32292 ( .A(n33256), .B(n33068), .Z(n33258) );
  XNOR U32293 ( .A(n33259), .B(n33260), .Z(n33068) );
  ANDN U32294 ( .B(n33261), .A(n33262), .Z(n33259) );
  XOR U32295 ( .A(n33260), .B(n33263), .Z(n33261) );
  XNOR U32296 ( .A(n33256), .B(n33070), .Z(n33257) );
  XOR U32297 ( .A(n33264), .B(n33265), .Z(n33070) );
  AND U32298 ( .A(n440), .B(n33266), .Z(n33264) );
  XOR U32299 ( .A(n33267), .B(n33265), .Z(n33266) );
  XOR U32300 ( .A(n33268), .B(n33269), .Z(n33256) );
  AND U32301 ( .A(n33270), .B(n33271), .Z(n33268) );
  XOR U32302 ( .A(n33269), .B(n33095), .Z(n33271) );
  XOR U32303 ( .A(n33262), .B(n33263), .Z(n33095) );
  XNOR U32304 ( .A(n33272), .B(n33273), .Z(n33263) );
  ANDN U32305 ( .B(n33274), .A(n33275), .Z(n33272) );
  XOR U32306 ( .A(n33276), .B(n33277), .Z(n33274) );
  XOR U32307 ( .A(n33278), .B(n33279), .Z(n33262) );
  XNOR U32308 ( .A(n33280), .B(n33281), .Z(n33279) );
  ANDN U32309 ( .B(n33282), .A(n33283), .Z(n33280) );
  XNOR U32310 ( .A(n33284), .B(n33285), .Z(n33282) );
  IV U32311 ( .A(n33260), .Z(n33278) );
  XOR U32312 ( .A(n33286), .B(n33287), .Z(n33260) );
  ANDN U32313 ( .B(n33288), .A(n33289), .Z(n33286) );
  XOR U32314 ( .A(n33287), .B(n33290), .Z(n33288) );
  XNOR U32315 ( .A(n33269), .B(n33097), .Z(n33270) );
  XOR U32316 ( .A(n33291), .B(n33292), .Z(n33097) );
  AND U32317 ( .A(n440), .B(n33293), .Z(n33291) );
  XOR U32318 ( .A(n33294), .B(n33292), .Z(n33293) );
  XNOR U32319 ( .A(n33295), .B(n33296), .Z(n33269) );
  AND U32320 ( .A(n33297), .B(n33298), .Z(n33295) );
  XNOR U32321 ( .A(n33296), .B(n33147), .Z(n33298) );
  XOR U32322 ( .A(n33289), .B(n33290), .Z(n33147) );
  XOR U32323 ( .A(n33299), .B(n33277), .Z(n33290) );
  XNOR U32324 ( .A(n33300), .B(n33301), .Z(n33277) );
  ANDN U32325 ( .B(n33302), .A(n33303), .Z(n33300) );
  XOR U32326 ( .A(n33304), .B(n33305), .Z(n33302) );
  IV U32327 ( .A(n33275), .Z(n33299) );
  XOR U32328 ( .A(n33273), .B(n33306), .Z(n33275) );
  XNOR U32329 ( .A(n33307), .B(n33308), .Z(n33306) );
  ANDN U32330 ( .B(n33309), .A(n33310), .Z(n33307) );
  XNOR U32331 ( .A(n33311), .B(n33312), .Z(n33309) );
  IV U32332 ( .A(n33276), .Z(n33273) );
  XOR U32333 ( .A(n33313), .B(n33314), .Z(n33276) );
  ANDN U32334 ( .B(n33315), .A(n33316), .Z(n33313) );
  XOR U32335 ( .A(n33314), .B(n33317), .Z(n33315) );
  XOR U32336 ( .A(n33318), .B(n33319), .Z(n33289) );
  XNOR U32337 ( .A(n33284), .B(n33320), .Z(n33319) );
  IV U32338 ( .A(n33287), .Z(n33320) );
  XOR U32339 ( .A(n33321), .B(n33322), .Z(n33287) );
  ANDN U32340 ( .B(n33323), .A(n33324), .Z(n33321) );
  XOR U32341 ( .A(n33322), .B(n33325), .Z(n33323) );
  XNOR U32342 ( .A(n33326), .B(n33327), .Z(n33284) );
  ANDN U32343 ( .B(n33328), .A(n33329), .Z(n33326) );
  XOR U32344 ( .A(n33327), .B(n33330), .Z(n33328) );
  IV U32345 ( .A(n33283), .Z(n33318) );
  XOR U32346 ( .A(n33281), .B(n33331), .Z(n33283) );
  XNOR U32347 ( .A(n33332), .B(n33333), .Z(n33331) );
  ANDN U32348 ( .B(n33334), .A(n33335), .Z(n33332) );
  XNOR U32349 ( .A(n33336), .B(n33337), .Z(n33334) );
  IV U32350 ( .A(n33285), .Z(n33281) );
  XOR U32351 ( .A(n33338), .B(n33339), .Z(n33285) );
  ANDN U32352 ( .B(n33340), .A(n33341), .Z(n33338) );
  XOR U32353 ( .A(n33342), .B(n33339), .Z(n33340) );
  XOR U32354 ( .A(n33296), .B(n33149), .Z(n33297) );
  XOR U32355 ( .A(n33343), .B(n33344), .Z(n33149) );
  AND U32356 ( .A(n440), .B(n33345), .Z(n33343) );
  XOR U32357 ( .A(n33346), .B(n33344), .Z(n33345) );
  XNOR U32358 ( .A(n33347), .B(n33348), .Z(n33296) );
  NAND U32359 ( .A(n33349), .B(n33350), .Z(n33348) );
  XOR U32360 ( .A(n33351), .B(n33248), .Z(n33350) );
  XOR U32361 ( .A(n33324), .B(n33325), .Z(n33248) );
  XOR U32362 ( .A(n33352), .B(n33317), .Z(n33325) );
  XOR U32363 ( .A(n33353), .B(n33305), .Z(n33317) );
  XOR U32364 ( .A(n33354), .B(n33355), .Z(n33305) );
  ANDN U32365 ( .B(n33356), .A(n33357), .Z(n33354) );
  XOR U32366 ( .A(n33355), .B(n33358), .Z(n33356) );
  IV U32367 ( .A(n33303), .Z(n33353) );
  XOR U32368 ( .A(n33301), .B(n33359), .Z(n33303) );
  XOR U32369 ( .A(n33360), .B(n33361), .Z(n33359) );
  ANDN U32370 ( .B(n33362), .A(n33363), .Z(n33360) );
  XOR U32371 ( .A(n33364), .B(n33361), .Z(n33362) );
  IV U32372 ( .A(n33304), .Z(n33301) );
  XOR U32373 ( .A(n33365), .B(n33366), .Z(n33304) );
  ANDN U32374 ( .B(n33367), .A(n33368), .Z(n33365) );
  XOR U32375 ( .A(n33366), .B(n33369), .Z(n33367) );
  IV U32376 ( .A(n33316), .Z(n33352) );
  XOR U32377 ( .A(n33370), .B(n33371), .Z(n33316) );
  XNOR U32378 ( .A(n33311), .B(n33372), .Z(n33371) );
  IV U32379 ( .A(n33314), .Z(n33372) );
  XOR U32380 ( .A(n33373), .B(n33374), .Z(n33314) );
  ANDN U32381 ( .B(n33375), .A(n33376), .Z(n33373) );
  XOR U32382 ( .A(n33374), .B(n33377), .Z(n33375) );
  XNOR U32383 ( .A(n33378), .B(n33379), .Z(n33311) );
  ANDN U32384 ( .B(n33380), .A(n33381), .Z(n33378) );
  XOR U32385 ( .A(n33379), .B(n33382), .Z(n33380) );
  IV U32386 ( .A(n33310), .Z(n33370) );
  XOR U32387 ( .A(n33308), .B(n33383), .Z(n33310) );
  XOR U32388 ( .A(n33384), .B(n33385), .Z(n33383) );
  ANDN U32389 ( .B(n33386), .A(n33387), .Z(n33384) );
  XOR U32390 ( .A(n33388), .B(n33385), .Z(n33386) );
  IV U32391 ( .A(n33312), .Z(n33308) );
  XOR U32392 ( .A(n33389), .B(n33390), .Z(n33312) );
  ANDN U32393 ( .B(n33391), .A(n33392), .Z(n33389) );
  XOR U32394 ( .A(n33393), .B(n33390), .Z(n33391) );
  XOR U32395 ( .A(n33394), .B(n33395), .Z(n33324) );
  XOR U32396 ( .A(n33342), .B(n33396), .Z(n33395) );
  IV U32397 ( .A(n33322), .Z(n33396) );
  XOR U32398 ( .A(n33397), .B(n33398), .Z(n33322) );
  ANDN U32399 ( .B(n33399), .A(n33400), .Z(n33397) );
  XOR U32400 ( .A(n33398), .B(n33401), .Z(n33399) );
  XOR U32401 ( .A(n33402), .B(n33330), .Z(n33342) );
  XOR U32402 ( .A(n33403), .B(n33404), .Z(n33330) );
  ANDN U32403 ( .B(n33405), .A(n33406), .Z(n33403) );
  XOR U32404 ( .A(n33404), .B(n33407), .Z(n33405) );
  IV U32405 ( .A(n33329), .Z(n33402) );
  XOR U32406 ( .A(n33408), .B(n33409), .Z(n33329) );
  XOR U32407 ( .A(n33410), .B(n33411), .Z(n33409) );
  ANDN U32408 ( .B(n33412), .A(n33413), .Z(n33410) );
  XOR U32409 ( .A(n33414), .B(n33411), .Z(n33412) );
  IV U32410 ( .A(n33327), .Z(n33408) );
  XOR U32411 ( .A(n33415), .B(n33416), .Z(n33327) );
  ANDN U32412 ( .B(n33417), .A(n33418), .Z(n33415) );
  XOR U32413 ( .A(n33416), .B(n33419), .Z(n33417) );
  IV U32414 ( .A(n33341), .Z(n33394) );
  XOR U32415 ( .A(n33420), .B(n33421), .Z(n33341) );
  XNOR U32416 ( .A(n33336), .B(n33422), .Z(n33421) );
  IV U32417 ( .A(n33339), .Z(n33422) );
  XOR U32418 ( .A(n33423), .B(n33424), .Z(n33339) );
  ANDN U32419 ( .B(n33425), .A(n33426), .Z(n33423) );
  XOR U32420 ( .A(n33427), .B(n33424), .Z(n33425) );
  XNOR U32421 ( .A(n33428), .B(n33429), .Z(n33336) );
  ANDN U32422 ( .B(n33430), .A(n33431), .Z(n33428) );
  XOR U32423 ( .A(n33429), .B(n33432), .Z(n33430) );
  IV U32424 ( .A(n33335), .Z(n33420) );
  XOR U32425 ( .A(n33333), .B(n33433), .Z(n33335) );
  XOR U32426 ( .A(n33434), .B(n33435), .Z(n33433) );
  ANDN U32427 ( .B(n33436), .A(n33437), .Z(n33434) );
  XOR U32428 ( .A(n33438), .B(n33435), .Z(n33436) );
  IV U32429 ( .A(n33337), .Z(n33333) );
  XOR U32430 ( .A(n33439), .B(n33440), .Z(n33337) );
  ANDN U32431 ( .B(n33441), .A(n33442), .Z(n33439) );
  XOR U32432 ( .A(n33443), .B(n33440), .Z(n33441) );
  IV U32433 ( .A(n33347), .Z(n33351) );
  XOR U32434 ( .A(n33347), .B(n33250), .Z(n33349) );
  XOR U32435 ( .A(n33444), .B(n33445), .Z(n33250) );
  AND U32436 ( .A(n440), .B(n33446), .Z(n33444) );
  XOR U32437 ( .A(n33447), .B(n33445), .Z(n33446) );
  NANDN U32438 ( .A(n33252), .B(n33254), .Z(n33347) );
  XOR U32439 ( .A(n33448), .B(n33449), .Z(n33254) );
  AND U32440 ( .A(n440), .B(n33450), .Z(n33448) );
  XOR U32441 ( .A(n33449), .B(n33451), .Z(n33450) );
  XNOR U32442 ( .A(n33452), .B(n33453), .Z(n440) );
  AND U32443 ( .A(n33454), .B(n33455), .Z(n33452) );
  XOR U32444 ( .A(n33453), .B(n33265), .Z(n33455) );
  XNOR U32445 ( .A(n33456), .B(n33457), .Z(n33265) );
  ANDN U32446 ( .B(n33458), .A(n33459), .Z(n33456) );
  XOR U32447 ( .A(n33457), .B(n33460), .Z(n33458) );
  XNOR U32448 ( .A(n33453), .B(n33267), .Z(n33454) );
  XOR U32449 ( .A(n33461), .B(n33462), .Z(n33267) );
  AND U32450 ( .A(n444), .B(n33463), .Z(n33461) );
  XOR U32451 ( .A(n33464), .B(n33462), .Z(n33463) );
  XOR U32452 ( .A(n33465), .B(n33466), .Z(n33453) );
  AND U32453 ( .A(n33467), .B(n33468), .Z(n33465) );
  XOR U32454 ( .A(n33466), .B(n33292), .Z(n33468) );
  XOR U32455 ( .A(n33459), .B(n33460), .Z(n33292) );
  XNOR U32456 ( .A(n33469), .B(n33470), .Z(n33460) );
  ANDN U32457 ( .B(n33471), .A(n33472), .Z(n33469) );
  XOR U32458 ( .A(n33473), .B(n33474), .Z(n33471) );
  XOR U32459 ( .A(n33475), .B(n33476), .Z(n33459) );
  XNOR U32460 ( .A(n33477), .B(n33478), .Z(n33476) );
  ANDN U32461 ( .B(n33479), .A(n33480), .Z(n33477) );
  XNOR U32462 ( .A(n33481), .B(n33482), .Z(n33479) );
  IV U32463 ( .A(n33457), .Z(n33475) );
  XOR U32464 ( .A(n33483), .B(n33484), .Z(n33457) );
  ANDN U32465 ( .B(n33485), .A(n33486), .Z(n33483) );
  XOR U32466 ( .A(n33484), .B(n33487), .Z(n33485) );
  XNOR U32467 ( .A(n33466), .B(n33294), .Z(n33467) );
  XOR U32468 ( .A(n33488), .B(n33489), .Z(n33294) );
  AND U32469 ( .A(n444), .B(n33490), .Z(n33488) );
  XOR U32470 ( .A(n33491), .B(n33489), .Z(n33490) );
  XNOR U32471 ( .A(n33492), .B(n33493), .Z(n33466) );
  AND U32472 ( .A(n33494), .B(n33495), .Z(n33492) );
  XNOR U32473 ( .A(n33493), .B(n33344), .Z(n33495) );
  XOR U32474 ( .A(n33486), .B(n33487), .Z(n33344) );
  XOR U32475 ( .A(n33496), .B(n33474), .Z(n33487) );
  XNOR U32476 ( .A(n33497), .B(n33498), .Z(n33474) );
  ANDN U32477 ( .B(n33499), .A(n33500), .Z(n33497) );
  XOR U32478 ( .A(n33501), .B(n33502), .Z(n33499) );
  IV U32479 ( .A(n33472), .Z(n33496) );
  XOR U32480 ( .A(n33470), .B(n33503), .Z(n33472) );
  XNOR U32481 ( .A(n33504), .B(n33505), .Z(n33503) );
  ANDN U32482 ( .B(n33506), .A(n33507), .Z(n33504) );
  XNOR U32483 ( .A(n33508), .B(n33509), .Z(n33506) );
  IV U32484 ( .A(n33473), .Z(n33470) );
  XOR U32485 ( .A(n33510), .B(n33511), .Z(n33473) );
  ANDN U32486 ( .B(n33512), .A(n33513), .Z(n33510) );
  XOR U32487 ( .A(n33511), .B(n33514), .Z(n33512) );
  XOR U32488 ( .A(n33515), .B(n33516), .Z(n33486) );
  XNOR U32489 ( .A(n33481), .B(n33517), .Z(n33516) );
  IV U32490 ( .A(n33484), .Z(n33517) );
  XOR U32491 ( .A(n33518), .B(n33519), .Z(n33484) );
  ANDN U32492 ( .B(n33520), .A(n33521), .Z(n33518) );
  XOR U32493 ( .A(n33519), .B(n33522), .Z(n33520) );
  XNOR U32494 ( .A(n33523), .B(n33524), .Z(n33481) );
  ANDN U32495 ( .B(n33525), .A(n33526), .Z(n33523) );
  XOR U32496 ( .A(n33524), .B(n33527), .Z(n33525) );
  IV U32497 ( .A(n33480), .Z(n33515) );
  XOR U32498 ( .A(n33478), .B(n33528), .Z(n33480) );
  XNOR U32499 ( .A(n33529), .B(n33530), .Z(n33528) );
  ANDN U32500 ( .B(n33531), .A(n33532), .Z(n33529) );
  XNOR U32501 ( .A(n33533), .B(n33534), .Z(n33531) );
  IV U32502 ( .A(n33482), .Z(n33478) );
  XOR U32503 ( .A(n33535), .B(n33536), .Z(n33482) );
  ANDN U32504 ( .B(n33537), .A(n33538), .Z(n33535) );
  XOR U32505 ( .A(n33539), .B(n33536), .Z(n33537) );
  XOR U32506 ( .A(n33493), .B(n33346), .Z(n33494) );
  XOR U32507 ( .A(n33540), .B(n33541), .Z(n33346) );
  AND U32508 ( .A(n444), .B(n33542), .Z(n33540) );
  XOR U32509 ( .A(n33543), .B(n33541), .Z(n33542) );
  XNOR U32510 ( .A(n33544), .B(n33545), .Z(n33493) );
  NAND U32511 ( .A(n33546), .B(n33547), .Z(n33545) );
  XOR U32512 ( .A(n33548), .B(n33445), .Z(n33547) );
  XOR U32513 ( .A(n33521), .B(n33522), .Z(n33445) );
  XOR U32514 ( .A(n33549), .B(n33514), .Z(n33522) );
  XOR U32515 ( .A(n33550), .B(n33502), .Z(n33514) );
  XOR U32516 ( .A(n33551), .B(n33552), .Z(n33502) );
  ANDN U32517 ( .B(n33553), .A(n33554), .Z(n33551) );
  XOR U32518 ( .A(n33552), .B(n33555), .Z(n33553) );
  IV U32519 ( .A(n33500), .Z(n33550) );
  XOR U32520 ( .A(n33498), .B(n33556), .Z(n33500) );
  XOR U32521 ( .A(n33557), .B(n33558), .Z(n33556) );
  ANDN U32522 ( .B(n33559), .A(n33560), .Z(n33557) );
  XOR U32523 ( .A(n33561), .B(n33558), .Z(n33559) );
  IV U32524 ( .A(n33501), .Z(n33498) );
  XOR U32525 ( .A(n33562), .B(n33563), .Z(n33501) );
  ANDN U32526 ( .B(n33564), .A(n33565), .Z(n33562) );
  XOR U32527 ( .A(n33563), .B(n33566), .Z(n33564) );
  IV U32528 ( .A(n33513), .Z(n33549) );
  XOR U32529 ( .A(n33567), .B(n33568), .Z(n33513) );
  XNOR U32530 ( .A(n33508), .B(n33569), .Z(n33568) );
  IV U32531 ( .A(n33511), .Z(n33569) );
  XOR U32532 ( .A(n33570), .B(n33571), .Z(n33511) );
  ANDN U32533 ( .B(n33572), .A(n33573), .Z(n33570) );
  XOR U32534 ( .A(n33571), .B(n33574), .Z(n33572) );
  XNOR U32535 ( .A(n33575), .B(n33576), .Z(n33508) );
  ANDN U32536 ( .B(n33577), .A(n33578), .Z(n33575) );
  XOR U32537 ( .A(n33576), .B(n33579), .Z(n33577) );
  IV U32538 ( .A(n33507), .Z(n33567) );
  XOR U32539 ( .A(n33505), .B(n33580), .Z(n33507) );
  XOR U32540 ( .A(n33581), .B(n33582), .Z(n33580) );
  ANDN U32541 ( .B(n33583), .A(n33584), .Z(n33581) );
  XOR U32542 ( .A(n33585), .B(n33582), .Z(n33583) );
  IV U32543 ( .A(n33509), .Z(n33505) );
  XOR U32544 ( .A(n33586), .B(n33587), .Z(n33509) );
  ANDN U32545 ( .B(n33588), .A(n33589), .Z(n33586) );
  XOR U32546 ( .A(n33590), .B(n33587), .Z(n33588) );
  XOR U32547 ( .A(n33591), .B(n33592), .Z(n33521) );
  XOR U32548 ( .A(n33539), .B(n33593), .Z(n33592) );
  IV U32549 ( .A(n33519), .Z(n33593) );
  XOR U32550 ( .A(n33594), .B(n33595), .Z(n33519) );
  ANDN U32551 ( .B(n33596), .A(n33597), .Z(n33594) );
  XOR U32552 ( .A(n33595), .B(n33598), .Z(n33596) );
  XOR U32553 ( .A(n33599), .B(n33527), .Z(n33539) );
  XOR U32554 ( .A(n33600), .B(n33601), .Z(n33527) );
  ANDN U32555 ( .B(n33602), .A(n33603), .Z(n33600) );
  XOR U32556 ( .A(n33601), .B(n33604), .Z(n33602) );
  IV U32557 ( .A(n33526), .Z(n33599) );
  XOR U32558 ( .A(n33605), .B(n33606), .Z(n33526) );
  XOR U32559 ( .A(n33607), .B(n33608), .Z(n33606) );
  ANDN U32560 ( .B(n33609), .A(n33610), .Z(n33607) );
  XOR U32561 ( .A(n33611), .B(n33608), .Z(n33609) );
  IV U32562 ( .A(n33524), .Z(n33605) );
  XOR U32563 ( .A(n33612), .B(n33613), .Z(n33524) );
  ANDN U32564 ( .B(n33614), .A(n33615), .Z(n33612) );
  XOR U32565 ( .A(n33613), .B(n33616), .Z(n33614) );
  IV U32566 ( .A(n33538), .Z(n33591) );
  XOR U32567 ( .A(n33617), .B(n33618), .Z(n33538) );
  XNOR U32568 ( .A(n33533), .B(n33619), .Z(n33618) );
  IV U32569 ( .A(n33536), .Z(n33619) );
  XOR U32570 ( .A(n33620), .B(n33621), .Z(n33536) );
  ANDN U32571 ( .B(n33622), .A(n33623), .Z(n33620) );
  XOR U32572 ( .A(n33624), .B(n33621), .Z(n33622) );
  XNOR U32573 ( .A(n33625), .B(n33626), .Z(n33533) );
  ANDN U32574 ( .B(n33627), .A(n33628), .Z(n33625) );
  XOR U32575 ( .A(n33626), .B(n33629), .Z(n33627) );
  IV U32576 ( .A(n33532), .Z(n33617) );
  XOR U32577 ( .A(n33530), .B(n33630), .Z(n33532) );
  XOR U32578 ( .A(n33631), .B(n33632), .Z(n33630) );
  ANDN U32579 ( .B(n33633), .A(n33634), .Z(n33631) );
  XOR U32580 ( .A(n33635), .B(n33632), .Z(n33633) );
  IV U32581 ( .A(n33534), .Z(n33530) );
  XOR U32582 ( .A(n33636), .B(n33637), .Z(n33534) );
  ANDN U32583 ( .B(n33638), .A(n33639), .Z(n33636) );
  XOR U32584 ( .A(n33640), .B(n33637), .Z(n33638) );
  IV U32585 ( .A(n33544), .Z(n33548) );
  XOR U32586 ( .A(n33544), .B(n33447), .Z(n33546) );
  XOR U32587 ( .A(n33641), .B(n33642), .Z(n33447) );
  AND U32588 ( .A(n444), .B(n33643), .Z(n33641) );
  XOR U32589 ( .A(n33644), .B(n33642), .Z(n33643) );
  NANDN U32590 ( .A(n33449), .B(n33451), .Z(n33544) );
  XOR U32591 ( .A(n33645), .B(n33646), .Z(n33451) );
  AND U32592 ( .A(n444), .B(n33647), .Z(n33645) );
  XOR U32593 ( .A(n33646), .B(n33648), .Z(n33647) );
  XNOR U32594 ( .A(n33649), .B(n33650), .Z(n444) );
  AND U32595 ( .A(n33651), .B(n33652), .Z(n33649) );
  XOR U32596 ( .A(n33650), .B(n33462), .Z(n33652) );
  XNOR U32597 ( .A(n33653), .B(n33654), .Z(n33462) );
  ANDN U32598 ( .B(n33655), .A(n33656), .Z(n33653) );
  XOR U32599 ( .A(n33654), .B(n33657), .Z(n33655) );
  XNOR U32600 ( .A(n33650), .B(n33464), .Z(n33651) );
  XOR U32601 ( .A(n33658), .B(n33659), .Z(n33464) );
  AND U32602 ( .A(n448), .B(n33660), .Z(n33658) );
  XOR U32603 ( .A(n33661), .B(n33659), .Z(n33660) );
  XOR U32604 ( .A(n33662), .B(n33663), .Z(n33650) );
  AND U32605 ( .A(n33664), .B(n33665), .Z(n33662) );
  XOR U32606 ( .A(n33663), .B(n33489), .Z(n33665) );
  XOR U32607 ( .A(n33656), .B(n33657), .Z(n33489) );
  XNOR U32608 ( .A(n33666), .B(n33667), .Z(n33657) );
  ANDN U32609 ( .B(n33668), .A(n33669), .Z(n33666) );
  XOR U32610 ( .A(n33670), .B(n33671), .Z(n33668) );
  XOR U32611 ( .A(n33672), .B(n33673), .Z(n33656) );
  XNOR U32612 ( .A(n33674), .B(n33675), .Z(n33673) );
  ANDN U32613 ( .B(n33676), .A(n33677), .Z(n33674) );
  XNOR U32614 ( .A(n33678), .B(n33679), .Z(n33676) );
  IV U32615 ( .A(n33654), .Z(n33672) );
  XOR U32616 ( .A(n33680), .B(n33681), .Z(n33654) );
  ANDN U32617 ( .B(n33682), .A(n33683), .Z(n33680) );
  XOR U32618 ( .A(n33681), .B(n33684), .Z(n33682) );
  XNOR U32619 ( .A(n33663), .B(n33491), .Z(n33664) );
  XOR U32620 ( .A(n33685), .B(n33686), .Z(n33491) );
  AND U32621 ( .A(n448), .B(n33687), .Z(n33685) );
  XOR U32622 ( .A(n33688), .B(n33686), .Z(n33687) );
  XNOR U32623 ( .A(n33689), .B(n33690), .Z(n33663) );
  AND U32624 ( .A(n33691), .B(n33692), .Z(n33689) );
  XNOR U32625 ( .A(n33690), .B(n33541), .Z(n33692) );
  XOR U32626 ( .A(n33683), .B(n33684), .Z(n33541) );
  XOR U32627 ( .A(n33693), .B(n33671), .Z(n33684) );
  XNOR U32628 ( .A(n33694), .B(n33695), .Z(n33671) );
  ANDN U32629 ( .B(n33696), .A(n33697), .Z(n33694) );
  XOR U32630 ( .A(n33698), .B(n33699), .Z(n33696) );
  IV U32631 ( .A(n33669), .Z(n33693) );
  XOR U32632 ( .A(n33667), .B(n33700), .Z(n33669) );
  XNOR U32633 ( .A(n33701), .B(n33702), .Z(n33700) );
  ANDN U32634 ( .B(n33703), .A(n33704), .Z(n33701) );
  XNOR U32635 ( .A(n33705), .B(n33706), .Z(n33703) );
  IV U32636 ( .A(n33670), .Z(n33667) );
  XOR U32637 ( .A(n33707), .B(n33708), .Z(n33670) );
  ANDN U32638 ( .B(n33709), .A(n33710), .Z(n33707) );
  XOR U32639 ( .A(n33708), .B(n33711), .Z(n33709) );
  XOR U32640 ( .A(n33712), .B(n33713), .Z(n33683) );
  XNOR U32641 ( .A(n33678), .B(n33714), .Z(n33713) );
  IV U32642 ( .A(n33681), .Z(n33714) );
  XOR U32643 ( .A(n33715), .B(n33716), .Z(n33681) );
  ANDN U32644 ( .B(n33717), .A(n33718), .Z(n33715) );
  XOR U32645 ( .A(n33716), .B(n33719), .Z(n33717) );
  XNOR U32646 ( .A(n33720), .B(n33721), .Z(n33678) );
  ANDN U32647 ( .B(n33722), .A(n33723), .Z(n33720) );
  XOR U32648 ( .A(n33721), .B(n33724), .Z(n33722) );
  IV U32649 ( .A(n33677), .Z(n33712) );
  XOR U32650 ( .A(n33675), .B(n33725), .Z(n33677) );
  XNOR U32651 ( .A(n33726), .B(n33727), .Z(n33725) );
  ANDN U32652 ( .B(n33728), .A(n33729), .Z(n33726) );
  XNOR U32653 ( .A(n33730), .B(n33731), .Z(n33728) );
  IV U32654 ( .A(n33679), .Z(n33675) );
  XOR U32655 ( .A(n33732), .B(n33733), .Z(n33679) );
  ANDN U32656 ( .B(n33734), .A(n33735), .Z(n33732) );
  XOR U32657 ( .A(n33736), .B(n33733), .Z(n33734) );
  XOR U32658 ( .A(n33690), .B(n33543), .Z(n33691) );
  XOR U32659 ( .A(n33737), .B(n33738), .Z(n33543) );
  AND U32660 ( .A(n448), .B(n33739), .Z(n33737) );
  XOR U32661 ( .A(n33740), .B(n33738), .Z(n33739) );
  XNOR U32662 ( .A(n33741), .B(n33742), .Z(n33690) );
  NAND U32663 ( .A(n33743), .B(n33744), .Z(n33742) );
  XOR U32664 ( .A(n33745), .B(n33642), .Z(n33744) );
  XOR U32665 ( .A(n33718), .B(n33719), .Z(n33642) );
  XOR U32666 ( .A(n33746), .B(n33711), .Z(n33719) );
  XOR U32667 ( .A(n33747), .B(n33699), .Z(n33711) );
  XOR U32668 ( .A(n33748), .B(n33749), .Z(n33699) );
  ANDN U32669 ( .B(n33750), .A(n33751), .Z(n33748) );
  XOR U32670 ( .A(n33749), .B(n33752), .Z(n33750) );
  IV U32671 ( .A(n33697), .Z(n33747) );
  XOR U32672 ( .A(n33695), .B(n33753), .Z(n33697) );
  XOR U32673 ( .A(n33754), .B(n33755), .Z(n33753) );
  ANDN U32674 ( .B(n33756), .A(n33757), .Z(n33754) );
  XOR U32675 ( .A(n33758), .B(n33755), .Z(n33756) );
  IV U32676 ( .A(n33698), .Z(n33695) );
  XOR U32677 ( .A(n33759), .B(n33760), .Z(n33698) );
  ANDN U32678 ( .B(n33761), .A(n33762), .Z(n33759) );
  XOR U32679 ( .A(n33760), .B(n33763), .Z(n33761) );
  IV U32680 ( .A(n33710), .Z(n33746) );
  XOR U32681 ( .A(n33764), .B(n33765), .Z(n33710) );
  XNOR U32682 ( .A(n33705), .B(n33766), .Z(n33765) );
  IV U32683 ( .A(n33708), .Z(n33766) );
  XOR U32684 ( .A(n33767), .B(n33768), .Z(n33708) );
  ANDN U32685 ( .B(n33769), .A(n33770), .Z(n33767) );
  XOR U32686 ( .A(n33768), .B(n33771), .Z(n33769) );
  XNOR U32687 ( .A(n33772), .B(n33773), .Z(n33705) );
  ANDN U32688 ( .B(n33774), .A(n33775), .Z(n33772) );
  XOR U32689 ( .A(n33773), .B(n33776), .Z(n33774) );
  IV U32690 ( .A(n33704), .Z(n33764) );
  XOR U32691 ( .A(n33702), .B(n33777), .Z(n33704) );
  XOR U32692 ( .A(n33778), .B(n33779), .Z(n33777) );
  ANDN U32693 ( .B(n33780), .A(n33781), .Z(n33778) );
  XOR U32694 ( .A(n33782), .B(n33779), .Z(n33780) );
  IV U32695 ( .A(n33706), .Z(n33702) );
  XOR U32696 ( .A(n33783), .B(n33784), .Z(n33706) );
  ANDN U32697 ( .B(n33785), .A(n33786), .Z(n33783) );
  XOR U32698 ( .A(n33787), .B(n33784), .Z(n33785) );
  XOR U32699 ( .A(n33788), .B(n33789), .Z(n33718) );
  XOR U32700 ( .A(n33736), .B(n33790), .Z(n33789) );
  IV U32701 ( .A(n33716), .Z(n33790) );
  XOR U32702 ( .A(n33791), .B(n33792), .Z(n33716) );
  ANDN U32703 ( .B(n33793), .A(n33794), .Z(n33791) );
  XOR U32704 ( .A(n33792), .B(n33795), .Z(n33793) );
  XOR U32705 ( .A(n33796), .B(n33724), .Z(n33736) );
  XOR U32706 ( .A(n33797), .B(n33798), .Z(n33724) );
  ANDN U32707 ( .B(n33799), .A(n33800), .Z(n33797) );
  XOR U32708 ( .A(n33798), .B(n33801), .Z(n33799) );
  IV U32709 ( .A(n33723), .Z(n33796) );
  XOR U32710 ( .A(n33802), .B(n33803), .Z(n33723) );
  XOR U32711 ( .A(n33804), .B(n33805), .Z(n33803) );
  ANDN U32712 ( .B(n33806), .A(n33807), .Z(n33804) );
  XOR U32713 ( .A(n33808), .B(n33805), .Z(n33806) );
  IV U32714 ( .A(n33721), .Z(n33802) );
  XOR U32715 ( .A(n33809), .B(n33810), .Z(n33721) );
  ANDN U32716 ( .B(n33811), .A(n33812), .Z(n33809) );
  XOR U32717 ( .A(n33810), .B(n33813), .Z(n33811) );
  IV U32718 ( .A(n33735), .Z(n33788) );
  XOR U32719 ( .A(n33814), .B(n33815), .Z(n33735) );
  XNOR U32720 ( .A(n33730), .B(n33816), .Z(n33815) );
  IV U32721 ( .A(n33733), .Z(n33816) );
  XOR U32722 ( .A(n33817), .B(n33818), .Z(n33733) );
  ANDN U32723 ( .B(n33819), .A(n33820), .Z(n33817) );
  XOR U32724 ( .A(n33821), .B(n33818), .Z(n33819) );
  XNOR U32725 ( .A(n33822), .B(n33823), .Z(n33730) );
  ANDN U32726 ( .B(n33824), .A(n33825), .Z(n33822) );
  XOR U32727 ( .A(n33823), .B(n33826), .Z(n33824) );
  IV U32728 ( .A(n33729), .Z(n33814) );
  XOR U32729 ( .A(n33727), .B(n33827), .Z(n33729) );
  XOR U32730 ( .A(n33828), .B(n33829), .Z(n33827) );
  ANDN U32731 ( .B(n33830), .A(n33831), .Z(n33828) );
  XOR U32732 ( .A(n33832), .B(n33829), .Z(n33830) );
  IV U32733 ( .A(n33731), .Z(n33727) );
  XOR U32734 ( .A(n33833), .B(n33834), .Z(n33731) );
  ANDN U32735 ( .B(n33835), .A(n33836), .Z(n33833) );
  XOR U32736 ( .A(n33837), .B(n33834), .Z(n33835) );
  IV U32737 ( .A(n33741), .Z(n33745) );
  XOR U32738 ( .A(n33741), .B(n33644), .Z(n33743) );
  XOR U32739 ( .A(n33838), .B(n33839), .Z(n33644) );
  AND U32740 ( .A(n448), .B(n33840), .Z(n33838) );
  XOR U32741 ( .A(n33841), .B(n33839), .Z(n33840) );
  NANDN U32742 ( .A(n33646), .B(n33648), .Z(n33741) );
  XOR U32743 ( .A(n33842), .B(n33843), .Z(n33648) );
  AND U32744 ( .A(n448), .B(n33844), .Z(n33842) );
  XOR U32745 ( .A(n33843), .B(n33845), .Z(n33844) );
  XNOR U32746 ( .A(n33846), .B(n33847), .Z(n448) );
  AND U32747 ( .A(n33848), .B(n33849), .Z(n33846) );
  XOR U32748 ( .A(n33847), .B(n33659), .Z(n33849) );
  XNOR U32749 ( .A(n33850), .B(n33851), .Z(n33659) );
  ANDN U32750 ( .B(n33852), .A(n33853), .Z(n33850) );
  XOR U32751 ( .A(n33851), .B(n33854), .Z(n33852) );
  XNOR U32752 ( .A(n33847), .B(n33661), .Z(n33848) );
  XOR U32753 ( .A(n33855), .B(n33856), .Z(n33661) );
  AND U32754 ( .A(n452), .B(n33857), .Z(n33855) );
  XOR U32755 ( .A(n33858), .B(n33856), .Z(n33857) );
  XOR U32756 ( .A(n33859), .B(n33860), .Z(n33847) );
  AND U32757 ( .A(n33861), .B(n33862), .Z(n33859) );
  XOR U32758 ( .A(n33860), .B(n33686), .Z(n33862) );
  XOR U32759 ( .A(n33853), .B(n33854), .Z(n33686) );
  XNOR U32760 ( .A(n33863), .B(n33864), .Z(n33854) );
  ANDN U32761 ( .B(n33865), .A(n33866), .Z(n33863) );
  XOR U32762 ( .A(n33867), .B(n33868), .Z(n33865) );
  XOR U32763 ( .A(n33869), .B(n33870), .Z(n33853) );
  XNOR U32764 ( .A(n33871), .B(n33872), .Z(n33870) );
  ANDN U32765 ( .B(n33873), .A(n33874), .Z(n33871) );
  XNOR U32766 ( .A(n33875), .B(n33876), .Z(n33873) );
  IV U32767 ( .A(n33851), .Z(n33869) );
  XOR U32768 ( .A(n33877), .B(n33878), .Z(n33851) );
  ANDN U32769 ( .B(n33879), .A(n33880), .Z(n33877) );
  XOR U32770 ( .A(n33878), .B(n33881), .Z(n33879) );
  XNOR U32771 ( .A(n33860), .B(n33688), .Z(n33861) );
  XOR U32772 ( .A(n33882), .B(n33883), .Z(n33688) );
  AND U32773 ( .A(n452), .B(n33884), .Z(n33882) );
  XOR U32774 ( .A(n33885), .B(n33883), .Z(n33884) );
  XNOR U32775 ( .A(n33886), .B(n33887), .Z(n33860) );
  AND U32776 ( .A(n33888), .B(n33889), .Z(n33886) );
  XNOR U32777 ( .A(n33887), .B(n33738), .Z(n33889) );
  XOR U32778 ( .A(n33880), .B(n33881), .Z(n33738) );
  XOR U32779 ( .A(n33890), .B(n33868), .Z(n33881) );
  XNOR U32780 ( .A(n33891), .B(n33892), .Z(n33868) );
  ANDN U32781 ( .B(n33893), .A(n33894), .Z(n33891) );
  XOR U32782 ( .A(n33895), .B(n33896), .Z(n33893) );
  IV U32783 ( .A(n33866), .Z(n33890) );
  XOR U32784 ( .A(n33864), .B(n33897), .Z(n33866) );
  XNOR U32785 ( .A(n33898), .B(n33899), .Z(n33897) );
  ANDN U32786 ( .B(n33900), .A(n33901), .Z(n33898) );
  XNOR U32787 ( .A(n33902), .B(n33903), .Z(n33900) );
  IV U32788 ( .A(n33867), .Z(n33864) );
  XOR U32789 ( .A(n33904), .B(n33905), .Z(n33867) );
  ANDN U32790 ( .B(n33906), .A(n33907), .Z(n33904) );
  XOR U32791 ( .A(n33905), .B(n33908), .Z(n33906) );
  XOR U32792 ( .A(n33909), .B(n33910), .Z(n33880) );
  XNOR U32793 ( .A(n33875), .B(n33911), .Z(n33910) );
  IV U32794 ( .A(n33878), .Z(n33911) );
  XOR U32795 ( .A(n33912), .B(n33913), .Z(n33878) );
  ANDN U32796 ( .B(n33914), .A(n33915), .Z(n33912) );
  XOR U32797 ( .A(n33913), .B(n33916), .Z(n33914) );
  XNOR U32798 ( .A(n33917), .B(n33918), .Z(n33875) );
  ANDN U32799 ( .B(n33919), .A(n33920), .Z(n33917) );
  XOR U32800 ( .A(n33918), .B(n33921), .Z(n33919) );
  IV U32801 ( .A(n33874), .Z(n33909) );
  XOR U32802 ( .A(n33872), .B(n33922), .Z(n33874) );
  XNOR U32803 ( .A(n33923), .B(n33924), .Z(n33922) );
  ANDN U32804 ( .B(n33925), .A(n33926), .Z(n33923) );
  XNOR U32805 ( .A(n33927), .B(n33928), .Z(n33925) );
  IV U32806 ( .A(n33876), .Z(n33872) );
  XOR U32807 ( .A(n33929), .B(n33930), .Z(n33876) );
  ANDN U32808 ( .B(n33931), .A(n33932), .Z(n33929) );
  XOR U32809 ( .A(n33933), .B(n33930), .Z(n33931) );
  XOR U32810 ( .A(n33887), .B(n33740), .Z(n33888) );
  XOR U32811 ( .A(n33934), .B(n33935), .Z(n33740) );
  AND U32812 ( .A(n452), .B(n33936), .Z(n33934) );
  XOR U32813 ( .A(n33937), .B(n33935), .Z(n33936) );
  XNOR U32814 ( .A(n33938), .B(n33939), .Z(n33887) );
  NAND U32815 ( .A(n33940), .B(n33941), .Z(n33939) );
  XOR U32816 ( .A(n33942), .B(n33839), .Z(n33941) );
  XOR U32817 ( .A(n33915), .B(n33916), .Z(n33839) );
  XOR U32818 ( .A(n33943), .B(n33908), .Z(n33916) );
  XOR U32819 ( .A(n33944), .B(n33896), .Z(n33908) );
  XOR U32820 ( .A(n33945), .B(n33946), .Z(n33896) );
  ANDN U32821 ( .B(n33947), .A(n33948), .Z(n33945) );
  XOR U32822 ( .A(n33946), .B(n33949), .Z(n33947) );
  IV U32823 ( .A(n33894), .Z(n33944) );
  XOR U32824 ( .A(n33892), .B(n33950), .Z(n33894) );
  XOR U32825 ( .A(n33951), .B(n33952), .Z(n33950) );
  ANDN U32826 ( .B(n33953), .A(n33954), .Z(n33951) );
  XOR U32827 ( .A(n33955), .B(n33952), .Z(n33953) );
  IV U32828 ( .A(n33895), .Z(n33892) );
  XOR U32829 ( .A(n33956), .B(n33957), .Z(n33895) );
  ANDN U32830 ( .B(n33958), .A(n33959), .Z(n33956) );
  XOR U32831 ( .A(n33957), .B(n33960), .Z(n33958) );
  IV U32832 ( .A(n33907), .Z(n33943) );
  XOR U32833 ( .A(n33961), .B(n33962), .Z(n33907) );
  XNOR U32834 ( .A(n33902), .B(n33963), .Z(n33962) );
  IV U32835 ( .A(n33905), .Z(n33963) );
  XOR U32836 ( .A(n33964), .B(n33965), .Z(n33905) );
  ANDN U32837 ( .B(n33966), .A(n33967), .Z(n33964) );
  XOR U32838 ( .A(n33965), .B(n33968), .Z(n33966) );
  XNOR U32839 ( .A(n33969), .B(n33970), .Z(n33902) );
  ANDN U32840 ( .B(n33971), .A(n33972), .Z(n33969) );
  XOR U32841 ( .A(n33970), .B(n33973), .Z(n33971) );
  IV U32842 ( .A(n33901), .Z(n33961) );
  XOR U32843 ( .A(n33899), .B(n33974), .Z(n33901) );
  XOR U32844 ( .A(n33975), .B(n33976), .Z(n33974) );
  ANDN U32845 ( .B(n33977), .A(n33978), .Z(n33975) );
  XOR U32846 ( .A(n33979), .B(n33976), .Z(n33977) );
  IV U32847 ( .A(n33903), .Z(n33899) );
  XOR U32848 ( .A(n33980), .B(n33981), .Z(n33903) );
  ANDN U32849 ( .B(n33982), .A(n33983), .Z(n33980) );
  XOR U32850 ( .A(n33984), .B(n33981), .Z(n33982) );
  XOR U32851 ( .A(n33985), .B(n33986), .Z(n33915) );
  XOR U32852 ( .A(n33933), .B(n33987), .Z(n33986) );
  IV U32853 ( .A(n33913), .Z(n33987) );
  XOR U32854 ( .A(n33988), .B(n33989), .Z(n33913) );
  ANDN U32855 ( .B(n33990), .A(n33991), .Z(n33988) );
  XOR U32856 ( .A(n33989), .B(n33992), .Z(n33990) );
  XOR U32857 ( .A(n33993), .B(n33921), .Z(n33933) );
  XOR U32858 ( .A(n33994), .B(n33995), .Z(n33921) );
  ANDN U32859 ( .B(n33996), .A(n33997), .Z(n33994) );
  XOR U32860 ( .A(n33995), .B(n33998), .Z(n33996) );
  IV U32861 ( .A(n33920), .Z(n33993) );
  XOR U32862 ( .A(n33999), .B(n34000), .Z(n33920) );
  XOR U32863 ( .A(n34001), .B(n34002), .Z(n34000) );
  ANDN U32864 ( .B(n34003), .A(n34004), .Z(n34001) );
  XOR U32865 ( .A(n34005), .B(n34002), .Z(n34003) );
  IV U32866 ( .A(n33918), .Z(n33999) );
  XOR U32867 ( .A(n34006), .B(n34007), .Z(n33918) );
  ANDN U32868 ( .B(n34008), .A(n34009), .Z(n34006) );
  XOR U32869 ( .A(n34007), .B(n34010), .Z(n34008) );
  IV U32870 ( .A(n33932), .Z(n33985) );
  XOR U32871 ( .A(n34011), .B(n34012), .Z(n33932) );
  XNOR U32872 ( .A(n33927), .B(n34013), .Z(n34012) );
  IV U32873 ( .A(n33930), .Z(n34013) );
  XOR U32874 ( .A(n34014), .B(n34015), .Z(n33930) );
  ANDN U32875 ( .B(n34016), .A(n34017), .Z(n34014) );
  XOR U32876 ( .A(n34018), .B(n34015), .Z(n34016) );
  XNOR U32877 ( .A(n34019), .B(n34020), .Z(n33927) );
  ANDN U32878 ( .B(n34021), .A(n34022), .Z(n34019) );
  XOR U32879 ( .A(n34020), .B(n34023), .Z(n34021) );
  IV U32880 ( .A(n33926), .Z(n34011) );
  XOR U32881 ( .A(n33924), .B(n34024), .Z(n33926) );
  XOR U32882 ( .A(n34025), .B(n34026), .Z(n34024) );
  ANDN U32883 ( .B(n34027), .A(n34028), .Z(n34025) );
  XOR U32884 ( .A(n34029), .B(n34026), .Z(n34027) );
  IV U32885 ( .A(n33928), .Z(n33924) );
  XOR U32886 ( .A(n34030), .B(n34031), .Z(n33928) );
  ANDN U32887 ( .B(n34032), .A(n34033), .Z(n34030) );
  XOR U32888 ( .A(n34034), .B(n34031), .Z(n34032) );
  IV U32889 ( .A(n33938), .Z(n33942) );
  XOR U32890 ( .A(n33938), .B(n33841), .Z(n33940) );
  XOR U32891 ( .A(n34035), .B(n34036), .Z(n33841) );
  AND U32892 ( .A(n452), .B(n34037), .Z(n34035) );
  XOR U32893 ( .A(n34038), .B(n34036), .Z(n34037) );
  NANDN U32894 ( .A(n33843), .B(n33845), .Z(n33938) );
  XOR U32895 ( .A(n34039), .B(n34040), .Z(n33845) );
  AND U32896 ( .A(n452), .B(n34041), .Z(n34039) );
  XOR U32897 ( .A(n34040), .B(n34042), .Z(n34041) );
  XNOR U32898 ( .A(n34043), .B(n34044), .Z(n452) );
  AND U32899 ( .A(n34045), .B(n34046), .Z(n34043) );
  XOR U32900 ( .A(n34044), .B(n33856), .Z(n34046) );
  XNOR U32901 ( .A(n34047), .B(n34048), .Z(n33856) );
  ANDN U32902 ( .B(n34049), .A(n34050), .Z(n34047) );
  XOR U32903 ( .A(n34048), .B(n34051), .Z(n34049) );
  XNOR U32904 ( .A(n34044), .B(n33858), .Z(n34045) );
  XOR U32905 ( .A(n34052), .B(n34053), .Z(n33858) );
  AND U32906 ( .A(n456), .B(n34054), .Z(n34052) );
  XOR U32907 ( .A(n34055), .B(n34053), .Z(n34054) );
  XOR U32908 ( .A(n34056), .B(n34057), .Z(n34044) );
  AND U32909 ( .A(n34058), .B(n34059), .Z(n34056) );
  XOR U32910 ( .A(n34057), .B(n33883), .Z(n34059) );
  XOR U32911 ( .A(n34050), .B(n34051), .Z(n33883) );
  XNOR U32912 ( .A(n34060), .B(n34061), .Z(n34051) );
  ANDN U32913 ( .B(n34062), .A(n34063), .Z(n34060) );
  XOR U32914 ( .A(n34064), .B(n34065), .Z(n34062) );
  XOR U32915 ( .A(n34066), .B(n34067), .Z(n34050) );
  XNOR U32916 ( .A(n34068), .B(n34069), .Z(n34067) );
  ANDN U32917 ( .B(n34070), .A(n34071), .Z(n34068) );
  XNOR U32918 ( .A(n34072), .B(n34073), .Z(n34070) );
  IV U32919 ( .A(n34048), .Z(n34066) );
  XOR U32920 ( .A(n34074), .B(n34075), .Z(n34048) );
  ANDN U32921 ( .B(n34076), .A(n34077), .Z(n34074) );
  XOR U32922 ( .A(n34075), .B(n34078), .Z(n34076) );
  XNOR U32923 ( .A(n34057), .B(n33885), .Z(n34058) );
  XOR U32924 ( .A(n34079), .B(n34080), .Z(n33885) );
  AND U32925 ( .A(n456), .B(n34081), .Z(n34079) );
  XOR U32926 ( .A(n34082), .B(n34080), .Z(n34081) );
  XNOR U32927 ( .A(n34083), .B(n34084), .Z(n34057) );
  AND U32928 ( .A(n34085), .B(n34086), .Z(n34083) );
  XNOR U32929 ( .A(n34084), .B(n33935), .Z(n34086) );
  XOR U32930 ( .A(n34077), .B(n34078), .Z(n33935) );
  XOR U32931 ( .A(n34087), .B(n34065), .Z(n34078) );
  XNOR U32932 ( .A(n34088), .B(n34089), .Z(n34065) );
  ANDN U32933 ( .B(n34090), .A(n34091), .Z(n34088) );
  XOR U32934 ( .A(n34092), .B(n34093), .Z(n34090) );
  IV U32935 ( .A(n34063), .Z(n34087) );
  XOR U32936 ( .A(n34061), .B(n34094), .Z(n34063) );
  XNOR U32937 ( .A(n34095), .B(n34096), .Z(n34094) );
  ANDN U32938 ( .B(n34097), .A(n34098), .Z(n34095) );
  XNOR U32939 ( .A(n34099), .B(n34100), .Z(n34097) );
  IV U32940 ( .A(n34064), .Z(n34061) );
  XOR U32941 ( .A(n34101), .B(n34102), .Z(n34064) );
  ANDN U32942 ( .B(n34103), .A(n34104), .Z(n34101) );
  XOR U32943 ( .A(n34102), .B(n34105), .Z(n34103) );
  XOR U32944 ( .A(n34106), .B(n34107), .Z(n34077) );
  XNOR U32945 ( .A(n34072), .B(n34108), .Z(n34107) );
  IV U32946 ( .A(n34075), .Z(n34108) );
  XOR U32947 ( .A(n34109), .B(n34110), .Z(n34075) );
  ANDN U32948 ( .B(n34111), .A(n34112), .Z(n34109) );
  XOR U32949 ( .A(n34110), .B(n34113), .Z(n34111) );
  XNOR U32950 ( .A(n34114), .B(n34115), .Z(n34072) );
  ANDN U32951 ( .B(n34116), .A(n34117), .Z(n34114) );
  XOR U32952 ( .A(n34115), .B(n34118), .Z(n34116) );
  IV U32953 ( .A(n34071), .Z(n34106) );
  XOR U32954 ( .A(n34069), .B(n34119), .Z(n34071) );
  XNOR U32955 ( .A(n34120), .B(n34121), .Z(n34119) );
  ANDN U32956 ( .B(n34122), .A(n34123), .Z(n34120) );
  XNOR U32957 ( .A(n34124), .B(n34125), .Z(n34122) );
  IV U32958 ( .A(n34073), .Z(n34069) );
  XOR U32959 ( .A(n34126), .B(n34127), .Z(n34073) );
  ANDN U32960 ( .B(n34128), .A(n34129), .Z(n34126) );
  XOR U32961 ( .A(n34130), .B(n34127), .Z(n34128) );
  XOR U32962 ( .A(n34084), .B(n33937), .Z(n34085) );
  XOR U32963 ( .A(n34131), .B(n34132), .Z(n33937) );
  AND U32964 ( .A(n456), .B(n34133), .Z(n34131) );
  XOR U32965 ( .A(n34134), .B(n34132), .Z(n34133) );
  XNOR U32966 ( .A(n34135), .B(n34136), .Z(n34084) );
  NAND U32967 ( .A(n34137), .B(n34138), .Z(n34136) );
  XOR U32968 ( .A(n34139), .B(n34036), .Z(n34138) );
  XOR U32969 ( .A(n34112), .B(n34113), .Z(n34036) );
  XOR U32970 ( .A(n34140), .B(n34105), .Z(n34113) );
  XOR U32971 ( .A(n34141), .B(n34093), .Z(n34105) );
  XOR U32972 ( .A(n34142), .B(n34143), .Z(n34093) );
  ANDN U32973 ( .B(n34144), .A(n34145), .Z(n34142) );
  XOR U32974 ( .A(n34143), .B(n34146), .Z(n34144) );
  IV U32975 ( .A(n34091), .Z(n34141) );
  XOR U32976 ( .A(n34089), .B(n34147), .Z(n34091) );
  XOR U32977 ( .A(n34148), .B(n34149), .Z(n34147) );
  ANDN U32978 ( .B(n34150), .A(n34151), .Z(n34148) );
  XOR U32979 ( .A(n34152), .B(n34149), .Z(n34150) );
  IV U32980 ( .A(n34092), .Z(n34089) );
  XOR U32981 ( .A(n34153), .B(n34154), .Z(n34092) );
  ANDN U32982 ( .B(n34155), .A(n34156), .Z(n34153) );
  XOR U32983 ( .A(n34154), .B(n34157), .Z(n34155) );
  IV U32984 ( .A(n34104), .Z(n34140) );
  XOR U32985 ( .A(n34158), .B(n34159), .Z(n34104) );
  XNOR U32986 ( .A(n34099), .B(n34160), .Z(n34159) );
  IV U32987 ( .A(n34102), .Z(n34160) );
  XOR U32988 ( .A(n34161), .B(n34162), .Z(n34102) );
  ANDN U32989 ( .B(n34163), .A(n34164), .Z(n34161) );
  XOR U32990 ( .A(n34162), .B(n34165), .Z(n34163) );
  XNOR U32991 ( .A(n34166), .B(n34167), .Z(n34099) );
  ANDN U32992 ( .B(n34168), .A(n34169), .Z(n34166) );
  XOR U32993 ( .A(n34167), .B(n34170), .Z(n34168) );
  IV U32994 ( .A(n34098), .Z(n34158) );
  XOR U32995 ( .A(n34096), .B(n34171), .Z(n34098) );
  XOR U32996 ( .A(n34172), .B(n34173), .Z(n34171) );
  ANDN U32997 ( .B(n34174), .A(n34175), .Z(n34172) );
  XOR U32998 ( .A(n34176), .B(n34173), .Z(n34174) );
  IV U32999 ( .A(n34100), .Z(n34096) );
  XOR U33000 ( .A(n34177), .B(n34178), .Z(n34100) );
  ANDN U33001 ( .B(n34179), .A(n34180), .Z(n34177) );
  XOR U33002 ( .A(n34181), .B(n34178), .Z(n34179) );
  XOR U33003 ( .A(n34182), .B(n34183), .Z(n34112) );
  XOR U33004 ( .A(n34130), .B(n34184), .Z(n34183) );
  IV U33005 ( .A(n34110), .Z(n34184) );
  XOR U33006 ( .A(n34185), .B(n34186), .Z(n34110) );
  ANDN U33007 ( .B(n34187), .A(n34188), .Z(n34185) );
  XOR U33008 ( .A(n34186), .B(n34189), .Z(n34187) );
  XOR U33009 ( .A(n34190), .B(n34118), .Z(n34130) );
  XOR U33010 ( .A(n34191), .B(n34192), .Z(n34118) );
  ANDN U33011 ( .B(n34193), .A(n34194), .Z(n34191) );
  XOR U33012 ( .A(n34192), .B(n34195), .Z(n34193) );
  IV U33013 ( .A(n34117), .Z(n34190) );
  XOR U33014 ( .A(n34196), .B(n34197), .Z(n34117) );
  XOR U33015 ( .A(n34198), .B(n34199), .Z(n34197) );
  ANDN U33016 ( .B(n34200), .A(n34201), .Z(n34198) );
  XOR U33017 ( .A(n34202), .B(n34199), .Z(n34200) );
  IV U33018 ( .A(n34115), .Z(n34196) );
  XOR U33019 ( .A(n34203), .B(n34204), .Z(n34115) );
  ANDN U33020 ( .B(n34205), .A(n34206), .Z(n34203) );
  XOR U33021 ( .A(n34204), .B(n34207), .Z(n34205) );
  IV U33022 ( .A(n34129), .Z(n34182) );
  XOR U33023 ( .A(n34208), .B(n34209), .Z(n34129) );
  XNOR U33024 ( .A(n34124), .B(n34210), .Z(n34209) );
  IV U33025 ( .A(n34127), .Z(n34210) );
  XOR U33026 ( .A(n34211), .B(n34212), .Z(n34127) );
  ANDN U33027 ( .B(n34213), .A(n34214), .Z(n34211) );
  XOR U33028 ( .A(n34215), .B(n34212), .Z(n34213) );
  XNOR U33029 ( .A(n34216), .B(n34217), .Z(n34124) );
  ANDN U33030 ( .B(n34218), .A(n34219), .Z(n34216) );
  XOR U33031 ( .A(n34217), .B(n34220), .Z(n34218) );
  IV U33032 ( .A(n34123), .Z(n34208) );
  XOR U33033 ( .A(n34121), .B(n34221), .Z(n34123) );
  XOR U33034 ( .A(n34222), .B(n34223), .Z(n34221) );
  ANDN U33035 ( .B(n34224), .A(n34225), .Z(n34222) );
  XOR U33036 ( .A(n34226), .B(n34223), .Z(n34224) );
  IV U33037 ( .A(n34125), .Z(n34121) );
  XOR U33038 ( .A(n34227), .B(n34228), .Z(n34125) );
  ANDN U33039 ( .B(n34229), .A(n34230), .Z(n34227) );
  XOR U33040 ( .A(n34231), .B(n34228), .Z(n34229) );
  IV U33041 ( .A(n34135), .Z(n34139) );
  XOR U33042 ( .A(n34135), .B(n34038), .Z(n34137) );
  XOR U33043 ( .A(n34232), .B(n34233), .Z(n34038) );
  AND U33044 ( .A(n456), .B(n34234), .Z(n34232) );
  XOR U33045 ( .A(n34235), .B(n34233), .Z(n34234) );
  NANDN U33046 ( .A(n34040), .B(n34042), .Z(n34135) );
  XOR U33047 ( .A(n34236), .B(n34237), .Z(n34042) );
  AND U33048 ( .A(n456), .B(n34238), .Z(n34236) );
  XOR U33049 ( .A(n34237), .B(n34239), .Z(n34238) );
  XNOR U33050 ( .A(n34240), .B(n34241), .Z(n456) );
  AND U33051 ( .A(n34242), .B(n34243), .Z(n34240) );
  XOR U33052 ( .A(n34241), .B(n34053), .Z(n34243) );
  XNOR U33053 ( .A(n34244), .B(n34245), .Z(n34053) );
  ANDN U33054 ( .B(n34246), .A(n34247), .Z(n34244) );
  XOR U33055 ( .A(n34245), .B(n34248), .Z(n34246) );
  XNOR U33056 ( .A(n34241), .B(n34055), .Z(n34242) );
  XOR U33057 ( .A(n34249), .B(n34250), .Z(n34055) );
  AND U33058 ( .A(n460), .B(n34251), .Z(n34249) );
  XOR U33059 ( .A(n34252), .B(n34250), .Z(n34251) );
  XOR U33060 ( .A(n34253), .B(n34254), .Z(n34241) );
  AND U33061 ( .A(n34255), .B(n34256), .Z(n34253) );
  XOR U33062 ( .A(n34254), .B(n34080), .Z(n34256) );
  XOR U33063 ( .A(n34247), .B(n34248), .Z(n34080) );
  XNOR U33064 ( .A(n34257), .B(n34258), .Z(n34248) );
  ANDN U33065 ( .B(n34259), .A(n34260), .Z(n34257) );
  XOR U33066 ( .A(n34261), .B(n34262), .Z(n34259) );
  XOR U33067 ( .A(n34263), .B(n34264), .Z(n34247) );
  XNOR U33068 ( .A(n34265), .B(n34266), .Z(n34264) );
  ANDN U33069 ( .B(n34267), .A(n34268), .Z(n34265) );
  XNOR U33070 ( .A(n34269), .B(n34270), .Z(n34267) );
  IV U33071 ( .A(n34245), .Z(n34263) );
  XOR U33072 ( .A(n34271), .B(n34272), .Z(n34245) );
  ANDN U33073 ( .B(n34273), .A(n34274), .Z(n34271) );
  XOR U33074 ( .A(n34272), .B(n34275), .Z(n34273) );
  XNOR U33075 ( .A(n34254), .B(n34082), .Z(n34255) );
  XOR U33076 ( .A(n34276), .B(n34277), .Z(n34082) );
  AND U33077 ( .A(n460), .B(n34278), .Z(n34276) );
  XOR U33078 ( .A(n34279), .B(n34277), .Z(n34278) );
  XNOR U33079 ( .A(n34280), .B(n34281), .Z(n34254) );
  AND U33080 ( .A(n34282), .B(n34283), .Z(n34280) );
  XNOR U33081 ( .A(n34281), .B(n34132), .Z(n34283) );
  XOR U33082 ( .A(n34274), .B(n34275), .Z(n34132) );
  XOR U33083 ( .A(n34284), .B(n34262), .Z(n34275) );
  XNOR U33084 ( .A(n34285), .B(n34286), .Z(n34262) );
  ANDN U33085 ( .B(n34287), .A(n34288), .Z(n34285) );
  XOR U33086 ( .A(n34289), .B(n34290), .Z(n34287) );
  IV U33087 ( .A(n34260), .Z(n34284) );
  XOR U33088 ( .A(n34258), .B(n34291), .Z(n34260) );
  XNOR U33089 ( .A(n34292), .B(n34293), .Z(n34291) );
  ANDN U33090 ( .B(n34294), .A(n34295), .Z(n34292) );
  XNOR U33091 ( .A(n34296), .B(n34297), .Z(n34294) );
  IV U33092 ( .A(n34261), .Z(n34258) );
  XOR U33093 ( .A(n34298), .B(n34299), .Z(n34261) );
  ANDN U33094 ( .B(n34300), .A(n34301), .Z(n34298) );
  XOR U33095 ( .A(n34299), .B(n34302), .Z(n34300) );
  XOR U33096 ( .A(n34303), .B(n34304), .Z(n34274) );
  XNOR U33097 ( .A(n34269), .B(n34305), .Z(n34304) );
  IV U33098 ( .A(n34272), .Z(n34305) );
  XOR U33099 ( .A(n34306), .B(n34307), .Z(n34272) );
  ANDN U33100 ( .B(n34308), .A(n34309), .Z(n34306) );
  XOR U33101 ( .A(n34307), .B(n34310), .Z(n34308) );
  XNOR U33102 ( .A(n34311), .B(n34312), .Z(n34269) );
  ANDN U33103 ( .B(n34313), .A(n34314), .Z(n34311) );
  XOR U33104 ( .A(n34312), .B(n34315), .Z(n34313) );
  IV U33105 ( .A(n34268), .Z(n34303) );
  XOR U33106 ( .A(n34266), .B(n34316), .Z(n34268) );
  XNOR U33107 ( .A(n34317), .B(n34318), .Z(n34316) );
  ANDN U33108 ( .B(n34319), .A(n34320), .Z(n34317) );
  XNOR U33109 ( .A(n34321), .B(n34322), .Z(n34319) );
  IV U33110 ( .A(n34270), .Z(n34266) );
  XOR U33111 ( .A(n34323), .B(n34324), .Z(n34270) );
  ANDN U33112 ( .B(n34325), .A(n34326), .Z(n34323) );
  XOR U33113 ( .A(n34327), .B(n34324), .Z(n34325) );
  XOR U33114 ( .A(n34281), .B(n34134), .Z(n34282) );
  XOR U33115 ( .A(n34328), .B(n34329), .Z(n34134) );
  AND U33116 ( .A(n460), .B(n34330), .Z(n34328) );
  XOR U33117 ( .A(n34331), .B(n34329), .Z(n34330) );
  XNOR U33118 ( .A(n34332), .B(n34333), .Z(n34281) );
  NAND U33119 ( .A(n34334), .B(n34335), .Z(n34333) );
  XOR U33120 ( .A(n34336), .B(n34233), .Z(n34335) );
  XOR U33121 ( .A(n34309), .B(n34310), .Z(n34233) );
  XOR U33122 ( .A(n34337), .B(n34302), .Z(n34310) );
  XOR U33123 ( .A(n34338), .B(n34290), .Z(n34302) );
  XOR U33124 ( .A(n34339), .B(n34340), .Z(n34290) );
  ANDN U33125 ( .B(n34341), .A(n34342), .Z(n34339) );
  XOR U33126 ( .A(n34340), .B(n34343), .Z(n34341) );
  IV U33127 ( .A(n34288), .Z(n34338) );
  XOR U33128 ( .A(n34286), .B(n34344), .Z(n34288) );
  XOR U33129 ( .A(n34345), .B(n34346), .Z(n34344) );
  ANDN U33130 ( .B(n34347), .A(n34348), .Z(n34345) );
  XOR U33131 ( .A(n34349), .B(n34346), .Z(n34347) );
  IV U33132 ( .A(n34289), .Z(n34286) );
  XOR U33133 ( .A(n34350), .B(n34351), .Z(n34289) );
  ANDN U33134 ( .B(n34352), .A(n34353), .Z(n34350) );
  XOR U33135 ( .A(n34351), .B(n34354), .Z(n34352) );
  IV U33136 ( .A(n34301), .Z(n34337) );
  XOR U33137 ( .A(n34355), .B(n34356), .Z(n34301) );
  XNOR U33138 ( .A(n34296), .B(n34357), .Z(n34356) );
  IV U33139 ( .A(n34299), .Z(n34357) );
  XOR U33140 ( .A(n34358), .B(n34359), .Z(n34299) );
  ANDN U33141 ( .B(n34360), .A(n34361), .Z(n34358) );
  XOR U33142 ( .A(n34359), .B(n34362), .Z(n34360) );
  XNOR U33143 ( .A(n34363), .B(n34364), .Z(n34296) );
  ANDN U33144 ( .B(n34365), .A(n34366), .Z(n34363) );
  XOR U33145 ( .A(n34364), .B(n34367), .Z(n34365) );
  IV U33146 ( .A(n34295), .Z(n34355) );
  XOR U33147 ( .A(n34293), .B(n34368), .Z(n34295) );
  XOR U33148 ( .A(n34369), .B(n34370), .Z(n34368) );
  ANDN U33149 ( .B(n34371), .A(n34372), .Z(n34369) );
  XOR U33150 ( .A(n34373), .B(n34370), .Z(n34371) );
  IV U33151 ( .A(n34297), .Z(n34293) );
  XOR U33152 ( .A(n34374), .B(n34375), .Z(n34297) );
  ANDN U33153 ( .B(n34376), .A(n34377), .Z(n34374) );
  XOR U33154 ( .A(n34378), .B(n34375), .Z(n34376) );
  XOR U33155 ( .A(n34379), .B(n34380), .Z(n34309) );
  XOR U33156 ( .A(n34327), .B(n34381), .Z(n34380) );
  IV U33157 ( .A(n34307), .Z(n34381) );
  XOR U33158 ( .A(n34382), .B(n34383), .Z(n34307) );
  ANDN U33159 ( .B(n34384), .A(n34385), .Z(n34382) );
  XOR U33160 ( .A(n34383), .B(n34386), .Z(n34384) );
  XOR U33161 ( .A(n34387), .B(n34315), .Z(n34327) );
  XOR U33162 ( .A(n34388), .B(n34389), .Z(n34315) );
  ANDN U33163 ( .B(n34390), .A(n34391), .Z(n34388) );
  XOR U33164 ( .A(n34389), .B(n34392), .Z(n34390) );
  IV U33165 ( .A(n34314), .Z(n34387) );
  XOR U33166 ( .A(n34393), .B(n34394), .Z(n34314) );
  XOR U33167 ( .A(n34395), .B(n34396), .Z(n34394) );
  ANDN U33168 ( .B(n34397), .A(n34398), .Z(n34395) );
  XOR U33169 ( .A(n34399), .B(n34396), .Z(n34397) );
  IV U33170 ( .A(n34312), .Z(n34393) );
  XOR U33171 ( .A(n34400), .B(n34401), .Z(n34312) );
  ANDN U33172 ( .B(n34402), .A(n34403), .Z(n34400) );
  XOR U33173 ( .A(n34401), .B(n34404), .Z(n34402) );
  IV U33174 ( .A(n34326), .Z(n34379) );
  XOR U33175 ( .A(n34405), .B(n34406), .Z(n34326) );
  XNOR U33176 ( .A(n34321), .B(n34407), .Z(n34406) );
  IV U33177 ( .A(n34324), .Z(n34407) );
  XOR U33178 ( .A(n34408), .B(n34409), .Z(n34324) );
  ANDN U33179 ( .B(n34410), .A(n34411), .Z(n34408) );
  XOR U33180 ( .A(n34412), .B(n34409), .Z(n34410) );
  XNOR U33181 ( .A(n34413), .B(n34414), .Z(n34321) );
  ANDN U33182 ( .B(n34415), .A(n34416), .Z(n34413) );
  XOR U33183 ( .A(n34414), .B(n34417), .Z(n34415) );
  IV U33184 ( .A(n34320), .Z(n34405) );
  XOR U33185 ( .A(n34318), .B(n34418), .Z(n34320) );
  XOR U33186 ( .A(n34419), .B(n34420), .Z(n34418) );
  ANDN U33187 ( .B(n34421), .A(n34422), .Z(n34419) );
  XOR U33188 ( .A(n34423), .B(n34420), .Z(n34421) );
  IV U33189 ( .A(n34322), .Z(n34318) );
  XOR U33190 ( .A(n34424), .B(n34425), .Z(n34322) );
  ANDN U33191 ( .B(n34426), .A(n34427), .Z(n34424) );
  XOR U33192 ( .A(n34428), .B(n34425), .Z(n34426) );
  IV U33193 ( .A(n34332), .Z(n34336) );
  XOR U33194 ( .A(n34332), .B(n34235), .Z(n34334) );
  XOR U33195 ( .A(n34429), .B(n34430), .Z(n34235) );
  AND U33196 ( .A(n460), .B(n34431), .Z(n34429) );
  XOR U33197 ( .A(n34432), .B(n34430), .Z(n34431) );
  NANDN U33198 ( .A(n34237), .B(n34239), .Z(n34332) );
  XOR U33199 ( .A(n34433), .B(n34434), .Z(n34239) );
  AND U33200 ( .A(n460), .B(n34435), .Z(n34433) );
  XOR U33201 ( .A(n34434), .B(n34436), .Z(n34435) );
  XNOR U33202 ( .A(n34437), .B(n34438), .Z(n460) );
  AND U33203 ( .A(n34439), .B(n34440), .Z(n34437) );
  XOR U33204 ( .A(n34438), .B(n34250), .Z(n34440) );
  XNOR U33205 ( .A(n34441), .B(n34442), .Z(n34250) );
  ANDN U33206 ( .B(n34443), .A(n34444), .Z(n34441) );
  XOR U33207 ( .A(n34442), .B(n34445), .Z(n34443) );
  XNOR U33208 ( .A(n34438), .B(n34252), .Z(n34439) );
  XOR U33209 ( .A(n34446), .B(n34447), .Z(n34252) );
  AND U33210 ( .A(n464), .B(n34448), .Z(n34446) );
  XOR U33211 ( .A(n34449), .B(n34447), .Z(n34448) );
  XOR U33212 ( .A(n34450), .B(n34451), .Z(n34438) );
  AND U33213 ( .A(n34452), .B(n34453), .Z(n34450) );
  XOR U33214 ( .A(n34451), .B(n34277), .Z(n34453) );
  XOR U33215 ( .A(n34444), .B(n34445), .Z(n34277) );
  XNOR U33216 ( .A(n34454), .B(n34455), .Z(n34445) );
  ANDN U33217 ( .B(n34456), .A(n34457), .Z(n34454) );
  XOR U33218 ( .A(n34458), .B(n34459), .Z(n34456) );
  XOR U33219 ( .A(n34460), .B(n34461), .Z(n34444) );
  XNOR U33220 ( .A(n34462), .B(n34463), .Z(n34461) );
  ANDN U33221 ( .B(n34464), .A(n34465), .Z(n34462) );
  XNOR U33222 ( .A(n34466), .B(n34467), .Z(n34464) );
  IV U33223 ( .A(n34442), .Z(n34460) );
  XOR U33224 ( .A(n34468), .B(n34469), .Z(n34442) );
  ANDN U33225 ( .B(n34470), .A(n34471), .Z(n34468) );
  XOR U33226 ( .A(n34469), .B(n34472), .Z(n34470) );
  XNOR U33227 ( .A(n34451), .B(n34279), .Z(n34452) );
  XOR U33228 ( .A(n34473), .B(n34474), .Z(n34279) );
  AND U33229 ( .A(n464), .B(n34475), .Z(n34473) );
  XOR U33230 ( .A(n34476), .B(n34474), .Z(n34475) );
  XNOR U33231 ( .A(n34477), .B(n34478), .Z(n34451) );
  AND U33232 ( .A(n34479), .B(n34480), .Z(n34477) );
  XNOR U33233 ( .A(n34478), .B(n34329), .Z(n34480) );
  XOR U33234 ( .A(n34471), .B(n34472), .Z(n34329) );
  XOR U33235 ( .A(n34481), .B(n34459), .Z(n34472) );
  XNOR U33236 ( .A(n34482), .B(n34483), .Z(n34459) );
  ANDN U33237 ( .B(n34484), .A(n34485), .Z(n34482) );
  XOR U33238 ( .A(n34486), .B(n34487), .Z(n34484) );
  IV U33239 ( .A(n34457), .Z(n34481) );
  XOR U33240 ( .A(n34455), .B(n34488), .Z(n34457) );
  XNOR U33241 ( .A(n34489), .B(n34490), .Z(n34488) );
  ANDN U33242 ( .B(n34491), .A(n34492), .Z(n34489) );
  XNOR U33243 ( .A(n34493), .B(n34494), .Z(n34491) );
  IV U33244 ( .A(n34458), .Z(n34455) );
  XOR U33245 ( .A(n34495), .B(n34496), .Z(n34458) );
  ANDN U33246 ( .B(n34497), .A(n34498), .Z(n34495) );
  XOR U33247 ( .A(n34496), .B(n34499), .Z(n34497) );
  XOR U33248 ( .A(n34500), .B(n34501), .Z(n34471) );
  XNOR U33249 ( .A(n34466), .B(n34502), .Z(n34501) );
  IV U33250 ( .A(n34469), .Z(n34502) );
  XOR U33251 ( .A(n34503), .B(n34504), .Z(n34469) );
  ANDN U33252 ( .B(n34505), .A(n34506), .Z(n34503) );
  XOR U33253 ( .A(n34504), .B(n34507), .Z(n34505) );
  XNOR U33254 ( .A(n34508), .B(n34509), .Z(n34466) );
  ANDN U33255 ( .B(n34510), .A(n34511), .Z(n34508) );
  XOR U33256 ( .A(n34509), .B(n34512), .Z(n34510) );
  IV U33257 ( .A(n34465), .Z(n34500) );
  XOR U33258 ( .A(n34463), .B(n34513), .Z(n34465) );
  XNOR U33259 ( .A(n34514), .B(n34515), .Z(n34513) );
  ANDN U33260 ( .B(n34516), .A(n34517), .Z(n34514) );
  XNOR U33261 ( .A(n34518), .B(n34519), .Z(n34516) );
  IV U33262 ( .A(n34467), .Z(n34463) );
  XOR U33263 ( .A(n34520), .B(n34521), .Z(n34467) );
  ANDN U33264 ( .B(n34522), .A(n34523), .Z(n34520) );
  XOR U33265 ( .A(n34524), .B(n34521), .Z(n34522) );
  XOR U33266 ( .A(n34478), .B(n34331), .Z(n34479) );
  XOR U33267 ( .A(n34525), .B(n34526), .Z(n34331) );
  AND U33268 ( .A(n464), .B(n34527), .Z(n34525) );
  XOR U33269 ( .A(n34528), .B(n34526), .Z(n34527) );
  XNOR U33270 ( .A(n34529), .B(n34530), .Z(n34478) );
  NAND U33271 ( .A(n34531), .B(n34532), .Z(n34530) );
  XOR U33272 ( .A(n34533), .B(n34430), .Z(n34532) );
  XOR U33273 ( .A(n34506), .B(n34507), .Z(n34430) );
  XOR U33274 ( .A(n34534), .B(n34499), .Z(n34507) );
  XOR U33275 ( .A(n34535), .B(n34487), .Z(n34499) );
  XOR U33276 ( .A(n34536), .B(n34537), .Z(n34487) );
  ANDN U33277 ( .B(n34538), .A(n34539), .Z(n34536) );
  XOR U33278 ( .A(n34537), .B(n34540), .Z(n34538) );
  IV U33279 ( .A(n34485), .Z(n34535) );
  XOR U33280 ( .A(n34483), .B(n34541), .Z(n34485) );
  XOR U33281 ( .A(n34542), .B(n34543), .Z(n34541) );
  ANDN U33282 ( .B(n34544), .A(n34545), .Z(n34542) );
  XOR U33283 ( .A(n34546), .B(n34543), .Z(n34544) );
  IV U33284 ( .A(n34486), .Z(n34483) );
  XOR U33285 ( .A(n34547), .B(n34548), .Z(n34486) );
  ANDN U33286 ( .B(n34549), .A(n34550), .Z(n34547) );
  XOR U33287 ( .A(n34548), .B(n34551), .Z(n34549) );
  IV U33288 ( .A(n34498), .Z(n34534) );
  XOR U33289 ( .A(n34552), .B(n34553), .Z(n34498) );
  XNOR U33290 ( .A(n34493), .B(n34554), .Z(n34553) );
  IV U33291 ( .A(n34496), .Z(n34554) );
  XOR U33292 ( .A(n34555), .B(n34556), .Z(n34496) );
  ANDN U33293 ( .B(n34557), .A(n34558), .Z(n34555) );
  XOR U33294 ( .A(n34556), .B(n34559), .Z(n34557) );
  XNOR U33295 ( .A(n34560), .B(n34561), .Z(n34493) );
  ANDN U33296 ( .B(n34562), .A(n34563), .Z(n34560) );
  XOR U33297 ( .A(n34561), .B(n34564), .Z(n34562) );
  IV U33298 ( .A(n34492), .Z(n34552) );
  XOR U33299 ( .A(n34490), .B(n34565), .Z(n34492) );
  XOR U33300 ( .A(n34566), .B(n34567), .Z(n34565) );
  ANDN U33301 ( .B(n34568), .A(n34569), .Z(n34566) );
  XOR U33302 ( .A(n34570), .B(n34567), .Z(n34568) );
  IV U33303 ( .A(n34494), .Z(n34490) );
  XOR U33304 ( .A(n34571), .B(n34572), .Z(n34494) );
  ANDN U33305 ( .B(n34573), .A(n34574), .Z(n34571) );
  XOR U33306 ( .A(n34575), .B(n34572), .Z(n34573) );
  XOR U33307 ( .A(n34576), .B(n34577), .Z(n34506) );
  XOR U33308 ( .A(n34524), .B(n34578), .Z(n34577) );
  IV U33309 ( .A(n34504), .Z(n34578) );
  XOR U33310 ( .A(n34579), .B(n34580), .Z(n34504) );
  ANDN U33311 ( .B(n34581), .A(n34582), .Z(n34579) );
  XOR U33312 ( .A(n34580), .B(n34583), .Z(n34581) );
  XOR U33313 ( .A(n34584), .B(n34512), .Z(n34524) );
  XOR U33314 ( .A(n34585), .B(n34586), .Z(n34512) );
  ANDN U33315 ( .B(n34587), .A(n34588), .Z(n34585) );
  XOR U33316 ( .A(n34586), .B(n34589), .Z(n34587) );
  IV U33317 ( .A(n34511), .Z(n34584) );
  XOR U33318 ( .A(n34590), .B(n34591), .Z(n34511) );
  XOR U33319 ( .A(n34592), .B(n34593), .Z(n34591) );
  ANDN U33320 ( .B(n34594), .A(n34595), .Z(n34592) );
  XOR U33321 ( .A(n34596), .B(n34593), .Z(n34594) );
  IV U33322 ( .A(n34509), .Z(n34590) );
  XOR U33323 ( .A(n34597), .B(n34598), .Z(n34509) );
  ANDN U33324 ( .B(n34599), .A(n34600), .Z(n34597) );
  XOR U33325 ( .A(n34598), .B(n34601), .Z(n34599) );
  IV U33326 ( .A(n34523), .Z(n34576) );
  XOR U33327 ( .A(n34602), .B(n34603), .Z(n34523) );
  XNOR U33328 ( .A(n34518), .B(n34604), .Z(n34603) );
  IV U33329 ( .A(n34521), .Z(n34604) );
  XOR U33330 ( .A(n34605), .B(n34606), .Z(n34521) );
  ANDN U33331 ( .B(n34607), .A(n34608), .Z(n34605) );
  XOR U33332 ( .A(n34609), .B(n34606), .Z(n34607) );
  XNOR U33333 ( .A(n34610), .B(n34611), .Z(n34518) );
  ANDN U33334 ( .B(n34612), .A(n34613), .Z(n34610) );
  XOR U33335 ( .A(n34611), .B(n34614), .Z(n34612) );
  IV U33336 ( .A(n34517), .Z(n34602) );
  XOR U33337 ( .A(n34515), .B(n34615), .Z(n34517) );
  XOR U33338 ( .A(n34616), .B(n34617), .Z(n34615) );
  ANDN U33339 ( .B(n34618), .A(n34619), .Z(n34616) );
  XOR U33340 ( .A(n34620), .B(n34617), .Z(n34618) );
  IV U33341 ( .A(n34519), .Z(n34515) );
  XOR U33342 ( .A(n34621), .B(n34622), .Z(n34519) );
  ANDN U33343 ( .B(n34623), .A(n34624), .Z(n34621) );
  XOR U33344 ( .A(n34625), .B(n34622), .Z(n34623) );
  IV U33345 ( .A(n34529), .Z(n34533) );
  XOR U33346 ( .A(n34529), .B(n34432), .Z(n34531) );
  XOR U33347 ( .A(n34626), .B(n34627), .Z(n34432) );
  AND U33348 ( .A(n464), .B(n34628), .Z(n34626) );
  XOR U33349 ( .A(n34629), .B(n34627), .Z(n34628) );
  NANDN U33350 ( .A(n34434), .B(n34436), .Z(n34529) );
  XOR U33351 ( .A(n34630), .B(n34631), .Z(n34436) );
  AND U33352 ( .A(n464), .B(n34632), .Z(n34630) );
  XOR U33353 ( .A(n34631), .B(n34633), .Z(n34632) );
  XNOR U33354 ( .A(n34634), .B(n34635), .Z(n464) );
  AND U33355 ( .A(n34636), .B(n34637), .Z(n34634) );
  XOR U33356 ( .A(n34635), .B(n34447), .Z(n34637) );
  XNOR U33357 ( .A(n34638), .B(n34639), .Z(n34447) );
  ANDN U33358 ( .B(n34640), .A(n34641), .Z(n34638) );
  XOR U33359 ( .A(n34639), .B(n34642), .Z(n34640) );
  XNOR U33360 ( .A(n34635), .B(n34449), .Z(n34636) );
  XOR U33361 ( .A(n34643), .B(n34644), .Z(n34449) );
  AND U33362 ( .A(n468), .B(n34645), .Z(n34643) );
  XOR U33363 ( .A(n34646), .B(n34644), .Z(n34645) );
  XOR U33364 ( .A(n34647), .B(n34648), .Z(n34635) );
  AND U33365 ( .A(n34649), .B(n34650), .Z(n34647) );
  XOR U33366 ( .A(n34648), .B(n34474), .Z(n34650) );
  XOR U33367 ( .A(n34641), .B(n34642), .Z(n34474) );
  XNOR U33368 ( .A(n34651), .B(n34652), .Z(n34642) );
  ANDN U33369 ( .B(n34653), .A(n34654), .Z(n34651) );
  XOR U33370 ( .A(n34655), .B(n34656), .Z(n34653) );
  XOR U33371 ( .A(n34657), .B(n34658), .Z(n34641) );
  XNOR U33372 ( .A(n34659), .B(n34660), .Z(n34658) );
  ANDN U33373 ( .B(n34661), .A(n34662), .Z(n34659) );
  XNOR U33374 ( .A(n34663), .B(n34664), .Z(n34661) );
  IV U33375 ( .A(n34639), .Z(n34657) );
  XOR U33376 ( .A(n34665), .B(n34666), .Z(n34639) );
  ANDN U33377 ( .B(n34667), .A(n34668), .Z(n34665) );
  XOR U33378 ( .A(n34666), .B(n34669), .Z(n34667) );
  XNOR U33379 ( .A(n34648), .B(n34476), .Z(n34649) );
  XOR U33380 ( .A(n34670), .B(n34671), .Z(n34476) );
  AND U33381 ( .A(n468), .B(n34672), .Z(n34670) );
  XOR U33382 ( .A(n34673), .B(n34671), .Z(n34672) );
  XNOR U33383 ( .A(n34674), .B(n34675), .Z(n34648) );
  AND U33384 ( .A(n34676), .B(n34677), .Z(n34674) );
  XNOR U33385 ( .A(n34675), .B(n34526), .Z(n34677) );
  XOR U33386 ( .A(n34668), .B(n34669), .Z(n34526) );
  XOR U33387 ( .A(n34678), .B(n34656), .Z(n34669) );
  XNOR U33388 ( .A(n34679), .B(n34680), .Z(n34656) );
  ANDN U33389 ( .B(n34681), .A(n34682), .Z(n34679) );
  XOR U33390 ( .A(n34683), .B(n34684), .Z(n34681) );
  IV U33391 ( .A(n34654), .Z(n34678) );
  XOR U33392 ( .A(n34652), .B(n34685), .Z(n34654) );
  XNOR U33393 ( .A(n34686), .B(n34687), .Z(n34685) );
  ANDN U33394 ( .B(n34688), .A(n34689), .Z(n34686) );
  XNOR U33395 ( .A(n34690), .B(n34691), .Z(n34688) );
  IV U33396 ( .A(n34655), .Z(n34652) );
  XOR U33397 ( .A(n34692), .B(n34693), .Z(n34655) );
  ANDN U33398 ( .B(n34694), .A(n34695), .Z(n34692) );
  XOR U33399 ( .A(n34693), .B(n34696), .Z(n34694) );
  XOR U33400 ( .A(n34697), .B(n34698), .Z(n34668) );
  XNOR U33401 ( .A(n34663), .B(n34699), .Z(n34698) );
  IV U33402 ( .A(n34666), .Z(n34699) );
  XOR U33403 ( .A(n34700), .B(n34701), .Z(n34666) );
  ANDN U33404 ( .B(n34702), .A(n34703), .Z(n34700) );
  XOR U33405 ( .A(n34701), .B(n34704), .Z(n34702) );
  XNOR U33406 ( .A(n34705), .B(n34706), .Z(n34663) );
  ANDN U33407 ( .B(n34707), .A(n34708), .Z(n34705) );
  XOR U33408 ( .A(n34706), .B(n34709), .Z(n34707) );
  IV U33409 ( .A(n34662), .Z(n34697) );
  XOR U33410 ( .A(n34660), .B(n34710), .Z(n34662) );
  XNOR U33411 ( .A(n34711), .B(n34712), .Z(n34710) );
  ANDN U33412 ( .B(n34713), .A(n34714), .Z(n34711) );
  XNOR U33413 ( .A(n34715), .B(n34716), .Z(n34713) );
  IV U33414 ( .A(n34664), .Z(n34660) );
  XOR U33415 ( .A(n34717), .B(n34718), .Z(n34664) );
  ANDN U33416 ( .B(n34719), .A(n34720), .Z(n34717) );
  XOR U33417 ( .A(n34721), .B(n34718), .Z(n34719) );
  XOR U33418 ( .A(n34675), .B(n34528), .Z(n34676) );
  XOR U33419 ( .A(n34722), .B(n34723), .Z(n34528) );
  AND U33420 ( .A(n468), .B(n34724), .Z(n34722) );
  XOR U33421 ( .A(n34725), .B(n34723), .Z(n34724) );
  XNOR U33422 ( .A(n34726), .B(n34727), .Z(n34675) );
  NAND U33423 ( .A(n34728), .B(n34729), .Z(n34727) );
  XOR U33424 ( .A(n34730), .B(n34627), .Z(n34729) );
  XOR U33425 ( .A(n34703), .B(n34704), .Z(n34627) );
  XOR U33426 ( .A(n34731), .B(n34696), .Z(n34704) );
  XOR U33427 ( .A(n34732), .B(n34684), .Z(n34696) );
  XOR U33428 ( .A(n34733), .B(n34734), .Z(n34684) );
  ANDN U33429 ( .B(n34735), .A(n34736), .Z(n34733) );
  XOR U33430 ( .A(n34734), .B(n34737), .Z(n34735) );
  IV U33431 ( .A(n34682), .Z(n34732) );
  XOR U33432 ( .A(n34680), .B(n34738), .Z(n34682) );
  XOR U33433 ( .A(n34739), .B(n34740), .Z(n34738) );
  ANDN U33434 ( .B(n34741), .A(n34742), .Z(n34739) );
  XOR U33435 ( .A(n34743), .B(n34740), .Z(n34741) );
  IV U33436 ( .A(n34683), .Z(n34680) );
  XOR U33437 ( .A(n34744), .B(n34745), .Z(n34683) );
  ANDN U33438 ( .B(n34746), .A(n34747), .Z(n34744) );
  XOR U33439 ( .A(n34745), .B(n34748), .Z(n34746) );
  IV U33440 ( .A(n34695), .Z(n34731) );
  XOR U33441 ( .A(n34749), .B(n34750), .Z(n34695) );
  XNOR U33442 ( .A(n34690), .B(n34751), .Z(n34750) );
  IV U33443 ( .A(n34693), .Z(n34751) );
  XOR U33444 ( .A(n34752), .B(n34753), .Z(n34693) );
  ANDN U33445 ( .B(n34754), .A(n34755), .Z(n34752) );
  XOR U33446 ( .A(n34753), .B(n34756), .Z(n34754) );
  XNOR U33447 ( .A(n34757), .B(n34758), .Z(n34690) );
  ANDN U33448 ( .B(n34759), .A(n34760), .Z(n34757) );
  XOR U33449 ( .A(n34758), .B(n34761), .Z(n34759) );
  IV U33450 ( .A(n34689), .Z(n34749) );
  XOR U33451 ( .A(n34687), .B(n34762), .Z(n34689) );
  XOR U33452 ( .A(n34763), .B(n34764), .Z(n34762) );
  ANDN U33453 ( .B(n34765), .A(n34766), .Z(n34763) );
  XOR U33454 ( .A(n34767), .B(n34764), .Z(n34765) );
  IV U33455 ( .A(n34691), .Z(n34687) );
  XOR U33456 ( .A(n34768), .B(n34769), .Z(n34691) );
  ANDN U33457 ( .B(n34770), .A(n34771), .Z(n34768) );
  XOR U33458 ( .A(n34772), .B(n34769), .Z(n34770) );
  XOR U33459 ( .A(n34773), .B(n34774), .Z(n34703) );
  XOR U33460 ( .A(n34721), .B(n34775), .Z(n34774) );
  IV U33461 ( .A(n34701), .Z(n34775) );
  XOR U33462 ( .A(n34776), .B(n34777), .Z(n34701) );
  ANDN U33463 ( .B(n34778), .A(n34779), .Z(n34776) );
  XOR U33464 ( .A(n34777), .B(n34780), .Z(n34778) );
  XOR U33465 ( .A(n34781), .B(n34709), .Z(n34721) );
  XOR U33466 ( .A(n34782), .B(n34783), .Z(n34709) );
  ANDN U33467 ( .B(n34784), .A(n34785), .Z(n34782) );
  XOR U33468 ( .A(n34783), .B(n34786), .Z(n34784) );
  IV U33469 ( .A(n34708), .Z(n34781) );
  XOR U33470 ( .A(n34787), .B(n34788), .Z(n34708) );
  XOR U33471 ( .A(n34789), .B(n34790), .Z(n34788) );
  ANDN U33472 ( .B(n34791), .A(n34792), .Z(n34789) );
  XOR U33473 ( .A(n34793), .B(n34790), .Z(n34791) );
  IV U33474 ( .A(n34706), .Z(n34787) );
  XOR U33475 ( .A(n34794), .B(n34795), .Z(n34706) );
  ANDN U33476 ( .B(n34796), .A(n34797), .Z(n34794) );
  XOR U33477 ( .A(n34795), .B(n34798), .Z(n34796) );
  IV U33478 ( .A(n34720), .Z(n34773) );
  XOR U33479 ( .A(n34799), .B(n34800), .Z(n34720) );
  XNOR U33480 ( .A(n34715), .B(n34801), .Z(n34800) );
  IV U33481 ( .A(n34718), .Z(n34801) );
  XOR U33482 ( .A(n34802), .B(n34803), .Z(n34718) );
  ANDN U33483 ( .B(n34804), .A(n34805), .Z(n34802) );
  XOR U33484 ( .A(n34806), .B(n34803), .Z(n34804) );
  XNOR U33485 ( .A(n34807), .B(n34808), .Z(n34715) );
  ANDN U33486 ( .B(n34809), .A(n34810), .Z(n34807) );
  XOR U33487 ( .A(n34808), .B(n34811), .Z(n34809) );
  IV U33488 ( .A(n34714), .Z(n34799) );
  XOR U33489 ( .A(n34712), .B(n34812), .Z(n34714) );
  XOR U33490 ( .A(n34813), .B(n34814), .Z(n34812) );
  ANDN U33491 ( .B(n34815), .A(n34816), .Z(n34813) );
  XOR U33492 ( .A(n34817), .B(n34814), .Z(n34815) );
  IV U33493 ( .A(n34716), .Z(n34712) );
  XOR U33494 ( .A(n34818), .B(n34819), .Z(n34716) );
  ANDN U33495 ( .B(n34820), .A(n34821), .Z(n34818) );
  XOR U33496 ( .A(n34822), .B(n34819), .Z(n34820) );
  IV U33497 ( .A(n34726), .Z(n34730) );
  XOR U33498 ( .A(n34726), .B(n34629), .Z(n34728) );
  XOR U33499 ( .A(n34823), .B(n34824), .Z(n34629) );
  AND U33500 ( .A(n468), .B(n34825), .Z(n34823) );
  XOR U33501 ( .A(n34826), .B(n34824), .Z(n34825) );
  NANDN U33502 ( .A(n34631), .B(n34633), .Z(n34726) );
  XOR U33503 ( .A(n34827), .B(n34828), .Z(n34633) );
  AND U33504 ( .A(n468), .B(n34829), .Z(n34827) );
  XOR U33505 ( .A(n34828), .B(n34830), .Z(n34829) );
  XNOR U33506 ( .A(n34831), .B(n34832), .Z(n468) );
  AND U33507 ( .A(n34833), .B(n34834), .Z(n34831) );
  XOR U33508 ( .A(n34832), .B(n34644), .Z(n34834) );
  XNOR U33509 ( .A(n34835), .B(n34836), .Z(n34644) );
  ANDN U33510 ( .B(n34837), .A(n34838), .Z(n34835) );
  XOR U33511 ( .A(n34836), .B(n34839), .Z(n34837) );
  XNOR U33512 ( .A(n34832), .B(n34646), .Z(n34833) );
  XOR U33513 ( .A(n34840), .B(n34841), .Z(n34646) );
  AND U33514 ( .A(n472), .B(n34842), .Z(n34840) );
  XOR U33515 ( .A(n34843), .B(n34841), .Z(n34842) );
  XOR U33516 ( .A(n34844), .B(n34845), .Z(n34832) );
  AND U33517 ( .A(n34846), .B(n34847), .Z(n34844) );
  XOR U33518 ( .A(n34845), .B(n34671), .Z(n34847) );
  XOR U33519 ( .A(n34838), .B(n34839), .Z(n34671) );
  XNOR U33520 ( .A(n34848), .B(n34849), .Z(n34839) );
  ANDN U33521 ( .B(n34850), .A(n34851), .Z(n34848) );
  XOR U33522 ( .A(n34852), .B(n34853), .Z(n34850) );
  XOR U33523 ( .A(n34854), .B(n34855), .Z(n34838) );
  XNOR U33524 ( .A(n34856), .B(n34857), .Z(n34855) );
  ANDN U33525 ( .B(n34858), .A(n34859), .Z(n34856) );
  XNOR U33526 ( .A(n34860), .B(n34861), .Z(n34858) );
  IV U33527 ( .A(n34836), .Z(n34854) );
  XOR U33528 ( .A(n34862), .B(n34863), .Z(n34836) );
  ANDN U33529 ( .B(n34864), .A(n34865), .Z(n34862) );
  XOR U33530 ( .A(n34863), .B(n34866), .Z(n34864) );
  XNOR U33531 ( .A(n34845), .B(n34673), .Z(n34846) );
  XOR U33532 ( .A(n34867), .B(n34868), .Z(n34673) );
  AND U33533 ( .A(n472), .B(n34869), .Z(n34867) );
  XOR U33534 ( .A(n34870), .B(n34868), .Z(n34869) );
  XNOR U33535 ( .A(n34871), .B(n34872), .Z(n34845) );
  AND U33536 ( .A(n34873), .B(n34874), .Z(n34871) );
  XNOR U33537 ( .A(n34872), .B(n34723), .Z(n34874) );
  XOR U33538 ( .A(n34865), .B(n34866), .Z(n34723) );
  XOR U33539 ( .A(n34875), .B(n34853), .Z(n34866) );
  XNOR U33540 ( .A(n34876), .B(n34877), .Z(n34853) );
  ANDN U33541 ( .B(n34878), .A(n34879), .Z(n34876) );
  XOR U33542 ( .A(n34880), .B(n34881), .Z(n34878) );
  IV U33543 ( .A(n34851), .Z(n34875) );
  XOR U33544 ( .A(n34849), .B(n34882), .Z(n34851) );
  XNOR U33545 ( .A(n34883), .B(n34884), .Z(n34882) );
  ANDN U33546 ( .B(n34885), .A(n34886), .Z(n34883) );
  XNOR U33547 ( .A(n34887), .B(n34888), .Z(n34885) );
  IV U33548 ( .A(n34852), .Z(n34849) );
  XOR U33549 ( .A(n34889), .B(n34890), .Z(n34852) );
  ANDN U33550 ( .B(n34891), .A(n34892), .Z(n34889) );
  XOR U33551 ( .A(n34890), .B(n34893), .Z(n34891) );
  XOR U33552 ( .A(n34894), .B(n34895), .Z(n34865) );
  XNOR U33553 ( .A(n34860), .B(n34896), .Z(n34895) );
  IV U33554 ( .A(n34863), .Z(n34896) );
  XOR U33555 ( .A(n34897), .B(n34898), .Z(n34863) );
  ANDN U33556 ( .B(n34899), .A(n34900), .Z(n34897) );
  XOR U33557 ( .A(n34898), .B(n34901), .Z(n34899) );
  XNOR U33558 ( .A(n34902), .B(n34903), .Z(n34860) );
  ANDN U33559 ( .B(n34904), .A(n34905), .Z(n34902) );
  XOR U33560 ( .A(n34903), .B(n34906), .Z(n34904) );
  IV U33561 ( .A(n34859), .Z(n34894) );
  XOR U33562 ( .A(n34857), .B(n34907), .Z(n34859) );
  XNOR U33563 ( .A(n34908), .B(n34909), .Z(n34907) );
  ANDN U33564 ( .B(n34910), .A(n34911), .Z(n34908) );
  XNOR U33565 ( .A(n34912), .B(n34913), .Z(n34910) );
  IV U33566 ( .A(n34861), .Z(n34857) );
  XOR U33567 ( .A(n34914), .B(n34915), .Z(n34861) );
  ANDN U33568 ( .B(n34916), .A(n34917), .Z(n34914) );
  XOR U33569 ( .A(n34918), .B(n34915), .Z(n34916) );
  XOR U33570 ( .A(n34872), .B(n34725), .Z(n34873) );
  XOR U33571 ( .A(n34919), .B(n34920), .Z(n34725) );
  AND U33572 ( .A(n472), .B(n34921), .Z(n34919) );
  XOR U33573 ( .A(n34922), .B(n34920), .Z(n34921) );
  XNOR U33574 ( .A(n34923), .B(n34924), .Z(n34872) );
  NAND U33575 ( .A(n34925), .B(n34926), .Z(n34924) );
  XOR U33576 ( .A(n34927), .B(n34824), .Z(n34926) );
  XOR U33577 ( .A(n34900), .B(n34901), .Z(n34824) );
  XOR U33578 ( .A(n34928), .B(n34893), .Z(n34901) );
  XOR U33579 ( .A(n34929), .B(n34881), .Z(n34893) );
  XOR U33580 ( .A(n34930), .B(n34931), .Z(n34881) );
  ANDN U33581 ( .B(n34932), .A(n34933), .Z(n34930) );
  XOR U33582 ( .A(n34931), .B(n34934), .Z(n34932) );
  IV U33583 ( .A(n34879), .Z(n34929) );
  XOR U33584 ( .A(n34877), .B(n34935), .Z(n34879) );
  XOR U33585 ( .A(n34936), .B(n34937), .Z(n34935) );
  ANDN U33586 ( .B(n34938), .A(n34939), .Z(n34936) );
  XOR U33587 ( .A(n34940), .B(n34937), .Z(n34938) );
  IV U33588 ( .A(n34880), .Z(n34877) );
  XOR U33589 ( .A(n34941), .B(n34942), .Z(n34880) );
  ANDN U33590 ( .B(n34943), .A(n34944), .Z(n34941) );
  XOR U33591 ( .A(n34942), .B(n34945), .Z(n34943) );
  IV U33592 ( .A(n34892), .Z(n34928) );
  XOR U33593 ( .A(n34946), .B(n34947), .Z(n34892) );
  XNOR U33594 ( .A(n34887), .B(n34948), .Z(n34947) );
  IV U33595 ( .A(n34890), .Z(n34948) );
  XOR U33596 ( .A(n34949), .B(n34950), .Z(n34890) );
  ANDN U33597 ( .B(n34951), .A(n34952), .Z(n34949) );
  XOR U33598 ( .A(n34950), .B(n34953), .Z(n34951) );
  XNOR U33599 ( .A(n34954), .B(n34955), .Z(n34887) );
  ANDN U33600 ( .B(n34956), .A(n34957), .Z(n34954) );
  XOR U33601 ( .A(n34955), .B(n34958), .Z(n34956) );
  IV U33602 ( .A(n34886), .Z(n34946) );
  XOR U33603 ( .A(n34884), .B(n34959), .Z(n34886) );
  XOR U33604 ( .A(n34960), .B(n34961), .Z(n34959) );
  ANDN U33605 ( .B(n34962), .A(n34963), .Z(n34960) );
  XOR U33606 ( .A(n34964), .B(n34961), .Z(n34962) );
  IV U33607 ( .A(n34888), .Z(n34884) );
  XOR U33608 ( .A(n34965), .B(n34966), .Z(n34888) );
  ANDN U33609 ( .B(n34967), .A(n34968), .Z(n34965) );
  XOR U33610 ( .A(n34969), .B(n34966), .Z(n34967) );
  XOR U33611 ( .A(n34970), .B(n34971), .Z(n34900) );
  XOR U33612 ( .A(n34918), .B(n34972), .Z(n34971) );
  IV U33613 ( .A(n34898), .Z(n34972) );
  XOR U33614 ( .A(n34973), .B(n34974), .Z(n34898) );
  ANDN U33615 ( .B(n34975), .A(n34976), .Z(n34973) );
  XOR U33616 ( .A(n34974), .B(n34977), .Z(n34975) );
  XOR U33617 ( .A(n34978), .B(n34906), .Z(n34918) );
  XOR U33618 ( .A(n34979), .B(n34980), .Z(n34906) );
  ANDN U33619 ( .B(n34981), .A(n34982), .Z(n34979) );
  XOR U33620 ( .A(n34980), .B(n34983), .Z(n34981) );
  IV U33621 ( .A(n34905), .Z(n34978) );
  XOR U33622 ( .A(n34984), .B(n34985), .Z(n34905) );
  XOR U33623 ( .A(n34986), .B(n34987), .Z(n34985) );
  ANDN U33624 ( .B(n34988), .A(n34989), .Z(n34986) );
  XOR U33625 ( .A(n34990), .B(n34987), .Z(n34988) );
  IV U33626 ( .A(n34903), .Z(n34984) );
  XOR U33627 ( .A(n34991), .B(n34992), .Z(n34903) );
  ANDN U33628 ( .B(n34993), .A(n34994), .Z(n34991) );
  XOR U33629 ( .A(n34992), .B(n34995), .Z(n34993) );
  IV U33630 ( .A(n34917), .Z(n34970) );
  XOR U33631 ( .A(n34996), .B(n34997), .Z(n34917) );
  XNOR U33632 ( .A(n34912), .B(n34998), .Z(n34997) );
  IV U33633 ( .A(n34915), .Z(n34998) );
  XOR U33634 ( .A(n34999), .B(n35000), .Z(n34915) );
  ANDN U33635 ( .B(n35001), .A(n35002), .Z(n34999) );
  XOR U33636 ( .A(n35003), .B(n35000), .Z(n35001) );
  XNOR U33637 ( .A(n35004), .B(n35005), .Z(n34912) );
  ANDN U33638 ( .B(n35006), .A(n35007), .Z(n35004) );
  XOR U33639 ( .A(n35005), .B(n35008), .Z(n35006) );
  IV U33640 ( .A(n34911), .Z(n34996) );
  XOR U33641 ( .A(n34909), .B(n35009), .Z(n34911) );
  XOR U33642 ( .A(n35010), .B(n35011), .Z(n35009) );
  ANDN U33643 ( .B(n35012), .A(n35013), .Z(n35010) );
  XOR U33644 ( .A(n35014), .B(n35011), .Z(n35012) );
  IV U33645 ( .A(n34913), .Z(n34909) );
  XOR U33646 ( .A(n35015), .B(n35016), .Z(n34913) );
  ANDN U33647 ( .B(n35017), .A(n35018), .Z(n35015) );
  XOR U33648 ( .A(n35019), .B(n35016), .Z(n35017) );
  IV U33649 ( .A(n34923), .Z(n34927) );
  XOR U33650 ( .A(n34923), .B(n34826), .Z(n34925) );
  XOR U33651 ( .A(n35020), .B(n35021), .Z(n34826) );
  AND U33652 ( .A(n472), .B(n35022), .Z(n35020) );
  XOR U33653 ( .A(n35023), .B(n35021), .Z(n35022) );
  NANDN U33654 ( .A(n34828), .B(n34830), .Z(n34923) );
  XOR U33655 ( .A(n35024), .B(n35025), .Z(n34830) );
  AND U33656 ( .A(n472), .B(n35026), .Z(n35024) );
  XOR U33657 ( .A(n35025), .B(n35027), .Z(n35026) );
  XNOR U33658 ( .A(n35028), .B(n35029), .Z(n472) );
  AND U33659 ( .A(n35030), .B(n35031), .Z(n35028) );
  XOR U33660 ( .A(n35029), .B(n34841), .Z(n35031) );
  XNOR U33661 ( .A(n35032), .B(n35033), .Z(n34841) );
  ANDN U33662 ( .B(n35034), .A(n35035), .Z(n35032) );
  XOR U33663 ( .A(n35033), .B(n35036), .Z(n35034) );
  XNOR U33664 ( .A(n35029), .B(n34843), .Z(n35030) );
  XOR U33665 ( .A(n35037), .B(n35038), .Z(n34843) );
  AND U33666 ( .A(n476), .B(n35039), .Z(n35037) );
  XOR U33667 ( .A(n35040), .B(n35038), .Z(n35039) );
  XOR U33668 ( .A(n35041), .B(n35042), .Z(n35029) );
  AND U33669 ( .A(n35043), .B(n35044), .Z(n35041) );
  XOR U33670 ( .A(n35042), .B(n34868), .Z(n35044) );
  XOR U33671 ( .A(n35035), .B(n35036), .Z(n34868) );
  XNOR U33672 ( .A(n35045), .B(n35046), .Z(n35036) );
  ANDN U33673 ( .B(n35047), .A(n35048), .Z(n35045) );
  XOR U33674 ( .A(n35049), .B(n35050), .Z(n35047) );
  XOR U33675 ( .A(n35051), .B(n35052), .Z(n35035) );
  XNOR U33676 ( .A(n35053), .B(n35054), .Z(n35052) );
  ANDN U33677 ( .B(n35055), .A(n35056), .Z(n35053) );
  XNOR U33678 ( .A(n35057), .B(n35058), .Z(n35055) );
  IV U33679 ( .A(n35033), .Z(n35051) );
  XOR U33680 ( .A(n35059), .B(n35060), .Z(n35033) );
  ANDN U33681 ( .B(n35061), .A(n35062), .Z(n35059) );
  XOR U33682 ( .A(n35060), .B(n35063), .Z(n35061) );
  XNOR U33683 ( .A(n35042), .B(n34870), .Z(n35043) );
  XOR U33684 ( .A(n35064), .B(n35065), .Z(n34870) );
  AND U33685 ( .A(n476), .B(n35066), .Z(n35064) );
  XOR U33686 ( .A(n35067), .B(n35065), .Z(n35066) );
  XNOR U33687 ( .A(n35068), .B(n35069), .Z(n35042) );
  AND U33688 ( .A(n35070), .B(n35071), .Z(n35068) );
  XNOR U33689 ( .A(n35069), .B(n34920), .Z(n35071) );
  XOR U33690 ( .A(n35062), .B(n35063), .Z(n34920) );
  XOR U33691 ( .A(n35072), .B(n35050), .Z(n35063) );
  XNOR U33692 ( .A(n35073), .B(n35074), .Z(n35050) );
  ANDN U33693 ( .B(n35075), .A(n35076), .Z(n35073) );
  XOR U33694 ( .A(n35077), .B(n35078), .Z(n35075) );
  IV U33695 ( .A(n35048), .Z(n35072) );
  XOR U33696 ( .A(n35046), .B(n35079), .Z(n35048) );
  XNOR U33697 ( .A(n35080), .B(n35081), .Z(n35079) );
  ANDN U33698 ( .B(n35082), .A(n35083), .Z(n35080) );
  XNOR U33699 ( .A(n35084), .B(n35085), .Z(n35082) );
  IV U33700 ( .A(n35049), .Z(n35046) );
  XOR U33701 ( .A(n35086), .B(n35087), .Z(n35049) );
  ANDN U33702 ( .B(n35088), .A(n35089), .Z(n35086) );
  XOR U33703 ( .A(n35087), .B(n35090), .Z(n35088) );
  XOR U33704 ( .A(n35091), .B(n35092), .Z(n35062) );
  XNOR U33705 ( .A(n35057), .B(n35093), .Z(n35092) );
  IV U33706 ( .A(n35060), .Z(n35093) );
  XOR U33707 ( .A(n35094), .B(n35095), .Z(n35060) );
  ANDN U33708 ( .B(n35096), .A(n35097), .Z(n35094) );
  XOR U33709 ( .A(n35095), .B(n35098), .Z(n35096) );
  XNOR U33710 ( .A(n35099), .B(n35100), .Z(n35057) );
  ANDN U33711 ( .B(n35101), .A(n35102), .Z(n35099) );
  XOR U33712 ( .A(n35100), .B(n35103), .Z(n35101) );
  IV U33713 ( .A(n35056), .Z(n35091) );
  XOR U33714 ( .A(n35054), .B(n35104), .Z(n35056) );
  XNOR U33715 ( .A(n35105), .B(n35106), .Z(n35104) );
  ANDN U33716 ( .B(n35107), .A(n35108), .Z(n35105) );
  XNOR U33717 ( .A(n35109), .B(n35110), .Z(n35107) );
  IV U33718 ( .A(n35058), .Z(n35054) );
  XOR U33719 ( .A(n35111), .B(n35112), .Z(n35058) );
  ANDN U33720 ( .B(n35113), .A(n35114), .Z(n35111) );
  XOR U33721 ( .A(n35115), .B(n35112), .Z(n35113) );
  XOR U33722 ( .A(n35069), .B(n34922), .Z(n35070) );
  XOR U33723 ( .A(n35116), .B(n35117), .Z(n34922) );
  AND U33724 ( .A(n476), .B(n35118), .Z(n35116) );
  XOR U33725 ( .A(n35119), .B(n35117), .Z(n35118) );
  XNOR U33726 ( .A(n35120), .B(n35121), .Z(n35069) );
  NAND U33727 ( .A(n35122), .B(n35123), .Z(n35121) );
  XOR U33728 ( .A(n35124), .B(n35021), .Z(n35123) );
  XOR U33729 ( .A(n35097), .B(n35098), .Z(n35021) );
  XOR U33730 ( .A(n35125), .B(n35090), .Z(n35098) );
  XOR U33731 ( .A(n35126), .B(n35078), .Z(n35090) );
  XOR U33732 ( .A(n35127), .B(n35128), .Z(n35078) );
  ANDN U33733 ( .B(n35129), .A(n35130), .Z(n35127) );
  XOR U33734 ( .A(n35128), .B(n35131), .Z(n35129) );
  IV U33735 ( .A(n35076), .Z(n35126) );
  XOR U33736 ( .A(n35074), .B(n35132), .Z(n35076) );
  XOR U33737 ( .A(n35133), .B(n35134), .Z(n35132) );
  ANDN U33738 ( .B(n35135), .A(n35136), .Z(n35133) );
  XOR U33739 ( .A(n35137), .B(n35134), .Z(n35135) );
  IV U33740 ( .A(n35077), .Z(n35074) );
  XOR U33741 ( .A(n35138), .B(n35139), .Z(n35077) );
  ANDN U33742 ( .B(n35140), .A(n35141), .Z(n35138) );
  XOR U33743 ( .A(n35139), .B(n35142), .Z(n35140) );
  IV U33744 ( .A(n35089), .Z(n35125) );
  XOR U33745 ( .A(n35143), .B(n35144), .Z(n35089) );
  XNOR U33746 ( .A(n35084), .B(n35145), .Z(n35144) );
  IV U33747 ( .A(n35087), .Z(n35145) );
  XOR U33748 ( .A(n35146), .B(n35147), .Z(n35087) );
  ANDN U33749 ( .B(n35148), .A(n35149), .Z(n35146) );
  XOR U33750 ( .A(n35147), .B(n35150), .Z(n35148) );
  XNOR U33751 ( .A(n35151), .B(n35152), .Z(n35084) );
  ANDN U33752 ( .B(n35153), .A(n35154), .Z(n35151) );
  XOR U33753 ( .A(n35152), .B(n35155), .Z(n35153) );
  IV U33754 ( .A(n35083), .Z(n35143) );
  XOR U33755 ( .A(n35081), .B(n35156), .Z(n35083) );
  XOR U33756 ( .A(n35157), .B(n35158), .Z(n35156) );
  ANDN U33757 ( .B(n35159), .A(n35160), .Z(n35157) );
  XOR U33758 ( .A(n35161), .B(n35158), .Z(n35159) );
  IV U33759 ( .A(n35085), .Z(n35081) );
  XOR U33760 ( .A(n35162), .B(n35163), .Z(n35085) );
  ANDN U33761 ( .B(n35164), .A(n35165), .Z(n35162) );
  XOR U33762 ( .A(n35166), .B(n35163), .Z(n35164) );
  XOR U33763 ( .A(n35167), .B(n35168), .Z(n35097) );
  XOR U33764 ( .A(n35115), .B(n35169), .Z(n35168) );
  IV U33765 ( .A(n35095), .Z(n35169) );
  XOR U33766 ( .A(n35170), .B(n35171), .Z(n35095) );
  ANDN U33767 ( .B(n35172), .A(n35173), .Z(n35170) );
  XOR U33768 ( .A(n35171), .B(n35174), .Z(n35172) );
  XOR U33769 ( .A(n35175), .B(n35103), .Z(n35115) );
  XOR U33770 ( .A(n35176), .B(n35177), .Z(n35103) );
  ANDN U33771 ( .B(n35178), .A(n35179), .Z(n35176) );
  XOR U33772 ( .A(n35177), .B(n35180), .Z(n35178) );
  IV U33773 ( .A(n35102), .Z(n35175) );
  XOR U33774 ( .A(n35181), .B(n35182), .Z(n35102) );
  XOR U33775 ( .A(n35183), .B(n35184), .Z(n35182) );
  ANDN U33776 ( .B(n35185), .A(n35186), .Z(n35183) );
  XOR U33777 ( .A(n35187), .B(n35184), .Z(n35185) );
  IV U33778 ( .A(n35100), .Z(n35181) );
  XOR U33779 ( .A(n35188), .B(n35189), .Z(n35100) );
  ANDN U33780 ( .B(n35190), .A(n35191), .Z(n35188) );
  XOR U33781 ( .A(n35189), .B(n35192), .Z(n35190) );
  IV U33782 ( .A(n35114), .Z(n35167) );
  XOR U33783 ( .A(n35193), .B(n35194), .Z(n35114) );
  XNOR U33784 ( .A(n35109), .B(n35195), .Z(n35194) );
  IV U33785 ( .A(n35112), .Z(n35195) );
  XOR U33786 ( .A(n35196), .B(n35197), .Z(n35112) );
  ANDN U33787 ( .B(n35198), .A(n35199), .Z(n35196) );
  XOR U33788 ( .A(n35200), .B(n35197), .Z(n35198) );
  XNOR U33789 ( .A(n35201), .B(n35202), .Z(n35109) );
  ANDN U33790 ( .B(n35203), .A(n35204), .Z(n35201) );
  XOR U33791 ( .A(n35202), .B(n35205), .Z(n35203) );
  IV U33792 ( .A(n35108), .Z(n35193) );
  XOR U33793 ( .A(n35106), .B(n35206), .Z(n35108) );
  XOR U33794 ( .A(n35207), .B(n35208), .Z(n35206) );
  ANDN U33795 ( .B(n35209), .A(n35210), .Z(n35207) );
  XOR U33796 ( .A(n35211), .B(n35208), .Z(n35209) );
  IV U33797 ( .A(n35110), .Z(n35106) );
  XOR U33798 ( .A(n35212), .B(n35213), .Z(n35110) );
  ANDN U33799 ( .B(n35214), .A(n35215), .Z(n35212) );
  XOR U33800 ( .A(n35216), .B(n35213), .Z(n35214) );
  IV U33801 ( .A(n35120), .Z(n35124) );
  XOR U33802 ( .A(n35120), .B(n35023), .Z(n35122) );
  XOR U33803 ( .A(n35217), .B(n35218), .Z(n35023) );
  AND U33804 ( .A(n476), .B(n35219), .Z(n35217) );
  XOR U33805 ( .A(n35220), .B(n35218), .Z(n35219) );
  NANDN U33806 ( .A(n35025), .B(n35027), .Z(n35120) );
  XOR U33807 ( .A(n35221), .B(n35222), .Z(n35027) );
  AND U33808 ( .A(n476), .B(n35223), .Z(n35221) );
  XOR U33809 ( .A(n35222), .B(n35224), .Z(n35223) );
  XNOR U33810 ( .A(n35225), .B(n35226), .Z(n476) );
  AND U33811 ( .A(n35227), .B(n35228), .Z(n35225) );
  XOR U33812 ( .A(n35226), .B(n35038), .Z(n35228) );
  XNOR U33813 ( .A(n35229), .B(n35230), .Z(n35038) );
  ANDN U33814 ( .B(n35231), .A(n35232), .Z(n35229) );
  XOR U33815 ( .A(n35230), .B(n35233), .Z(n35231) );
  XNOR U33816 ( .A(n35226), .B(n35040), .Z(n35227) );
  XOR U33817 ( .A(n35234), .B(n35235), .Z(n35040) );
  AND U33818 ( .A(n480), .B(n35236), .Z(n35234) );
  XOR U33819 ( .A(n35237), .B(n35235), .Z(n35236) );
  XOR U33820 ( .A(n35238), .B(n35239), .Z(n35226) );
  AND U33821 ( .A(n35240), .B(n35241), .Z(n35238) );
  XOR U33822 ( .A(n35239), .B(n35065), .Z(n35241) );
  XOR U33823 ( .A(n35232), .B(n35233), .Z(n35065) );
  XNOR U33824 ( .A(n35242), .B(n35243), .Z(n35233) );
  ANDN U33825 ( .B(n35244), .A(n35245), .Z(n35242) );
  XOR U33826 ( .A(n35246), .B(n35247), .Z(n35244) );
  XOR U33827 ( .A(n35248), .B(n35249), .Z(n35232) );
  XNOR U33828 ( .A(n35250), .B(n35251), .Z(n35249) );
  ANDN U33829 ( .B(n35252), .A(n35253), .Z(n35250) );
  XNOR U33830 ( .A(n35254), .B(n35255), .Z(n35252) );
  IV U33831 ( .A(n35230), .Z(n35248) );
  XOR U33832 ( .A(n35256), .B(n35257), .Z(n35230) );
  ANDN U33833 ( .B(n35258), .A(n35259), .Z(n35256) );
  XOR U33834 ( .A(n35257), .B(n35260), .Z(n35258) );
  XNOR U33835 ( .A(n35239), .B(n35067), .Z(n35240) );
  XOR U33836 ( .A(n35261), .B(n35262), .Z(n35067) );
  AND U33837 ( .A(n480), .B(n35263), .Z(n35261) );
  XOR U33838 ( .A(n35264), .B(n35262), .Z(n35263) );
  XNOR U33839 ( .A(n35265), .B(n35266), .Z(n35239) );
  AND U33840 ( .A(n35267), .B(n35268), .Z(n35265) );
  XNOR U33841 ( .A(n35266), .B(n35117), .Z(n35268) );
  XOR U33842 ( .A(n35259), .B(n35260), .Z(n35117) );
  XOR U33843 ( .A(n35269), .B(n35247), .Z(n35260) );
  XNOR U33844 ( .A(n35270), .B(n35271), .Z(n35247) );
  ANDN U33845 ( .B(n35272), .A(n35273), .Z(n35270) );
  XOR U33846 ( .A(n35274), .B(n35275), .Z(n35272) );
  IV U33847 ( .A(n35245), .Z(n35269) );
  XOR U33848 ( .A(n35243), .B(n35276), .Z(n35245) );
  XNOR U33849 ( .A(n35277), .B(n35278), .Z(n35276) );
  ANDN U33850 ( .B(n35279), .A(n35280), .Z(n35277) );
  XNOR U33851 ( .A(n35281), .B(n35282), .Z(n35279) );
  IV U33852 ( .A(n35246), .Z(n35243) );
  XOR U33853 ( .A(n35283), .B(n35284), .Z(n35246) );
  ANDN U33854 ( .B(n35285), .A(n35286), .Z(n35283) );
  XOR U33855 ( .A(n35284), .B(n35287), .Z(n35285) );
  XOR U33856 ( .A(n35288), .B(n35289), .Z(n35259) );
  XNOR U33857 ( .A(n35254), .B(n35290), .Z(n35289) );
  IV U33858 ( .A(n35257), .Z(n35290) );
  XOR U33859 ( .A(n35291), .B(n35292), .Z(n35257) );
  ANDN U33860 ( .B(n35293), .A(n35294), .Z(n35291) );
  XOR U33861 ( .A(n35292), .B(n35295), .Z(n35293) );
  XNOR U33862 ( .A(n35296), .B(n35297), .Z(n35254) );
  ANDN U33863 ( .B(n35298), .A(n35299), .Z(n35296) );
  XOR U33864 ( .A(n35297), .B(n35300), .Z(n35298) );
  IV U33865 ( .A(n35253), .Z(n35288) );
  XOR U33866 ( .A(n35251), .B(n35301), .Z(n35253) );
  XNOR U33867 ( .A(n35302), .B(n35303), .Z(n35301) );
  ANDN U33868 ( .B(n35304), .A(n35305), .Z(n35302) );
  XNOR U33869 ( .A(n35306), .B(n35307), .Z(n35304) );
  IV U33870 ( .A(n35255), .Z(n35251) );
  XOR U33871 ( .A(n35308), .B(n35309), .Z(n35255) );
  ANDN U33872 ( .B(n35310), .A(n35311), .Z(n35308) );
  XOR U33873 ( .A(n35312), .B(n35309), .Z(n35310) );
  XOR U33874 ( .A(n35266), .B(n35119), .Z(n35267) );
  XOR U33875 ( .A(n35313), .B(n35314), .Z(n35119) );
  AND U33876 ( .A(n480), .B(n35315), .Z(n35313) );
  XOR U33877 ( .A(n35316), .B(n35314), .Z(n35315) );
  XNOR U33878 ( .A(n35317), .B(n35318), .Z(n35266) );
  NAND U33879 ( .A(n35319), .B(n35320), .Z(n35318) );
  XOR U33880 ( .A(n35321), .B(n35218), .Z(n35320) );
  XOR U33881 ( .A(n35294), .B(n35295), .Z(n35218) );
  XOR U33882 ( .A(n35322), .B(n35287), .Z(n35295) );
  XOR U33883 ( .A(n35323), .B(n35275), .Z(n35287) );
  XOR U33884 ( .A(n35324), .B(n35325), .Z(n35275) );
  ANDN U33885 ( .B(n35326), .A(n35327), .Z(n35324) );
  XOR U33886 ( .A(n35325), .B(n35328), .Z(n35326) );
  IV U33887 ( .A(n35273), .Z(n35323) );
  XOR U33888 ( .A(n35271), .B(n35329), .Z(n35273) );
  XOR U33889 ( .A(n35330), .B(n35331), .Z(n35329) );
  ANDN U33890 ( .B(n35332), .A(n35333), .Z(n35330) );
  XOR U33891 ( .A(n35334), .B(n35331), .Z(n35332) );
  IV U33892 ( .A(n35274), .Z(n35271) );
  XOR U33893 ( .A(n35335), .B(n35336), .Z(n35274) );
  ANDN U33894 ( .B(n35337), .A(n35338), .Z(n35335) );
  XOR U33895 ( .A(n35336), .B(n35339), .Z(n35337) );
  IV U33896 ( .A(n35286), .Z(n35322) );
  XOR U33897 ( .A(n35340), .B(n35341), .Z(n35286) );
  XNOR U33898 ( .A(n35281), .B(n35342), .Z(n35341) );
  IV U33899 ( .A(n35284), .Z(n35342) );
  XOR U33900 ( .A(n35343), .B(n35344), .Z(n35284) );
  ANDN U33901 ( .B(n35345), .A(n35346), .Z(n35343) );
  XOR U33902 ( .A(n35344), .B(n35347), .Z(n35345) );
  XNOR U33903 ( .A(n35348), .B(n35349), .Z(n35281) );
  ANDN U33904 ( .B(n35350), .A(n35351), .Z(n35348) );
  XOR U33905 ( .A(n35349), .B(n35352), .Z(n35350) );
  IV U33906 ( .A(n35280), .Z(n35340) );
  XOR U33907 ( .A(n35278), .B(n35353), .Z(n35280) );
  XOR U33908 ( .A(n35354), .B(n35355), .Z(n35353) );
  ANDN U33909 ( .B(n35356), .A(n35357), .Z(n35354) );
  XOR U33910 ( .A(n35358), .B(n35355), .Z(n35356) );
  IV U33911 ( .A(n35282), .Z(n35278) );
  XOR U33912 ( .A(n35359), .B(n35360), .Z(n35282) );
  ANDN U33913 ( .B(n35361), .A(n35362), .Z(n35359) );
  XOR U33914 ( .A(n35363), .B(n35360), .Z(n35361) );
  XOR U33915 ( .A(n35364), .B(n35365), .Z(n35294) );
  XOR U33916 ( .A(n35312), .B(n35366), .Z(n35365) );
  IV U33917 ( .A(n35292), .Z(n35366) );
  XOR U33918 ( .A(n35367), .B(n35368), .Z(n35292) );
  ANDN U33919 ( .B(n35369), .A(n35370), .Z(n35367) );
  XOR U33920 ( .A(n35368), .B(n35371), .Z(n35369) );
  XOR U33921 ( .A(n35372), .B(n35300), .Z(n35312) );
  XOR U33922 ( .A(n35373), .B(n35374), .Z(n35300) );
  ANDN U33923 ( .B(n35375), .A(n35376), .Z(n35373) );
  XOR U33924 ( .A(n35374), .B(n35377), .Z(n35375) );
  IV U33925 ( .A(n35299), .Z(n35372) );
  XOR U33926 ( .A(n35378), .B(n35379), .Z(n35299) );
  XOR U33927 ( .A(n35380), .B(n35381), .Z(n35379) );
  ANDN U33928 ( .B(n35382), .A(n35383), .Z(n35380) );
  XOR U33929 ( .A(n35384), .B(n35381), .Z(n35382) );
  IV U33930 ( .A(n35297), .Z(n35378) );
  XOR U33931 ( .A(n35385), .B(n35386), .Z(n35297) );
  ANDN U33932 ( .B(n35387), .A(n35388), .Z(n35385) );
  XOR U33933 ( .A(n35386), .B(n35389), .Z(n35387) );
  IV U33934 ( .A(n35311), .Z(n35364) );
  XOR U33935 ( .A(n35390), .B(n35391), .Z(n35311) );
  XNOR U33936 ( .A(n35306), .B(n35392), .Z(n35391) );
  IV U33937 ( .A(n35309), .Z(n35392) );
  XOR U33938 ( .A(n35393), .B(n35394), .Z(n35309) );
  ANDN U33939 ( .B(n35395), .A(n35396), .Z(n35393) );
  XOR U33940 ( .A(n35397), .B(n35394), .Z(n35395) );
  XNOR U33941 ( .A(n35398), .B(n35399), .Z(n35306) );
  ANDN U33942 ( .B(n35400), .A(n35401), .Z(n35398) );
  XOR U33943 ( .A(n35399), .B(n35402), .Z(n35400) );
  IV U33944 ( .A(n35305), .Z(n35390) );
  XOR U33945 ( .A(n35303), .B(n35403), .Z(n35305) );
  XOR U33946 ( .A(n35404), .B(n35405), .Z(n35403) );
  ANDN U33947 ( .B(n35406), .A(n35407), .Z(n35404) );
  XOR U33948 ( .A(n35408), .B(n35405), .Z(n35406) );
  IV U33949 ( .A(n35307), .Z(n35303) );
  XOR U33950 ( .A(n35409), .B(n35410), .Z(n35307) );
  ANDN U33951 ( .B(n35411), .A(n35412), .Z(n35409) );
  XOR U33952 ( .A(n35413), .B(n35410), .Z(n35411) );
  IV U33953 ( .A(n35317), .Z(n35321) );
  XOR U33954 ( .A(n35317), .B(n35220), .Z(n35319) );
  XOR U33955 ( .A(n35414), .B(n35415), .Z(n35220) );
  AND U33956 ( .A(n480), .B(n35416), .Z(n35414) );
  XOR U33957 ( .A(n35417), .B(n35415), .Z(n35416) );
  NANDN U33958 ( .A(n35222), .B(n35224), .Z(n35317) );
  XOR U33959 ( .A(n35418), .B(n35419), .Z(n35224) );
  AND U33960 ( .A(n480), .B(n35420), .Z(n35418) );
  XOR U33961 ( .A(n35419), .B(n35421), .Z(n35420) );
  XNOR U33962 ( .A(n35422), .B(n35423), .Z(n480) );
  AND U33963 ( .A(n35424), .B(n35425), .Z(n35422) );
  XOR U33964 ( .A(n35423), .B(n35235), .Z(n35425) );
  XNOR U33965 ( .A(n35426), .B(n35427), .Z(n35235) );
  ANDN U33966 ( .B(n35428), .A(n35429), .Z(n35426) );
  XOR U33967 ( .A(n35427), .B(n35430), .Z(n35428) );
  XNOR U33968 ( .A(n35423), .B(n35237), .Z(n35424) );
  XOR U33969 ( .A(n35431), .B(n35432), .Z(n35237) );
  AND U33970 ( .A(n484), .B(n35433), .Z(n35431) );
  XOR U33971 ( .A(n35434), .B(n35432), .Z(n35433) );
  XOR U33972 ( .A(n35435), .B(n35436), .Z(n35423) );
  AND U33973 ( .A(n35437), .B(n35438), .Z(n35435) );
  XOR U33974 ( .A(n35436), .B(n35262), .Z(n35438) );
  XOR U33975 ( .A(n35429), .B(n35430), .Z(n35262) );
  XNOR U33976 ( .A(n35439), .B(n35440), .Z(n35430) );
  ANDN U33977 ( .B(n35441), .A(n35442), .Z(n35439) );
  XOR U33978 ( .A(n35443), .B(n35444), .Z(n35441) );
  XOR U33979 ( .A(n35445), .B(n35446), .Z(n35429) );
  XNOR U33980 ( .A(n35447), .B(n35448), .Z(n35446) );
  ANDN U33981 ( .B(n35449), .A(n35450), .Z(n35447) );
  XNOR U33982 ( .A(n35451), .B(n35452), .Z(n35449) );
  IV U33983 ( .A(n35427), .Z(n35445) );
  XOR U33984 ( .A(n35453), .B(n35454), .Z(n35427) );
  ANDN U33985 ( .B(n35455), .A(n35456), .Z(n35453) );
  XOR U33986 ( .A(n35454), .B(n35457), .Z(n35455) );
  XNOR U33987 ( .A(n35436), .B(n35264), .Z(n35437) );
  XOR U33988 ( .A(n35458), .B(n35459), .Z(n35264) );
  AND U33989 ( .A(n484), .B(n35460), .Z(n35458) );
  XOR U33990 ( .A(n35461), .B(n35459), .Z(n35460) );
  XNOR U33991 ( .A(n35462), .B(n35463), .Z(n35436) );
  AND U33992 ( .A(n35464), .B(n35465), .Z(n35462) );
  XNOR U33993 ( .A(n35463), .B(n35314), .Z(n35465) );
  XOR U33994 ( .A(n35456), .B(n35457), .Z(n35314) );
  XOR U33995 ( .A(n35466), .B(n35444), .Z(n35457) );
  XNOR U33996 ( .A(n35467), .B(n35468), .Z(n35444) );
  ANDN U33997 ( .B(n35469), .A(n35470), .Z(n35467) );
  XOR U33998 ( .A(n35471), .B(n35472), .Z(n35469) );
  IV U33999 ( .A(n35442), .Z(n35466) );
  XOR U34000 ( .A(n35440), .B(n35473), .Z(n35442) );
  XNOR U34001 ( .A(n35474), .B(n35475), .Z(n35473) );
  ANDN U34002 ( .B(n35476), .A(n35477), .Z(n35474) );
  XNOR U34003 ( .A(n35478), .B(n35479), .Z(n35476) );
  IV U34004 ( .A(n35443), .Z(n35440) );
  XOR U34005 ( .A(n35480), .B(n35481), .Z(n35443) );
  ANDN U34006 ( .B(n35482), .A(n35483), .Z(n35480) );
  XOR U34007 ( .A(n35481), .B(n35484), .Z(n35482) );
  XOR U34008 ( .A(n35485), .B(n35486), .Z(n35456) );
  XNOR U34009 ( .A(n35451), .B(n35487), .Z(n35486) );
  IV U34010 ( .A(n35454), .Z(n35487) );
  XOR U34011 ( .A(n35488), .B(n35489), .Z(n35454) );
  ANDN U34012 ( .B(n35490), .A(n35491), .Z(n35488) );
  XOR U34013 ( .A(n35489), .B(n35492), .Z(n35490) );
  XNOR U34014 ( .A(n35493), .B(n35494), .Z(n35451) );
  ANDN U34015 ( .B(n35495), .A(n35496), .Z(n35493) );
  XOR U34016 ( .A(n35494), .B(n35497), .Z(n35495) );
  IV U34017 ( .A(n35450), .Z(n35485) );
  XOR U34018 ( .A(n35448), .B(n35498), .Z(n35450) );
  XNOR U34019 ( .A(n35499), .B(n35500), .Z(n35498) );
  ANDN U34020 ( .B(n35501), .A(n35502), .Z(n35499) );
  XNOR U34021 ( .A(n35503), .B(n35504), .Z(n35501) );
  IV U34022 ( .A(n35452), .Z(n35448) );
  XOR U34023 ( .A(n35505), .B(n35506), .Z(n35452) );
  ANDN U34024 ( .B(n35507), .A(n35508), .Z(n35505) );
  XOR U34025 ( .A(n35509), .B(n35506), .Z(n35507) );
  XOR U34026 ( .A(n35463), .B(n35316), .Z(n35464) );
  XOR U34027 ( .A(n35510), .B(n35511), .Z(n35316) );
  AND U34028 ( .A(n484), .B(n35512), .Z(n35510) );
  XOR U34029 ( .A(n35513), .B(n35511), .Z(n35512) );
  XNOR U34030 ( .A(n35514), .B(n35515), .Z(n35463) );
  NAND U34031 ( .A(n35516), .B(n35517), .Z(n35515) );
  XOR U34032 ( .A(n35518), .B(n35415), .Z(n35517) );
  XOR U34033 ( .A(n35491), .B(n35492), .Z(n35415) );
  XOR U34034 ( .A(n35519), .B(n35484), .Z(n35492) );
  XOR U34035 ( .A(n35520), .B(n35472), .Z(n35484) );
  XOR U34036 ( .A(n35521), .B(n35522), .Z(n35472) );
  ANDN U34037 ( .B(n35523), .A(n35524), .Z(n35521) );
  XOR U34038 ( .A(n35522), .B(n35525), .Z(n35523) );
  IV U34039 ( .A(n35470), .Z(n35520) );
  XOR U34040 ( .A(n35468), .B(n35526), .Z(n35470) );
  XOR U34041 ( .A(n35527), .B(n35528), .Z(n35526) );
  ANDN U34042 ( .B(n35529), .A(n35530), .Z(n35527) );
  XOR U34043 ( .A(n35531), .B(n35528), .Z(n35529) );
  IV U34044 ( .A(n35471), .Z(n35468) );
  XOR U34045 ( .A(n35532), .B(n35533), .Z(n35471) );
  ANDN U34046 ( .B(n35534), .A(n35535), .Z(n35532) );
  XOR U34047 ( .A(n35533), .B(n35536), .Z(n35534) );
  IV U34048 ( .A(n35483), .Z(n35519) );
  XOR U34049 ( .A(n35537), .B(n35538), .Z(n35483) );
  XNOR U34050 ( .A(n35478), .B(n35539), .Z(n35538) );
  IV U34051 ( .A(n35481), .Z(n35539) );
  XOR U34052 ( .A(n35540), .B(n35541), .Z(n35481) );
  ANDN U34053 ( .B(n35542), .A(n35543), .Z(n35540) );
  XOR U34054 ( .A(n35541), .B(n35544), .Z(n35542) );
  XNOR U34055 ( .A(n35545), .B(n35546), .Z(n35478) );
  ANDN U34056 ( .B(n35547), .A(n35548), .Z(n35545) );
  XOR U34057 ( .A(n35546), .B(n35549), .Z(n35547) );
  IV U34058 ( .A(n35477), .Z(n35537) );
  XOR U34059 ( .A(n35475), .B(n35550), .Z(n35477) );
  XOR U34060 ( .A(n35551), .B(n35552), .Z(n35550) );
  ANDN U34061 ( .B(n35553), .A(n35554), .Z(n35551) );
  XOR U34062 ( .A(n35555), .B(n35552), .Z(n35553) );
  IV U34063 ( .A(n35479), .Z(n35475) );
  XOR U34064 ( .A(n35556), .B(n35557), .Z(n35479) );
  ANDN U34065 ( .B(n35558), .A(n35559), .Z(n35556) );
  XOR U34066 ( .A(n35560), .B(n35557), .Z(n35558) );
  XOR U34067 ( .A(n35561), .B(n35562), .Z(n35491) );
  XOR U34068 ( .A(n35509), .B(n35563), .Z(n35562) );
  IV U34069 ( .A(n35489), .Z(n35563) );
  XOR U34070 ( .A(n35564), .B(n35565), .Z(n35489) );
  ANDN U34071 ( .B(n35566), .A(n35567), .Z(n35564) );
  XOR U34072 ( .A(n35565), .B(n35568), .Z(n35566) );
  XOR U34073 ( .A(n35569), .B(n35497), .Z(n35509) );
  XOR U34074 ( .A(n35570), .B(n35571), .Z(n35497) );
  ANDN U34075 ( .B(n35572), .A(n35573), .Z(n35570) );
  XOR U34076 ( .A(n35571), .B(n35574), .Z(n35572) );
  IV U34077 ( .A(n35496), .Z(n35569) );
  XOR U34078 ( .A(n35575), .B(n35576), .Z(n35496) );
  XOR U34079 ( .A(n35577), .B(n35578), .Z(n35576) );
  ANDN U34080 ( .B(n35579), .A(n35580), .Z(n35577) );
  XOR U34081 ( .A(n35581), .B(n35578), .Z(n35579) );
  IV U34082 ( .A(n35494), .Z(n35575) );
  XOR U34083 ( .A(n35582), .B(n35583), .Z(n35494) );
  ANDN U34084 ( .B(n35584), .A(n35585), .Z(n35582) );
  XOR U34085 ( .A(n35583), .B(n35586), .Z(n35584) );
  IV U34086 ( .A(n35508), .Z(n35561) );
  XOR U34087 ( .A(n35587), .B(n35588), .Z(n35508) );
  XNOR U34088 ( .A(n35503), .B(n35589), .Z(n35588) );
  IV U34089 ( .A(n35506), .Z(n35589) );
  XOR U34090 ( .A(n35590), .B(n35591), .Z(n35506) );
  ANDN U34091 ( .B(n35592), .A(n35593), .Z(n35590) );
  XOR U34092 ( .A(n35594), .B(n35591), .Z(n35592) );
  XNOR U34093 ( .A(n35595), .B(n35596), .Z(n35503) );
  ANDN U34094 ( .B(n35597), .A(n35598), .Z(n35595) );
  XOR U34095 ( .A(n35596), .B(n35599), .Z(n35597) );
  IV U34096 ( .A(n35502), .Z(n35587) );
  XOR U34097 ( .A(n35500), .B(n35600), .Z(n35502) );
  XOR U34098 ( .A(n35601), .B(n35602), .Z(n35600) );
  ANDN U34099 ( .B(n35603), .A(n35604), .Z(n35601) );
  XOR U34100 ( .A(n35605), .B(n35602), .Z(n35603) );
  IV U34101 ( .A(n35504), .Z(n35500) );
  XOR U34102 ( .A(n35606), .B(n35607), .Z(n35504) );
  ANDN U34103 ( .B(n35608), .A(n35609), .Z(n35606) );
  XOR U34104 ( .A(n35610), .B(n35607), .Z(n35608) );
  IV U34105 ( .A(n35514), .Z(n35518) );
  XOR U34106 ( .A(n35514), .B(n35417), .Z(n35516) );
  XOR U34107 ( .A(n35611), .B(n35612), .Z(n35417) );
  AND U34108 ( .A(n484), .B(n35613), .Z(n35611) );
  XOR U34109 ( .A(n35614), .B(n35612), .Z(n35613) );
  NANDN U34110 ( .A(n35419), .B(n35421), .Z(n35514) );
  XOR U34111 ( .A(n35615), .B(n35616), .Z(n35421) );
  AND U34112 ( .A(n484), .B(n35617), .Z(n35615) );
  XOR U34113 ( .A(n35616), .B(n35618), .Z(n35617) );
  XNOR U34114 ( .A(n35619), .B(n35620), .Z(n484) );
  AND U34115 ( .A(n35621), .B(n35622), .Z(n35619) );
  XOR U34116 ( .A(n35620), .B(n35432), .Z(n35622) );
  XNOR U34117 ( .A(n35623), .B(n35624), .Z(n35432) );
  ANDN U34118 ( .B(n35625), .A(n35626), .Z(n35623) );
  XOR U34119 ( .A(n35624), .B(n35627), .Z(n35625) );
  XNOR U34120 ( .A(n35620), .B(n35434), .Z(n35621) );
  XOR U34121 ( .A(n35628), .B(n35629), .Z(n35434) );
  AND U34122 ( .A(n488), .B(n35630), .Z(n35628) );
  XOR U34123 ( .A(n35631), .B(n35629), .Z(n35630) );
  XOR U34124 ( .A(n35632), .B(n35633), .Z(n35620) );
  AND U34125 ( .A(n35634), .B(n35635), .Z(n35632) );
  XOR U34126 ( .A(n35633), .B(n35459), .Z(n35635) );
  XOR U34127 ( .A(n35626), .B(n35627), .Z(n35459) );
  XNOR U34128 ( .A(n35636), .B(n35637), .Z(n35627) );
  ANDN U34129 ( .B(n35638), .A(n35639), .Z(n35636) );
  XOR U34130 ( .A(n35640), .B(n35641), .Z(n35638) );
  XOR U34131 ( .A(n35642), .B(n35643), .Z(n35626) );
  XNOR U34132 ( .A(n35644), .B(n35645), .Z(n35643) );
  ANDN U34133 ( .B(n35646), .A(n35647), .Z(n35644) );
  XNOR U34134 ( .A(n35648), .B(n35649), .Z(n35646) );
  IV U34135 ( .A(n35624), .Z(n35642) );
  XOR U34136 ( .A(n35650), .B(n35651), .Z(n35624) );
  ANDN U34137 ( .B(n35652), .A(n35653), .Z(n35650) );
  XOR U34138 ( .A(n35651), .B(n35654), .Z(n35652) );
  XNOR U34139 ( .A(n35633), .B(n35461), .Z(n35634) );
  XOR U34140 ( .A(n35655), .B(n35656), .Z(n35461) );
  AND U34141 ( .A(n488), .B(n35657), .Z(n35655) );
  XOR U34142 ( .A(n35658), .B(n35656), .Z(n35657) );
  XNOR U34143 ( .A(n35659), .B(n35660), .Z(n35633) );
  AND U34144 ( .A(n35661), .B(n35662), .Z(n35659) );
  XNOR U34145 ( .A(n35660), .B(n35511), .Z(n35662) );
  XOR U34146 ( .A(n35653), .B(n35654), .Z(n35511) );
  XOR U34147 ( .A(n35663), .B(n35641), .Z(n35654) );
  XNOR U34148 ( .A(n35664), .B(n35665), .Z(n35641) );
  ANDN U34149 ( .B(n35666), .A(n35667), .Z(n35664) );
  XOR U34150 ( .A(n35668), .B(n35669), .Z(n35666) );
  IV U34151 ( .A(n35639), .Z(n35663) );
  XOR U34152 ( .A(n35637), .B(n35670), .Z(n35639) );
  XNOR U34153 ( .A(n35671), .B(n35672), .Z(n35670) );
  ANDN U34154 ( .B(n35673), .A(n35674), .Z(n35671) );
  XNOR U34155 ( .A(n35675), .B(n35676), .Z(n35673) );
  IV U34156 ( .A(n35640), .Z(n35637) );
  XOR U34157 ( .A(n35677), .B(n35678), .Z(n35640) );
  ANDN U34158 ( .B(n35679), .A(n35680), .Z(n35677) );
  XOR U34159 ( .A(n35678), .B(n35681), .Z(n35679) );
  XOR U34160 ( .A(n35682), .B(n35683), .Z(n35653) );
  XNOR U34161 ( .A(n35648), .B(n35684), .Z(n35683) );
  IV U34162 ( .A(n35651), .Z(n35684) );
  XOR U34163 ( .A(n35685), .B(n35686), .Z(n35651) );
  ANDN U34164 ( .B(n35687), .A(n35688), .Z(n35685) );
  XOR U34165 ( .A(n35686), .B(n35689), .Z(n35687) );
  XNOR U34166 ( .A(n35690), .B(n35691), .Z(n35648) );
  ANDN U34167 ( .B(n35692), .A(n35693), .Z(n35690) );
  XOR U34168 ( .A(n35691), .B(n35694), .Z(n35692) );
  IV U34169 ( .A(n35647), .Z(n35682) );
  XOR U34170 ( .A(n35645), .B(n35695), .Z(n35647) );
  XNOR U34171 ( .A(n35696), .B(n35697), .Z(n35695) );
  ANDN U34172 ( .B(n35698), .A(n35699), .Z(n35696) );
  XNOR U34173 ( .A(n35700), .B(n35701), .Z(n35698) );
  IV U34174 ( .A(n35649), .Z(n35645) );
  XOR U34175 ( .A(n35702), .B(n35703), .Z(n35649) );
  ANDN U34176 ( .B(n35704), .A(n35705), .Z(n35702) );
  XOR U34177 ( .A(n35706), .B(n35703), .Z(n35704) );
  XOR U34178 ( .A(n35660), .B(n35513), .Z(n35661) );
  XOR U34179 ( .A(n35707), .B(n35708), .Z(n35513) );
  AND U34180 ( .A(n488), .B(n35709), .Z(n35707) );
  XOR U34181 ( .A(n35710), .B(n35708), .Z(n35709) );
  XNOR U34182 ( .A(n35711), .B(n35712), .Z(n35660) );
  NAND U34183 ( .A(n35713), .B(n35714), .Z(n35712) );
  XOR U34184 ( .A(n35715), .B(n35612), .Z(n35714) );
  XOR U34185 ( .A(n35688), .B(n35689), .Z(n35612) );
  XOR U34186 ( .A(n35716), .B(n35681), .Z(n35689) );
  XOR U34187 ( .A(n35717), .B(n35669), .Z(n35681) );
  XOR U34188 ( .A(n35718), .B(n35719), .Z(n35669) );
  ANDN U34189 ( .B(n35720), .A(n35721), .Z(n35718) );
  XOR U34190 ( .A(n35719), .B(n35722), .Z(n35720) );
  IV U34191 ( .A(n35667), .Z(n35717) );
  XOR U34192 ( .A(n35665), .B(n35723), .Z(n35667) );
  XOR U34193 ( .A(n35724), .B(n35725), .Z(n35723) );
  ANDN U34194 ( .B(n35726), .A(n35727), .Z(n35724) );
  XOR U34195 ( .A(n35728), .B(n35725), .Z(n35726) );
  IV U34196 ( .A(n35668), .Z(n35665) );
  XOR U34197 ( .A(n35729), .B(n35730), .Z(n35668) );
  ANDN U34198 ( .B(n35731), .A(n35732), .Z(n35729) );
  XOR U34199 ( .A(n35730), .B(n35733), .Z(n35731) );
  IV U34200 ( .A(n35680), .Z(n35716) );
  XOR U34201 ( .A(n35734), .B(n35735), .Z(n35680) );
  XNOR U34202 ( .A(n35675), .B(n35736), .Z(n35735) );
  IV U34203 ( .A(n35678), .Z(n35736) );
  XOR U34204 ( .A(n35737), .B(n35738), .Z(n35678) );
  ANDN U34205 ( .B(n35739), .A(n35740), .Z(n35737) );
  XOR U34206 ( .A(n35738), .B(n35741), .Z(n35739) );
  XNOR U34207 ( .A(n35742), .B(n35743), .Z(n35675) );
  ANDN U34208 ( .B(n35744), .A(n35745), .Z(n35742) );
  XOR U34209 ( .A(n35743), .B(n35746), .Z(n35744) );
  IV U34210 ( .A(n35674), .Z(n35734) );
  XOR U34211 ( .A(n35672), .B(n35747), .Z(n35674) );
  XOR U34212 ( .A(n35748), .B(n35749), .Z(n35747) );
  ANDN U34213 ( .B(n35750), .A(n35751), .Z(n35748) );
  XOR U34214 ( .A(n35752), .B(n35749), .Z(n35750) );
  IV U34215 ( .A(n35676), .Z(n35672) );
  XOR U34216 ( .A(n35753), .B(n35754), .Z(n35676) );
  ANDN U34217 ( .B(n35755), .A(n35756), .Z(n35753) );
  XOR U34218 ( .A(n35757), .B(n35754), .Z(n35755) );
  XOR U34219 ( .A(n35758), .B(n35759), .Z(n35688) );
  XOR U34220 ( .A(n35706), .B(n35760), .Z(n35759) );
  IV U34221 ( .A(n35686), .Z(n35760) );
  XOR U34222 ( .A(n35761), .B(n35762), .Z(n35686) );
  ANDN U34223 ( .B(n35763), .A(n35764), .Z(n35761) );
  XOR U34224 ( .A(n35762), .B(n35765), .Z(n35763) );
  XOR U34225 ( .A(n35766), .B(n35694), .Z(n35706) );
  XOR U34226 ( .A(n35767), .B(n35768), .Z(n35694) );
  ANDN U34227 ( .B(n35769), .A(n35770), .Z(n35767) );
  XOR U34228 ( .A(n35768), .B(n35771), .Z(n35769) );
  IV U34229 ( .A(n35693), .Z(n35766) );
  XOR U34230 ( .A(n35772), .B(n35773), .Z(n35693) );
  XOR U34231 ( .A(n35774), .B(n35775), .Z(n35773) );
  ANDN U34232 ( .B(n35776), .A(n35777), .Z(n35774) );
  XOR U34233 ( .A(n35778), .B(n35775), .Z(n35776) );
  IV U34234 ( .A(n35691), .Z(n35772) );
  XOR U34235 ( .A(n35779), .B(n35780), .Z(n35691) );
  ANDN U34236 ( .B(n35781), .A(n35782), .Z(n35779) );
  XOR U34237 ( .A(n35780), .B(n35783), .Z(n35781) );
  IV U34238 ( .A(n35705), .Z(n35758) );
  XOR U34239 ( .A(n35784), .B(n35785), .Z(n35705) );
  XNOR U34240 ( .A(n35700), .B(n35786), .Z(n35785) );
  IV U34241 ( .A(n35703), .Z(n35786) );
  XOR U34242 ( .A(n35787), .B(n35788), .Z(n35703) );
  ANDN U34243 ( .B(n35789), .A(n35790), .Z(n35787) );
  XOR U34244 ( .A(n35791), .B(n35788), .Z(n35789) );
  XNOR U34245 ( .A(n35792), .B(n35793), .Z(n35700) );
  ANDN U34246 ( .B(n35794), .A(n35795), .Z(n35792) );
  XOR U34247 ( .A(n35793), .B(n35796), .Z(n35794) );
  IV U34248 ( .A(n35699), .Z(n35784) );
  XOR U34249 ( .A(n35697), .B(n35797), .Z(n35699) );
  XOR U34250 ( .A(n35798), .B(n35799), .Z(n35797) );
  ANDN U34251 ( .B(n35800), .A(n35801), .Z(n35798) );
  XOR U34252 ( .A(n35802), .B(n35799), .Z(n35800) );
  IV U34253 ( .A(n35701), .Z(n35697) );
  XOR U34254 ( .A(n35803), .B(n35804), .Z(n35701) );
  ANDN U34255 ( .B(n35805), .A(n35806), .Z(n35803) );
  XOR U34256 ( .A(n35807), .B(n35804), .Z(n35805) );
  IV U34257 ( .A(n35711), .Z(n35715) );
  XOR U34258 ( .A(n35711), .B(n35614), .Z(n35713) );
  XOR U34259 ( .A(n35808), .B(n35809), .Z(n35614) );
  AND U34260 ( .A(n488), .B(n35810), .Z(n35808) );
  XOR U34261 ( .A(n35811), .B(n35809), .Z(n35810) );
  NANDN U34262 ( .A(n35616), .B(n35618), .Z(n35711) );
  XOR U34263 ( .A(n35812), .B(n35813), .Z(n35618) );
  AND U34264 ( .A(n488), .B(n35814), .Z(n35812) );
  XOR U34265 ( .A(n35813), .B(n35815), .Z(n35814) );
  XNOR U34266 ( .A(n35816), .B(n35817), .Z(n488) );
  AND U34267 ( .A(n35818), .B(n35819), .Z(n35816) );
  XOR U34268 ( .A(n35817), .B(n35629), .Z(n35819) );
  XNOR U34269 ( .A(n35820), .B(n35821), .Z(n35629) );
  ANDN U34270 ( .B(n35822), .A(n35823), .Z(n35820) );
  XOR U34271 ( .A(n35821), .B(n35824), .Z(n35822) );
  XNOR U34272 ( .A(n35817), .B(n35631), .Z(n35818) );
  XOR U34273 ( .A(n35825), .B(n35826), .Z(n35631) );
  AND U34274 ( .A(n492), .B(n35827), .Z(n35825) );
  XOR U34275 ( .A(n35828), .B(n35826), .Z(n35827) );
  XOR U34276 ( .A(n35829), .B(n35830), .Z(n35817) );
  AND U34277 ( .A(n35831), .B(n35832), .Z(n35829) );
  XOR U34278 ( .A(n35830), .B(n35656), .Z(n35832) );
  XOR U34279 ( .A(n35823), .B(n35824), .Z(n35656) );
  XNOR U34280 ( .A(n35833), .B(n35834), .Z(n35824) );
  ANDN U34281 ( .B(n35835), .A(n35836), .Z(n35833) );
  XOR U34282 ( .A(n35837), .B(n35838), .Z(n35835) );
  XOR U34283 ( .A(n35839), .B(n35840), .Z(n35823) );
  XNOR U34284 ( .A(n35841), .B(n35842), .Z(n35840) );
  ANDN U34285 ( .B(n35843), .A(n35844), .Z(n35841) );
  XNOR U34286 ( .A(n35845), .B(n35846), .Z(n35843) );
  IV U34287 ( .A(n35821), .Z(n35839) );
  XOR U34288 ( .A(n35847), .B(n35848), .Z(n35821) );
  ANDN U34289 ( .B(n35849), .A(n35850), .Z(n35847) );
  XOR U34290 ( .A(n35848), .B(n35851), .Z(n35849) );
  XNOR U34291 ( .A(n35830), .B(n35658), .Z(n35831) );
  XOR U34292 ( .A(n35852), .B(n35853), .Z(n35658) );
  AND U34293 ( .A(n492), .B(n35854), .Z(n35852) );
  XOR U34294 ( .A(n35855), .B(n35853), .Z(n35854) );
  XNOR U34295 ( .A(n35856), .B(n35857), .Z(n35830) );
  AND U34296 ( .A(n35858), .B(n35859), .Z(n35856) );
  XNOR U34297 ( .A(n35857), .B(n35708), .Z(n35859) );
  XOR U34298 ( .A(n35850), .B(n35851), .Z(n35708) );
  XOR U34299 ( .A(n35860), .B(n35838), .Z(n35851) );
  XNOR U34300 ( .A(n35861), .B(n35862), .Z(n35838) );
  ANDN U34301 ( .B(n35863), .A(n35864), .Z(n35861) );
  XOR U34302 ( .A(n35865), .B(n35866), .Z(n35863) );
  IV U34303 ( .A(n35836), .Z(n35860) );
  XOR U34304 ( .A(n35834), .B(n35867), .Z(n35836) );
  XNOR U34305 ( .A(n35868), .B(n35869), .Z(n35867) );
  ANDN U34306 ( .B(n35870), .A(n35871), .Z(n35868) );
  XNOR U34307 ( .A(n35872), .B(n35873), .Z(n35870) );
  IV U34308 ( .A(n35837), .Z(n35834) );
  XOR U34309 ( .A(n35874), .B(n35875), .Z(n35837) );
  ANDN U34310 ( .B(n35876), .A(n35877), .Z(n35874) );
  XOR U34311 ( .A(n35875), .B(n35878), .Z(n35876) );
  XOR U34312 ( .A(n35879), .B(n35880), .Z(n35850) );
  XNOR U34313 ( .A(n35845), .B(n35881), .Z(n35880) );
  IV U34314 ( .A(n35848), .Z(n35881) );
  XOR U34315 ( .A(n35882), .B(n35883), .Z(n35848) );
  ANDN U34316 ( .B(n35884), .A(n35885), .Z(n35882) );
  XOR U34317 ( .A(n35883), .B(n35886), .Z(n35884) );
  XNOR U34318 ( .A(n35887), .B(n35888), .Z(n35845) );
  ANDN U34319 ( .B(n35889), .A(n35890), .Z(n35887) );
  XOR U34320 ( .A(n35888), .B(n35891), .Z(n35889) );
  IV U34321 ( .A(n35844), .Z(n35879) );
  XOR U34322 ( .A(n35842), .B(n35892), .Z(n35844) );
  XNOR U34323 ( .A(n35893), .B(n35894), .Z(n35892) );
  ANDN U34324 ( .B(n35895), .A(n35896), .Z(n35893) );
  XNOR U34325 ( .A(n35897), .B(n35898), .Z(n35895) );
  IV U34326 ( .A(n35846), .Z(n35842) );
  XOR U34327 ( .A(n35899), .B(n35900), .Z(n35846) );
  ANDN U34328 ( .B(n35901), .A(n35902), .Z(n35899) );
  XOR U34329 ( .A(n35903), .B(n35900), .Z(n35901) );
  XOR U34330 ( .A(n35857), .B(n35710), .Z(n35858) );
  XOR U34331 ( .A(n35904), .B(n35905), .Z(n35710) );
  AND U34332 ( .A(n492), .B(n35906), .Z(n35904) );
  XOR U34333 ( .A(n35907), .B(n35905), .Z(n35906) );
  XNOR U34334 ( .A(n35908), .B(n35909), .Z(n35857) );
  NAND U34335 ( .A(n35910), .B(n35911), .Z(n35909) );
  XOR U34336 ( .A(n35912), .B(n35809), .Z(n35911) );
  XOR U34337 ( .A(n35885), .B(n35886), .Z(n35809) );
  XOR U34338 ( .A(n35913), .B(n35878), .Z(n35886) );
  XOR U34339 ( .A(n35914), .B(n35866), .Z(n35878) );
  XOR U34340 ( .A(n35915), .B(n35916), .Z(n35866) );
  ANDN U34341 ( .B(n35917), .A(n35918), .Z(n35915) );
  XOR U34342 ( .A(n35916), .B(n35919), .Z(n35917) );
  IV U34343 ( .A(n35864), .Z(n35914) );
  XOR U34344 ( .A(n35862), .B(n35920), .Z(n35864) );
  XOR U34345 ( .A(n35921), .B(n35922), .Z(n35920) );
  ANDN U34346 ( .B(n35923), .A(n35924), .Z(n35921) );
  XOR U34347 ( .A(n35925), .B(n35922), .Z(n35923) );
  IV U34348 ( .A(n35865), .Z(n35862) );
  XOR U34349 ( .A(n35926), .B(n35927), .Z(n35865) );
  ANDN U34350 ( .B(n35928), .A(n35929), .Z(n35926) );
  XOR U34351 ( .A(n35927), .B(n35930), .Z(n35928) );
  IV U34352 ( .A(n35877), .Z(n35913) );
  XOR U34353 ( .A(n35931), .B(n35932), .Z(n35877) );
  XNOR U34354 ( .A(n35872), .B(n35933), .Z(n35932) );
  IV U34355 ( .A(n35875), .Z(n35933) );
  XOR U34356 ( .A(n35934), .B(n35935), .Z(n35875) );
  ANDN U34357 ( .B(n35936), .A(n35937), .Z(n35934) );
  XOR U34358 ( .A(n35935), .B(n35938), .Z(n35936) );
  XNOR U34359 ( .A(n35939), .B(n35940), .Z(n35872) );
  ANDN U34360 ( .B(n35941), .A(n35942), .Z(n35939) );
  XOR U34361 ( .A(n35940), .B(n35943), .Z(n35941) );
  IV U34362 ( .A(n35871), .Z(n35931) );
  XOR U34363 ( .A(n35869), .B(n35944), .Z(n35871) );
  XOR U34364 ( .A(n35945), .B(n35946), .Z(n35944) );
  ANDN U34365 ( .B(n35947), .A(n35948), .Z(n35945) );
  XOR U34366 ( .A(n35949), .B(n35946), .Z(n35947) );
  IV U34367 ( .A(n35873), .Z(n35869) );
  XOR U34368 ( .A(n35950), .B(n35951), .Z(n35873) );
  ANDN U34369 ( .B(n35952), .A(n35953), .Z(n35950) );
  XOR U34370 ( .A(n35954), .B(n35951), .Z(n35952) );
  XOR U34371 ( .A(n35955), .B(n35956), .Z(n35885) );
  XOR U34372 ( .A(n35903), .B(n35957), .Z(n35956) );
  IV U34373 ( .A(n35883), .Z(n35957) );
  XOR U34374 ( .A(n35958), .B(n35959), .Z(n35883) );
  ANDN U34375 ( .B(n35960), .A(n35961), .Z(n35958) );
  XOR U34376 ( .A(n35959), .B(n35962), .Z(n35960) );
  XOR U34377 ( .A(n35963), .B(n35891), .Z(n35903) );
  XOR U34378 ( .A(n35964), .B(n35965), .Z(n35891) );
  ANDN U34379 ( .B(n35966), .A(n35967), .Z(n35964) );
  XOR U34380 ( .A(n35965), .B(n35968), .Z(n35966) );
  IV U34381 ( .A(n35890), .Z(n35963) );
  XOR U34382 ( .A(n35969), .B(n35970), .Z(n35890) );
  XOR U34383 ( .A(n35971), .B(n35972), .Z(n35970) );
  ANDN U34384 ( .B(n35973), .A(n35974), .Z(n35971) );
  XOR U34385 ( .A(n35975), .B(n35972), .Z(n35973) );
  IV U34386 ( .A(n35888), .Z(n35969) );
  XOR U34387 ( .A(n35976), .B(n35977), .Z(n35888) );
  ANDN U34388 ( .B(n35978), .A(n35979), .Z(n35976) );
  XOR U34389 ( .A(n35977), .B(n35980), .Z(n35978) );
  IV U34390 ( .A(n35902), .Z(n35955) );
  XOR U34391 ( .A(n35981), .B(n35982), .Z(n35902) );
  XNOR U34392 ( .A(n35897), .B(n35983), .Z(n35982) );
  IV U34393 ( .A(n35900), .Z(n35983) );
  XOR U34394 ( .A(n35984), .B(n35985), .Z(n35900) );
  ANDN U34395 ( .B(n35986), .A(n35987), .Z(n35984) );
  XOR U34396 ( .A(n35988), .B(n35985), .Z(n35986) );
  XNOR U34397 ( .A(n35989), .B(n35990), .Z(n35897) );
  ANDN U34398 ( .B(n35991), .A(n35992), .Z(n35989) );
  XOR U34399 ( .A(n35990), .B(n35993), .Z(n35991) );
  IV U34400 ( .A(n35896), .Z(n35981) );
  XOR U34401 ( .A(n35894), .B(n35994), .Z(n35896) );
  XOR U34402 ( .A(n35995), .B(n35996), .Z(n35994) );
  ANDN U34403 ( .B(n35997), .A(n35998), .Z(n35995) );
  XOR U34404 ( .A(n35999), .B(n35996), .Z(n35997) );
  IV U34405 ( .A(n35898), .Z(n35894) );
  XOR U34406 ( .A(n36000), .B(n36001), .Z(n35898) );
  ANDN U34407 ( .B(n36002), .A(n36003), .Z(n36000) );
  XOR U34408 ( .A(n36004), .B(n36001), .Z(n36002) );
  IV U34409 ( .A(n35908), .Z(n35912) );
  XOR U34410 ( .A(n35908), .B(n35811), .Z(n35910) );
  XOR U34411 ( .A(n36005), .B(n36006), .Z(n35811) );
  AND U34412 ( .A(n492), .B(n36007), .Z(n36005) );
  XOR U34413 ( .A(n36008), .B(n36006), .Z(n36007) );
  NANDN U34414 ( .A(n35813), .B(n35815), .Z(n35908) );
  XOR U34415 ( .A(n36009), .B(n36010), .Z(n35815) );
  AND U34416 ( .A(n492), .B(n36011), .Z(n36009) );
  XOR U34417 ( .A(n36010), .B(n36012), .Z(n36011) );
  XNOR U34418 ( .A(n36013), .B(n36014), .Z(n492) );
  AND U34419 ( .A(n36015), .B(n36016), .Z(n36013) );
  XOR U34420 ( .A(n36014), .B(n35826), .Z(n36016) );
  XNOR U34421 ( .A(n36017), .B(n36018), .Z(n35826) );
  ANDN U34422 ( .B(n36019), .A(n36020), .Z(n36017) );
  XOR U34423 ( .A(n36018), .B(n36021), .Z(n36019) );
  XNOR U34424 ( .A(n36014), .B(n35828), .Z(n36015) );
  XOR U34425 ( .A(n36022), .B(n36023), .Z(n35828) );
  AND U34426 ( .A(n496), .B(n36024), .Z(n36022) );
  XOR U34427 ( .A(n36025), .B(n36023), .Z(n36024) );
  XOR U34428 ( .A(n36026), .B(n36027), .Z(n36014) );
  AND U34429 ( .A(n36028), .B(n36029), .Z(n36026) );
  XOR U34430 ( .A(n36027), .B(n35853), .Z(n36029) );
  XOR U34431 ( .A(n36020), .B(n36021), .Z(n35853) );
  XNOR U34432 ( .A(n36030), .B(n36031), .Z(n36021) );
  ANDN U34433 ( .B(n36032), .A(n36033), .Z(n36030) );
  XOR U34434 ( .A(n36034), .B(n36035), .Z(n36032) );
  XOR U34435 ( .A(n36036), .B(n36037), .Z(n36020) );
  XNOR U34436 ( .A(n36038), .B(n36039), .Z(n36037) );
  ANDN U34437 ( .B(n36040), .A(n36041), .Z(n36038) );
  XNOR U34438 ( .A(n36042), .B(n36043), .Z(n36040) );
  IV U34439 ( .A(n36018), .Z(n36036) );
  XOR U34440 ( .A(n36044), .B(n36045), .Z(n36018) );
  ANDN U34441 ( .B(n36046), .A(n36047), .Z(n36044) );
  XOR U34442 ( .A(n36045), .B(n36048), .Z(n36046) );
  XNOR U34443 ( .A(n36027), .B(n35855), .Z(n36028) );
  XOR U34444 ( .A(n36049), .B(n36050), .Z(n35855) );
  AND U34445 ( .A(n496), .B(n36051), .Z(n36049) );
  XOR U34446 ( .A(n36052), .B(n36050), .Z(n36051) );
  XNOR U34447 ( .A(n36053), .B(n36054), .Z(n36027) );
  AND U34448 ( .A(n36055), .B(n36056), .Z(n36053) );
  XNOR U34449 ( .A(n36054), .B(n35905), .Z(n36056) );
  XOR U34450 ( .A(n36047), .B(n36048), .Z(n35905) );
  XOR U34451 ( .A(n36057), .B(n36035), .Z(n36048) );
  XNOR U34452 ( .A(n36058), .B(n36059), .Z(n36035) );
  ANDN U34453 ( .B(n36060), .A(n36061), .Z(n36058) );
  XOR U34454 ( .A(n36062), .B(n36063), .Z(n36060) );
  IV U34455 ( .A(n36033), .Z(n36057) );
  XOR U34456 ( .A(n36031), .B(n36064), .Z(n36033) );
  XNOR U34457 ( .A(n36065), .B(n36066), .Z(n36064) );
  ANDN U34458 ( .B(n36067), .A(n36068), .Z(n36065) );
  XNOR U34459 ( .A(n36069), .B(n36070), .Z(n36067) );
  IV U34460 ( .A(n36034), .Z(n36031) );
  XOR U34461 ( .A(n36071), .B(n36072), .Z(n36034) );
  ANDN U34462 ( .B(n36073), .A(n36074), .Z(n36071) );
  XOR U34463 ( .A(n36072), .B(n36075), .Z(n36073) );
  XOR U34464 ( .A(n36076), .B(n36077), .Z(n36047) );
  XNOR U34465 ( .A(n36042), .B(n36078), .Z(n36077) );
  IV U34466 ( .A(n36045), .Z(n36078) );
  XOR U34467 ( .A(n36079), .B(n36080), .Z(n36045) );
  ANDN U34468 ( .B(n36081), .A(n36082), .Z(n36079) );
  XOR U34469 ( .A(n36080), .B(n36083), .Z(n36081) );
  XNOR U34470 ( .A(n36084), .B(n36085), .Z(n36042) );
  ANDN U34471 ( .B(n36086), .A(n36087), .Z(n36084) );
  XOR U34472 ( .A(n36085), .B(n36088), .Z(n36086) );
  IV U34473 ( .A(n36041), .Z(n36076) );
  XOR U34474 ( .A(n36039), .B(n36089), .Z(n36041) );
  XNOR U34475 ( .A(n36090), .B(n36091), .Z(n36089) );
  ANDN U34476 ( .B(n36092), .A(n36093), .Z(n36090) );
  XNOR U34477 ( .A(n36094), .B(n36095), .Z(n36092) );
  IV U34478 ( .A(n36043), .Z(n36039) );
  XOR U34479 ( .A(n36096), .B(n36097), .Z(n36043) );
  ANDN U34480 ( .B(n36098), .A(n36099), .Z(n36096) );
  XOR U34481 ( .A(n36100), .B(n36097), .Z(n36098) );
  XOR U34482 ( .A(n36054), .B(n35907), .Z(n36055) );
  XOR U34483 ( .A(n36101), .B(n36102), .Z(n35907) );
  AND U34484 ( .A(n496), .B(n36103), .Z(n36101) );
  XOR U34485 ( .A(n36104), .B(n36102), .Z(n36103) );
  XNOR U34486 ( .A(n36105), .B(n36106), .Z(n36054) );
  NAND U34487 ( .A(n36107), .B(n36108), .Z(n36106) );
  XOR U34488 ( .A(n36109), .B(n36006), .Z(n36108) );
  XOR U34489 ( .A(n36082), .B(n36083), .Z(n36006) );
  XOR U34490 ( .A(n36110), .B(n36075), .Z(n36083) );
  XOR U34491 ( .A(n36111), .B(n36063), .Z(n36075) );
  XOR U34492 ( .A(n36112), .B(n36113), .Z(n36063) );
  ANDN U34493 ( .B(n36114), .A(n36115), .Z(n36112) );
  XOR U34494 ( .A(n36113), .B(n36116), .Z(n36114) );
  IV U34495 ( .A(n36061), .Z(n36111) );
  XOR U34496 ( .A(n36059), .B(n36117), .Z(n36061) );
  XOR U34497 ( .A(n36118), .B(n36119), .Z(n36117) );
  ANDN U34498 ( .B(n36120), .A(n36121), .Z(n36118) );
  XOR U34499 ( .A(n36122), .B(n36119), .Z(n36120) );
  IV U34500 ( .A(n36062), .Z(n36059) );
  XOR U34501 ( .A(n36123), .B(n36124), .Z(n36062) );
  ANDN U34502 ( .B(n36125), .A(n36126), .Z(n36123) );
  XOR U34503 ( .A(n36124), .B(n36127), .Z(n36125) );
  IV U34504 ( .A(n36074), .Z(n36110) );
  XOR U34505 ( .A(n36128), .B(n36129), .Z(n36074) );
  XNOR U34506 ( .A(n36069), .B(n36130), .Z(n36129) );
  IV U34507 ( .A(n36072), .Z(n36130) );
  XOR U34508 ( .A(n36131), .B(n36132), .Z(n36072) );
  ANDN U34509 ( .B(n36133), .A(n36134), .Z(n36131) );
  XOR U34510 ( .A(n36132), .B(n36135), .Z(n36133) );
  XNOR U34511 ( .A(n36136), .B(n36137), .Z(n36069) );
  ANDN U34512 ( .B(n36138), .A(n36139), .Z(n36136) );
  XOR U34513 ( .A(n36137), .B(n36140), .Z(n36138) );
  IV U34514 ( .A(n36068), .Z(n36128) );
  XOR U34515 ( .A(n36066), .B(n36141), .Z(n36068) );
  XOR U34516 ( .A(n36142), .B(n36143), .Z(n36141) );
  ANDN U34517 ( .B(n36144), .A(n36145), .Z(n36142) );
  XOR U34518 ( .A(n36146), .B(n36143), .Z(n36144) );
  IV U34519 ( .A(n36070), .Z(n36066) );
  XOR U34520 ( .A(n36147), .B(n36148), .Z(n36070) );
  ANDN U34521 ( .B(n36149), .A(n36150), .Z(n36147) );
  XOR U34522 ( .A(n36151), .B(n36148), .Z(n36149) );
  XOR U34523 ( .A(n36152), .B(n36153), .Z(n36082) );
  XOR U34524 ( .A(n36100), .B(n36154), .Z(n36153) );
  IV U34525 ( .A(n36080), .Z(n36154) );
  XOR U34526 ( .A(n36155), .B(n36156), .Z(n36080) );
  ANDN U34527 ( .B(n36157), .A(n36158), .Z(n36155) );
  XOR U34528 ( .A(n36156), .B(n36159), .Z(n36157) );
  XOR U34529 ( .A(n36160), .B(n36088), .Z(n36100) );
  XOR U34530 ( .A(n36161), .B(n36162), .Z(n36088) );
  ANDN U34531 ( .B(n36163), .A(n36164), .Z(n36161) );
  XOR U34532 ( .A(n36162), .B(n36165), .Z(n36163) );
  IV U34533 ( .A(n36087), .Z(n36160) );
  XOR U34534 ( .A(n36166), .B(n36167), .Z(n36087) );
  XOR U34535 ( .A(n36168), .B(n36169), .Z(n36167) );
  ANDN U34536 ( .B(n36170), .A(n36171), .Z(n36168) );
  XOR U34537 ( .A(n36172), .B(n36169), .Z(n36170) );
  IV U34538 ( .A(n36085), .Z(n36166) );
  XOR U34539 ( .A(n36173), .B(n36174), .Z(n36085) );
  ANDN U34540 ( .B(n36175), .A(n36176), .Z(n36173) );
  XOR U34541 ( .A(n36174), .B(n36177), .Z(n36175) );
  IV U34542 ( .A(n36099), .Z(n36152) );
  XOR U34543 ( .A(n36178), .B(n36179), .Z(n36099) );
  XNOR U34544 ( .A(n36094), .B(n36180), .Z(n36179) );
  IV U34545 ( .A(n36097), .Z(n36180) );
  XOR U34546 ( .A(n36181), .B(n36182), .Z(n36097) );
  ANDN U34547 ( .B(n36183), .A(n36184), .Z(n36181) );
  XOR U34548 ( .A(n36185), .B(n36182), .Z(n36183) );
  XNOR U34549 ( .A(n36186), .B(n36187), .Z(n36094) );
  ANDN U34550 ( .B(n36188), .A(n36189), .Z(n36186) );
  XOR U34551 ( .A(n36187), .B(n36190), .Z(n36188) );
  IV U34552 ( .A(n36093), .Z(n36178) );
  XOR U34553 ( .A(n36091), .B(n36191), .Z(n36093) );
  XOR U34554 ( .A(n36192), .B(n36193), .Z(n36191) );
  ANDN U34555 ( .B(n36194), .A(n36195), .Z(n36192) );
  XOR U34556 ( .A(n36196), .B(n36193), .Z(n36194) );
  IV U34557 ( .A(n36095), .Z(n36091) );
  XOR U34558 ( .A(n36197), .B(n36198), .Z(n36095) );
  ANDN U34559 ( .B(n36199), .A(n36200), .Z(n36197) );
  XOR U34560 ( .A(n36201), .B(n36198), .Z(n36199) );
  IV U34561 ( .A(n36105), .Z(n36109) );
  XOR U34562 ( .A(n36105), .B(n36008), .Z(n36107) );
  XOR U34563 ( .A(n36202), .B(n36203), .Z(n36008) );
  AND U34564 ( .A(n496), .B(n36204), .Z(n36202) );
  XOR U34565 ( .A(n36205), .B(n36203), .Z(n36204) );
  NANDN U34566 ( .A(n36010), .B(n36012), .Z(n36105) );
  XOR U34567 ( .A(n36206), .B(n36207), .Z(n36012) );
  AND U34568 ( .A(n496), .B(n36208), .Z(n36206) );
  XOR U34569 ( .A(n36207), .B(n36209), .Z(n36208) );
  XNOR U34570 ( .A(n36210), .B(n36211), .Z(n496) );
  AND U34571 ( .A(n36212), .B(n36213), .Z(n36210) );
  XOR U34572 ( .A(n36211), .B(n36023), .Z(n36213) );
  XNOR U34573 ( .A(n36214), .B(n36215), .Z(n36023) );
  ANDN U34574 ( .B(n36216), .A(n36217), .Z(n36214) );
  XOR U34575 ( .A(n36215), .B(n36218), .Z(n36216) );
  XNOR U34576 ( .A(n36211), .B(n36025), .Z(n36212) );
  XOR U34577 ( .A(n36219), .B(n36220), .Z(n36025) );
  AND U34578 ( .A(n500), .B(n36221), .Z(n36219) );
  XOR U34579 ( .A(n36222), .B(n36220), .Z(n36221) );
  XOR U34580 ( .A(n36223), .B(n36224), .Z(n36211) );
  AND U34581 ( .A(n36225), .B(n36226), .Z(n36223) );
  XOR U34582 ( .A(n36224), .B(n36050), .Z(n36226) );
  XOR U34583 ( .A(n36217), .B(n36218), .Z(n36050) );
  XNOR U34584 ( .A(n36227), .B(n36228), .Z(n36218) );
  ANDN U34585 ( .B(n36229), .A(n36230), .Z(n36227) );
  XOR U34586 ( .A(n36231), .B(n36232), .Z(n36229) );
  XOR U34587 ( .A(n36233), .B(n36234), .Z(n36217) );
  XNOR U34588 ( .A(n36235), .B(n36236), .Z(n36234) );
  ANDN U34589 ( .B(n36237), .A(n36238), .Z(n36235) );
  XNOR U34590 ( .A(n36239), .B(n36240), .Z(n36237) );
  IV U34591 ( .A(n36215), .Z(n36233) );
  XOR U34592 ( .A(n36241), .B(n36242), .Z(n36215) );
  ANDN U34593 ( .B(n36243), .A(n36244), .Z(n36241) );
  XOR U34594 ( .A(n36242), .B(n36245), .Z(n36243) );
  XNOR U34595 ( .A(n36224), .B(n36052), .Z(n36225) );
  XOR U34596 ( .A(n36246), .B(n36247), .Z(n36052) );
  AND U34597 ( .A(n500), .B(n36248), .Z(n36246) );
  XOR U34598 ( .A(n36249), .B(n36247), .Z(n36248) );
  XNOR U34599 ( .A(n36250), .B(n36251), .Z(n36224) );
  AND U34600 ( .A(n36252), .B(n36253), .Z(n36250) );
  XNOR U34601 ( .A(n36251), .B(n36102), .Z(n36253) );
  XOR U34602 ( .A(n36244), .B(n36245), .Z(n36102) );
  XOR U34603 ( .A(n36254), .B(n36232), .Z(n36245) );
  XNOR U34604 ( .A(n36255), .B(n36256), .Z(n36232) );
  ANDN U34605 ( .B(n36257), .A(n36258), .Z(n36255) );
  XOR U34606 ( .A(n36259), .B(n36260), .Z(n36257) );
  IV U34607 ( .A(n36230), .Z(n36254) );
  XOR U34608 ( .A(n36228), .B(n36261), .Z(n36230) );
  XNOR U34609 ( .A(n36262), .B(n36263), .Z(n36261) );
  ANDN U34610 ( .B(n36264), .A(n36265), .Z(n36262) );
  XNOR U34611 ( .A(n36266), .B(n36267), .Z(n36264) );
  IV U34612 ( .A(n36231), .Z(n36228) );
  XOR U34613 ( .A(n36268), .B(n36269), .Z(n36231) );
  ANDN U34614 ( .B(n36270), .A(n36271), .Z(n36268) );
  XOR U34615 ( .A(n36269), .B(n36272), .Z(n36270) );
  XOR U34616 ( .A(n36273), .B(n36274), .Z(n36244) );
  XNOR U34617 ( .A(n36239), .B(n36275), .Z(n36274) );
  IV U34618 ( .A(n36242), .Z(n36275) );
  XOR U34619 ( .A(n36276), .B(n36277), .Z(n36242) );
  ANDN U34620 ( .B(n36278), .A(n36279), .Z(n36276) );
  XOR U34621 ( .A(n36277), .B(n36280), .Z(n36278) );
  XNOR U34622 ( .A(n36281), .B(n36282), .Z(n36239) );
  ANDN U34623 ( .B(n36283), .A(n36284), .Z(n36281) );
  XOR U34624 ( .A(n36282), .B(n36285), .Z(n36283) );
  IV U34625 ( .A(n36238), .Z(n36273) );
  XOR U34626 ( .A(n36236), .B(n36286), .Z(n36238) );
  XNOR U34627 ( .A(n36287), .B(n36288), .Z(n36286) );
  ANDN U34628 ( .B(n36289), .A(n36290), .Z(n36287) );
  XNOR U34629 ( .A(n36291), .B(n36292), .Z(n36289) );
  IV U34630 ( .A(n36240), .Z(n36236) );
  XOR U34631 ( .A(n36293), .B(n36294), .Z(n36240) );
  ANDN U34632 ( .B(n36295), .A(n36296), .Z(n36293) );
  XOR U34633 ( .A(n36297), .B(n36294), .Z(n36295) );
  XOR U34634 ( .A(n36251), .B(n36104), .Z(n36252) );
  XOR U34635 ( .A(n36298), .B(n36299), .Z(n36104) );
  AND U34636 ( .A(n500), .B(n36300), .Z(n36298) );
  XOR U34637 ( .A(n36301), .B(n36299), .Z(n36300) );
  XNOR U34638 ( .A(n36302), .B(n36303), .Z(n36251) );
  NAND U34639 ( .A(n36304), .B(n36305), .Z(n36303) );
  XOR U34640 ( .A(n36306), .B(n36203), .Z(n36305) );
  XOR U34641 ( .A(n36279), .B(n36280), .Z(n36203) );
  XOR U34642 ( .A(n36307), .B(n36272), .Z(n36280) );
  XOR U34643 ( .A(n36308), .B(n36260), .Z(n36272) );
  XOR U34644 ( .A(n36309), .B(n36310), .Z(n36260) );
  ANDN U34645 ( .B(n36311), .A(n36312), .Z(n36309) );
  XOR U34646 ( .A(n36310), .B(n36313), .Z(n36311) );
  IV U34647 ( .A(n36258), .Z(n36308) );
  XOR U34648 ( .A(n36256), .B(n36314), .Z(n36258) );
  XOR U34649 ( .A(n36315), .B(n36316), .Z(n36314) );
  ANDN U34650 ( .B(n36317), .A(n36318), .Z(n36315) );
  XOR U34651 ( .A(n36319), .B(n36316), .Z(n36317) );
  IV U34652 ( .A(n36259), .Z(n36256) );
  XOR U34653 ( .A(n36320), .B(n36321), .Z(n36259) );
  ANDN U34654 ( .B(n36322), .A(n36323), .Z(n36320) );
  XOR U34655 ( .A(n36321), .B(n36324), .Z(n36322) );
  IV U34656 ( .A(n36271), .Z(n36307) );
  XOR U34657 ( .A(n36325), .B(n36326), .Z(n36271) );
  XNOR U34658 ( .A(n36266), .B(n36327), .Z(n36326) );
  IV U34659 ( .A(n36269), .Z(n36327) );
  XOR U34660 ( .A(n36328), .B(n36329), .Z(n36269) );
  ANDN U34661 ( .B(n36330), .A(n36331), .Z(n36328) );
  XOR U34662 ( .A(n36329), .B(n36332), .Z(n36330) );
  XNOR U34663 ( .A(n36333), .B(n36334), .Z(n36266) );
  ANDN U34664 ( .B(n36335), .A(n36336), .Z(n36333) );
  XOR U34665 ( .A(n36334), .B(n36337), .Z(n36335) );
  IV U34666 ( .A(n36265), .Z(n36325) );
  XOR U34667 ( .A(n36263), .B(n36338), .Z(n36265) );
  XOR U34668 ( .A(n36339), .B(n36340), .Z(n36338) );
  ANDN U34669 ( .B(n36341), .A(n36342), .Z(n36339) );
  XOR U34670 ( .A(n36343), .B(n36340), .Z(n36341) );
  IV U34671 ( .A(n36267), .Z(n36263) );
  XOR U34672 ( .A(n36344), .B(n36345), .Z(n36267) );
  ANDN U34673 ( .B(n36346), .A(n36347), .Z(n36344) );
  XOR U34674 ( .A(n36348), .B(n36345), .Z(n36346) );
  XOR U34675 ( .A(n36349), .B(n36350), .Z(n36279) );
  XOR U34676 ( .A(n36297), .B(n36351), .Z(n36350) );
  IV U34677 ( .A(n36277), .Z(n36351) );
  XOR U34678 ( .A(n36352), .B(n36353), .Z(n36277) );
  ANDN U34679 ( .B(n36354), .A(n36355), .Z(n36352) );
  XOR U34680 ( .A(n36353), .B(n36356), .Z(n36354) );
  XOR U34681 ( .A(n36357), .B(n36285), .Z(n36297) );
  XOR U34682 ( .A(n36358), .B(n36359), .Z(n36285) );
  ANDN U34683 ( .B(n36360), .A(n36361), .Z(n36358) );
  XOR U34684 ( .A(n36359), .B(n36362), .Z(n36360) );
  IV U34685 ( .A(n36284), .Z(n36357) );
  XOR U34686 ( .A(n36363), .B(n36364), .Z(n36284) );
  XOR U34687 ( .A(n36365), .B(n36366), .Z(n36364) );
  ANDN U34688 ( .B(n36367), .A(n36368), .Z(n36365) );
  XOR U34689 ( .A(n36369), .B(n36366), .Z(n36367) );
  IV U34690 ( .A(n36282), .Z(n36363) );
  XOR U34691 ( .A(n36370), .B(n36371), .Z(n36282) );
  ANDN U34692 ( .B(n36372), .A(n36373), .Z(n36370) );
  XOR U34693 ( .A(n36371), .B(n36374), .Z(n36372) );
  IV U34694 ( .A(n36296), .Z(n36349) );
  XOR U34695 ( .A(n36375), .B(n36376), .Z(n36296) );
  XNOR U34696 ( .A(n36291), .B(n36377), .Z(n36376) );
  IV U34697 ( .A(n36294), .Z(n36377) );
  XOR U34698 ( .A(n36378), .B(n36379), .Z(n36294) );
  ANDN U34699 ( .B(n36380), .A(n36381), .Z(n36378) );
  XOR U34700 ( .A(n36382), .B(n36379), .Z(n36380) );
  XNOR U34701 ( .A(n36383), .B(n36384), .Z(n36291) );
  ANDN U34702 ( .B(n36385), .A(n36386), .Z(n36383) );
  XOR U34703 ( .A(n36384), .B(n36387), .Z(n36385) );
  IV U34704 ( .A(n36290), .Z(n36375) );
  XOR U34705 ( .A(n36288), .B(n36388), .Z(n36290) );
  XOR U34706 ( .A(n36389), .B(n36390), .Z(n36388) );
  ANDN U34707 ( .B(n36391), .A(n36392), .Z(n36389) );
  XOR U34708 ( .A(n36393), .B(n36390), .Z(n36391) );
  IV U34709 ( .A(n36292), .Z(n36288) );
  XOR U34710 ( .A(n36394), .B(n36395), .Z(n36292) );
  ANDN U34711 ( .B(n36396), .A(n36397), .Z(n36394) );
  XOR U34712 ( .A(n36398), .B(n36395), .Z(n36396) );
  IV U34713 ( .A(n36302), .Z(n36306) );
  XOR U34714 ( .A(n36302), .B(n36205), .Z(n36304) );
  XOR U34715 ( .A(n36399), .B(n36400), .Z(n36205) );
  AND U34716 ( .A(n500), .B(n36401), .Z(n36399) );
  XOR U34717 ( .A(n36402), .B(n36400), .Z(n36401) );
  NANDN U34718 ( .A(n36207), .B(n36209), .Z(n36302) );
  XOR U34719 ( .A(n36403), .B(n36404), .Z(n36209) );
  AND U34720 ( .A(n500), .B(n36405), .Z(n36403) );
  XOR U34721 ( .A(n36404), .B(n36406), .Z(n36405) );
  XNOR U34722 ( .A(n36407), .B(n36408), .Z(n500) );
  AND U34723 ( .A(n36409), .B(n36410), .Z(n36407) );
  XOR U34724 ( .A(n36408), .B(n36220), .Z(n36410) );
  XNOR U34725 ( .A(n36411), .B(n36412), .Z(n36220) );
  ANDN U34726 ( .B(n36413), .A(n36414), .Z(n36411) );
  XOR U34727 ( .A(n36412), .B(n36415), .Z(n36413) );
  XNOR U34728 ( .A(n36408), .B(n36222), .Z(n36409) );
  XOR U34729 ( .A(n36416), .B(n36417), .Z(n36222) );
  AND U34730 ( .A(n504), .B(n36418), .Z(n36416) );
  XOR U34731 ( .A(n36419), .B(n36417), .Z(n36418) );
  XOR U34732 ( .A(n36420), .B(n36421), .Z(n36408) );
  AND U34733 ( .A(n36422), .B(n36423), .Z(n36420) );
  XOR U34734 ( .A(n36421), .B(n36247), .Z(n36423) );
  XOR U34735 ( .A(n36414), .B(n36415), .Z(n36247) );
  XNOR U34736 ( .A(n36424), .B(n36425), .Z(n36415) );
  ANDN U34737 ( .B(n36426), .A(n36427), .Z(n36424) );
  XOR U34738 ( .A(n36428), .B(n36429), .Z(n36426) );
  XOR U34739 ( .A(n36430), .B(n36431), .Z(n36414) );
  XNOR U34740 ( .A(n36432), .B(n36433), .Z(n36431) );
  ANDN U34741 ( .B(n36434), .A(n36435), .Z(n36432) );
  XNOR U34742 ( .A(n36436), .B(n36437), .Z(n36434) );
  IV U34743 ( .A(n36412), .Z(n36430) );
  XOR U34744 ( .A(n36438), .B(n36439), .Z(n36412) );
  ANDN U34745 ( .B(n36440), .A(n36441), .Z(n36438) );
  XOR U34746 ( .A(n36439), .B(n36442), .Z(n36440) );
  XNOR U34747 ( .A(n36421), .B(n36249), .Z(n36422) );
  XOR U34748 ( .A(n36443), .B(n36444), .Z(n36249) );
  AND U34749 ( .A(n504), .B(n36445), .Z(n36443) );
  XOR U34750 ( .A(n36446), .B(n36444), .Z(n36445) );
  XNOR U34751 ( .A(n36447), .B(n36448), .Z(n36421) );
  AND U34752 ( .A(n36449), .B(n36450), .Z(n36447) );
  XNOR U34753 ( .A(n36448), .B(n36299), .Z(n36450) );
  XOR U34754 ( .A(n36441), .B(n36442), .Z(n36299) );
  XOR U34755 ( .A(n36451), .B(n36429), .Z(n36442) );
  XNOR U34756 ( .A(n36452), .B(n36453), .Z(n36429) );
  ANDN U34757 ( .B(n36454), .A(n36455), .Z(n36452) );
  XOR U34758 ( .A(n36456), .B(n36457), .Z(n36454) );
  IV U34759 ( .A(n36427), .Z(n36451) );
  XOR U34760 ( .A(n36425), .B(n36458), .Z(n36427) );
  XNOR U34761 ( .A(n36459), .B(n36460), .Z(n36458) );
  ANDN U34762 ( .B(n36461), .A(n36462), .Z(n36459) );
  XNOR U34763 ( .A(n36463), .B(n36464), .Z(n36461) );
  IV U34764 ( .A(n36428), .Z(n36425) );
  XOR U34765 ( .A(n36465), .B(n36466), .Z(n36428) );
  ANDN U34766 ( .B(n36467), .A(n36468), .Z(n36465) );
  XOR U34767 ( .A(n36466), .B(n36469), .Z(n36467) );
  XOR U34768 ( .A(n36470), .B(n36471), .Z(n36441) );
  XNOR U34769 ( .A(n36436), .B(n36472), .Z(n36471) );
  IV U34770 ( .A(n36439), .Z(n36472) );
  XOR U34771 ( .A(n36473), .B(n36474), .Z(n36439) );
  ANDN U34772 ( .B(n36475), .A(n36476), .Z(n36473) );
  XOR U34773 ( .A(n36474), .B(n36477), .Z(n36475) );
  XNOR U34774 ( .A(n36478), .B(n36479), .Z(n36436) );
  ANDN U34775 ( .B(n36480), .A(n36481), .Z(n36478) );
  XOR U34776 ( .A(n36479), .B(n36482), .Z(n36480) );
  IV U34777 ( .A(n36435), .Z(n36470) );
  XOR U34778 ( .A(n36433), .B(n36483), .Z(n36435) );
  XNOR U34779 ( .A(n36484), .B(n36485), .Z(n36483) );
  ANDN U34780 ( .B(n36486), .A(n36487), .Z(n36484) );
  XNOR U34781 ( .A(n36488), .B(n36489), .Z(n36486) );
  IV U34782 ( .A(n36437), .Z(n36433) );
  XOR U34783 ( .A(n36490), .B(n36491), .Z(n36437) );
  ANDN U34784 ( .B(n36492), .A(n36493), .Z(n36490) );
  XOR U34785 ( .A(n36494), .B(n36491), .Z(n36492) );
  XOR U34786 ( .A(n36448), .B(n36301), .Z(n36449) );
  XOR U34787 ( .A(n36495), .B(n36496), .Z(n36301) );
  AND U34788 ( .A(n504), .B(n36497), .Z(n36495) );
  XOR U34789 ( .A(n36498), .B(n36496), .Z(n36497) );
  XNOR U34790 ( .A(n36499), .B(n36500), .Z(n36448) );
  NAND U34791 ( .A(n36501), .B(n36502), .Z(n36500) );
  XOR U34792 ( .A(n36503), .B(n36400), .Z(n36502) );
  XOR U34793 ( .A(n36476), .B(n36477), .Z(n36400) );
  XOR U34794 ( .A(n36504), .B(n36469), .Z(n36477) );
  XOR U34795 ( .A(n36505), .B(n36457), .Z(n36469) );
  XOR U34796 ( .A(n36506), .B(n36507), .Z(n36457) );
  ANDN U34797 ( .B(n36508), .A(n36509), .Z(n36506) );
  XOR U34798 ( .A(n36507), .B(n36510), .Z(n36508) );
  IV U34799 ( .A(n36455), .Z(n36505) );
  XOR U34800 ( .A(n36453), .B(n36511), .Z(n36455) );
  XOR U34801 ( .A(n36512), .B(n36513), .Z(n36511) );
  ANDN U34802 ( .B(n36514), .A(n36515), .Z(n36512) );
  XOR U34803 ( .A(n36516), .B(n36513), .Z(n36514) );
  IV U34804 ( .A(n36456), .Z(n36453) );
  XOR U34805 ( .A(n36517), .B(n36518), .Z(n36456) );
  ANDN U34806 ( .B(n36519), .A(n36520), .Z(n36517) );
  XOR U34807 ( .A(n36518), .B(n36521), .Z(n36519) );
  IV U34808 ( .A(n36468), .Z(n36504) );
  XOR U34809 ( .A(n36522), .B(n36523), .Z(n36468) );
  XNOR U34810 ( .A(n36463), .B(n36524), .Z(n36523) );
  IV U34811 ( .A(n36466), .Z(n36524) );
  XOR U34812 ( .A(n36525), .B(n36526), .Z(n36466) );
  ANDN U34813 ( .B(n36527), .A(n36528), .Z(n36525) );
  XOR U34814 ( .A(n36526), .B(n36529), .Z(n36527) );
  XNOR U34815 ( .A(n36530), .B(n36531), .Z(n36463) );
  ANDN U34816 ( .B(n36532), .A(n36533), .Z(n36530) );
  XOR U34817 ( .A(n36531), .B(n36534), .Z(n36532) );
  IV U34818 ( .A(n36462), .Z(n36522) );
  XOR U34819 ( .A(n36460), .B(n36535), .Z(n36462) );
  XOR U34820 ( .A(n36536), .B(n36537), .Z(n36535) );
  ANDN U34821 ( .B(n36538), .A(n36539), .Z(n36536) );
  XOR U34822 ( .A(n36540), .B(n36537), .Z(n36538) );
  IV U34823 ( .A(n36464), .Z(n36460) );
  XOR U34824 ( .A(n36541), .B(n36542), .Z(n36464) );
  ANDN U34825 ( .B(n36543), .A(n36544), .Z(n36541) );
  XOR U34826 ( .A(n36545), .B(n36542), .Z(n36543) );
  XOR U34827 ( .A(n36546), .B(n36547), .Z(n36476) );
  XOR U34828 ( .A(n36494), .B(n36548), .Z(n36547) );
  IV U34829 ( .A(n36474), .Z(n36548) );
  XOR U34830 ( .A(n36549), .B(n36550), .Z(n36474) );
  ANDN U34831 ( .B(n36551), .A(n36552), .Z(n36549) );
  XOR U34832 ( .A(n36550), .B(n36553), .Z(n36551) );
  XOR U34833 ( .A(n36554), .B(n36482), .Z(n36494) );
  XOR U34834 ( .A(n36555), .B(n36556), .Z(n36482) );
  ANDN U34835 ( .B(n36557), .A(n36558), .Z(n36555) );
  XOR U34836 ( .A(n36556), .B(n36559), .Z(n36557) );
  IV U34837 ( .A(n36481), .Z(n36554) );
  XOR U34838 ( .A(n36560), .B(n36561), .Z(n36481) );
  XOR U34839 ( .A(n36562), .B(n36563), .Z(n36561) );
  ANDN U34840 ( .B(n36564), .A(n36565), .Z(n36562) );
  XOR U34841 ( .A(n36566), .B(n36563), .Z(n36564) );
  IV U34842 ( .A(n36479), .Z(n36560) );
  XOR U34843 ( .A(n36567), .B(n36568), .Z(n36479) );
  ANDN U34844 ( .B(n36569), .A(n36570), .Z(n36567) );
  XOR U34845 ( .A(n36568), .B(n36571), .Z(n36569) );
  IV U34846 ( .A(n36493), .Z(n36546) );
  XOR U34847 ( .A(n36572), .B(n36573), .Z(n36493) );
  XNOR U34848 ( .A(n36488), .B(n36574), .Z(n36573) );
  IV U34849 ( .A(n36491), .Z(n36574) );
  XOR U34850 ( .A(n36575), .B(n36576), .Z(n36491) );
  ANDN U34851 ( .B(n36577), .A(n36578), .Z(n36575) );
  XOR U34852 ( .A(n36579), .B(n36576), .Z(n36577) );
  XNOR U34853 ( .A(n36580), .B(n36581), .Z(n36488) );
  ANDN U34854 ( .B(n36582), .A(n36583), .Z(n36580) );
  XOR U34855 ( .A(n36581), .B(n36584), .Z(n36582) );
  IV U34856 ( .A(n36487), .Z(n36572) );
  XOR U34857 ( .A(n36485), .B(n36585), .Z(n36487) );
  XOR U34858 ( .A(n36586), .B(n36587), .Z(n36585) );
  ANDN U34859 ( .B(n36588), .A(n36589), .Z(n36586) );
  XOR U34860 ( .A(n36590), .B(n36587), .Z(n36588) );
  IV U34861 ( .A(n36489), .Z(n36485) );
  XOR U34862 ( .A(n36591), .B(n36592), .Z(n36489) );
  ANDN U34863 ( .B(n36593), .A(n36594), .Z(n36591) );
  XOR U34864 ( .A(n36595), .B(n36592), .Z(n36593) );
  IV U34865 ( .A(n36499), .Z(n36503) );
  XOR U34866 ( .A(n36499), .B(n36402), .Z(n36501) );
  XOR U34867 ( .A(n36596), .B(n36597), .Z(n36402) );
  AND U34868 ( .A(n504), .B(n36598), .Z(n36596) );
  XOR U34869 ( .A(n36599), .B(n36597), .Z(n36598) );
  NANDN U34870 ( .A(n36404), .B(n36406), .Z(n36499) );
  XOR U34871 ( .A(n36600), .B(n36601), .Z(n36406) );
  AND U34872 ( .A(n504), .B(n36602), .Z(n36600) );
  XOR U34873 ( .A(n36601), .B(n36603), .Z(n36602) );
  XNOR U34874 ( .A(n36604), .B(n36605), .Z(n504) );
  AND U34875 ( .A(n36606), .B(n36607), .Z(n36604) );
  XOR U34876 ( .A(n36605), .B(n36417), .Z(n36607) );
  XNOR U34877 ( .A(n36608), .B(n36609), .Z(n36417) );
  ANDN U34878 ( .B(n36610), .A(n36611), .Z(n36608) );
  XOR U34879 ( .A(n36609), .B(n36612), .Z(n36610) );
  XNOR U34880 ( .A(n36605), .B(n36419), .Z(n36606) );
  XOR U34881 ( .A(n36613), .B(n36614), .Z(n36419) );
  AND U34882 ( .A(n508), .B(n36615), .Z(n36613) );
  XOR U34883 ( .A(n36616), .B(n36614), .Z(n36615) );
  XOR U34884 ( .A(n36617), .B(n36618), .Z(n36605) );
  AND U34885 ( .A(n36619), .B(n36620), .Z(n36617) );
  XOR U34886 ( .A(n36618), .B(n36444), .Z(n36620) );
  XOR U34887 ( .A(n36611), .B(n36612), .Z(n36444) );
  XNOR U34888 ( .A(n36621), .B(n36622), .Z(n36612) );
  ANDN U34889 ( .B(n36623), .A(n36624), .Z(n36621) );
  XOR U34890 ( .A(n36625), .B(n36626), .Z(n36623) );
  XOR U34891 ( .A(n36627), .B(n36628), .Z(n36611) );
  XNOR U34892 ( .A(n36629), .B(n36630), .Z(n36628) );
  ANDN U34893 ( .B(n36631), .A(n36632), .Z(n36629) );
  XNOR U34894 ( .A(n36633), .B(n36634), .Z(n36631) );
  IV U34895 ( .A(n36609), .Z(n36627) );
  XOR U34896 ( .A(n36635), .B(n36636), .Z(n36609) );
  ANDN U34897 ( .B(n36637), .A(n36638), .Z(n36635) );
  XOR U34898 ( .A(n36636), .B(n36639), .Z(n36637) );
  XNOR U34899 ( .A(n36618), .B(n36446), .Z(n36619) );
  XOR U34900 ( .A(n36640), .B(n36641), .Z(n36446) );
  AND U34901 ( .A(n508), .B(n36642), .Z(n36640) );
  XNOR U34902 ( .A(n36643), .B(n36641), .Z(n36642) );
  XNOR U34903 ( .A(n36644), .B(n36645), .Z(n36618) );
  AND U34904 ( .A(n36646), .B(n36647), .Z(n36644) );
  XNOR U34905 ( .A(n36645), .B(n36496), .Z(n36647) );
  XOR U34906 ( .A(n36638), .B(n36639), .Z(n36496) );
  XOR U34907 ( .A(n36648), .B(n36626), .Z(n36639) );
  XNOR U34908 ( .A(n36649), .B(n36650), .Z(n36626) );
  ANDN U34909 ( .B(n36651), .A(n36652), .Z(n36649) );
  XOR U34910 ( .A(n36653), .B(n36654), .Z(n36651) );
  IV U34911 ( .A(n36624), .Z(n36648) );
  XOR U34912 ( .A(n36622), .B(n36655), .Z(n36624) );
  XNOR U34913 ( .A(n36656), .B(n36657), .Z(n36655) );
  ANDN U34914 ( .B(n36658), .A(n36659), .Z(n36656) );
  XNOR U34915 ( .A(n36660), .B(n36661), .Z(n36658) );
  IV U34916 ( .A(n36625), .Z(n36622) );
  XOR U34917 ( .A(n36662), .B(n36663), .Z(n36625) );
  ANDN U34918 ( .B(n36664), .A(n36665), .Z(n36662) );
  XOR U34919 ( .A(n36663), .B(n36666), .Z(n36664) );
  XOR U34920 ( .A(n36667), .B(n36668), .Z(n36638) );
  XNOR U34921 ( .A(n36633), .B(n36669), .Z(n36668) );
  IV U34922 ( .A(n36636), .Z(n36669) );
  XOR U34923 ( .A(n36670), .B(n36671), .Z(n36636) );
  ANDN U34924 ( .B(n36672), .A(n36673), .Z(n36670) );
  XOR U34925 ( .A(n36671), .B(n36674), .Z(n36672) );
  XNOR U34926 ( .A(n36675), .B(n36676), .Z(n36633) );
  ANDN U34927 ( .B(n36677), .A(n36678), .Z(n36675) );
  XOR U34928 ( .A(n36676), .B(n36679), .Z(n36677) );
  IV U34929 ( .A(n36632), .Z(n36667) );
  XOR U34930 ( .A(n36630), .B(n36680), .Z(n36632) );
  XNOR U34931 ( .A(n36681), .B(n36682), .Z(n36680) );
  ANDN U34932 ( .B(n36683), .A(n36684), .Z(n36681) );
  XNOR U34933 ( .A(n36685), .B(n36686), .Z(n36683) );
  IV U34934 ( .A(n36634), .Z(n36630) );
  XOR U34935 ( .A(n36687), .B(n36688), .Z(n36634) );
  ANDN U34936 ( .B(n36689), .A(n36690), .Z(n36687) );
  XOR U34937 ( .A(n36691), .B(n36688), .Z(n36689) );
  XOR U34938 ( .A(n36645), .B(n36498), .Z(n36646) );
  XOR U34939 ( .A(n36692), .B(n36693), .Z(n36498) );
  AND U34940 ( .A(n508), .B(n36694), .Z(n36692) );
  XNOR U34941 ( .A(n36695), .B(n36693), .Z(n36694) );
  XNOR U34942 ( .A(n36696), .B(n36697), .Z(n36645) );
  NAND U34943 ( .A(n36698), .B(n36699), .Z(n36697) );
  XOR U34944 ( .A(n36700), .B(n36597), .Z(n36699) );
  XOR U34945 ( .A(n36673), .B(n36674), .Z(n36597) );
  XOR U34946 ( .A(n36701), .B(n36666), .Z(n36674) );
  XOR U34947 ( .A(n36702), .B(n36654), .Z(n36666) );
  XOR U34948 ( .A(n36703), .B(n36704), .Z(n36654) );
  ANDN U34949 ( .B(n36705), .A(n36706), .Z(n36703) );
  XOR U34950 ( .A(n36704), .B(n36707), .Z(n36705) );
  IV U34951 ( .A(n36652), .Z(n36702) );
  XOR U34952 ( .A(n36650), .B(n36708), .Z(n36652) );
  XOR U34953 ( .A(n36709), .B(n36710), .Z(n36708) );
  ANDN U34954 ( .B(n36711), .A(n36712), .Z(n36709) );
  XOR U34955 ( .A(n36713), .B(n36710), .Z(n36711) );
  IV U34956 ( .A(n36653), .Z(n36650) );
  XOR U34957 ( .A(n36714), .B(n36715), .Z(n36653) );
  ANDN U34958 ( .B(n36716), .A(n36717), .Z(n36714) );
  XOR U34959 ( .A(n36715), .B(n36718), .Z(n36716) );
  IV U34960 ( .A(n36665), .Z(n36701) );
  XOR U34961 ( .A(n36719), .B(n36720), .Z(n36665) );
  XNOR U34962 ( .A(n36660), .B(n36721), .Z(n36720) );
  IV U34963 ( .A(n36663), .Z(n36721) );
  XOR U34964 ( .A(n36722), .B(n36723), .Z(n36663) );
  ANDN U34965 ( .B(n36724), .A(n36725), .Z(n36722) );
  XOR U34966 ( .A(n36723), .B(n36726), .Z(n36724) );
  XNOR U34967 ( .A(n36727), .B(n36728), .Z(n36660) );
  ANDN U34968 ( .B(n36729), .A(n36730), .Z(n36727) );
  XOR U34969 ( .A(n36728), .B(n36731), .Z(n36729) );
  IV U34970 ( .A(n36659), .Z(n36719) );
  XOR U34971 ( .A(n36657), .B(n36732), .Z(n36659) );
  XOR U34972 ( .A(n36733), .B(n36734), .Z(n36732) );
  ANDN U34973 ( .B(n36735), .A(n36736), .Z(n36733) );
  XOR U34974 ( .A(n36737), .B(n36734), .Z(n36735) );
  IV U34975 ( .A(n36661), .Z(n36657) );
  XOR U34976 ( .A(n36738), .B(n36739), .Z(n36661) );
  ANDN U34977 ( .B(n36740), .A(n36741), .Z(n36738) );
  XOR U34978 ( .A(n36742), .B(n36739), .Z(n36740) );
  XOR U34979 ( .A(n36743), .B(n36744), .Z(n36673) );
  XOR U34980 ( .A(n36691), .B(n36745), .Z(n36744) );
  IV U34981 ( .A(n36671), .Z(n36745) );
  XOR U34982 ( .A(n36746), .B(n36747), .Z(n36671) );
  ANDN U34983 ( .B(n36748), .A(n36749), .Z(n36746) );
  XOR U34984 ( .A(n36747), .B(n36750), .Z(n36748) );
  XOR U34985 ( .A(n36751), .B(n36679), .Z(n36691) );
  XOR U34986 ( .A(n36752), .B(n36753), .Z(n36679) );
  ANDN U34987 ( .B(n36754), .A(n36755), .Z(n36752) );
  XOR U34988 ( .A(n36753), .B(n36756), .Z(n36754) );
  IV U34989 ( .A(n36678), .Z(n36751) );
  XOR U34990 ( .A(n36757), .B(n36758), .Z(n36678) );
  XOR U34991 ( .A(n36759), .B(n36760), .Z(n36758) );
  ANDN U34992 ( .B(n36761), .A(n36762), .Z(n36759) );
  XOR U34993 ( .A(n36763), .B(n36760), .Z(n36761) );
  IV U34994 ( .A(n36676), .Z(n36757) );
  XOR U34995 ( .A(n36764), .B(n36765), .Z(n36676) );
  ANDN U34996 ( .B(n36766), .A(n36767), .Z(n36764) );
  XOR U34997 ( .A(n36765), .B(n36768), .Z(n36766) );
  IV U34998 ( .A(n36690), .Z(n36743) );
  XOR U34999 ( .A(n36769), .B(n36770), .Z(n36690) );
  XNOR U35000 ( .A(n36685), .B(n36771), .Z(n36770) );
  IV U35001 ( .A(n36688), .Z(n36771) );
  XOR U35002 ( .A(n36772), .B(n36773), .Z(n36688) );
  ANDN U35003 ( .B(n36774), .A(n36775), .Z(n36772) );
  XOR U35004 ( .A(n36776), .B(n36773), .Z(n36774) );
  XNOR U35005 ( .A(n36777), .B(n36778), .Z(n36685) );
  ANDN U35006 ( .B(n36779), .A(n36780), .Z(n36777) );
  XOR U35007 ( .A(n36778), .B(n36781), .Z(n36779) );
  IV U35008 ( .A(n36684), .Z(n36769) );
  XOR U35009 ( .A(n36682), .B(n36782), .Z(n36684) );
  XOR U35010 ( .A(n36783), .B(n36784), .Z(n36782) );
  ANDN U35011 ( .B(n36785), .A(n36786), .Z(n36783) );
  XOR U35012 ( .A(n36787), .B(n36784), .Z(n36785) );
  IV U35013 ( .A(n36686), .Z(n36682) );
  XOR U35014 ( .A(n36788), .B(n36789), .Z(n36686) );
  ANDN U35015 ( .B(n36790), .A(n36791), .Z(n36788) );
  XOR U35016 ( .A(n36792), .B(n36789), .Z(n36790) );
  IV U35017 ( .A(n36696), .Z(n36700) );
  XOR U35018 ( .A(n36696), .B(n36599), .Z(n36698) );
  XOR U35019 ( .A(n36793), .B(n36794), .Z(n36599) );
  AND U35020 ( .A(n508), .B(n36795), .Z(n36793) );
  XNOR U35021 ( .A(n36796), .B(n36794), .Z(n36795) );
  NANDN U35022 ( .A(n36601), .B(n36603), .Z(n36696) );
  XOR U35023 ( .A(n36797), .B(n36798), .Z(n36603) );
  AND U35024 ( .A(n508), .B(n36799), .Z(n36797) );
  XOR U35025 ( .A(n36798), .B(n36800), .Z(n36799) );
  XNOR U35026 ( .A(n36801), .B(n36802), .Z(n508) );
  AND U35027 ( .A(n36803), .B(n36804), .Z(n36801) );
  XOR U35028 ( .A(n36802), .B(n36614), .Z(n36804) );
  XNOR U35029 ( .A(n36805), .B(n36806), .Z(n36614) );
  ANDN U35030 ( .B(n36807), .A(n36808), .Z(n36805) );
  XOR U35031 ( .A(n36806), .B(n36809), .Z(n36807) );
  XNOR U35032 ( .A(n36802), .B(n36616), .Z(n36803) );
  XNOR U35033 ( .A(n36810), .B(n36811), .Z(n36616) );
  ANDN U35034 ( .B(n36812), .A(n36813), .Z(n36810) );
  XOR U35035 ( .A(n36811), .B(n36814), .Z(n36812) );
  XOR U35036 ( .A(n36815), .B(n36816), .Z(n36802) );
  AND U35037 ( .A(n36817), .B(n36818), .Z(n36815) );
  XOR U35038 ( .A(n36816), .B(n36641), .Z(n36818) );
  XOR U35039 ( .A(n36808), .B(n36809), .Z(n36641) );
  XNOR U35040 ( .A(n36819), .B(n36820), .Z(n36809) );
  ANDN U35041 ( .B(n36821), .A(n36822), .Z(n36819) );
  XOR U35042 ( .A(n36823), .B(n36824), .Z(n36821) );
  XOR U35043 ( .A(n36825), .B(n36826), .Z(n36808) );
  XNOR U35044 ( .A(n36827), .B(n36828), .Z(n36826) );
  ANDN U35045 ( .B(n36829), .A(n36830), .Z(n36827) );
  XNOR U35046 ( .A(n36831), .B(n36832), .Z(n36829) );
  IV U35047 ( .A(n36806), .Z(n36825) );
  XOR U35048 ( .A(n36833), .B(n36834), .Z(n36806) );
  ANDN U35049 ( .B(n36835), .A(n36836), .Z(n36833) );
  XOR U35050 ( .A(n36834), .B(n36837), .Z(n36835) );
  XOR U35051 ( .A(n36816), .B(n36643), .Z(n36817) );
  XOR U35052 ( .A(n36838), .B(n36814), .Z(n36643) );
  XNOR U35053 ( .A(n36839), .B(n36840), .Z(n36814) );
  ANDN U35054 ( .B(n36841), .A(n36842), .Z(n36839) );
  XOR U35055 ( .A(n36843), .B(n36844), .Z(n36841) );
  IV U35056 ( .A(n36813), .Z(n36838) );
  XOR U35057 ( .A(n36845), .B(n36846), .Z(n36813) );
  XNOR U35058 ( .A(n36847), .B(n36848), .Z(n36846) );
  ANDN U35059 ( .B(n36849), .A(n36850), .Z(n36847) );
  XNOR U35060 ( .A(n36851), .B(n36852), .Z(n36849) );
  IV U35061 ( .A(n36811), .Z(n36845) );
  XOR U35062 ( .A(n36853), .B(n36854), .Z(n36811) );
  ANDN U35063 ( .B(n36855), .A(n36856), .Z(n36853) );
  XOR U35064 ( .A(n36854), .B(n36857), .Z(n36855) );
  XNOR U35065 ( .A(n36858), .B(n36859), .Z(n36816) );
  AND U35066 ( .A(n36860), .B(n36861), .Z(n36858) );
  XNOR U35067 ( .A(n36859), .B(n36693), .Z(n36861) );
  XOR U35068 ( .A(n36836), .B(n36837), .Z(n36693) );
  XOR U35069 ( .A(n36862), .B(n36824), .Z(n36837) );
  XNOR U35070 ( .A(n36863), .B(n36864), .Z(n36824) );
  ANDN U35071 ( .B(n36865), .A(n36866), .Z(n36863) );
  XOR U35072 ( .A(n36867), .B(n36868), .Z(n36865) );
  IV U35073 ( .A(n36822), .Z(n36862) );
  XOR U35074 ( .A(n36820), .B(n36869), .Z(n36822) );
  XNOR U35075 ( .A(n36870), .B(n36871), .Z(n36869) );
  ANDN U35076 ( .B(n36872), .A(n36873), .Z(n36870) );
  XNOR U35077 ( .A(n36874), .B(n36875), .Z(n36872) );
  IV U35078 ( .A(n36823), .Z(n36820) );
  XOR U35079 ( .A(n36876), .B(n36877), .Z(n36823) );
  ANDN U35080 ( .B(n36878), .A(n36879), .Z(n36876) );
  XOR U35081 ( .A(n36877), .B(n36880), .Z(n36878) );
  XOR U35082 ( .A(n36881), .B(n36882), .Z(n36836) );
  XNOR U35083 ( .A(n36831), .B(n36883), .Z(n36882) );
  IV U35084 ( .A(n36834), .Z(n36883) );
  XOR U35085 ( .A(n36884), .B(n36885), .Z(n36834) );
  ANDN U35086 ( .B(n36886), .A(n36887), .Z(n36884) );
  XOR U35087 ( .A(n36885), .B(n36888), .Z(n36886) );
  XNOR U35088 ( .A(n36889), .B(n36890), .Z(n36831) );
  ANDN U35089 ( .B(n36891), .A(n36892), .Z(n36889) );
  XOR U35090 ( .A(n36890), .B(n36893), .Z(n36891) );
  IV U35091 ( .A(n36830), .Z(n36881) );
  XOR U35092 ( .A(n36828), .B(n36894), .Z(n36830) );
  XNOR U35093 ( .A(n36895), .B(n36896), .Z(n36894) );
  ANDN U35094 ( .B(n36897), .A(n36898), .Z(n36895) );
  XNOR U35095 ( .A(n36899), .B(n36900), .Z(n36897) );
  IV U35096 ( .A(n36832), .Z(n36828) );
  XOR U35097 ( .A(n36901), .B(n36902), .Z(n36832) );
  ANDN U35098 ( .B(n36903), .A(n36904), .Z(n36901) );
  XOR U35099 ( .A(n36905), .B(n36902), .Z(n36903) );
  XNOR U35100 ( .A(n36859), .B(n36695), .Z(n36860) );
  XOR U35101 ( .A(n36906), .B(n36857), .Z(n36695) );
  XOR U35102 ( .A(n36907), .B(n36844), .Z(n36857) );
  XNOR U35103 ( .A(n36908), .B(n36909), .Z(n36844) );
  ANDN U35104 ( .B(n36910), .A(n36911), .Z(n36908) );
  XOR U35105 ( .A(n36912), .B(n36913), .Z(n36910) );
  IV U35106 ( .A(n36842), .Z(n36907) );
  XOR U35107 ( .A(n36840), .B(n36914), .Z(n36842) );
  XNOR U35108 ( .A(n36915), .B(n36916), .Z(n36914) );
  ANDN U35109 ( .B(n36917), .A(n36918), .Z(n36915) );
  XNOR U35110 ( .A(n36919), .B(n36920), .Z(n36917) );
  IV U35111 ( .A(n36843), .Z(n36840) );
  XOR U35112 ( .A(n36921), .B(n36922), .Z(n36843) );
  ANDN U35113 ( .B(n36923), .A(n36924), .Z(n36921) );
  XOR U35114 ( .A(n36922), .B(n36925), .Z(n36923) );
  IV U35115 ( .A(n36856), .Z(n36906) );
  XOR U35116 ( .A(n36926), .B(n36927), .Z(n36856) );
  XNOR U35117 ( .A(n36851), .B(n36928), .Z(n36927) );
  IV U35118 ( .A(n36854), .Z(n36928) );
  XOR U35119 ( .A(n36929), .B(n36930), .Z(n36854) );
  ANDN U35120 ( .B(n36931), .A(n36932), .Z(n36929) );
  XOR U35121 ( .A(n36930), .B(n36933), .Z(n36931) );
  XNOR U35122 ( .A(n36934), .B(n36935), .Z(n36851) );
  ANDN U35123 ( .B(n36936), .A(n36937), .Z(n36934) );
  XOR U35124 ( .A(n36935), .B(n36938), .Z(n36936) );
  IV U35125 ( .A(n36850), .Z(n36926) );
  XOR U35126 ( .A(n36848), .B(n36939), .Z(n36850) );
  XNOR U35127 ( .A(n36940), .B(n36941), .Z(n36939) );
  ANDN U35128 ( .B(n36942), .A(n36943), .Z(n36940) );
  XNOR U35129 ( .A(n36944), .B(n36945), .Z(n36942) );
  IV U35130 ( .A(n36852), .Z(n36848) );
  XOR U35131 ( .A(n36946), .B(n36947), .Z(n36852) );
  ANDN U35132 ( .B(n36948), .A(n36949), .Z(n36946) );
  XOR U35133 ( .A(n36950), .B(n36947), .Z(n36948) );
  XNOR U35134 ( .A(n36951), .B(n36952), .Z(n36859) );
  NAND U35135 ( .A(n36953), .B(n36954), .Z(n36952) );
  XOR U35136 ( .A(n36955), .B(n36794), .Z(n36954) );
  XOR U35137 ( .A(n36887), .B(n36888), .Z(n36794) );
  XOR U35138 ( .A(n36956), .B(n36880), .Z(n36888) );
  XOR U35139 ( .A(n36957), .B(n36868), .Z(n36880) );
  XOR U35140 ( .A(n36958), .B(n36959), .Z(n36868) );
  ANDN U35141 ( .B(n36960), .A(n36961), .Z(n36958) );
  XOR U35142 ( .A(n36959), .B(n36962), .Z(n36960) );
  IV U35143 ( .A(n36866), .Z(n36957) );
  XOR U35144 ( .A(n36864), .B(n36963), .Z(n36866) );
  XOR U35145 ( .A(n36964), .B(n36965), .Z(n36963) );
  ANDN U35146 ( .B(n36966), .A(n36967), .Z(n36964) );
  XOR U35147 ( .A(n36968), .B(n36965), .Z(n36966) );
  IV U35148 ( .A(n36867), .Z(n36864) );
  XOR U35149 ( .A(n36969), .B(n36970), .Z(n36867) );
  ANDN U35150 ( .B(n36971), .A(n36972), .Z(n36969) );
  XOR U35151 ( .A(n36970), .B(n36973), .Z(n36971) );
  IV U35152 ( .A(n36879), .Z(n36956) );
  XOR U35153 ( .A(n36974), .B(n36975), .Z(n36879) );
  XNOR U35154 ( .A(n36874), .B(n36976), .Z(n36975) );
  IV U35155 ( .A(n36877), .Z(n36976) );
  XOR U35156 ( .A(n36977), .B(n36978), .Z(n36877) );
  ANDN U35157 ( .B(n36979), .A(n36980), .Z(n36977) );
  XOR U35158 ( .A(n36978), .B(n36981), .Z(n36979) );
  XNOR U35159 ( .A(n36982), .B(n36983), .Z(n36874) );
  ANDN U35160 ( .B(n36984), .A(n36985), .Z(n36982) );
  XOR U35161 ( .A(n36983), .B(n36986), .Z(n36984) );
  IV U35162 ( .A(n36873), .Z(n36974) );
  XOR U35163 ( .A(n36871), .B(n36987), .Z(n36873) );
  XOR U35164 ( .A(n36988), .B(n36989), .Z(n36987) );
  ANDN U35165 ( .B(n36990), .A(n36991), .Z(n36988) );
  XOR U35166 ( .A(n36992), .B(n36989), .Z(n36990) );
  IV U35167 ( .A(n36875), .Z(n36871) );
  XOR U35168 ( .A(n36993), .B(n36994), .Z(n36875) );
  ANDN U35169 ( .B(n36995), .A(n36996), .Z(n36993) );
  XOR U35170 ( .A(n36997), .B(n36994), .Z(n36995) );
  XOR U35171 ( .A(n36998), .B(n36999), .Z(n36887) );
  XOR U35172 ( .A(n36905), .B(n37000), .Z(n36999) );
  IV U35173 ( .A(n36885), .Z(n37000) );
  XOR U35174 ( .A(n37001), .B(n37002), .Z(n36885) );
  ANDN U35175 ( .B(n37003), .A(n37004), .Z(n37001) );
  XOR U35176 ( .A(n37002), .B(n37005), .Z(n37003) );
  XOR U35177 ( .A(n37006), .B(n36893), .Z(n36905) );
  XOR U35178 ( .A(n37007), .B(n37008), .Z(n36893) );
  ANDN U35179 ( .B(n37009), .A(n37010), .Z(n37007) );
  XOR U35180 ( .A(n37008), .B(n37011), .Z(n37009) );
  IV U35181 ( .A(n36892), .Z(n37006) );
  XOR U35182 ( .A(n37012), .B(n37013), .Z(n36892) );
  XOR U35183 ( .A(n37014), .B(n37015), .Z(n37013) );
  ANDN U35184 ( .B(n37016), .A(n37017), .Z(n37014) );
  XOR U35185 ( .A(n37018), .B(n37015), .Z(n37016) );
  IV U35186 ( .A(n36890), .Z(n37012) );
  XOR U35187 ( .A(n37019), .B(n37020), .Z(n36890) );
  ANDN U35188 ( .B(n37021), .A(n37022), .Z(n37019) );
  XOR U35189 ( .A(n37020), .B(n37023), .Z(n37021) );
  IV U35190 ( .A(n36904), .Z(n36998) );
  XOR U35191 ( .A(n37024), .B(n37025), .Z(n36904) );
  XNOR U35192 ( .A(n36899), .B(n37026), .Z(n37025) );
  IV U35193 ( .A(n36902), .Z(n37026) );
  XOR U35194 ( .A(n37027), .B(n37028), .Z(n36902) );
  ANDN U35195 ( .B(n37029), .A(n37030), .Z(n37027) );
  XOR U35196 ( .A(n37031), .B(n37028), .Z(n37029) );
  XNOR U35197 ( .A(n37032), .B(n37033), .Z(n36899) );
  ANDN U35198 ( .B(n37034), .A(n37035), .Z(n37032) );
  XOR U35199 ( .A(n37033), .B(n37036), .Z(n37034) );
  IV U35200 ( .A(n36898), .Z(n37024) );
  XOR U35201 ( .A(n36896), .B(n37037), .Z(n36898) );
  XOR U35202 ( .A(n37038), .B(n37039), .Z(n37037) );
  ANDN U35203 ( .B(n37040), .A(n37041), .Z(n37038) );
  XOR U35204 ( .A(n37042), .B(n37039), .Z(n37040) );
  IV U35205 ( .A(n36900), .Z(n36896) );
  XOR U35206 ( .A(n37043), .B(n37044), .Z(n36900) );
  ANDN U35207 ( .B(n37045), .A(n37046), .Z(n37043) );
  XOR U35208 ( .A(n37047), .B(n37044), .Z(n37045) );
  IV U35209 ( .A(n36951), .Z(n36955) );
  XNOR U35210 ( .A(n36951), .B(n36796), .Z(n36953) );
  XOR U35211 ( .A(n37048), .B(n36933), .Z(n36796) );
  XOR U35212 ( .A(n37049), .B(n36925), .Z(n36933) );
  XOR U35213 ( .A(n37050), .B(n36913), .Z(n36925) );
  XOR U35214 ( .A(n37051), .B(n37052), .Z(n36913) );
  ANDN U35215 ( .B(n37053), .A(n37054), .Z(n37051) );
  XOR U35216 ( .A(n37052), .B(n37055), .Z(n37053) );
  IV U35217 ( .A(n36911), .Z(n37050) );
  XOR U35218 ( .A(n36909), .B(n37056), .Z(n36911) );
  XOR U35219 ( .A(n37057), .B(n37058), .Z(n37056) );
  ANDN U35220 ( .B(n37059), .A(n37060), .Z(n37057) );
  XOR U35221 ( .A(n37061), .B(n37058), .Z(n37059) );
  IV U35222 ( .A(n36912), .Z(n36909) );
  XOR U35223 ( .A(n37062), .B(n37063), .Z(n36912) );
  ANDN U35224 ( .B(n37064), .A(n37065), .Z(n37062) );
  XOR U35225 ( .A(n37063), .B(n37066), .Z(n37064) );
  IV U35226 ( .A(n36924), .Z(n37049) );
  XOR U35227 ( .A(n37067), .B(n37068), .Z(n36924) );
  XNOR U35228 ( .A(n36919), .B(n37069), .Z(n37068) );
  IV U35229 ( .A(n36922), .Z(n37069) );
  XOR U35230 ( .A(n37070), .B(n37071), .Z(n36922) );
  ANDN U35231 ( .B(n37072), .A(n37073), .Z(n37070) );
  XOR U35232 ( .A(n37071), .B(n37074), .Z(n37072) );
  XNOR U35233 ( .A(n37075), .B(n37076), .Z(n36919) );
  ANDN U35234 ( .B(n37077), .A(n37078), .Z(n37075) );
  XOR U35235 ( .A(n37076), .B(n37079), .Z(n37077) );
  IV U35236 ( .A(n36918), .Z(n37067) );
  XOR U35237 ( .A(n36916), .B(n37080), .Z(n36918) );
  XOR U35238 ( .A(n37081), .B(n37082), .Z(n37080) );
  ANDN U35239 ( .B(n37083), .A(n37084), .Z(n37081) );
  XOR U35240 ( .A(n37085), .B(n37082), .Z(n37083) );
  IV U35241 ( .A(n36920), .Z(n36916) );
  XOR U35242 ( .A(n37086), .B(n37087), .Z(n36920) );
  ANDN U35243 ( .B(n37088), .A(n37089), .Z(n37086) );
  XOR U35244 ( .A(n37090), .B(n37087), .Z(n37088) );
  IV U35245 ( .A(n36932), .Z(n37048) );
  XOR U35246 ( .A(n37091), .B(n37092), .Z(n36932) );
  XOR U35247 ( .A(n36950), .B(n37093), .Z(n37092) );
  IV U35248 ( .A(n36930), .Z(n37093) );
  XNOR U35249 ( .A(n37094), .B(n37095), .Z(n36930) );
  ANDN U35250 ( .B(n37096), .A(n37097), .Z(n37094) );
  XNOR U35251 ( .A(n37095), .B(n37098), .Z(n37096) );
  XOR U35252 ( .A(n37099), .B(n36938), .Z(n36950) );
  XOR U35253 ( .A(n37100), .B(n37101), .Z(n36938) );
  ANDN U35254 ( .B(n37102), .A(n37103), .Z(n37100) );
  XOR U35255 ( .A(n37101), .B(n37104), .Z(n37102) );
  IV U35256 ( .A(n36937), .Z(n37099) );
  XOR U35257 ( .A(n37105), .B(n37106), .Z(n36937) );
  XOR U35258 ( .A(n37107), .B(n37108), .Z(n37106) );
  ANDN U35259 ( .B(n37109), .A(n37110), .Z(n37107) );
  XOR U35260 ( .A(n37111), .B(n37108), .Z(n37109) );
  IV U35261 ( .A(n36935), .Z(n37105) );
  XNOR U35262 ( .A(n37112), .B(n37113), .Z(n36935) );
  ANDN U35263 ( .B(n37114), .A(n37115), .Z(n37112) );
  XNOR U35264 ( .A(n37113), .B(n37116), .Z(n37114) );
  IV U35265 ( .A(n36949), .Z(n37091) );
  XOR U35266 ( .A(n37117), .B(n37118), .Z(n36949) );
  XNOR U35267 ( .A(n36944), .B(n37119), .Z(n37118) );
  IV U35268 ( .A(n36947), .Z(n37119) );
  XOR U35269 ( .A(n37120), .B(n37121), .Z(n36947) );
  ANDN U35270 ( .B(n37122), .A(n37123), .Z(n37120) );
  XOR U35271 ( .A(n37124), .B(n37121), .Z(n37122) );
  XNOR U35272 ( .A(n37125), .B(n37126), .Z(n36944) );
  ANDN U35273 ( .B(n37127), .A(n37128), .Z(n37125) );
  XOR U35274 ( .A(n37126), .B(n37129), .Z(n37127) );
  IV U35275 ( .A(n36943), .Z(n37117) );
  XOR U35276 ( .A(n36941), .B(n37130), .Z(n36943) );
  XOR U35277 ( .A(n37131), .B(n37132), .Z(n37130) );
  ANDN U35278 ( .B(n37133), .A(n37134), .Z(n37131) );
  XOR U35279 ( .A(n37135), .B(n37132), .Z(n37133) );
  IV U35280 ( .A(n36945), .Z(n36941) );
  XOR U35281 ( .A(n37136), .B(n37137), .Z(n36945) );
  ANDN U35282 ( .B(n37138), .A(n37139), .Z(n37136) );
  XOR U35283 ( .A(n37140), .B(n37137), .Z(n37138) );
  NANDN U35284 ( .A(n36798), .B(n36800), .Z(n36951) );
  XOR U35285 ( .A(n37141), .B(n37098), .Z(n36800) );
  XOR U35286 ( .A(n37142), .B(n37074), .Z(n37098) );
  XOR U35287 ( .A(n37143), .B(n37066), .Z(n37074) );
  XOR U35288 ( .A(n37144), .B(n37055), .Z(n37066) );
  XNOR U35289 ( .A(q[30]), .B(DB[30]), .Z(n37055) );
  IV U35290 ( .A(n37054), .Z(n37144) );
  XNOR U35291 ( .A(n37052), .B(n37145), .Z(n37054) );
  XNOR U35292 ( .A(q[29]), .B(DB[29]), .Z(n37145) );
  XNOR U35293 ( .A(q[28]), .B(DB[28]), .Z(n37052) );
  IV U35294 ( .A(n37065), .Z(n37143) );
  XOR U35295 ( .A(n37146), .B(n37147), .Z(n37065) );
  XNOR U35296 ( .A(n37061), .B(n37063), .Z(n37147) );
  XNOR U35297 ( .A(q[24]), .B(DB[24]), .Z(n37063) );
  XNOR U35298 ( .A(q[27]), .B(DB[27]), .Z(n37061) );
  IV U35299 ( .A(n37060), .Z(n37146) );
  XNOR U35300 ( .A(n37058), .B(n37148), .Z(n37060) );
  XNOR U35301 ( .A(q[26]), .B(DB[26]), .Z(n37148) );
  XNOR U35302 ( .A(q[25]), .B(DB[25]), .Z(n37058) );
  IV U35303 ( .A(n37073), .Z(n37142) );
  XOR U35304 ( .A(n37149), .B(n37150), .Z(n37073) );
  XNOR U35305 ( .A(n37090), .B(n37071), .Z(n37150) );
  XNOR U35306 ( .A(q[16]), .B(DB[16]), .Z(n37071) );
  XOR U35307 ( .A(n37151), .B(n37079), .Z(n37090) );
  XNOR U35308 ( .A(q[23]), .B(DB[23]), .Z(n37079) );
  IV U35309 ( .A(n37078), .Z(n37151) );
  XNOR U35310 ( .A(n37076), .B(n37152), .Z(n37078) );
  XNOR U35311 ( .A(q[22]), .B(DB[22]), .Z(n37152) );
  XNOR U35312 ( .A(q[21]), .B(DB[21]), .Z(n37076) );
  IV U35313 ( .A(n37089), .Z(n37149) );
  XOR U35314 ( .A(n37153), .B(n37154), .Z(n37089) );
  XNOR U35315 ( .A(n37085), .B(n37087), .Z(n37154) );
  XNOR U35316 ( .A(q[17]), .B(DB[17]), .Z(n37087) );
  XNOR U35317 ( .A(q[20]), .B(DB[20]), .Z(n37085) );
  IV U35318 ( .A(n37084), .Z(n37153) );
  XNOR U35319 ( .A(n37082), .B(n37155), .Z(n37084) );
  XNOR U35320 ( .A(q[19]), .B(DB[19]), .Z(n37155) );
  XNOR U35321 ( .A(q[18]), .B(DB[18]), .Z(n37082) );
  IV U35322 ( .A(n37097), .Z(n37141) );
  XOR U35323 ( .A(n37156), .B(n37157), .Z(n37097) );
  XOR U35324 ( .A(n37095), .B(n37124), .Z(n37157) );
  XOR U35325 ( .A(n37158), .B(n37116), .Z(n37124) );
  XOR U35326 ( .A(n37159), .B(n37104), .Z(n37116) );
  XNOR U35327 ( .A(q[15]), .B(DB[15]), .Z(n37104) );
  IV U35328 ( .A(n37103), .Z(n37159) );
  XNOR U35329 ( .A(n37101), .B(n37160), .Z(n37103) );
  XNOR U35330 ( .A(q[14]), .B(DB[14]), .Z(n37160) );
  XNOR U35331 ( .A(q[13]), .B(DB[13]), .Z(n37101) );
  IV U35332 ( .A(n37115), .Z(n37158) );
  XOR U35333 ( .A(n37161), .B(n37162), .Z(n37115) );
  XOR U35334 ( .A(n37113), .B(n37111), .Z(n37162) );
  XNOR U35335 ( .A(q[12]), .B(DB[12]), .Z(n37111) );
  XOR U35336 ( .A(q[9]), .B(DB[9]), .Z(n37113) );
  IV U35337 ( .A(n37110), .Z(n37161) );
  XNOR U35338 ( .A(n37108), .B(n37163), .Z(n37110) );
  XNOR U35339 ( .A(q[11]), .B(DB[11]), .Z(n37163) );
  XNOR U35340 ( .A(q[10]), .B(DB[10]), .Z(n37108) );
  XOR U35341 ( .A(q[0]), .B(DB[0]), .Z(n37095) );
  IV U35342 ( .A(n37123), .Z(n37156) );
  XOR U35343 ( .A(n37164), .B(n37165), .Z(n37123) );
  XNOR U35344 ( .A(n37140), .B(n37121), .Z(n37165) );
  XNOR U35345 ( .A(q[1]), .B(DB[1]), .Z(n37121) );
  XOR U35346 ( .A(n37166), .B(n37129), .Z(n37140) );
  XNOR U35347 ( .A(q[8]), .B(DB[8]), .Z(n37129) );
  IV U35348 ( .A(n37128), .Z(n37166) );
  XNOR U35349 ( .A(n37126), .B(n37167), .Z(n37128) );
  XNOR U35350 ( .A(q[7]), .B(DB[7]), .Z(n37167) );
  XNOR U35351 ( .A(q[6]), .B(DB[6]), .Z(n37126) );
  IV U35352 ( .A(n37139), .Z(n37164) );
  XOR U35353 ( .A(n37168), .B(n37169), .Z(n37139) );
  XNOR U35354 ( .A(n37135), .B(n37137), .Z(n37169) );
  XNOR U35355 ( .A(q[2]), .B(DB[2]), .Z(n37137) );
  XNOR U35356 ( .A(q[5]), .B(DB[5]), .Z(n37135) );
  IV U35357 ( .A(n37134), .Z(n37168) );
  XNOR U35358 ( .A(n37132), .B(n37170), .Z(n37134) );
  XNOR U35359 ( .A(q[4]), .B(DB[4]), .Z(n37170) );
  XNOR U35360 ( .A(q[3]), .B(DB[3]), .Z(n37132) );
  XOR U35361 ( .A(n37171), .B(n37005), .Z(n36798) );
  XOR U35362 ( .A(n37172), .B(n36981), .Z(n37005) );
  XOR U35363 ( .A(n37173), .B(n36973), .Z(n36981) );
  XOR U35364 ( .A(n37174), .B(n36962), .Z(n36973) );
  XNOR U35365 ( .A(q[30]), .B(DB[61]), .Z(n36962) );
  IV U35366 ( .A(n36961), .Z(n37174) );
  XNOR U35367 ( .A(n36959), .B(n37175), .Z(n36961) );
  XNOR U35368 ( .A(q[29]), .B(DB[60]), .Z(n37175) );
  XNOR U35369 ( .A(q[28]), .B(DB[59]), .Z(n36959) );
  IV U35370 ( .A(n36972), .Z(n37173) );
  XOR U35371 ( .A(n37176), .B(n37177), .Z(n36972) );
  XNOR U35372 ( .A(n36968), .B(n36970), .Z(n37177) );
  XNOR U35373 ( .A(q[24]), .B(DB[55]), .Z(n36970) );
  XNOR U35374 ( .A(q[27]), .B(DB[58]), .Z(n36968) );
  IV U35375 ( .A(n36967), .Z(n37176) );
  XNOR U35376 ( .A(n36965), .B(n37178), .Z(n36967) );
  XNOR U35377 ( .A(q[26]), .B(DB[57]), .Z(n37178) );
  XNOR U35378 ( .A(q[25]), .B(DB[56]), .Z(n36965) );
  IV U35379 ( .A(n36980), .Z(n37172) );
  XOR U35380 ( .A(n37179), .B(n37180), .Z(n36980) );
  XNOR U35381 ( .A(n36997), .B(n36978), .Z(n37180) );
  XNOR U35382 ( .A(q[16]), .B(DB[47]), .Z(n36978) );
  XOR U35383 ( .A(n37181), .B(n36986), .Z(n36997) );
  XNOR U35384 ( .A(q[23]), .B(DB[54]), .Z(n36986) );
  IV U35385 ( .A(n36985), .Z(n37181) );
  XNOR U35386 ( .A(n36983), .B(n37182), .Z(n36985) );
  XNOR U35387 ( .A(q[22]), .B(DB[53]), .Z(n37182) );
  XNOR U35388 ( .A(q[21]), .B(DB[52]), .Z(n36983) );
  IV U35389 ( .A(n36996), .Z(n37179) );
  XOR U35390 ( .A(n37183), .B(n37184), .Z(n36996) );
  XNOR U35391 ( .A(n36992), .B(n36994), .Z(n37184) );
  XNOR U35392 ( .A(q[17]), .B(DB[48]), .Z(n36994) );
  XNOR U35393 ( .A(q[20]), .B(DB[51]), .Z(n36992) );
  IV U35394 ( .A(n36991), .Z(n37183) );
  XNOR U35395 ( .A(n36989), .B(n37185), .Z(n36991) );
  XNOR U35396 ( .A(q[19]), .B(DB[50]), .Z(n37185) );
  XNOR U35397 ( .A(q[18]), .B(DB[49]), .Z(n36989) );
  IV U35398 ( .A(n37004), .Z(n37171) );
  XOR U35399 ( .A(n37186), .B(n37187), .Z(n37004) );
  XNOR U35400 ( .A(n37031), .B(n37002), .Z(n37187) );
  XNOR U35401 ( .A(q[0]), .B(DB[31]), .Z(n37002) );
  XOR U35402 ( .A(n37188), .B(n37023), .Z(n37031) );
  XOR U35403 ( .A(n37189), .B(n37011), .Z(n37023) );
  XNOR U35404 ( .A(q[15]), .B(DB[46]), .Z(n37011) );
  IV U35405 ( .A(n37010), .Z(n37189) );
  XNOR U35406 ( .A(n37008), .B(n37190), .Z(n37010) );
  XNOR U35407 ( .A(q[14]), .B(DB[45]), .Z(n37190) );
  XNOR U35408 ( .A(q[13]), .B(DB[44]), .Z(n37008) );
  IV U35409 ( .A(n37022), .Z(n37188) );
  XOR U35410 ( .A(n37191), .B(n37192), .Z(n37022) );
  XNOR U35411 ( .A(n37018), .B(n37020), .Z(n37192) );
  XNOR U35412 ( .A(q[9]), .B(DB[40]), .Z(n37020) );
  XNOR U35413 ( .A(q[12]), .B(DB[43]), .Z(n37018) );
  IV U35414 ( .A(n37017), .Z(n37191) );
  XNOR U35415 ( .A(n37015), .B(n37193), .Z(n37017) );
  XNOR U35416 ( .A(q[11]), .B(DB[42]), .Z(n37193) );
  XNOR U35417 ( .A(q[10]), .B(DB[41]), .Z(n37015) );
  IV U35418 ( .A(n37030), .Z(n37186) );
  XOR U35419 ( .A(n37194), .B(n37195), .Z(n37030) );
  XNOR U35420 ( .A(n37047), .B(n37028), .Z(n37195) );
  XNOR U35421 ( .A(q[1]), .B(DB[32]), .Z(n37028) );
  XOR U35422 ( .A(n37196), .B(n37036), .Z(n37047) );
  XNOR U35423 ( .A(q[8]), .B(DB[39]), .Z(n37036) );
  IV U35424 ( .A(n37035), .Z(n37196) );
  XNOR U35425 ( .A(n37033), .B(n37197), .Z(n37035) );
  XNOR U35426 ( .A(q[7]), .B(DB[38]), .Z(n37197) );
  XNOR U35427 ( .A(q[6]), .B(DB[37]), .Z(n37033) );
  IV U35428 ( .A(n37046), .Z(n37194) );
  XOR U35429 ( .A(n37198), .B(n37199), .Z(n37046) );
  XNOR U35430 ( .A(n37042), .B(n37044), .Z(n37199) );
  XNOR U35431 ( .A(q[2]), .B(DB[33]), .Z(n37044) );
  XNOR U35432 ( .A(q[5]), .B(DB[36]), .Z(n37042) );
  IV U35433 ( .A(n37041), .Z(n37198) );
  XNOR U35434 ( .A(n37039), .B(n37200), .Z(n37041) );
  XNOR U35435 ( .A(q[4]), .B(DB[35]), .Z(n37200) );
  XNOR U35436 ( .A(q[3]), .B(DB[34]), .Z(n37039) );
  XOR U35437 ( .A(n37201), .B(n36750), .Z(n36601) );
  XOR U35438 ( .A(n37202), .B(n36726), .Z(n36750) );
  XOR U35439 ( .A(n37203), .B(n36718), .Z(n36726) );
  XOR U35440 ( .A(n37204), .B(n36707), .Z(n36718) );
  XNOR U35441 ( .A(q[30]), .B(DB[92]), .Z(n36707) );
  IV U35442 ( .A(n36706), .Z(n37204) );
  XNOR U35443 ( .A(n36704), .B(n37205), .Z(n36706) );
  XNOR U35444 ( .A(q[29]), .B(DB[91]), .Z(n37205) );
  XNOR U35445 ( .A(q[28]), .B(DB[90]), .Z(n36704) );
  IV U35446 ( .A(n36717), .Z(n37203) );
  XOR U35447 ( .A(n37206), .B(n37207), .Z(n36717) );
  XNOR U35448 ( .A(n36713), .B(n36715), .Z(n37207) );
  XNOR U35449 ( .A(q[24]), .B(DB[86]), .Z(n36715) );
  XNOR U35450 ( .A(q[27]), .B(DB[89]), .Z(n36713) );
  IV U35451 ( .A(n36712), .Z(n37206) );
  XNOR U35452 ( .A(n36710), .B(n37208), .Z(n36712) );
  XNOR U35453 ( .A(q[26]), .B(DB[88]), .Z(n37208) );
  XNOR U35454 ( .A(q[25]), .B(DB[87]), .Z(n36710) );
  IV U35455 ( .A(n36725), .Z(n37202) );
  XOR U35456 ( .A(n37209), .B(n37210), .Z(n36725) );
  XNOR U35457 ( .A(n36742), .B(n36723), .Z(n37210) );
  XNOR U35458 ( .A(q[16]), .B(DB[78]), .Z(n36723) );
  XOR U35459 ( .A(n37211), .B(n36731), .Z(n36742) );
  XNOR U35460 ( .A(q[23]), .B(DB[85]), .Z(n36731) );
  IV U35461 ( .A(n36730), .Z(n37211) );
  XNOR U35462 ( .A(n36728), .B(n37212), .Z(n36730) );
  XNOR U35463 ( .A(q[22]), .B(DB[84]), .Z(n37212) );
  XNOR U35464 ( .A(q[21]), .B(DB[83]), .Z(n36728) );
  IV U35465 ( .A(n36741), .Z(n37209) );
  XOR U35466 ( .A(n37213), .B(n37214), .Z(n36741) );
  XNOR U35467 ( .A(n36737), .B(n36739), .Z(n37214) );
  XNOR U35468 ( .A(q[17]), .B(DB[79]), .Z(n36739) );
  XNOR U35469 ( .A(q[20]), .B(DB[82]), .Z(n36737) );
  IV U35470 ( .A(n36736), .Z(n37213) );
  XNOR U35471 ( .A(n36734), .B(n37215), .Z(n36736) );
  XNOR U35472 ( .A(q[19]), .B(DB[81]), .Z(n37215) );
  XNOR U35473 ( .A(q[18]), .B(DB[80]), .Z(n36734) );
  IV U35474 ( .A(n36749), .Z(n37201) );
  XOR U35475 ( .A(n37216), .B(n37217), .Z(n36749) );
  XNOR U35476 ( .A(n36776), .B(n36747), .Z(n37217) );
  XNOR U35477 ( .A(q[0]), .B(DB[62]), .Z(n36747) );
  XOR U35478 ( .A(n37218), .B(n36768), .Z(n36776) );
  XOR U35479 ( .A(n37219), .B(n36756), .Z(n36768) );
  XNOR U35480 ( .A(q[15]), .B(DB[77]), .Z(n36756) );
  IV U35481 ( .A(n36755), .Z(n37219) );
  XNOR U35482 ( .A(n36753), .B(n37220), .Z(n36755) );
  XNOR U35483 ( .A(q[14]), .B(DB[76]), .Z(n37220) );
  XNOR U35484 ( .A(q[13]), .B(DB[75]), .Z(n36753) );
  IV U35485 ( .A(n36767), .Z(n37218) );
  XOR U35486 ( .A(n37221), .B(n37222), .Z(n36767) );
  XNOR U35487 ( .A(n36763), .B(n36765), .Z(n37222) );
  XNOR U35488 ( .A(q[9]), .B(DB[71]), .Z(n36765) );
  XNOR U35489 ( .A(q[12]), .B(DB[74]), .Z(n36763) );
  IV U35490 ( .A(n36762), .Z(n37221) );
  XNOR U35491 ( .A(n36760), .B(n37223), .Z(n36762) );
  XNOR U35492 ( .A(q[11]), .B(DB[73]), .Z(n37223) );
  XNOR U35493 ( .A(q[10]), .B(DB[72]), .Z(n36760) );
  IV U35494 ( .A(n36775), .Z(n37216) );
  XOR U35495 ( .A(n37224), .B(n37225), .Z(n36775) );
  XNOR U35496 ( .A(n36792), .B(n36773), .Z(n37225) );
  XNOR U35497 ( .A(q[1]), .B(DB[63]), .Z(n36773) );
  XOR U35498 ( .A(n37226), .B(n36781), .Z(n36792) );
  XNOR U35499 ( .A(q[8]), .B(DB[70]), .Z(n36781) );
  IV U35500 ( .A(n36780), .Z(n37226) );
  XNOR U35501 ( .A(n36778), .B(n37227), .Z(n36780) );
  XNOR U35502 ( .A(q[7]), .B(DB[69]), .Z(n37227) );
  XNOR U35503 ( .A(q[6]), .B(DB[68]), .Z(n36778) );
  IV U35504 ( .A(n36791), .Z(n37224) );
  XOR U35505 ( .A(n37228), .B(n37229), .Z(n36791) );
  XNOR U35506 ( .A(n36787), .B(n36789), .Z(n37229) );
  XNOR U35507 ( .A(q[2]), .B(DB[64]), .Z(n36789) );
  XNOR U35508 ( .A(q[5]), .B(DB[67]), .Z(n36787) );
  IV U35509 ( .A(n36786), .Z(n37228) );
  XNOR U35510 ( .A(n36784), .B(n37230), .Z(n36786) );
  XNOR U35511 ( .A(q[4]), .B(DB[66]), .Z(n37230) );
  XNOR U35512 ( .A(q[3]), .B(DB[65]), .Z(n36784) );
  XOR U35513 ( .A(n37231), .B(n36553), .Z(n36404) );
  XOR U35514 ( .A(n37232), .B(n36529), .Z(n36553) );
  XOR U35515 ( .A(n37233), .B(n36521), .Z(n36529) );
  XOR U35516 ( .A(n37234), .B(n36510), .Z(n36521) );
  XNOR U35517 ( .A(q[30]), .B(DB[123]), .Z(n36510) );
  IV U35518 ( .A(n36509), .Z(n37234) );
  XNOR U35519 ( .A(n36507), .B(n37235), .Z(n36509) );
  XNOR U35520 ( .A(q[29]), .B(DB[122]), .Z(n37235) );
  XNOR U35521 ( .A(q[28]), .B(DB[121]), .Z(n36507) );
  IV U35522 ( .A(n36520), .Z(n37233) );
  XOR U35523 ( .A(n37236), .B(n37237), .Z(n36520) );
  XNOR U35524 ( .A(n36516), .B(n36518), .Z(n37237) );
  XNOR U35525 ( .A(q[24]), .B(DB[117]), .Z(n36518) );
  XNOR U35526 ( .A(q[27]), .B(DB[120]), .Z(n36516) );
  IV U35527 ( .A(n36515), .Z(n37236) );
  XNOR U35528 ( .A(n36513), .B(n37238), .Z(n36515) );
  XNOR U35529 ( .A(q[26]), .B(DB[119]), .Z(n37238) );
  XNOR U35530 ( .A(q[25]), .B(DB[118]), .Z(n36513) );
  IV U35531 ( .A(n36528), .Z(n37232) );
  XOR U35532 ( .A(n37239), .B(n37240), .Z(n36528) );
  XNOR U35533 ( .A(n36545), .B(n36526), .Z(n37240) );
  XNOR U35534 ( .A(q[16]), .B(DB[109]), .Z(n36526) );
  XOR U35535 ( .A(n37241), .B(n36534), .Z(n36545) );
  XNOR U35536 ( .A(q[23]), .B(DB[116]), .Z(n36534) );
  IV U35537 ( .A(n36533), .Z(n37241) );
  XNOR U35538 ( .A(n36531), .B(n37242), .Z(n36533) );
  XNOR U35539 ( .A(q[22]), .B(DB[115]), .Z(n37242) );
  XNOR U35540 ( .A(q[21]), .B(DB[114]), .Z(n36531) );
  IV U35541 ( .A(n36544), .Z(n37239) );
  XOR U35542 ( .A(n37243), .B(n37244), .Z(n36544) );
  XNOR U35543 ( .A(n36540), .B(n36542), .Z(n37244) );
  XNOR U35544 ( .A(q[17]), .B(DB[110]), .Z(n36542) );
  XNOR U35545 ( .A(q[20]), .B(DB[113]), .Z(n36540) );
  IV U35546 ( .A(n36539), .Z(n37243) );
  XNOR U35547 ( .A(n36537), .B(n37245), .Z(n36539) );
  XNOR U35548 ( .A(q[19]), .B(DB[112]), .Z(n37245) );
  XNOR U35549 ( .A(q[18]), .B(DB[111]), .Z(n36537) );
  IV U35550 ( .A(n36552), .Z(n37231) );
  XOR U35551 ( .A(n37246), .B(n37247), .Z(n36552) );
  XNOR U35552 ( .A(n36579), .B(n36550), .Z(n37247) );
  XNOR U35553 ( .A(q[0]), .B(DB[93]), .Z(n36550) );
  XOR U35554 ( .A(n37248), .B(n36571), .Z(n36579) );
  XOR U35555 ( .A(n37249), .B(n36559), .Z(n36571) );
  XNOR U35556 ( .A(q[15]), .B(DB[108]), .Z(n36559) );
  IV U35557 ( .A(n36558), .Z(n37249) );
  XNOR U35558 ( .A(n36556), .B(n37250), .Z(n36558) );
  XNOR U35559 ( .A(q[14]), .B(DB[107]), .Z(n37250) );
  XNOR U35560 ( .A(q[13]), .B(DB[106]), .Z(n36556) );
  IV U35561 ( .A(n36570), .Z(n37248) );
  XOR U35562 ( .A(n37251), .B(n37252), .Z(n36570) );
  XNOR U35563 ( .A(n36566), .B(n36568), .Z(n37252) );
  XNOR U35564 ( .A(q[9]), .B(DB[102]), .Z(n36568) );
  XNOR U35565 ( .A(q[12]), .B(DB[105]), .Z(n36566) );
  IV U35566 ( .A(n36565), .Z(n37251) );
  XNOR U35567 ( .A(n36563), .B(n37253), .Z(n36565) );
  XNOR U35568 ( .A(q[11]), .B(DB[104]), .Z(n37253) );
  XNOR U35569 ( .A(q[10]), .B(DB[103]), .Z(n36563) );
  IV U35570 ( .A(n36578), .Z(n37246) );
  XOR U35571 ( .A(n37254), .B(n37255), .Z(n36578) );
  XNOR U35572 ( .A(n36595), .B(n36576), .Z(n37255) );
  XNOR U35573 ( .A(q[1]), .B(DB[94]), .Z(n36576) );
  XOR U35574 ( .A(n37256), .B(n36584), .Z(n36595) );
  XNOR U35575 ( .A(q[8]), .B(DB[101]), .Z(n36584) );
  IV U35576 ( .A(n36583), .Z(n37256) );
  XNOR U35577 ( .A(n36581), .B(n37257), .Z(n36583) );
  XNOR U35578 ( .A(q[7]), .B(DB[100]), .Z(n37257) );
  XNOR U35579 ( .A(q[6]), .B(DB[99]), .Z(n36581) );
  IV U35580 ( .A(n36594), .Z(n37254) );
  XOR U35581 ( .A(n37258), .B(n37259), .Z(n36594) );
  XNOR U35582 ( .A(n36590), .B(n36592), .Z(n37259) );
  XNOR U35583 ( .A(q[2]), .B(DB[95]), .Z(n36592) );
  XNOR U35584 ( .A(q[5]), .B(DB[98]), .Z(n36590) );
  IV U35585 ( .A(n36589), .Z(n37258) );
  XNOR U35586 ( .A(n36587), .B(n37260), .Z(n36589) );
  XNOR U35587 ( .A(q[4]), .B(DB[97]), .Z(n37260) );
  XNOR U35588 ( .A(q[3]), .B(DB[96]), .Z(n36587) );
  XOR U35589 ( .A(n37261), .B(n36356), .Z(n36207) );
  XOR U35590 ( .A(n37262), .B(n36332), .Z(n36356) );
  XOR U35591 ( .A(n37263), .B(n36324), .Z(n36332) );
  XOR U35592 ( .A(n37264), .B(n36313), .Z(n36324) );
  XNOR U35593 ( .A(q[30]), .B(DB[154]), .Z(n36313) );
  IV U35594 ( .A(n36312), .Z(n37264) );
  XNOR U35595 ( .A(n36310), .B(n37265), .Z(n36312) );
  XNOR U35596 ( .A(q[29]), .B(DB[153]), .Z(n37265) );
  XNOR U35597 ( .A(q[28]), .B(DB[152]), .Z(n36310) );
  IV U35598 ( .A(n36323), .Z(n37263) );
  XOR U35599 ( .A(n37266), .B(n37267), .Z(n36323) );
  XNOR U35600 ( .A(n36319), .B(n36321), .Z(n37267) );
  XNOR U35601 ( .A(q[24]), .B(DB[148]), .Z(n36321) );
  XNOR U35602 ( .A(q[27]), .B(DB[151]), .Z(n36319) );
  IV U35603 ( .A(n36318), .Z(n37266) );
  XNOR U35604 ( .A(n36316), .B(n37268), .Z(n36318) );
  XNOR U35605 ( .A(q[26]), .B(DB[150]), .Z(n37268) );
  XNOR U35606 ( .A(q[25]), .B(DB[149]), .Z(n36316) );
  IV U35607 ( .A(n36331), .Z(n37262) );
  XOR U35608 ( .A(n37269), .B(n37270), .Z(n36331) );
  XNOR U35609 ( .A(n36348), .B(n36329), .Z(n37270) );
  XNOR U35610 ( .A(q[16]), .B(DB[140]), .Z(n36329) );
  XOR U35611 ( .A(n37271), .B(n36337), .Z(n36348) );
  XNOR U35612 ( .A(q[23]), .B(DB[147]), .Z(n36337) );
  IV U35613 ( .A(n36336), .Z(n37271) );
  XNOR U35614 ( .A(n36334), .B(n37272), .Z(n36336) );
  XNOR U35615 ( .A(q[22]), .B(DB[146]), .Z(n37272) );
  XNOR U35616 ( .A(q[21]), .B(DB[145]), .Z(n36334) );
  IV U35617 ( .A(n36347), .Z(n37269) );
  XOR U35618 ( .A(n37273), .B(n37274), .Z(n36347) );
  XNOR U35619 ( .A(n36343), .B(n36345), .Z(n37274) );
  XNOR U35620 ( .A(q[17]), .B(DB[141]), .Z(n36345) );
  XNOR U35621 ( .A(q[20]), .B(DB[144]), .Z(n36343) );
  IV U35622 ( .A(n36342), .Z(n37273) );
  XNOR U35623 ( .A(n36340), .B(n37275), .Z(n36342) );
  XNOR U35624 ( .A(q[19]), .B(DB[143]), .Z(n37275) );
  XNOR U35625 ( .A(q[18]), .B(DB[142]), .Z(n36340) );
  IV U35626 ( .A(n36355), .Z(n37261) );
  XOR U35627 ( .A(n37276), .B(n37277), .Z(n36355) );
  XNOR U35628 ( .A(n36382), .B(n36353), .Z(n37277) );
  XNOR U35629 ( .A(q[0]), .B(DB[124]), .Z(n36353) );
  XOR U35630 ( .A(n37278), .B(n36374), .Z(n36382) );
  XOR U35631 ( .A(n37279), .B(n36362), .Z(n36374) );
  XNOR U35632 ( .A(q[15]), .B(DB[139]), .Z(n36362) );
  IV U35633 ( .A(n36361), .Z(n37279) );
  XNOR U35634 ( .A(n36359), .B(n37280), .Z(n36361) );
  XNOR U35635 ( .A(q[14]), .B(DB[138]), .Z(n37280) );
  XNOR U35636 ( .A(q[13]), .B(DB[137]), .Z(n36359) );
  IV U35637 ( .A(n36373), .Z(n37278) );
  XOR U35638 ( .A(n37281), .B(n37282), .Z(n36373) );
  XNOR U35639 ( .A(n36369), .B(n36371), .Z(n37282) );
  XNOR U35640 ( .A(q[9]), .B(DB[133]), .Z(n36371) );
  XNOR U35641 ( .A(q[12]), .B(DB[136]), .Z(n36369) );
  IV U35642 ( .A(n36368), .Z(n37281) );
  XNOR U35643 ( .A(n36366), .B(n37283), .Z(n36368) );
  XNOR U35644 ( .A(q[11]), .B(DB[135]), .Z(n37283) );
  XNOR U35645 ( .A(q[10]), .B(DB[134]), .Z(n36366) );
  IV U35646 ( .A(n36381), .Z(n37276) );
  XOR U35647 ( .A(n37284), .B(n37285), .Z(n36381) );
  XNOR U35648 ( .A(n36398), .B(n36379), .Z(n37285) );
  XNOR U35649 ( .A(q[1]), .B(DB[125]), .Z(n36379) );
  XOR U35650 ( .A(n37286), .B(n36387), .Z(n36398) );
  XNOR U35651 ( .A(q[8]), .B(DB[132]), .Z(n36387) );
  IV U35652 ( .A(n36386), .Z(n37286) );
  XNOR U35653 ( .A(n36384), .B(n37287), .Z(n36386) );
  XNOR U35654 ( .A(q[7]), .B(DB[131]), .Z(n37287) );
  XNOR U35655 ( .A(q[6]), .B(DB[130]), .Z(n36384) );
  IV U35656 ( .A(n36397), .Z(n37284) );
  XOR U35657 ( .A(n37288), .B(n37289), .Z(n36397) );
  XNOR U35658 ( .A(n36393), .B(n36395), .Z(n37289) );
  XNOR U35659 ( .A(q[2]), .B(DB[126]), .Z(n36395) );
  XNOR U35660 ( .A(q[5]), .B(DB[129]), .Z(n36393) );
  IV U35661 ( .A(n36392), .Z(n37288) );
  XNOR U35662 ( .A(n36390), .B(n37290), .Z(n36392) );
  XNOR U35663 ( .A(q[4]), .B(DB[128]), .Z(n37290) );
  XNOR U35664 ( .A(q[3]), .B(DB[127]), .Z(n36390) );
  XOR U35665 ( .A(n37291), .B(n36159), .Z(n36010) );
  XOR U35666 ( .A(n37292), .B(n36135), .Z(n36159) );
  XOR U35667 ( .A(n37293), .B(n36127), .Z(n36135) );
  XOR U35668 ( .A(n37294), .B(n36116), .Z(n36127) );
  XNOR U35669 ( .A(q[30]), .B(DB[185]), .Z(n36116) );
  IV U35670 ( .A(n36115), .Z(n37294) );
  XNOR U35671 ( .A(n36113), .B(n37295), .Z(n36115) );
  XNOR U35672 ( .A(q[29]), .B(DB[184]), .Z(n37295) );
  XNOR U35673 ( .A(q[28]), .B(DB[183]), .Z(n36113) );
  IV U35674 ( .A(n36126), .Z(n37293) );
  XOR U35675 ( .A(n37296), .B(n37297), .Z(n36126) );
  XNOR U35676 ( .A(n36122), .B(n36124), .Z(n37297) );
  XNOR U35677 ( .A(q[24]), .B(DB[179]), .Z(n36124) );
  XNOR U35678 ( .A(q[27]), .B(DB[182]), .Z(n36122) );
  IV U35679 ( .A(n36121), .Z(n37296) );
  XNOR U35680 ( .A(n36119), .B(n37298), .Z(n36121) );
  XNOR U35681 ( .A(q[26]), .B(DB[181]), .Z(n37298) );
  XNOR U35682 ( .A(q[25]), .B(DB[180]), .Z(n36119) );
  IV U35683 ( .A(n36134), .Z(n37292) );
  XOR U35684 ( .A(n37299), .B(n37300), .Z(n36134) );
  XNOR U35685 ( .A(n36151), .B(n36132), .Z(n37300) );
  XNOR U35686 ( .A(q[16]), .B(DB[171]), .Z(n36132) );
  XOR U35687 ( .A(n37301), .B(n36140), .Z(n36151) );
  XNOR U35688 ( .A(q[23]), .B(DB[178]), .Z(n36140) );
  IV U35689 ( .A(n36139), .Z(n37301) );
  XNOR U35690 ( .A(n36137), .B(n37302), .Z(n36139) );
  XNOR U35691 ( .A(q[22]), .B(DB[177]), .Z(n37302) );
  XNOR U35692 ( .A(q[21]), .B(DB[176]), .Z(n36137) );
  IV U35693 ( .A(n36150), .Z(n37299) );
  XOR U35694 ( .A(n37303), .B(n37304), .Z(n36150) );
  XNOR U35695 ( .A(n36146), .B(n36148), .Z(n37304) );
  XNOR U35696 ( .A(q[17]), .B(DB[172]), .Z(n36148) );
  XNOR U35697 ( .A(q[20]), .B(DB[175]), .Z(n36146) );
  IV U35698 ( .A(n36145), .Z(n37303) );
  XNOR U35699 ( .A(n36143), .B(n37305), .Z(n36145) );
  XNOR U35700 ( .A(q[19]), .B(DB[174]), .Z(n37305) );
  XNOR U35701 ( .A(q[18]), .B(DB[173]), .Z(n36143) );
  IV U35702 ( .A(n36158), .Z(n37291) );
  XOR U35703 ( .A(n37306), .B(n37307), .Z(n36158) );
  XNOR U35704 ( .A(n36185), .B(n36156), .Z(n37307) );
  XNOR U35705 ( .A(q[0]), .B(DB[155]), .Z(n36156) );
  XOR U35706 ( .A(n37308), .B(n36177), .Z(n36185) );
  XOR U35707 ( .A(n37309), .B(n36165), .Z(n36177) );
  XNOR U35708 ( .A(q[15]), .B(DB[170]), .Z(n36165) );
  IV U35709 ( .A(n36164), .Z(n37309) );
  XNOR U35710 ( .A(n36162), .B(n37310), .Z(n36164) );
  XNOR U35711 ( .A(q[14]), .B(DB[169]), .Z(n37310) );
  XNOR U35712 ( .A(q[13]), .B(DB[168]), .Z(n36162) );
  IV U35713 ( .A(n36176), .Z(n37308) );
  XOR U35714 ( .A(n37311), .B(n37312), .Z(n36176) );
  XNOR U35715 ( .A(n36172), .B(n36174), .Z(n37312) );
  XNOR U35716 ( .A(q[9]), .B(DB[164]), .Z(n36174) );
  XNOR U35717 ( .A(q[12]), .B(DB[167]), .Z(n36172) );
  IV U35718 ( .A(n36171), .Z(n37311) );
  XNOR U35719 ( .A(n36169), .B(n37313), .Z(n36171) );
  XNOR U35720 ( .A(q[11]), .B(DB[166]), .Z(n37313) );
  XNOR U35721 ( .A(q[10]), .B(DB[165]), .Z(n36169) );
  IV U35722 ( .A(n36184), .Z(n37306) );
  XOR U35723 ( .A(n37314), .B(n37315), .Z(n36184) );
  XNOR U35724 ( .A(n36201), .B(n36182), .Z(n37315) );
  XNOR U35725 ( .A(q[1]), .B(DB[156]), .Z(n36182) );
  XOR U35726 ( .A(n37316), .B(n36190), .Z(n36201) );
  XNOR U35727 ( .A(q[8]), .B(DB[163]), .Z(n36190) );
  IV U35728 ( .A(n36189), .Z(n37316) );
  XNOR U35729 ( .A(n36187), .B(n37317), .Z(n36189) );
  XNOR U35730 ( .A(q[7]), .B(DB[162]), .Z(n37317) );
  XNOR U35731 ( .A(q[6]), .B(DB[161]), .Z(n36187) );
  IV U35732 ( .A(n36200), .Z(n37314) );
  XOR U35733 ( .A(n37318), .B(n37319), .Z(n36200) );
  XNOR U35734 ( .A(n36196), .B(n36198), .Z(n37319) );
  XNOR U35735 ( .A(q[2]), .B(DB[157]), .Z(n36198) );
  XNOR U35736 ( .A(q[5]), .B(DB[160]), .Z(n36196) );
  IV U35737 ( .A(n36195), .Z(n37318) );
  XNOR U35738 ( .A(n36193), .B(n37320), .Z(n36195) );
  XNOR U35739 ( .A(q[4]), .B(DB[159]), .Z(n37320) );
  XNOR U35740 ( .A(q[3]), .B(DB[158]), .Z(n36193) );
  XOR U35741 ( .A(n37321), .B(n35962), .Z(n35813) );
  XOR U35742 ( .A(n37322), .B(n35938), .Z(n35962) );
  XOR U35743 ( .A(n37323), .B(n35930), .Z(n35938) );
  XOR U35744 ( .A(n37324), .B(n35919), .Z(n35930) );
  XNOR U35745 ( .A(q[30]), .B(DB[216]), .Z(n35919) );
  IV U35746 ( .A(n35918), .Z(n37324) );
  XNOR U35747 ( .A(n35916), .B(n37325), .Z(n35918) );
  XNOR U35748 ( .A(q[29]), .B(DB[215]), .Z(n37325) );
  XNOR U35749 ( .A(q[28]), .B(DB[214]), .Z(n35916) );
  IV U35750 ( .A(n35929), .Z(n37323) );
  XOR U35751 ( .A(n37326), .B(n37327), .Z(n35929) );
  XNOR U35752 ( .A(n35925), .B(n35927), .Z(n37327) );
  XNOR U35753 ( .A(q[24]), .B(DB[210]), .Z(n35927) );
  XNOR U35754 ( .A(q[27]), .B(DB[213]), .Z(n35925) );
  IV U35755 ( .A(n35924), .Z(n37326) );
  XNOR U35756 ( .A(n35922), .B(n37328), .Z(n35924) );
  XNOR U35757 ( .A(q[26]), .B(DB[212]), .Z(n37328) );
  XNOR U35758 ( .A(q[25]), .B(DB[211]), .Z(n35922) );
  IV U35759 ( .A(n35937), .Z(n37322) );
  XOR U35760 ( .A(n37329), .B(n37330), .Z(n35937) );
  XNOR U35761 ( .A(n35954), .B(n35935), .Z(n37330) );
  XNOR U35762 ( .A(q[16]), .B(DB[202]), .Z(n35935) );
  XOR U35763 ( .A(n37331), .B(n35943), .Z(n35954) );
  XNOR U35764 ( .A(q[23]), .B(DB[209]), .Z(n35943) );
  IV U35765 ( .A(n35942), .Z(n37331) );
  XNOR U35766 ( .A(n35940), .B(n37332), .Z(n35942) );
  XNOR U35767 ( .A(q[22]), .B(DB[208]), .Z(n37332) );
  XNOR U35768 ( .A(q[21]), .B(DB[207]), .Z(n35940) );
  IV U35769 ( .A(n35953), .Z(n37329) );
  XOR U35770 ( .A(n37333), .B(n37334), .Z(n35953) );
  XNOR U35771 ( .A(n35949), .B(n35951), .Z(n37334) );
  XNOR U35772 ( .A(q[17]), .B(DB[203]), .Z(n35951) );
  XNOR U35773 ( .A(q[20]), .B(DB[206]), .Z(n35949) );
  IV U35774 ( .A(n35948), .Z(n37333) );
  XNOR U35775 ( .A(n35946), .B(n37335), .Z(n35948) );
  XNOR U35776 ( .A(q[19]), .B(DB[205]), .Z(n37335) );
  XNOR U35777 ( .A(q[18]), .B(DB[204]), .Z(n35946) );
  IV U35778 ( .A(n35961), .Z(n37321) );
  XOR U35779 ( .A(n37336), .B(n37337), .Z(n35961) );
  XNOR U35780 ( .A(n35988), .B(n35959), .Z(n37337) );
  XNOR U35781 ( .A(q[0]), .B(DB[186]), .Z(n35959) );
  XOR U35782 ( .A(n37338), .B(n35980), .Z(n35988) );
  XOR U35783 ( .A(n37339), .B(n35968), .Z(n35980) );
  XNOR U35784 ( .A(q[15]), .B(DB[201]), .Z(n35968) );
  IV U35785 ( .A(n35967), .Z(n37339) );
  XNOR U35786 ( .A(n35965), .B(n37340), .Z(n35967) );
  XNOR U35787 ( .A(q[14]), .B(DB[200]), .Z(n37340) );
  XNOR U35788 ( .A(q[13]), .B(DB[199]), .Z(n35965) );
  IV U35789 ( .A(n35979), .Z(n37338) );
  XOR U35790 ( .A(n37341), .B(n37342), .Z(n35979) );
  XNOR U35791 ( .A(n35975), .B(n35977), .Z(n37342) );
  XNOR U35792 ( .A(q[9]), .B(DB[195]), .Z(n35977) );
  XNOR U35793 ( .A(q[12]), .B(DB[198]), .Z(n35975) );
  IV U35794 ( .A(n35974), .Z(n37341) );
  XNOR U35795 ( .A(n35972), .B(n37343), .Z(n35974) );
  XNOR U35796 ( .A(q[11]), .B(DB[197]), .Z(n37343) );
  XNOR U35797 ( .A(q[10]), .B(DB[196]), .Z(n35972) );
  IV U35798 ( .A(n35987), .Z(n37336) );
  XOR U35799 ( .A(n37344), .B(n37345), .Z(n35987) );
  XNOR U35800 ( .A(n36004), .B(n35985), .Z(n37345) );
  XNOR U35801 ( .A(q[1]), .B(DB[187]), .Z(n35985) );
  XOR U35802 ( .A(n37346), .B(n35993), .Z(n36004) );
  XNOR U35803 ( .A(q[8]), .B(DB[194]), .Z(n35993) );
  IV U35804 ( .A(n35992), .Z(n37346) );
  XNOR U35805 ( .A(n35990), .B(n37347), .Z(n35992) );
  XNOR U35806 ( .A(q[7]), .B(DB[193]), .Z(n37347) );
  XNOR U35807 ( .A(q[6]), .B(DB[192]), .Z(n35990) );
  IV U35808 ( .A(n36003), .Z(n37344) );
  XOR U35809 ( .A(n37348), .B(n37349), .Z(n36003) );
  XNOR U35810 ( .A(n35999), .B(n36001), .Z(n37349) );
  XNOR U35811 ( .A(q[2]), .B(DB[188]), .Z(n36001) );
  XNOR U35812 ( .A(q[5]), .B(DB[191]), .Z(n35999) );
  IV U35813 ( .A(n35998), .Z(n37348) );
  XNOR U35814 ( .A(n35996), .B(n37350), .Z(n35998) );
  XNOR U35815 ( .A(q[4]), .B(DB[190]), .Z(n37350) );
  XNOR U35816 ( .A(q[3]), .B(DB[189]), .Z(n35996) );
  XOR U35817 ( .A(n37351), .B(n35765), .Z(n35616) );
  XOR U35818 ( .A(n37352), .B(n35741), .Z(n35765) );
  XOR U35819 ( .A(n37353), .B(n35733), .Z(n35741) );
  XOR U35820 ( .A(n37354), .B(n35722), .Z(n35733) );
  XNOR U35821 ( .A(q[30]), .B(DB[247]), .Z(n35722) );
  IV U35822 ( .A(n35721), .Z(n37354) );
  XNOR U35823 ( .A(n35719), .B(n37355), .Z(n35721) );
  XNOR U35824 ( .A(q[29]), .B(DB[246]), .Z(n37355) );
  XNOR U35825 ( .A(q[28]), .B(DB[245]), .Z(n35719) );
  IV U35826 ( .A(n35732), .Z(n37353) );
  XOR U35827 ( .A(n37356), .B(n37357), .Z(n35732) );
  XNOR U35828 ( .A(n35728), .B(n35730), .Z(n37357) );
  XNOR U35829 ( .A(q[24]), .B(DB[241]), .Z(n35730) );
  XNOR U35830 ( .A(q[27]), .B(DB[244]), .Z(n35728) );
  IV U35831 ( .A(n35727), .Z(n37356) );
  XNOR U35832 ( .A(n35725), .B(n37358), .Z(n35727) );
  XNOR U35833 ( .A(q[26]), .B(DB[243]), .Z(n37358) );
  XNOR U35834 ( .A(q[25]), .B(DB[242]), .Z(n35725) );
  IV U35835 ( .A(n35740), .Z(n37352) );
  XOR U35836 ( .A(n37359), .B(n37360), .Z(n35740) );
  XNOR U35837 ( .A(n35757), .B(n35738), .Z(n37360) );
  XNOR U35838 ( .A(q[16]), .B(DB[233]), .Z(n35738) );
  XOR U35839 ( .A(n37361), .B(n35746), .Z(n35757) );
  XNOR U35840 ( .A(q[23]), .B(DB[240]), .Z(n35746) );
  IV U35841 ( .A(n35745), .Z(n37361) );
  XNOR U35842 ( .A(n35743), .B(n37362), .Z(n35745) );
  XNOR U35843 ( .A(q[22]), .B(DB[239]), .Z(n37362) );
  XNOR U35844 ( .A(q[21]), .B(DB[238]), .Z(n35743) );
  IV U35845 ( .A(n35756), .Z(n37359) );
  XOR U35846 ( .A(n37363), .B(n37364), .Z(n35756) );
  XNOR U35847 ( .A(n35752), .B(n35754), .Z(n37364) );
  XNOR U35848 ( .A(q[17]), .B(DB[234]), .Z(n35754) );
  XNOR U35849 ( .A(q[20]), .B(DB[237]), .Z(n35752) );
  IV U35850 ( .A(n35751), .Z(n37363) );
  XNOR U35851 ( .A(n35749), .B(n37365), .Z(n35751) );
  XNOR U35852 ( .A(q[19]), .B(DB[236]), .Z(n37365) );
  XNOR U35853 ( .A(q[18]), .B(DB[235]), .Z(n35749) );
  IV U35854 ( .A(n35764), .Z(n37351) );
  XOR U35855 ( .A(n37366), .B(n37367), .Z(n35764) );
  XNOR U35856 ( .A(n35791), .B(n35762), .Z(n37367) );
  XNOR U35857 ( .A(q[0]), .B(DB[217]), .Z(n35762) );
  XOR U35858 ( .A(n37368), .B(n35783), .Z(n35791) );
  XOR U35859 ( .A(n37369), .B(n35771), .Z(n35783) );
  XNOR U35860 ( .A(q[15]), .B(DB[232]), .Z(n35771) );
  IV U35861 ( .A(n35770), .Z(n37369) );
  XNOR U35862 ( .A(n35768), .B(n37370), .Z(n35770) );
  XNOR U35863 ( .A(q[14]), .B(DB[231]), .Z(n37370) );
  XNOR U35864 ( .A(q[13]), .B(DB[230]), .Z(n35768) );
  IV U35865 ( .A(n35782), .Z(n37368) );
  XOR U35866 ( .A(n37371), .B(n37372), .Z(n35782) );
  XNOR U35867 ( .A(n35778), .B(n35780), .Z(n37372) );
  XNOR U35868 ( .A(q[9]), .B(DB[226]), .Z(n35780) );
  XNOR U35869 ( .A(q[12]), .B(DB[229]), .Z(n35778) );
  IV U35870 ( .A(n35777), .Z(n37371) );
  XNOR U35871 ( .A(n35775), .B(n37373), .Z(n35777) );
  XNOR U35872 ( .A(q[11]), .B(DB[228]), .Z(n37373) );
  XNOR U35873 ( .A(q[10]), .B(DB[227]), .Z(n35775) );
  IV U35874 ( .A(n35790), .Z(n37366) );
  XOR U35875 ( .A(n37374), .B(n37375), .Z(n35790) );
  XNOR U35876 ( .A(n35807), .B(n35788), .Z(n37375) );
  XNOR U35877 ( .A(q[1]), .B(DB[218]), .Z(n35788) );
  XOR U35878 ( .A(n37376), .B(n35796), .Z(n35807) );
  XNOR U35879 ( .A(q[8]), .B(DB[225]), .Z(n35796) );
  IV U35880 ( .A(n35795), .Z(n37376) );
  XNOR U35881 ( .A(n35793), .B(n37377), .Z(n35795) );
  XNOR U35882 ( .A(q[7]), .B(DB[224]), .Z(n37377) );
  XNOR U35883 ( .A(q[6]), .B(DB[223]), .Z(n35793) );
  IV U35884 ( .A(n35806), .Z(n37374) );
  XOR U35885 ( .A(n37378), .B(n37379), .Z(n35806) );
  XNOR U35886 ( .A(n35802), .B(n35804), .Z(n37379) );
  XNOR U35887 ( .A(q[2]), .B(DB[219]), .Z(n35804) );
  XNOR U35888 ( .A(q[5]), .B(DB[222]), .Z(n35802) );
  IV U35889 ( .A(n35801), .Z(n37378) );
  XNOR U35890 ( .A(n35799), .B(n37380), .Z(n35801) );
  XNOR U35891 ( .A(q[4]), .B(DB[221]), .Z(n37380) );
  XNOR U35892 ( .A(q[3]), .B(DB[220]), .Z(n35799) );
  XOR U35893 ( .A(n37381), .B(n35568), .Z(n35419) );
  XOR U35894 ( .A(n37382), .B(n35544), .Z(n35568) );
  XOR U35895 ( .A(n37383), .B(n35536), .Z(n35544) );
  XOR U35896 ( .A(n37384), .B(n35525), .Z(n35536) );
  XNOR U35897 ( .A(q[30]), .B(DB[278]), .Z(n35525) );
  IV U35898 ( .A(n35524), .Z(n37384) );
  XNOR U35899 ( .A(n35522), .B(n37385), .Z(n35524) );
  XNOR U35900 ( .A(q[29]), .B(DB[277]), .Z(n37385) );
  XNOR U35901 ( .A(q[28]), .B(DB[276]), .Z(n35522) );
  IV U35902 ( .A(n35535), .Z(n37383) );
  XOR U35903 ( .A(n37386), .B(n37387), .Z(n35535) );
  XNOR U35904 ( .A(n35531), .B(n35533), .Z(n37387) );
  XNOR U35905 ( .A(q[24]), .B(DB[272]), .Z(n35533) );
  XNOR U35906 ( .A(q[27]), .B(DB[275]), .Z(n35531) );
  IV U35907 ( .A(n35530), .Z(n37386) );
  XNOR U35908 ( .A(n35528), .B(n37388), .Z(n35530) );
  XNOR U35909 ( .A(q[26]), .B(DB[274]), .Z(n37388) );
  XNOR U35910 ( .A(q[25]), .B(DB[273]), .Z(n35528) );
  IV U35911 ( .A(n35543), .Z(n37382) );
  XOR U35912 ( .A(n37389), .B(n37390), .Z(n35543) );
  XNOR U35913 ( .A(n35560), .B(n35541), .Z(n37390) );
  XNOR U35914 ( .A(q[16]), .B(DB[264]), .Z(n35541) );
  XOR U35915 ( .A(n37391), .B(n35549), .Z(n35560) );
  XNOR U35916 ( .A(q[23]), .B(DB[271]), .Z(n35549) );
  IV U35917 ( .A(n35548), .Z(n37391) );
  XNOR U35918 ( .A(n35546), .B(n37392), .Z(n35548) );
  XNOR U35919 ( .A(q[22]), .B(DB[270]), .Z(n37392) );
  XNOR U35920 ( .A(q[21]), .B(DB[269]), .Z(n35546) );
  IV U35921 ( .A(n35559), .Z(n37389) );
  XOR U35922 ( .A(n37393), .B(n37394), .Z(n35559) );
  XNOR U35923 ( .A(n35555), .B(n35557), .Z(n37394) );
  XNOR U35924 ( .A(q[17]), .B(DB[265]), .Z(n35557) );
  XNOR U35925 ( .A(q[20]), .B(DB[268]), .Z(n35555) );
  IV U35926 ( .A(n35554), .Z(n37393) );
  XNOR U35927 ( .A(n35552), .B(n37395), .Z(n35554) );
  XNOR U35928 ( .A(q[19]), .B(DB[267]), .Z(n37395) );
  XNOR U35929 ( .A(q[18]), .B(DB[266]), .Z(n35552) );
  IV U35930 ( .A(n35567), .Z(n37381) );
  XOR U35931 ( .A(n37396), .B(n37397), .Z(n35567) );
  XNOR U35932 ( .A(n35594), .B(n35565), .Z(n37397) );
  XNOR U35933 ( .A(q[0]), .B(DB[248]), .Z(n35565) );
  XOR U35934 ( .A(n37398), .B(n35586), .Z(n35594) );
  XOR U35935 ( .A(n37399), .B(n35574), .Z(n35586) );
  XNOR U35936 ( .A(q[15]), .B(DB[263]), .Z(n35574) );
  IV U35937 ( .A(n35573), .Z(n37399) );
  XNOR U35938 ( .A(n35571), .B(n37400), .Z(n35573) );
  XNOR U35939 ( .A(q[14]), .B(DB[262]), .Z(n37400) );
  XNOR U35940 ( .A(q[13]), .B(DB[261]), .Z(n35571) );
  IV U35941 ( .A(n35585), .Z(n37398) );
  XOR U35942 ( .A(n37401), .B(n37402), .Z(n35585) );
  XNOR U35943 ( .A(n35581), .B(n35583), .Z(n37402) );
  XNOR U35944 ( .A(q[9]), .B(DB[257]), .Z(n35583) );
  XNOR U35945 ( .A(q[12]), .B(DB[260]), .Z(n35581) );
  IV U35946 ( .A(n35580), .Z(n37401) );
  XNOR U35947 ( .A(n35578), .B(n37403), .Z(n35580) );
  XNOR U35948 ( .A(q[11]), .B(DB[259]), .Z(n37403) );
  XNOR U35949 ( .A(q[10]), .B(DB[258]), .Z(n35578) );
  IV U35950 ( .A(n35593), .Z(n37396) );
  XOR U35951 ( .A(n37404), .B(n37405), .Z(n35593) );
  XNOR U35952 ( .A(n35610), .B(n35591), .Z(n37405) );
  XNOR U35953 ( .A(q[1]), .B(DB[249]), .Z(n35591) );
  XOR U35954 ( .A(n37406), .B(n35599), .Z(n35610) );
  XNOR U35955 ( .A(q[8]), .B(DB[256]), .Z(n35599) );
  IV U35956 ( .A(n35598), .Z(n37406) );
  XNOR U35957 ( .A(n35596), .B(n37407), .Z(n35598) );
  XNOR U35958 ( .A(q[7]), .B(DB[255]), .Z(n37407) );
  XNOR U35959 ( .A(q[6]), .B(DB[254]), .Z(n35596) );
  IV U35960 ( .A(n35609), .Z(n37404) );
  XOR U35961 ( .A(n37408), .B(n37409), .Z(n35609) );
  XNOR U35962 ( .A(n35605), .B(n35607), .Z(n37409) );
  XNOR U35963 ( .A(q[2]), .B(DB[250]), .Z(n35607) );
  XNOR U35964 ( .A(q[5]), .B(DB[253]), .Z(n35605) );
  IV U35965 ( .A(n35604), .Z(n37408) );
  XNOR U35966 ( .A(n35602), .B(n37410), .Z(n35604) );
  XNOR U35967 ( .A(q[4]), .B(DB[252]), .Z(n37410) );
  XNOR U35968 ( .A(q[3]), .B(DB[251]), .Z(n35602) );
  XOR U35969 ( .A(n37411), .B(n35371), .Z(n35222) );
  XOR U35970 ( .A(n37412), .B(n35347), .Z(n35371) );
  XOR U35971 ( .A(n37413), .B(n35339), .Z(n35347) );
  XOR U35972 ( .A(n37414), .B(n35328), .Z(n35339) );
  XNOR U35973 ( .A(q[30]), .B(DB[309]), .Z(n35328) );
  IV U35974 ( .A(n35327), .Z(n37414) );
  XNOR U35975 ( .A(n35325), .B(n37415), .Z(n35327) );
  XNOR U35976 ( .A(q[29]), .B(DB[308]), .Z(n37415) );
  XNOR U35977 ( .A(q[28]), .B(DB[307]), .Z(n35325) );
  IV U35978 ( .A(n35338), .Z(n37413) );
  XOR U35979 ( .A(n37416), .B(n37417), .Z(n35338) );
  XNOR U35980 ( .A(n35334), .B(n35336), .Z(n37417) );
  XNOR U35981 ( .A(q[24]), .B(DB[303]), .Z(n35336) );
  XNOR U35982 ( .A(q[27]), .B(DB[306]), .Z(n35334) );
  IV U35983 ( .A(n35333), .Z(n37416) );
  XNOR U35984 ( .A(n35331), .B(n37418), .Z(n35333) );
  XNOR U35985 ( .A(q[26]), .B(DB[305]), .Z(n37418) );
  XNOR U35986 ( .A(q[25]), .B(DB[304]), .Z(n35331) );
  IV U35987 ( .A(n35346), .Z(n37412) );
  XOR U35988 ( .A(n37419), .B(n37420), .Z(n35346) );
  XNOR U35989 ( .A(n35363), .B(n35344), .Z(n37420) );
  XNOR U35990 ( .A(q[16]), .B(DB[295]), .Z(n35344) );
  XOR U35991 ( .A(n37421), .B(n35352), .Z(n35363) );
  XNOR U35992 ( .A(q[23]), .B(DB[302]), .Z(n35352) );
  IV U35993 ( .A(n35351), .Z(n37421) );
  XNOR U35994 ( .A(n35349), .B(n37422), .Z(n35351) );
  XNOR U35995 ( .A(q[22]), .B(DB[301]), .Z(n37422) );
  XNOR U35996 ( .A(q[21]), .B(DB[300]), .Z(n35349) );
  IV U35997 ( .A(n35362), .Z(n37419) );
  XOR U35998 ( .A(n37423), .B(n37424), .Z(n35362) );
  XNOR U35999 ( .A(n35358), .B(n35360), .Z(n37424) );
  XNOR U36000 ( .A(q[17]), .B(DB[296]), .Z(n35360) );
  XNOR U36001 ( .A(q[20]), .B(DB[299]), .Z(n35358) );
  IV U36002 ( .A(n35357), .Z(n37423) );
  XNOR U36003 ( .A(n35355), .B(n37425), .Z(n35357) );
  XNOR U36004 ( .A(q[19]), .B(DB[298]), .Z(n37425) );
  XNOR U36005 ( .A(q[18]), .B(DB[297]), .Z(n35355) );
  IV U36006 ( .A(n35370), .Z(n37411) );
  XOR U36007 ( .A(n37426), .B(n37427), .Z(n35370) );
  XNOR U36008 ( .A(n35397), .B(n35368), .Z(n37427) );
  XNOR U36009 ( .A(q[0]), .B(DB[279]), .Z(n35368) );
  XOR U36010 ( .A(n37428), .B(n35389), .Z(n35397) );
  XOR U36011 ( .A(n37429), .B(n35377), .Z(n35389) );
  XNOR U36012 ( .A(q[15]), .B(DB[294]), .Z(n35377) );
  IV U36013 ( .A(n35376), .Z(n37429) );
  XNOR U36014 ( .A(n35374), .B(n37430), .Z(n35376) );
  XNOR U36015 ( .A(q[14]), .B(DB[293]), .Z(n37430) );
  XNOR U36016 ( .A(q[13]), .B(DB[292]), .Z(n35374) );
  IV U36017 ( .A(n35388), .Z(n37428) );
  XOR U36018 ( .A(n37431), .B(n37432), .Z(n35388) );
  XNOR U36019 ( .A(n35384), .B(n35386), .Z(n37432) );
  XNOR U36020 ( .A(q[9]), .B(DB[288]), .Z(n35386) );
  XNOR U36021 ( .A(q[12]), .B(DB[291]), .Z(n35384) );
  IV U36022 ( .A(n35383), .Z(n37431) );
  XNOR U36023 ( .A(n35381), .B(n37433), .Z(n35383) );
  XNOR U36024 ( .A(q[11]), .B(DB[290]), .Z(n37433) );
  XNOR U36025 ( .A(q[10]), .B(DB[289]), .Z(n35381) );
  IV U36026 ( .A(n35396), .Z(n37426) );
  XOR U36027 ( .A(n37434), .B(n37435), .Z(n35396) );
  XNOR U36028 ( .A(n35413), .B(n35394), .Z(n37435) );
  XNOR U36029 ( .A(q[1]), .B(DB[280]), .Z(n35394) );
  XOR U36030 ( .A(n37436), .B(n35402), .Z(n35413) );
  XNOR U36031 ( .A(q[8]), .B(DB[287]), .Z(n35402) );
  IV U36032 ( .A(n35401), .Z(n37436) );
  XNOR U36033 ( .A(n35399), .B(n37437), .Z(n35401) );
  XNOR U36034 ( .A(q[7]), .B(DB[286]), .Z(n37437) );
  XNOR U36035 ( .A(q[6]), .B(DB[285]), .Z(n35399) );
  IV U36036 ( .A(n35412), .Z(n37434) );
  XOR U36037 ( .A(n37438), .B(n37439), .Z(n35412) );
  XNOR U36038 ( .A(n35408), .B(n35410), .Z(n37439) );
  XNOR U36039 ( .A(q[2]), .B(DB[281]), .Z(n35410) );
  XNOR U36040 ( .A(q[5]), .B(DB[284]), .Z(n35408) );
  IV U36041 ( .A(n35407), .Z(n37438) );
  XNOR U36042 ( .A(n35405), .B(n37440), .Z(n35407) );
  XNOR U36043 ( .A(q[4]), .B(DB[283]), .Z(n37440) );
  XNOR U36044 ( .A(q[3]), .B(DB[282]), .Z(n35405) );
  XOR U36045 ( .A(n37441), .B(n35174), .Z(n35025) );
  XOR U36046 ( .A(n37442), .B(n35150), .Z(n35174) );
  XOR U36047 ( .A(n37443), .B(n35142), .Z(n35150) );
  XOR U36048 ( .A(n37444), .B(n35131), .Z(n35142) );
  XNOR U36049 ( .A(q[30]), .B(DB[340]), .Z(n35131) );
  IV U36050 ( .A(n35130), .Z(n37444) );
  XNOR U36051 ( .A(n35128), .B(n37445), .Z(n35130) );
  XNOR U36052 ( .A(q[29]), .B(DB[339]), .Z(n37445) );
  XNOR U36053 ( .A(q[28]), .B(DB[338]), .Z(n35128) );
  IV U36054 ( .A(n35141), .Z(n37443) );
  XOR U36055 ( .A(n37446), .B(n37447), .Z(n35141) );
  XNOR U36056 ( .A(n35137), .B(n35139), .Z(n37447) );
  XNOR U36057 ( .A(q[24]), .B(DB[334]), .Z(n35139) );
  XNOR U36058 ( .A(q[27]), .B(DB[337]), .Z(n35137) );
  IV U36059 ( .A(n35136), .Z(n37446) );
  XNOR U36060 ( .A(n35134), .B(n37448), .Z(n35136) );
  XNOR U36061 ( .A(q[26]), .B(DB[336]), .Z(n37448) );
  XNOR U36062 ( .A(q[25]), .B(DB[335]), .Z(n35134) );
  IV U36063 ( .A(n35149), .Z(n37442) );
  XOR U36064 ( .A(n37449), .B(n37450), .Z(n35149) );
  XNOR U36065 ( .A(n35166), .B(n35147), .Z(n37450) );
  XNOR U36066 ( .A(q[16]), .B(DB[326]), .Z(n35147) );
  XOR U36067 ( .A(n37451), .B(n35155), .Z(n35166) );
  XNOR U36068 ( .A(q[23]), .B(DB[333]), .Z(n35155) );
  IV U36069 ( .A(n35154), .Z(n37451) );
  XNOR U36070 ( .A(n35152), .B(n37452), .Z(n35154) );
  XNOR U36071 ( .A(q[22]), .B(DB[332]), .Z(n37452) );
  XNOR U36072 ( .A(q[21]), .B(DB[331]), .Z(n35152) );
  IV U36073 ( .A(n35165), .Z(n37449) );
  XOR U36074 ( .A(n37453), .B(n37454), .Z(n35165) );
  XNOR U36075 ( .A(n35161), .B(n35163), .Z(n37454) );
  XNOR U36076 ( .A(q[17]), .B(DB[327]), .Z(n35163) );
  XNOR U36077 ( .A(q[20]), .B(DB[330]), .Z(n35161) );
  IV U36078 ( .A(n35160), .Z(n37453) );
  XNOR U36079 ( .A(n35158), .B(n37455), .Z(n35160) );
  XNOR U36080 ( .A(q[19]), .B(DB[329]), .Z(n37455) );
  XNOR U36081 ( .A(q[18]), .B(DB[328]), .Z(n35158) );
  IV U36082 ( .A(n35173), .Z(n37441) );
  XOR U36083 ( .A(n37456), .B(n37457), .Z(n35173) );
  XNOR U36084 ( .A(n35200), .B(n35171), .Z(n37457) );
  XNOR U36085 ( .A(q[0]), .B(DB[310]), .Z(n35171) );
  XOR U36086 ( .A(n37458), .B(n35192), .Z(n35200) );
  XOR U36087 ( .A(n37459), .B(n35180), .Z(n35192) );
  XNOR U36088 ( .A(q[15]), .B(DB[325]), .Z(n35180) );
  IV U36089 ( .A(n35179), .Z(n37459) );
  XNOR U36090 ( .A(n35177), .B(n37460), .Z(n35179) );
  XNOR U36091 ( .A(q[14]), .B(DB[324]), .Z(n37460) );
  XNOR U36092 ( .A(q[13]), .B(DB[323]), .Z(n35177) );
  IV U36093 ( .A(n35191), .Z(n37458) );
  XOR U36094 ( .A(n37461), .B(n37462), .Z(n35191) );
  XNOR U36095 ( .A(n35187), .B(n35189), .Z(n37462) );
  XNOR U36096 ( .A(q[9]), .B(DB[319]), .Z(n35189) );
  XNOR U36097 ( .A(q[12]), .B(DB[322]), .Z(n35187) );
  IV U36098 ( .A(n35186), .Z(n37461) );
  XNOR U36099 ( .A(n35184), .B(n37463), .Z(n35186) );
  XNOR U36100 ( .A(q[11]), .B(DB[321]), .Z(n37463) );
  XNOR U36101 ( .A(q[10]), .B(DB[320]), .Z(n35184) );
  IV U36102 ( .A(n35199), .Z(n37456) );
  XOR U36103 ( .A(n37464), .B(n37465), .Z(n35199) );
  XNOR U36104 ( .A(n35216), .B(n35197), .Z(n37465) );
  XNOR U36105 ( .A(q[1]), .B(DB[311]), .Z(n35197) );
  XOR U36106 ( .A(n37466), .B(n35205), .Z(n35216) );
  XNOR U36107 ( .A(q[8]), .B(DB[318]), .Z(n35205) );
  IV U36108 ( .A(n35204), .Z(n37466) );
  XNOR U36109 ( .A(n35202), .B(n37467), .Z(n35204) );
  XNOR U36110 ( .A(q[7]), .B(DB[317]), .Z(n37467) );
  XNOR U36111 ( .A(q[6]), .B(DB[316]), .Z(n35202) );
  IV U36112 ( .A(n35215), .Z(n37464) );
  XOR U36113 ( .A(n37468), .B(n37469), .Z(n35215) );
  XNOR U36114 ( .A(n35211), .B(n35213), .Z(n37469) );
  XNOR U36115 ( .A(q[2]), .B(DB[312]), .Z(n35213) );
  XNOR U36116 ( .A(q[5]), .B(DB[315]), .Z(n35211) );
  IV U36117 ( .A(n35210), .Z(n37468) );
  XNOR U36118 ( .A(n35208), .B(n37470), .Z(n35210) );
  XNOR U36119 ( .A(q[4]), .B(DB[314]), .Z(n37470) );
  XNOR U36120 ( .A(q[3]), .B(DB[313]), .Z(n35208) );
  XOR U36121 ( .A(n37471), .B(n34977), .Z(n34828) );
  XOR U36122 ( .A(n37472), .B(n34953), .Z(n34977) );
  XOR U36123 ( .A(n37473), .B(n34945), .Z(n34953) );
  XOR U36124 ( .A(n37474), .B(n34934), .Z(n34945) );
  XNOR U36125 ( .A(q[30]), .B(DB[371]), .Z(n34934) );
  IV U36126 ( .A(n34933), .Z(n37474) );
  XNOR U36127 ( .A(n34931), .B(n37475), .Z(n34933) );
  XNOR U36128 ( .A(q[29]), .B(DB[370]), .Z(n37475) );
  XNOR U36129 ( .A(q[28]), .B(DB[369]), .Z(n34931) );
  IV U36130 ( .A(n34944), .Z(n37473) );
  XOR U36131 ( .A(n37476), .B(n37477), .Z(n34944) );
  XNOR U36132 ( .A(n34940), .B(n34942), .Z(n37477) );
  XNOR U36133 ( .A(q[24]), .B(DB[365]), .Z(n34942) );
  XNOR U36134 ( .A(q[27]), .B(DB[368]), .Z(n34940) );
  IV U36135 ( .A(n34939), .Z(n37476) );
  XNOR U36136 ( .A(n34937), .B(n37478), .Z(n34939) );
  XNOR U36137 ( .A(q[26]), .B(DB[367]), .Z(n37478) );
  XNOR U36138 ( .A(q[25]), .B(DB[366]), .Z(n34937) );
  IV U36139 ( .A(n34952), .Z(n37472) );
  XOR U36140 ( .A(n37479), .B(n37480), .Z(n34952) );
  XNOR U36141 ( .A(n34969), .B(n34950), .Z(n37480) );
  XNOR U36142 ( .A(q[16]), .B(DB[357]), .Z(n34950) );
  XOR U36143 ( .A(n37481), .B(n34958), .Z(n34969) );
  XNOR U36144 ( .A(q[23]), .B(DB[364]), .Z(n34958) );
  IV U36145 ( .A(n34957), .Z(n37481) );
  XNOR U36146 ( .A(n34955), .B(n37482), .Z(n34957) );
  XNOR U36147 ( .A(q[22]), .B(DB[363]), .Z(n37482) );
  XNOR U36148 ( .A(q[21]), .B(DB[362]), .Z(n34955) );
  IV U36149 ( .A(n34968), .Z(n37479) );
  XOR U36150 ( .A(n37483), .B(n37484), .Z(n34968) );
  XNOR U36151 ( .A(n34964), .B(n34966), .Z(n37484) );
  XNOR U36152 ( .A(q[17]), .B(DB[358]), .Z(n34966) );
  XNOR U36153 ( .A(q[20]), .B(DB[361]), .Z(n34964) );
  IV U36154 ( .A(n34963), .Z(n37483) );
  XNOR U36155 ( .A(n34961), .B(n37485), .Z(n34963) );
  XNOR U36156 ( .A(q[19]), .B(DB[360]), .Z(n37485) );
  XNOR U36157 ( .A(q[18]), .B(DB[359]), .Z(n34961) );
  IV U36158 ( .A(n34976), .Z(n37471) );
  XOR U36159 ( .A(n37486), .B(n37487), .Z(n34976) );
  XNOR U36160 ( .A(n35003), .B(n34974), .Z(n37487) );
  XNOR U36161 ( .A(q[0]), .B(DB[341]), .Z(n34974) );
  XOR U36162 ( .A(n37488), .B(n34995), .Z(n35003) );
  XOR U36163 ( .A(n37489), .B(n34983), .Z(n34995) );
  XNOR U36164 ( .A(q[15]), .B(DB[356]), .Z(n34983) );
  IV U36165 ( .A(n34982), .Z(n37489) );
  XNOR U36166 ( .A(n34980), .B(n37490), .Z(n34982) );
  XNOR U36167 ( .A(q[14]), .B(DB[355]), .Z(n37490) );
  XNOR U36168 ( .A(q[13]), .B(DB[354]), .Z(n34980) );
  IV U36169 ( .A(n34994), .Z(n37488) );
  XOR U36170 ( .A(n37491), .B(n37492), .Z(n34994) );
  XNOR U36171 ( .A(n34990), .B(n34992), .Z(n37492) );
  XNOR U36172 ( .A(q[9]), .B(DB[350]), .Z(n34992) );
  XNOR U36173 ( .A(q[12]), .B(DB[353]), .Z(n34990) );
  IV U36174 ( .A(n34989), .Z(n37491) );
  XNOR U36175 ( .A(n34987), .B(n37493), .Z(n34989) );
  XNOR U36176 ( .A(q[11]), .B(DB[352]), .Z(n37493) );
  XNOR U36177 ( .A(q[10]), .B(DB[351]), .Z(n34987) );
  IV U36178 ( .A(n35002), .Z(n37486) );
  XOR U36179 ( .A(n37494), .B(n37495), .Z(n35002) );
  XNOR U36180 ( .A(n35019), .B(n35000), .Z(n37495) );
  XNOR U36181 ( .A(q[1]), .B(DB[342]), .Z(n35000) );
  XOR U36182 ( .A(n37496), .B(n35008), .Z(n35019) );
  XNOR U36183 ( .A(q[8]), .B(DB[349]), .Z(n35008) );
  IV U36184 ( .A(n35007), .Z(n37496) );
  XNOR U36185 ( .A(n35005), .B(n37497), .Z(n35007) );
  XNOR U36186 ( .A(q[7]), .B(DB[348]), .Z(n37497) );
  XNOR U36187 ( .A(q[6]), .B(DB[347]), .Z(n35005) );
  IV U36188 ( .A(n35018), .Z(n37494) );
  XOR U36189 ( .A(n37498), .B(n37499), .Z(n35018) );
  XNOR U36190 ( .A(n35014), .B(n35016), .Z(n37499) );
  XNOR U36191 ( .A(q[2]), .B(DB[343]), .Z(n35016) );
  XNOR U36192 ( .A(q[5]), .B(DB[346]), .Z(n35014) );
  IV U36193 ( .A(n35013), .Z(n37498) );
  XNOR U36194 ( .A(n35011), .B(n37500), .Z(n35013) );
  XNOR U36195 ( .A(q[4]), .B(DB[345]), .Z(n37500) );
  XNOR U36196 ( .A(q[3]), .B(DB[344]), .Z(n35011) );
  XOR U36197 ( .A(n37501), .B(n34780), .Z(n34631) );
  XOR U36198 ( .A(n37502), .B(n34756), .Z(n34780) );
  XOR U36199 ( .A(n37503), .B(n34748), .Z(n34756) );
  XOR U36200 ( .A(n37504), .B(n34737), .Z(n34748) );
  XNOR U36201 ( .A(q[30]), .B(DB[402]), .Z(n34737) );
  IV U36202 ( .A(n34736), .Z(n37504) );
  XNOR U36203 ( .A(n34734), .B(n37505), .Z(n34736) );
  XNOR U36204 ( .A(q[29]), .B(DB[401]), .Z(n37505) );
  XNOR U36205 ( .A(q[28]), .B(DB[400]), .Z(n34734) );
  IV U36206 ( .A(n34747), .Z(n37503) );
  XOR U36207 ( .A(n37506), .B(n37507), .Z(n34747) );
  XNOR U36208 ( .A(n34743), .B(n34745), .Z(n37507) );
  XNOR U36209 ( .A(q[24]), .B(DB[396]), .Z(n34745) );
  XNOR U36210 ( .A(q[27]), .B(DB[399]), .Z(n34743) );
  IV U36211 ( .A(n34742), .Z(n37506) );
  XNOR U36212 ( .A(n34740), .B(n37508), .Z(n34742) );
  XNOR U36213 ( .A(q[26]), .B(DB[398]), .Z(n37508) );
  XNOR U36214 ( .A(q[25]), .B(DB[397]), .Z(n34740) );
  IV U36215 ( .A(n34755), .Z(n37502) );
  XOR U36216 ( .A(n37509), .B(n37510), .Z(n34755) );
  XNOR U36217 ( .A(n34772), .B(n34753), .Z(n37510) );
  XNOR U36218 ( .A(q[16]), .B(DB[388]), .Z(n34753) );
  XOR U36219 ( .A(n37511), .B(n34761), .Z(n34772) );
  XNOR U36220 ( .A(q[23]), .B(DB[395]), .Z(n34761) );
  IV U36221 ( .A(n34760), .Z(n37511) );
  XNOR U36222 ( .A(n34758), .B(n37512), .Z(n34760) );
  XNOR U36223 ( .A(q[22]), .B(DB[394]), .Z(n37512) );
  XNOR U36224 ( .A(q[21]), .B(DB[393]), .Z(n34758) );
  IV U36225 ( .A(n34771), .Z(n37509) );
  XOR U36226 ( .A(n37513), .B(n37514), .Z(n34771) );
  XNOR U36227 ( .A(n34767), .B(n34769), .Z(n37514) );
  XNOR U36228 ( .A(q[17]), .B(DB[389]), .Z(n34769) );
  XNOR U36229 ( .A(q[20]), .B(DB[392]), .Z(n34767) );
  IV U36230 ( .A(n34766), .Z(n37513) );
  XNOR U36231 ( .A(n34764), .B(n37515), .Z(n34766) );
  XNOR U36232 ( .A(q[19]), .B(DB[391]), .Z(n37515) );
  XNOR U36233 ( .A(q[18]), .B(DB[390]), .Z(n34764) );
  IV U36234 ( .A(n34779), .Z(n37501) );
  XOR U36235 ( .A(n37516), .B(n37517), .Z(n34779) );
  XNOR U36236 ( .A(n34806), .B(n34777), .Z(n37517) );
  XNOR U36237 ( .A(q[0]), .B(DB[372]), .Z(n34777) );
  XOR U36238 ( .A(n37518), .B(n34798), .Z(n34806) );
  XOR U36239 ( .A(n37519), .B(n34786), .Z(n34798) );
  XNOR U36240 ( .A(q[15]), .B(DB[387]), .Z(n34786) );
  IV U36241 ( .A(n34785), .Z(n37519) );
  XNOR U36242 ( .A(n34783), .B(n37520), .Z(n34785) );
  XNOR U36243 ( .A(q[14]), .B(DB[386]), .Z(n37520) );
  XNOR U36244 ( .A(q[13]), .B(DB[385]), .Z(n34783) );
  IV U36245 ( .A(n34797), .Z(n37518) );
  XOR U36246 ( .A(n37521), .B(n37522), .Z(n34797) );
  XNOR U36247 ( .A(n34793), .B(n34795), .Z(n37522) );
  XNOR U36248 ( .A(q[9]), .B(DB[381]), .Z(n34795) );
  XNOR U36249 ( .A(q[12]), .B(DB[384]), .Z(n34793) );
  IV U36250 ( .A(n34792), .Z(n37521) );
  XNOR U36251 ( .A(n34790), .B(n37523), .Z(n34792) );
  XNOR U36252 ( .A(q[11]), .B(DB[383]), .Z(n37523) );
  XNOR U36253 ( .A(q[10]), .B(DB[382]), .Z(n34790) );
  IV U36254 ( .A(n34805), .Z(n37516) );
  XOR U36255 ( .A(n37524), .B(n37525), .Z(n34805) );
  XNOR U36256 ( .A(n34822), .B(n34803), .Z(n37525) );
  XNOR U36257 ( .A(q[1]), .B(DB[373]), .Z(n34803) );
  XOR U36258 ( .A(n37526), .B(n34811), .Z(n34822) );
  XNOR U36259 ( .A(q[8]), .B(DB[380]), .Z(n34811) );
  IV U36260 ( .A(n34810), .Z(n37526) );
  XNOR U36261 ( .A(n34808), .B(n37527), .Z(n34810) );
  XNOR U36262 ( .A(q[7]), .B(DB[379]), .Z(n37527) );
  XNOR U36263 ( .A(q[6]), .B(DB[378]), .Z(n34808) );
  IV U36264 ( .A(n34821), .Z(n37524) );
  XOR U36265 ( .A(n37528), .B(n37529), .Z(n34821) );
  XNOR U36266 ( .A(n34817), .B(n34819), .Z(n37529) );
  XNOR U36267 ( .A(q[2]), .B(DB[374]), .Z(n34819) );
  XNOR U36268 ( .A(q[5]), .B(DB[377]), .Z(n34817) );
  IV U36269 ( .A(n34816), .Z(n37528) );
  XNOR U36270 ( .A(n34814), .B(n37530), .Z(n34816) );
  XNOR U36271 ( .A(q[4]), .B(DB[376]), .Z(n37530) );
  XNOR U36272 ( .A(q[3]), .B(DB[375]), .Z(n34814) );
  XOR U36273 ( .A(n37531), .B(n34583), .Z(n34434) );
  XOR U36274 ( .A(n37532), .B(n34559), .Z(n34583) );
  XOR U36275 ( .A(n37533), .B(n34551), .Z(n34559) );
  XOR U36276 ( .A(n37534), .B(n34540), .Z(n34551) );
  XNOR U36277 ( .A(q[30]), .B(DB[433]), .Z(n34540) );
  IV U36278 ( .A(n34539), .Z(n37534) );
  XNOR U36279 ( .A(n34537), .B(n37535), .Z(n34539) );
  XNOR U36280 ( .A(q[29]), .B(DB[432]), .Z(n37535) );
  XNOR U36281 ( .A(q[28]), .B(DB[431]), .Z(n34537) );
  IV U36282 ( .A(n34550), .Z(n37533) );
  XOR U36283 ( .A(n37536), .B(n37537), .Z(n34550) );
  XNOR U36284 ( .A(n34546), .B(n34548), .Z(n37537) );
  XNOR U36285 ( .A(q[24]), .B(DB[427]), .Z(n34548) );
  XNOR U36286 ( .A(q[27]), .B(DB[430]), .Z(n34546) );
  IV U36287 ( .A(n34545), .Z(n37536) );
  XNOR U36288 ( .A(n34543), .B(n37538), .Z(n34545) );
  XNOR U36289 ( .A(q[26]), .B(DB[429]), .Z(n37538) );
  XNOR U36290 ( .A(q[25]), .B(DB[428]), .Z(n34543) );
  IV U36291 ( .A(n34558), .Z(n37532) );
  XOR U36292 ( .A(n37539), .B(n37540), .Z(n34558) );
  XNOR U36293 ( .A(n34575), .B(n34556), .Z(n37540) );
  XNOR U36294 ( .A(q[16]), .B(DB[419]), .Z(n34556) );
  XOR U36295 ( .A(n37541), .B(n34564), .Z(n34575) );
  XNOR U36296 ( .A(q[23]), .B(DB[426]), .Z(n34564) );
  IV U36297 ( .A(n34563), .Z(n37541) );
  XNOR U36298 ( .A(n34561), .B(n37542), .Z(n34563) );
  XNOR U36299 ( .A(q[22]), .B(DB[425]), .Z(n37542) );
  XNOR U36300 ( .A(q[21]), .B(DB[424]), .Z(n34561) );
  IV U36301 ( .A(n34574), .Z(n37539) );
  XOR U36302 ( .A(n37543), .B(n37544), .Z(n34574) );
  XNOR U36303 ( .A(n34570), .B(n34572), .Z(n37544) );
  XNOR U36304 ( .A(q[17]), .B(DB[420]), .Z(n34572) );
  XNOR U36305 ( .A(q[20]), .B(DB[423]), .Z(n34570) );
  IV U36306 ( .A(n34569), .Z(n37543) );
  XNOR U36307 ( .A(n34567), .B(n37545), .Z(n34569) );
  XNOR U36308 ( .A(q[19]), .B(DB[422]), .Z(n37545) );
  XNOR U36309 ( .A(q[18]), .B(DB[421]), .Z(n34567) );
  IV U36310 ( .A(n34582), .Z(n37531) );
  XOR U36311 ( .A(n37546), .B(n37547), .Z(n34582) );
  XNOR U36312 ( .A(n34609), .B(n34580), .Z(n37547) );
  XNOR U36313 ( .A(q[0]), .B(DB[403]), .Z(n34580) );
  XOR U36314 ( .A(n37548), .B(n34601), .Z(n34609) );
  XOR U36315 ( .A(n37549), .B(n34589), .Z(n34601) );
  XNOR U36316 ( .A(q[15]), .B(DB[418]), .Z(n34589) );
  IV U36317 ( .A(n34588), .Z(n37549) );
  XNOR U36318 ( .A(n34586), .B(n37550), .Z(n34588) );
  XNOR U36319 ( .A(q[14]), .B(DB[417]), .Z(n37550) );
  XNOR U36320 ( .A(q[13]), .B(DB[416]), .Z(n34586) );
  IV U36321 ( .A(n34600), .Z(n37548) );
  XOR U36322 ( .A(n37551), .B(n37552), .Z(n34600) );
  XNOR U36323 ( .A(n34596), .B(n34598), .Z(n37552) );
  XNOR U36324 ( .A(q[9]), .B(DB[412]), .Z(n34598) );
  XNOR U36325 ( .A(q[12]), .B(DB[415]), .Z(n34596) );
  IV U36326 ( .A(n34595), .Z(n37551) );
  XNOR U36327 ( .A(n34593), .B(n37553), .Z(n34595) );
  XNOR U36328 ( .A(q[11]), .B(DB[414]), .Z(n37553) );
  XNOR U36329 ( .A(q[10]), .B(DB[413]), .Z(n34593) );
  IV U36330 ( .A(n34608), .Z(n37546) );
  XOR U36331 ( .A(n37554), .B(n37555), .Z(n34608) );
  XNOR U36332 ( .A(n34625), .B(n34606), .Z(n37555) );
  XNOR U36333 ( .A(q[1]), .B(DB[404]), .Z(n34606) );
  XOR U36334 ( .A(n37556), .B(n34614), .Z(n34625) );
  XNOR U36335 ( .A(q[8]), .B(DB[411]), .Z(n34614) );
  IV U36336 ( .A(n34613), .Z(n37556) );
  XNOR U36337 ( .A(n34611), .B(n37557), .Z(n34613) );
  XNOR U36338 ( .A(q[7]), .B(DB[410]), .Z(n37557) );
  XNOR U36339 ( .A(q[6]), .B(DB[409]), .Z(n34611) );
  IV U36340 ( .A(n34624), .Z(n37554) );
  XOR U36341 ( .A(n37558), .B(n37559), .Z(n34624) );
  XNOR U36342 ( .A(n34620), .B(n34622), .Z(n37559) );
  XNOR U36343 ( .A(q[2]), .B(DB[405]), .Z(n34622) );
  XNOR U36344 ( .A(q[5]), .B(DB[408]), .Z(n34620) );
  IV U36345 ( .A(n34619), .Z(n37558) );
  XNOR U36346 ( .A(n34617), .B(n37560), .Z(n34619) );
  XNOR U36347 ( .A(q[4]), .B(DB[407]), .Z(n37560) );
  XNOR U36348 ( .A(q[3]), .B(DB[406]), .Z(n34617) );
  XOR U36349 ( .A(n37561), .B(n34386), .Z(n34237) );
  XOR U36350 ( .A(n37562), .B(n34362), .Z(n34386) );
  XOR U36351 ( .A(n37563), .B(n34354), .Z(n34362) );
  XOR U36352 ( .A(n37564), .B(n34343), .Z(n34354) );
  XNOR U36353 ( .A(q[30]), .B(DB[464]), .Z(n34343) );
  IV U36354 ( .A(n34342), .Z(n37564) );
  XNOR U36355 ( .A(n34340), .B(n37565), .Z(n34342) );
  XNOR U36356 ( .A(q[29]), .B(DB[463]), .Z(n37565) );
  XNOR U36357 ( .A(q[28]), .B(DB[462]), .Z(n34340) );
  IV U36358 ( .A(n34353), .Z(n37563) );
  XOR U36359 ( .A(n37566), .B(n37567), .Z(n34353) );
  XNOR U36360 ( .A(n34349), .B(n34351), .Z(n37567) );
  XNOR U36361 ( .A(q[24]), .B(DB[458]), .Z(n34351) );
  XNOR U36362 ( .A(q[27]), .B(DB[461]), .Z(n34349) );
  IV U36363 ( .A(n34348), .Z(n37566) );
  XNOR U36364 ( .A(n34346), .B(n37568), .Z(n34348) );
  XNOR U36365 ( .A(q[26]), .B(DB[460]), .Z(n37568) );
  XNOR U36366 ( .A(q[25]), .B(DB[459]), .Z(n34346) );
  IV U36367 ( .A(n34361), .Z(n37562) );
  XOR U36368 ( .A(n37569), .B(n37570), .Z(n34361) );
  XNOR U36369 ( .A(n34378), .B(n34359), .Z(n37570) );
  XNOR U36370 ( .A(q[16]), .B(DB[450]), .Z(n34359) );
  XOR U36371 ( .A(n37571), .B(n34367), .Z(n34378) );
  XNOR U36372 ( .A(q[23]), .B(DB[457]), .Z(n34367) );
  IV U36373 ( .A(n34366), .Z(n37571) );
  XNOR U36374 ( .A(n34364), .B(n37572), .Z(n34366) );
  XNOR U36375 ( .A(q[22]), .B(DB[456]), .Z(n37572) );
  XNOR U36376 ( .A(q[21]), .B(DB[455]), .Z(n34364) );
  IV U36377 ( .A(n34377), .Z(n37569) );
  XOR U36378 ( .A(n37573), .B(n37574), .Z(n34377) );
  XNOR U36379 ( .A(n34373), .B(n34375), .Z(n37574) );
  XNOR U36380 ( .A(q[17]), .B(DB[451]), .Z(n34375) );
  XNOR U36381 ( .A(q[20]), .B(DB[454]), .Z(n34373) );
  IV U36382 ( .A(n34372), .Z(n37573) );
  XNOR U36383 ( .A(n34370), .B(n37575), .Z(n34372) );
  XNOR U36384 ( .A(q[19]), .B(DB[453]), .Z(n37575) );
  XNOR U36385 ( .A(q[18]), .B(DB[452]), .Z(n34370) );
  IV U36386 ( .A(n34385), .Z(n37561) );
  XOR U36387 ( .A(n37576), .B(n37577), .Z(n34385) );
  XNOR U36388 ( .A(n34412), .B(n34383), .Z(n37577) );
  XNOR U36389 ( .A(q[0]), .B(DB[434]), .Z(n34383) );
  XOR U36390 ( .A(n37578), .B(n34404), .Z(n34412) );
  XOR U36391 ( .A(n37579), .B(n34392), .Z(n34404) );
  XNOR U36392 ( .A(q[15]), .B(DB[449]), .Z(n34392) );
  IV U36393 ( .A(n34391), .Z(n37579) );
  XNOR U36394 ( .A(n34389), .B(n37580), .Z(n34391) );
  XNOR U36395 ( .A(q[14]), .B(DB[448]), .Z(n37580) );
  XNOR U36396 ( .A(q[13]), .B(DB[447]), .Z(n34389) );
  IV U36397 ( .A(n34403), .Z(n37578) );
  XOR U36398 ( .A(n37581), .B(n37582), .Z(n34403) );
  XNOR U36399 ( .A(n34399), .B(n34401), .Z(n37582) );
  XNOR U36400 ( .A(q[9]), .B(DB[443]), .Z(n34401) );
  XNOR U36401 ( .A(q[12]), .B(DB[446]), .Z(n34399) );
  IV U36402 ( .A(n34398), .Z(n37581) );
  XNOR U36403 ( .A(n34396), .B(n37583), .Z(n34398) );
  XNOR U36404 ( .A(q[11]), .B(DB[445]), .Z(n37583) );
  XNOR U36405 ( .A(q[10]), .B(DB[444]), .Z(n34396) );
  IV U36406 ( .A(n34411), .Z(n37576) );
  XOR U36407 ( .A(n37584), .B(n37585), .Z(n34411) );
  XNOR U36408 ( .A(n34428), .B(n34409), .Z(n37585) );
  XNOR U36409 ( .A(q[1]), .B(DB[435]), .Z(n34409) );
  XOR U36410 ( .A(n37586), .B(n34417), .Z(n34428) );
  XNOR U36411 ( .A(q[8]), .B(DB[442]), .Z(n34417) );
  IV U36412 ( .A(n34416), .Z(n37586) );
  XNOR U36413 ( .A(n34414), .B(n37587), .Z(n34416) );
  XNOR U36414 ( .A(q[7]), .B(DB[441]), .Z(n37587) );
  XNOR U36415 ( .A(q[6]), .B(DB[440]), .Z(n34414) );
  IV U36416 ( .A(n34427), .Z(n37584) );
  XOR U36417 ( .A(n37588), .B(n37589), .Z(n34427) );
  XNOR U36418 ( .A(n34423), .B(n34425), .Z(n37589) );
  XNOR U36419 ( .A(q[2]), .B(DB[436]), .Z(n34425) );
  XNOR U36420 ( .A(q[5]), .B(DB[439]), .Z(n34423) );
  IV U36421 ( .A(n34422), .Z(n37588) );
  XNOR U36422 ( .A(n34420), .B(n37590), .Z(n34422) );
  XNOR U36423 ( .A(q[4]), .B(DB[438]), .Z(n37590) );
  XNOR U36424 ( .A(q[3]), .B(DB[437]), .Z(n34420) );
  XOR U36425 ( .A(n37591), .B(n34189), .Z(n34040) );
  XOR U36426 ( .A(n37592), .B(n34165), .Z(n34189) );
  XOR U36427 ( .A(n37593), .B(n34157), .Z(n34165) );
  XOR U36428 ( .A(n37594), .B(n34146), .Z(n34157) );
  XNOR U36429 ( .A(q[30]), .B(DB[495]), .Z(n34146) );
  IV U36430 ( .A(n34145), .Z(n37594) );
  XNOR U36431 ( .A(n34143), .B(n37595), .Z(n34145) );
  XNOR U36432 ( .A(q[29]), .B(DB[494]), .Z(n37595) );
  XNOR U36433 ( .A(q[28]), .B(DB[493]), .Z(n34143) );
  IV U36434 ( .A(n34156), .Z(n37593) );
  XOR U36435 ( .A(n37596), .B(n37597), .Z(n34156) );
  XNOR U36436 ( .A(n34152), .B(n34154), .Z(n37597) );
  XNOR U36437 ( .A(q[24]), .B(DB[489]), .Z(n34154) );
  XNOR U36438 ( .A(q[27]), .B(DB[492]), .Z(n34152) );
  IV U36439 ( .A(n34151), .Z(n37596) );
  XNOR U36440 ( .A(n34149), .B(n37598), .Z(n34151) );
  XNOR U36441 ( .A(q[26]), .B(DB[491]), .Z(n37598) );
  XNOR U36442 ( .A(q[25]), .B(DB[490]), .Z(n34149) );
  IV U36443 ( .A(n34164), .Z(n37592) );
  XOR U36444 ( .A(n37599), .B(n37600), .Z(n34164) );
  XNOR U36445 ( .A(n34181), .B(n34162), .Z(n37600) );
  XNOR U36446 ( .A(q[16]), .B(DB[481]), .Z(n34162) );
  XOR U36447 ( .A(n37601), .B(n34170), .Z(n34181) );
  XNOR U36448 ( .A(q[23]), .B(DB[488]), .Z(n34170) );
  IV U36449 ( .A(n34169), .Z(n37601) );
  XNOR U36450 ( .A(n34167), .B(n37602), .Z(n34169) );
  XNOR U36451 ( .A(q[22]), .B(DB[487]), .Z(n37602) );
  XNOR U36452 ( .A(q[21]), .B(DB[486]), .Z(n34167) );
  IV U36453 ( .A(n34180), .Z(n37599) );
  XOR U36454 ( .A(n37603), .B(n37604), .Z(n34180) );
  XNOR U36455 ( .A(n34176), .B(n34178), .Z(n37604) );
  XNOR U36456 ( .A(q[17]), .B(DB[482]), .Z(n34178) );
  XNOR U36457 ( .A(q[20]), .B(DB[485]), .Z(n34176) );
  IV U36458 ( .A(n34175), .Z(n37603) );
  XNOR U36459 ( .A(n34173), .B(n37605), .Z(n34175) );
  XNOR U36460 ( .A(q[19]), .B(DB[484]), .Z(n37605) );
  XNOR U36461 ( .A(q[18]), .B(DB[483]), .Z(n34173) );
  IV U36462 ( .A(n34188), .Z(n37591) );
  XOR U36463 ( .A(n37606), .B(n37607), .Z(n34188) );
  XNOR U36464 ( .A(n34215), .B(n34186), .Z(n37607) );
  XNOR U36465 ( .A(q[0]), .B(DB[465]), .Z(n34186) );
  XOR U36466 ( .A(n37608), .B(n34207), .Z(n34215) );
  XOR U36467 ( .A(n37609), .B(n34195), .Z(n34207) );
  XNOR U36468 ( .A(q[15]), .B(DB[480]), .Z(n34195) );
  IV U36469 ( .A(n34194), .Z(n37609) );
  XNOR U36470 ( .A(n34192), .B(n37610), .Z(n34194) );
  XNOR U36471 ( .A(q[14]), .B(DB[479]), .Z(n37610) );
  XNOR U36472 ( .A(q[13]), .B(DB[478]), .Z(n34192) );
  IV U36473 ( .A(n34206), .Z(n37608) );
  XOR U36474 ( .A(n37611), .B(n37612), .Z(n34206) );
  XNOR U36475 ( .A(n34202), .B(n34204), .Z(n37612) );
  XNOR U36476 ( .A(q[9]), .B(DB[474]), .Z(n34204) );
  XNOR U36477 ( .A(q[12]), .B(DB[477]), .Z(n34202) );
  IV U36478 ( .A(n34201), .Z(n37611) );
  XNOR U36479 ( .A(n34199), .B(n37613), .Z(n34201) );
  XNOR U36480 ( .A(q[11]), .B(DB[476]), .Z(n37613) );
  XNOR U36481 ( .A(q[10]), .B(DB[475]), .Z(n34199) );
  IV U36482 ( .A(n34214), .Z(n37606) );
  XOR U36483 ( .A(n37614), .B(n37615), .Z(n34214) );
  XNOR U36484 ( .A(n34231), .B(n34212), .Z(n37615) );
  XNOR U36485 ( .A(q[1]), .B(DB[466]), .Z(n34212) );
  XOR U36486 ( .A(n37616), .B(n34220), .Z(n34231) );
  XNOR U36487 ( .A(q[8]), .B(DB[473]), .Z(n34220) );
  IV U36488 ( .A(n34219), .Z(n37616) );
  XNOR U36489 ( .A(n34217), .B(n37617), .Z(n34219) );
  XNOR U36490 ( .A(q[7]), .B(DB[472]), .Z(n37617) );
  XNOR U36491 ( .A(q[6]), .B(DB[471]), .Z(n34217) );
  IV U36492 ( .A(n34230), .Z(n37614) );
  XOR U36493 ( .A(n37618), .B(n37619), .Z(n34230) );
  XNOR U36494 ( .A(n34226), .B(n34228), .Z(n37619) );
  XNOR U36495 ( .A(q[2]), .B(DB[467]), .Z(n34228) );
  XNOR U36496 ( .A(q[5]), .B(DB[470]), .Z(n34226) );
  IV U36497 ( .A(n34225), .Z(n37618) );
  XNOR U36498 ( .A(n34223), .B(n37620), .Z(n34225) );
  XNOR U36499 ( .A(q[4]), .B(DB[469]), .Z(n37620) );
  XNOR U36500 ( .A(q[3]), .B(DB[468]), .Z(n34223) );
  XOR U36501 ( .A(n37621), .B(n33992), .Z(n33843) );
  XOR U36502 ( .A(n37622), .B(n33968), .Z(n33992) );
  XOR U36503 ( .A(n37623), .B(n33960), .Z(n33968) );
  XOR U36504 ( .A(n37624), .B(n33949), .Z(n33960) );
  XNOR U36505 ( .A(q[30]), .B(DB[526]), .Z(n33949) );
  IV U36506 ( .A(n33948), .Z(n37624) );
  XNOR U36507 ( .A(n33946), .B(n37625), .Z(n33948) );
  XNOR U36508 ( .A(q[29]), .B(DB[525]), .Z(n37625) );
  XNOR U36509 ( .A(q[28]), .B(DB[524]), .Z(n33946) );
  IV U36510 ( .A(n33959), .Z(n37623) );
  XOR U36511 ( .A(n37626), .B(n37627), .Z(n33959) );
  XNOR U36512 ( .A(n33955), .B(n33957), .Z(n37627) );
  XNOR U36513 ( .A(q[24]), .B(DB[520]), .Z(n33957) );
  XNOR U36514 ( .A(q[27]), .B(DB[523]), .Z(n33955) );
  IV U36515 ( .A(n33954), .Z(n37626) );
  XNOR U36516 ( .A(n33952), .B(n37628), .Z(n33954) );
  XNOR U36517 ( .A(q[26]), .B(DB[522]), .Z(n37628) );
  XNOR U36518 ( .A(q[25]), .B(DB[521]), .Z(n33952) );
  IV U36519 ( .A(n33967), .Z(n37622) );
  XOR U36520 ( .A(n37629), .B(n37630), .Z(n33967) );
  XNOR U36521 ( .A(n33984), .B(n33965), .Z(n37630) );
  XNOR U36522 ( .A(q[16]), .B(DB[512]), .Z(n33965) );
  XOR U36523 ( .A(n37631), .B(n33973), .Z(n33984) );
  XNOR U36524 ( .A(q[23]), .B(DB[519]), .Z(n33973) );
  IV U36525 ( .A(n33972), .Z(n37631) );
  XNOR U36526 ( .A(n33970), .B(n37632), .Z(n33972) );
  XNOR U36527 ( .A(q[22]), .B(DB[518]), .Z(n37632) );
  XNOR U36528 ( .A(q[21]), .B(DB[517]), .Z(n33970) );
  IV U36529 ( .A(n33983), .Z(n37629) );
  XOR U36530 ( .A(n37633), .B(n37634), .Z(n33983) );
  XNOR U36531 ( .A(n33979), .B(n33981), .Z(n37634) );
  XNOR U36532 ( .A(q[17]), .B(DB[513]), .Z(n33981) );
  XNOR U36533 ( .A(q[20]), .B(DB[516]), .Z(n33979) );
  IV U36534 ( .A(n33978), .Z(n37633) );
  XNOR U36535 ( .A(n33976), .B(n37635), .Z(n33978) );
  XNOR U36536 ( .A(q[19]), .B(DB[515]), .Z(n37635) );
  XNOR U36537 ( .A(q[18]), .B(DB[514]), .Z(n33976) );
  IV U36538 ( .A(n33991), .Z(n37621) );
  XOR U36539 ( .A(n37636), .B(n37637), .Z(n33991) );
  XNOR U36540 ( .A(n34018), .B(n33989), .Z(n37637) );
  XNOR U36541 ( .A(q[0]), .B(DB[496]), .Z(n33989) );
  XOR U36542 ( .A(n37638), .B(n34010), .Z(n34018) );
  XOR U36543 ( .A(n37639), .B(n33998), .Z(n34010) );
  XNOR U36544 ( .A(q[15]), .B(DB[511]), .Z(n33998) );
  IV U36545 ( .A(n33997), .Z(n37639) );
  XNOR U36546 ( .A(n33995), .B(n37640), .Z(n33997) );
  XNOR U36547 ( .A(q[14]), .B(DB[510]), .Z(n37640) );
  XNOR U36548 ( .A(q[13]), .B(DB[509]), .Z(n33995) );
  IV U36549 ( .A(n34009), .Z(n37638) );
  XOR U36550 ( .A(n37641), .B(n37642), .Z(n34009) );
  XNOR U36551 ( .A(n34005), .B(n34007), .Z(n37642) );
  XNOR U36552 ( .A(q[9]), .B(DB[505]), .Z(n34007) );
  XNOR U36553 ( .A(q[12]), .B(DB[508]), .Z(n34005) );
  IV U36554 ( .A(n34004), .Z(n37641) );
  XNOR U36555 ( .A(n34002), .B(n37643), .Z(n34004) );
  XNOR U36556 ( .A(q[11]), .B(DB[507]), .Z(n37643) );
  XNOR U36557 ( .A(q[10]), .B(DB[506]), .Z(n34002) );
  IV U36558 ( .A(n34017), .Z(n37636) );
  XOR U36559 ( .A(n37644), .B(n37645), .Z(n34017) );
  XNOR U36560 ( .A(n34034), .B(n34015), .Z(n37645) );
  XNOR U36561 ( .A(q[1]), .B(DB[497]), .Z(n34015) );
  XOR U36562 ( .A(n37646), .B(n34023), .Z(n34034) );
  XNOR U36563 ( .A(q[8]), .B(DB[504]), .Z(n34023) );
  IV U36564 ( .A(n34022), .Z(n37646) );
  XNOR U36565 ( .A(n34020), .B(n37647), .Z(n34022) );
  XNOR U36566 ( .A(q[7]), .B(DB[503]), .Z(n37647) );
  XNOR U36567 ( .A(q[6]), .B(DB[502]), .Z(n34020) );
  IV U36568 ( .A(n34033), .Z(n37644) );
  XOR U36569 ( .A(n37648), .B(n37649), .Z(n34033) );
  XNOR U36570 ( .A(n34029), .B(n34031), .Z(n37649) );
  XNOR U36571 ( .A(q[2]), .B(DB[498]), .Z(n34031) );
  XNOR U36572 ( .A(q[5]), .B(DB[501]), .Z(n34029) );
  IV U36573 ( .A(n34028), .Z(n37648) );
  XNOR U36574 ( .A(n34026), .B(n37650), .Z(n34028) );
  XNOR U36575 ( .A(q[4]), .B(DB[500]), .Z(n37650) );
  XNOR U36576 ( .A(q[3]), .B(DB[499]), .Z(n34026) );
  XOR U36577 ( .A(n37651), .B(n33795), .Z(n33646) );
  XOR U36578 ( .A(n37652), .B(n33771), .Z(n33795) );
  XOR U36579 ( .A(n37653), .B(n33763), .Z(n33771) );
  XOR U36580 ( .A(n37654), .B(n33752), .Z(n33763) );
  XNOR U36581 ( .A(q[30]), .B(DB[557]), .Z(n33752) );
  IV U36582 ( .A(n33751), .Z(n37654) );
  XNOR U36583 ( .A(n33749), .B(n37655), .Z(n33751) );
  XNOR U36584 ( .A(q[29]), .B(DB[556]), .Z(n37655) );
  XNOR U36585 ( .A(q[28]), .B(DB[555]), .Z(n33749) );
  IV U36586 ( .A(n33762), .Z(n37653) );
  XOR U36587 ( .A(n37656), .B(n37657), .Z(n33762) );
  XNOR U36588 ( .A(n33758), .B(n33760), .Z(n37657) );
  XNOR U36589 ( .A(q[24]), .B(DB[551]), .Z(n33760) );
  XNOR U36590 ( .A(q[27]), .B(DB[554]), .Z(n33758) );
  IV U36591 ( .A(n33757), .Z(n37656) );
  XNOR U36592 ( .A(n33755), .B(n37658), .Z(n33757) );
  XNOR U36593 ( .A(q[26]), .B(DB[553]), .Z(n37658) );
  XNOR U36594 ( .A(q[25]), .B(DB[552]), .Z(n33755) );
  IV U36595 ( .A(n33770), .Z(n37652) );
  XOR U36596 ( .A(n37659), .B(n37660), .Z(n33770) );
  XNOR U36597 ( .A(n33787), .B(n33768), .Z(n37660) );
  XNOR U36598 ( .A(q[16]), .B(DB[543]), .Z(n33768) );
  XOR U36599 ( .A(n37661), .B(n33776), .Z(n33787) );
  XNOR U36600 ( .A(q[23]), .B(DB[550]), .Z(n33776) );
  IV U36601 ( .A(n33775), .Z(n37661) );
  XNOR U36602 ( .A(n33773), .B(n37662), .Z(n33775) );
  XNOR U36603 ( .A(q[22]), .B(DB[549]), .Z(n37662) );
  XNOR U36604 ( .A(q[21]), .B(DB[548]), .Z(n33773) );
  IV U36605 ( .A(n33786), .Z(n37659) );
  XOR U36606 ( .A(n37663), .B(n37664), .Z(n33786) );
  XNOR U36607 ( .A(n33782), .B(n33784), .Z(n37664) );
  XNOR U36608 ( .A(q[17]), .B(DB[544]), .Z(n33784) );
  XNOR U36609 ( .A(q[20]), .B(DB[547]), .Z(n33782) );
  IV U36610 ( .A(n33781), .Z(n37663) );
  XNOR U36611 ( .A(n33779), .B(n37665), .Z(n33781) );
  XNOR U36612 ( .A(q[19]), .B(DB[546]), .Z(n37665) );
  XNOR U36613 ( .A(q[18]), .B(DB[545]), .Z(n33779) );
  IV U36614 ( .A(n33794), .Z(n37651) );
  XOR U36615 ( .A(n37666), .B(n37667), .Z(n33794) );
  XNOR U36616 ( .A(n33821), .B(n33792), .Z(n37667) );
  XNOR U36617 ( .A(q[0]), .B(DB[527]), .Z(n33792) );
  XOR U36618 ( .A(n37668), .B(n33813), .Z(n33821) );
  XOR U36619 ( .A(n37669), .B(n33801), .Z(n33813) );
  XNOR U36620 ( .A(q[15]), .B(DB[542]), .Z(n33801) );
  IV U36621 ( .A(n33800), .Z(n37669) );
  XNOR U36622 ( .A(n33798), .B(n37670), .Z(n33800) );
  XNOR U36623 ( .A(q[14]), .B(DB[541]), .Z(n37670) );
  XNOR U36624 ( .A(q[13]), .B(DB[540]), .Z(n33798) );
  IV U36625 ( .A(n33812), .Z(n37668) );
  XOR U36626 ( .A(n37671), .B(n37672), .Z(n33812) );
  XNOR U36627 ( .A(n33808), .B(n33810), .Z(n37672) );
  XNOR U36628 ( .A(q[9]), .B(DB[536]), .Z(n33810) );
  XNOR U36629 ( .A(q[12]), .B(DB[539]), .Z(n33808) );
  IV U36630 ( .A(n33807), .Z(n37671) );
  XNOR U36631 ( .A(n33805), .B(n37673), .Z(n33807) );
  XNOR U36632 ( .A(q[11]), .B(DB[538]), .Z(n37673) );
  XNOR U36633 ( .A(q[10]), .B(DB[537]), .Z(n33805) );
  IV U36634 ( .A(n33820), .Z(n37666) );
  XOR U36635 ( .A(n37674), .B(n37675), .Z(n33820) );
  XNOR U36636 ( .A(n33837), .B(n33818), .Z(n37675) );
  XNOR U36637 ( .A(q[1]), .B(DB[528]), .Z(n33818) );
  XOR U36638 ( .A(n37676), .B(n33826), .Z(n33837) );
  XNOR U36639 ( .A(q[8]), .B(DB[535]), .Z(n33826) );
  IV U36640 ( .A(n33825), .Z(n37676) );
  XNOR U36641 ( .A(n33823), .B(n37677), .Z(n33825) );
  XNOR U36642 ( .A(q[7]), .B(DB[534]), .Z(n37677) );
  XNOR U36643 ( .A(q[6]), .B(DB[533]), .Z(n33823) );
  IV U36644 ( .A(n33836), .Z(n37674) );
  XOR U36645 ( .A(n37678), .B(n37679), .Z(n33836) );
  XNOR U36646 ( .A(n33832), .B(n33834), .Z(n37679) );
  XNOR U36647 ( .A(q[2]), .B(DB[529]), .Z(n33834) );
  XNOR U36648 ( .A(q[5]), .B(DB[532]), .Z(n33832) );
  IV U36649 ( .A(n33831), .Z(n37678) );
  XNOR U36650 ( .A(n33829), .B(n37680), .Z(n33831) );
  XNOR U36651 ( .A(q[4]), .B(DB[531]), .Z(n37680) );
  XNOR U36652 ( .A(q[3]), .B(DB[530]), .Z(n33829) );
  XOR U36653 ( .A(n37681), .B(n33598), .Z(n33449) );
  XOR U36654 ( .A(n37682), .B(n33574), .Z(n33598) );
  XOR U36655 ( .A(n37683), .B(n33566), .Z(n33574) );
  XOR U36656 ( .A(n37684), .B(n33555), .Z(n33566) );
  XNOR U36657 ( .A(q[30]), .B(DB[588]), .Z(n33555) );
  IV U36658 ( .A(n33554), .Z(n37684) );
  XNOR U36659 ( .A(n33552), .B(n37685), .Z(n33554) );
  XNOR U36660 ( .A(q[29]), .B(DB[587]), .Z(n37685) );
  XNOR U36661 ( .A(q[28]), .B(DB[586]), .Z(n33552) );
  IV U36662 ( .A(n33565), .Z(n37683) );
  XOR U36663 ( .A(n37686), .B(n37687), .Z(n33565) );
  XNOR U36664 ( .A(n33561), .B(n33563), .Z(n37687) );
  XNOR U36665 ( .A(q[24]), .B(DB[582]), .Z(n33563) );
  XNOR U36666 ( .A(q[27]), .B(DB[585]), .Z(n33561) );
  IV U36667 ( .A(n33560), .Z(n37686) );
  XNOR U36668 ( .A(n33558), .B(n37688), .Z(n33560) );
  XNOR U36669 ( .A(q[26]), .B(DB[584]), .Z(n37688) );
  XNOR U36670 ( .A(q[25]), .B(DB[583]), .Z(n33558) );
  IV U36671 ( .A(n33573), .Z(n37682) );
  XOR U36672 ( .A(n37689), .B(n37690), .Z(n33573) );
  XNOR U36673 ( .A(n33590), .B(n33571), .Z(n37690) );
  XNOR U36674 ( .A(q[16]), .B(DB[574]), .Z(n33571) );
  XOR U36675 ( .A(n37691), .B(n33579), .Z(n33590) );
  XNOR U36676 ( .A(q[23]), .B(DB[581]), .Z(n33579) );
  IV U36677 ( .A(n33578), .Z(n37691) );
  XNOR U36678 ( .A(n33576), .B(n37692), .Z(n33578) );
  XNOR U36679 ( .A(q[22]), .B(DB[580]), .Z(n37692) );
  XNOR U36680 ( .A(q[21]), .B(DB[579]), .Z(n33576) );
  IV U36681 ( .A(n33589), .Z(n37689) );
  XOR U36682 ( .A(n37693), .B(n37694), .Z(n33589) );
  XNOR U36683 ( .A(n33585), .B(n33587), .Z(n37694) );
  XNOR U36684 ( .A(q[17]), .B(DB[575]), .Z(n33587) );
  XNOR U36685 ( .A(q[20]), .B(DB[578]), .Z(n33585) );
  IV U36686 ( .A(n33584), .Z(n37693) );
  XNOR U36687 ( .A(n33582), .B(n37695), .Z(n33584) );
  XNOR U36688 ( .A(q[19]), .B(DB[577]), .Z(n37695) );
  XNOR U36689 ( .A(q[18]), .B(DB[576]), .Z(n33582) );
  IV U36690 ( .A(n33597), .Z(n37681) );
  XOR U36691 ( .A(n37696), .B(n37697), .Z(n33597) );
  XNOR U36692 ( .A(n33624), .B(n33595), .Z(n37697) );
  XNOR U36693 ( .A(q[0]), .B(DB[558]), .Z(n33595) );
  XOR U36694 ( .A(n37698), .B(n33616), .Z(n33624) );
  XOR U36695 ( .A(n37699), .B(n33604), .Z(n33616) );
  XNOR U36696 ( .A(q[15]), .B(DB[573]), .Z(n33604) );
  IV U36697 ( .A(n33603), .Z(n37699) );
  XNOR U36698 ( .A(n33601), .B(n37700), .Z(n33603) );
  XNOR U36699 ( .A(q[14]), .B(DB[572]), .Z(n37700) );
  XNOR U36700 ( .A(q[13]), .B(DB[571]), .Z(n33601) );
  IV U36701 ( .A(n33615), .Z(n37698) );
  XOR U36702 ( .A(n37701), .B(n37702), .Z(n33615) );
  XNOR U36703 ( .A(n33611), .B(n33613), .Z(n37702) );
  XNOR U36704 ( .A(q[9]), .B(DB[567]), .Z(n33613) );
  XNOR U36705 ( .A(q[12]), .B(DB[570]), .Z(n33611) );
  IV U36706 ( .A(n33610), .Z(n37701) );
  XNOR U36707 ( .A(n33608), .B(n37703), .Z(n33610) );
  XNOR U36708 ( .A(q[11]), .B(DB[569]), .Z(n37703) );
  XNOR U36709 ( .A(q[10]), .B(DB[568]), .Z(n33608) );
  IV U36710 ( .A(n33623), .Z(n37696) );
  XOR U36711 ( .A(n37704), .B(n37705), .Z(n33623) );
  XNOR U36712 ( .A(n33640), .B(n33621), .Z(n37705) );
  XNOR U36713 ( .A(q[1]), .B(DB[559]), .Z(n33621) );
  XOR U36714 ( .A(n37706), .B(n33629), .Z(n33640) );
  XNOR U36715 ( .A(q[8]), .B(DB[566]), .Z(n33629) );
  IV U36716 ( .A(n33628), .Z(n37706) );
  XNOR U36717 ( .A(n33626), .B(n37707), .Z(n33628) );
  XNOR U36718 ( .A(q[7]), .B(DB[565]), .Z(n37707) );
  XNOR U36719 ( .A(q[6]), .B(DB[564]), .Z(n33626) );
  IV U36720 ( .A(n33639), .Z(n37704) );
  XOR U36721 ( .A(n37708), .B(n37709), .Z(n33639) );
  XNOR U36722 ( .A(n33635), .B(n33637), .Z(n37709) );
  XNOR U36723 ( .A(q[2]), .B(DB[560]), .Z(n33637) );
  XNOR U36724 ( .A(q[5]), .B(DB[563]), .Z(n33635) );
  IV U36725 ( .A(n33634), .Z(n37708) );
  XNOR U36726 ( .A(n33632), .B(n37710), .Z(n33634) );
  XNOR U36727 ( .A(q[4]), .B(DB[562]), .Z(n37710) );
  XNOR U36728 ( .A(q[3]), .B(DB[561]), .Z(n33632) );
  XOR U36729 ( .A(n37711), .B(n33401), .Z(n33252) );
  XOR U36730 ( .A(n37712), .B(n33377), .Z(n33401) );
  XOR U36731 ( .A(n37713), .B(n33369), .Z(n33377) );
  XOR U36732 ( .A(n37714), .B(n33358), .Z(n33369) );
  XNOR U36733 ( .A(q[30]), .B(DB[619]), .Z(n33358) );
  IV U36734 ( .A(n33357), .Z(n37714) );
  XNOR U36735 ( .A(n33355), .B(n37715), .Z(n33357) );
  XNOR U36736 ( .A(q[29]), .B(DB[618]), .Z(n37715) );
  XNOR U36737 ( .A(q[28]), .B(DB[617]), .Z(n33355) );
  IV U36738 ( .A(n33368), .Z(n37713) );
  XOR U36739 ( .A(n37716), .B(n37717), .Z(n33368) );
  XNOR U36740 ( .A(n33364), .B(n33366), .Z(n37717) );
  XNOR U36741 ( .A(q[24]), .B(DB[613]), .Z(n33366) );
  XNOR U36742 ( .A(q[27]), .B(DB[616]), .Z(n33364) );
  IV U36743 ( .A(n33363), .Z(n37716) );
  XNOR U36744 ( .A(n33361), .B(n37718), .Z(n33363) );
  XNOR U36745 ( .A(q[26]), .B(DB[615]), .Z(n37718) );
  XNOR U36746 ( .A(q[25]), .B(DB[614]), .Z(n33361) );
  IV U36747 ( .A(n33376), .Z(n37712) );
  XOR U36748 ( .A(n37719), .B(n37720), .Z(n33376) );
  XNOR U36749 ( .A(n33393), .B(n33374), .Z(n37720) );
  XNOR U36750 ( .A(q[16]), .B(DB[605]), .Z(n33374) );
  XOR U36751 ( .A(n37721), .B(n33382), .Z(n33393) );
  XNOR U36752 ( .A(q[23]), .B(DB[612]), .Z(n33382) );
  IV U36753 ( .A(n33381), .Z(n37721) );
  XNOR U36754 ( .A(n33379), .B(n37722), .Z(n33381) );
  XNOR U36755 ( .A(q[22]), .B(DB[611]), .Z(n37722) );
  XNOR U36756 ( .A(q[21]), .B(DB[610]), .Z(n33379) );
  IV U36757 ( .A(n33392), .Z(n37719) );
  XOR U36758 ( .A(n37723), .B(n37724), .Z(n33392) );
  XNOR U36759 ( .A(n33388), .B(n33390), .Z(n37724) );
  XNOR U36760 ( .A(q[17]), .B(DB[606]), .Z(n33390) );
  XNOR U36761 ( .A(q[20]), .B(DB[609]), .Z(n33388) );
  IV U36762 ( .A(n33387), .Z(n37723) );
  XNOR U36763 ( .A(n33385), .B(n37725), .Z(n33387) );
  XNOR U36764 ( .A(q[19]), .B(DB[608]), .Z(n37725) );
  XNOR U36765 ( .A(q[18]), .B(DB[607]), .Z(n33385) );
  IV U36766 ( .A(n33400), .Z(n37711) );
  XOR U36767 ( .A(n37726), .B(n37727), .Z(n33400) );
  XNOR U36768 ( .A(n33427), .B(n33398), .Z(n37727) );
  XNOR U36769 ( .A(q[0]), .B(DB[589]), .Z(n33398) );
  XOR U36770 ( .A(n37728), .B(n33419), .Z(n33427) );
  XOR U36771 ( .A(n37729), .B(n33407), .Z(n33419) );
  XNOR U36772 ( .A(q[15]), .B(DB[604]), .Z(n33407) );
  IV U36773 ( .A(n33406), .Z(n37729) );
  XNOR U36774 ( .A(n33404), .B(n37730), .Z(n33406) );
  XNOR U36775 ( .A(q[14]), .B(DB[603]), .Z(n37730) );
  XNOR U36776 ( .A(q[13]), .B(DB[602]), .Z(n33404) );
  IV U36777 ( .A(n33418), .Z(n37728) );
  XOR U36778 ( .A(n37731), .B(n37732), .Z(n33418) );
  XNOR U36779 ( .A(n33414), .B(n33416), .Z(n37732) );
  XNOR U36780 ( .A(q[9]), .B(DB[598]), .Z(n33416) );
  XNOR U36781 ( .A(q[12]), .B(DB[601]), .Z(n33414) );
  IV U36782 ( .A(n33413), .Z(n37731) );
  XNOR U36783 ( .A(n33411), .B(n37733), .Z(n33413) );
  XNOR U36784 ( .A(q[11]), .B(DB[600]), .Z(n37733) );
  XNOR U36785 ( .A(q[10]), .B(DB[599]), .Z(n33411) );
  IV U36786 ( .A(n33426), .Z(n37726) );
  XOR U36787 ( .A(n37734), .B(n37735), .Z(n33426) );
  XNOR U36788 ( .A(n33443), .B(n33424), .Z(n37735) );
  XNOR U36789 ( .A(q[1]), .B(DB[590]), .Z(n33424) );
  XOR U36790 ( .A(n37736), .B(n33432), .Z(n33443) );
  XNOR U36791 ( .A(q[8]), .B(DB[597]), .Z(n33432) );
  IV U36792 ( .A(n33431), .Z(n37736) );
  XNOR U36793 ( .A(n33429), .B(n37737), .Z(n33431) );
  XNOR U36794 ( .A(q[7]), .B(DB[596]), .Z(n37737) );
  XNOR U36795 ( .A(q[6]), .B(DB[595]), .Z(n33429) );
  IV U36796 ( .A(n33442), .Z(n37734) );
  XOR U36797 ( .A(n37738), .B(n37739), .Z(n33442) );
  XNOR U36798 ( .A(n33438), .B(n33440), .Z(n37739) );
  XNOR U36799 ( .A(q[2]), .B(DB[591]), .Z(n33440) );
  XNOR U36800 ( .A(q[5]), .B(DB[594]), .Z(n33438) );
  IV U36801 ( .A(n33437), .Z(n37738) );
  XNOR U36802 ( .A(n33435), .B(n37740), .Z(n33437) );
  XNOR U36803 ( .A(q[4]), .B(DB[593]), .Z(n37740) );
  XNOR U36804 ( .A(q[3]), .B(DB[592]), .Z(n33435) );
  XOR U36805 ( .A(n37741), .B(n33204), .Z(n33055) );
  XOR U36806 ( .A(n37742), .B(n33180), .Z(n33204) );
  XOR U36807 ( .A(n37743), .B(n33172), .Z(n33180) );
  XOR U36808 ( .A(n37744), .B(n33161), .Z(n33172) );
  XNOR U36809 ( .A(q[30]), .B(DB[650]), .Z(n33161) );
  IV U36810 ( .A(n33160), .Z(n37744) );
  XNOR U36811 ( .A(n33158), .B(n37745), .Z(n33160) );
  XNOR U36812 ( .A(q[29]), .B(DB[649]), .Z(n37745) );
  XNOR U36813 ( .A(q[28]), .B(DB[648]), .Z(n33158) );
  IV U36814 ( .A(n33171), .Z(n37743) );
  XOR U36815 ( .A(n37746), .B(n37747), .Z(n33171) );
  XNOR U36816 ( .A(n33167), .B(n33169), .Z(n37747) );
  XNOR U36817 ( .A(q[24]), .B(DB[644]), .Z(n33169) );
  XNOR U36818 ( .A(q[27]), .B(DB[647]), .Z(n33167) );
  IV U36819 ( .A(n33166), .Z(n37746) );
  XNOR U36820 ( .A(n33164), .B(n37748), .Z(n33166) );
  XNOR U36821 ( .A(q[26]), .B(DB[646]), .Z(n37748) );
  XNOR U36822 ( .A(q[25]), .B(DB[645]), .Z(n33164) );
  IV U36823 ( .A(n33179), .Z(n37742) );
  XOR U36824 ( .A(n37749), .B(n37750), .Z(n33179) );
  XNOR U36825 ( .A(n33196), .B(n33177), .Z(n37750) );
  XNOR U36826 ( .A(q[16]), .B(DB[636]), .Z(n33177) );
  XOR U36827 ( .A(n37751), .B(n33185), .Z(n33196) );
  XNOR U36828 ( .A(q[23]), .B(DB[643]), .Z(n33185) );
  IV U36829 ( .A(n33184), .Z(n37751) );
  XNOR U36830 ( .A(n33182), .B(n37752), .Z(n33184) );
  XNOR U36831 ( .A(q[22]), .B(DB[642]), .Z(n37752) );
  XNOR U36832 ( .A(q[21]), .B(DB[641]), .Z(n33182) );
  IV U36833 ( .A(n33195), .Z(n37749) );
  XOR U36834 ( .A(n37753), .B(n37754), .Z(n33195) );
  XNOR U36835 ( .A(n33191), .B(n33193), .Z(n37754) );
  XNOR U36836 ( .A(q[17]), .B(DB[637]), .Z(n33193) );
  XNOR U36837 ( .A(q[20]), .B(DB[640]), .Z(n33191) );
  IV U36838 ( .A(n33190), .Z(n37753) );
  XNOR U36839 ( .A(n33188), .B(n37755), .Z(n33190) );
  XNOR U36840 ( .A(q[19]), .B(DB[639]), .Z(n37755) );
  XNOR U36841 ( .A(q[18]), .B(DB[638]), .Z(n33188) );
  IV U36842 ( .A(n33203), .Z(n37741) );
  XOR U36843 ( .A(n37756), .B(n37757), .Z(n33203) );
  XNOR U36844 ( .A(n33230), .B(n33201), .Z(n37757) );
  XNOR U36845 ( .A(q[0]), .B(DB[620]), .Z(n33201) );
  XOR U36846 ( .A(n37758), .B(n33222), .Z(n33230) );
  XOR U36847 ( .A(n37759), .B(n33210), .Z(n33222) );
  XNOR U36848 ( .A(q[15]), .B(DB[635]), .Z(n33210) );
  IV U36849 ( .A(n33209), .Z(n37759) );
  XNOR U36850 ( .A(n33207), .B(n37760), .Z(n33209) );
  XNOR U36851 ( .A(q[14]), .B(DB[634]), .Z(n37760) );
  XNOR U36852 ( .A(q[13]), .B(DB[633]), .Z(n33207) );
  IV U36853 ( .A(n33221), .Z(n37758) );
  XOR U36854 ( .A(n37761), .B(n37762), .Z(n33221) );
  XNOR U36855 ( .A(n33217), .B(n33219), .Z(n37762) );
  XNOR U36856 ( .A(q[9]), .B(DB[629]), .Z(n33219) );
  XNOR U36857 ( .A(q[12]), .B(DB[632]), .Z(n33217) );
  IV U36858 ( .A(n33216), .Z(n37761) );
  XNOR U36859 ( .A(n33214), .B(n37763), .Z(n33216) );
  XNOR U36860 ( .A(q[11]), .B(DB[631]), .Z(n37763) );
  XNOR U36861 ( .A(q[10]), .B(DB[630]), .Z(n33214) );
  IV U36862 ( .A(n33229), .Z(n37756) );
  XOR U36863 ( .A(n37764), .B(n37765), .Z(n33229) );
  XNOR U36864 ( .A(n33246), .B(n33227), .Z(n37765) );
  XNOR U36865 ( .A(q[1]), .B(DB[621]), .Z(n33227) );
  XOR U36866 ( .A(n37766), .B(n33235), .Z(n33246) );
  XNOR U36867 ( .A(q[8]), .B(DB[628]), .Z(n33235) );
  IV U36868 ( .A(n33234), .Z(n37766) );
  XNOR U36869 ( .A(n33232), .B(n37767), .Z(n33234) );
  XNOR U36870 ( .A(q[7]), .B(DB[627]), .Z(n37767) );
  XNOR U36871 ( .A(q[6]), .B(DB[626]), .Z(n33232) );
  IV U36872 ( .A(n33245), .Z(n37764) );
  XOR U36873 ( .A(n37768), .B(n37769), .Z(n33245) );
  XNOR U36874 ( .A(n33241), .B(n33243), .Z(n37769) );
  XNOR U36875 ( .A(q[2]), .B(DB[622]), .Z(n33243) );
  XNOR U36876 ( .A(q[5]), .B(DB[625]), .Z(n33241) );
  IV U36877 ( .A(n33240), .Z(n37768) );
  XNOR U36878 ( .A(n33238), .B(n37770), .Z(n33240) );
  XNOR U36879 ( .A(q[4]), .B(DB[624]), .Z(n37770) );
  XNOR U36880 ( .A(q[3]), .B(DB[623]), .Z(n33238) );
  XOR U36881 ( .A(n37771), .B(n33007), .Z(n32858) );
  XOR U36882 ( .A(n37772), .B(n32983), .Z(n33007) );
  XOR U36883 ( .A(n37773), .B(n32975), .Z(n32983) );
  XOR U36884 ( .A(n37774), .B(n32964), .Z(n32975) );
  XNOR U36885 ( .A(q[30]), .B(DB[681]), .Z(n32964) );
  IV U36886 ( .A(n32963), .Z(n37774) );
  XNOR U36887 ( .A(n32961), .B(n37775), .Z(n32963) );
  XNOR U36888 ( .A(q[29]), .B(DB[680]), .Z(n37775) );
  XNOR U36889 ( .A(q[28]), .B(DB[679]), .Z(n32961) );
  IV U36890 ( .A(n32974), .Z(n37773) );
  XOR U36891 ( .A(n37776), .B(n37777), .Z(n32974) );
  XNOR U36892 ( .A(n32970), .B(n32972), .Z(n37777) );
  XNOR U36893 ( .A(q[24]), .B(DB[675]), .Z(n32972) );
  XNOR U36894 ( .A(q[27]), .B(DB[678]), .Z(n32970) );
  IV U36895 ( .A(n32969), .Z(n37776) );
  XNOR U36896 ( .A(n32967), .B(n37778), .Z(n32969) );
  XNOR U36897 ( .A(q[26]), .B(DB[677]), .Z(n37778) );
  XNOR U36898 ( .A(q[25]), .B(DB[676]), .Z(n32967) );
  IV U36899 ( .A(n32982), .Z(n37772) );
  XOR U36900 ( .A(n37779), .B(n37780), .Z(n32982) );
  XNOR U36901 ( .A(n32999), .B(n32980), .Z(n37780) );
  XNOR U36902 ( .A(q[16]), .B(DB[667]), .Z(n32980) );
  XOR U36903 ( .A(n37781), .B(n32988), .Z(n32999) );
  XNOR U36904 ( .A(q[23]), .B(DB[674]), .Z(n32988) );
  IV U36905 ( .A(n32987), .Z(n37781) );
  XNOR U36906 ( .A(n32985), .B(n37782), .Z(n32987) );
  XNOR U36907 ( .A(q[22]), .B(DB[673]), .Z(n37782) );
  XNOR U36908 ( .A(q[21]), .B(DB[672]), .Z(n32985) );
  IV U36909 ( .A(n32998), .Z(n37779) );
  XOR U36910 ( .A(n37783), .B(n37784), .Z(n32998) );
  XNOR U36911 ( .A(n32994), .B(n32996), .Z(n37784) );
  XNOR U36912 ( .A(q[17]), .B(DB[668]), .Z(n32996) );
  XNOR U36913 ( .A(q[20]), .B(DB[671]), .Z(n32994) );
  IV U36914 ( .A(n32993), .Z(n37783) );
  XNOR U36915 ( .A(n32991), .B(n37785), .Z(n32993) );
  XNOR U36916 ( .A(q[19]), .B(DB[670]), .Z(n37785) );
  XNOR U36917 ( .A(q[18]), .B(DB[669]), .Z(n32991) );
  IV U36918 ( .A(n33006), .Z(n37771) );
  XOR U36919 ( .A(n37786), .B(n37787), .Z(n33006) );
  XNOR U36920 ( .A(n33033), .B(n33004), .Z(n37787) );
  XNOR U36921 ( .A(q[0]), .B(DB[651]), .Z(n33004) );
  XOR U36922 ( .A(n37788), .B(n33025), .Z(n33033) );
  XOR U36923 ( .A(n37789), .B(n33013), .Z(n33025) );
  XNOR U36924 ( .A(q[15]), .B(DB[666]), .Z(n33013) );
  IV U36925 ( .A(n33012), .Z(n37789) );
  XNOR U36926 ( .A(n33010), .B(n37790), .Z(n33012) );
  XNOR U36927 ( .A(q[14]), .B(DB[665]), .Z(n37790) );
  XNOR U36928 ( .A(q[13]), .B(DB[664]), .Z(n33010) );
  IV U36929 ( .A(n33024), .Z(n37788) );
  XOR U36930 ( .A(n37791), .B(n37792), .Z(n33024) );
  XNOR U36931 ( .A(n33020), .B(n33022), .Z(n37792) );
  XNOR U36932 ( .A(q[9]), .B(DB[660]), .Z(n33022) );
  XNOR U36933 ( .A(q[12]), .B(DB[663]), .Z(n33020) );
  IV U36934 ( .A(n33019), .Z(n37791) );
  XNOR U36935 ( .A(n33017), .B(n37793), .Z(n33019) );
  XNOR U36936 ( .A(q[11]), .B(DB[662]), .Z(n37793) );
  XNOR U36937 ( .A(q[10]), .B(DB[661]), .Z(n33017) );
  IV U36938 ( .A(n33032), .Z(n37786) );
  XOR U36939 ( .A(n37794), .B(n37795), .Z(n33032) );
  XNOR U36940 ( .A(n33049), .B(n33030), .Z(n37795) );
  XNOR U36941 ( .A(q[1]), .B(DB[652]), .Z(n33030) );
  XOR U36942 ( .A(n37796), .B(n33038), .Z(n33049) );
  XNOR U36943 ( .A(q[8]), .B(DB[659]), .Z(n33038) );
  IV U36944 ( .A(n33037), .Z(n37796) );
  XNOR U36945 ( .A(n33035), .B(n37797), .Z(n33037) );
  XNOR U36946 ( .A(q[7]), .B(DB[658]), .Z(n37797) );
  XNOR U36947 ( .A(q[6]), .B(DB[657]), .Z(n33035) );
  IV U36948 ( .A(n33048), .Z(n37794) );
  XOR U36949 ( .A(n37798), .B(n37799), .Z(n33048) );
  XNOR U36950 ( .A(n33044), .B(n33046), .Z(n37799) );
  XNOR U36951 ( .A(q[2]), .B(DB[653]), .Z(n33046) );
  XNOR U36952 ( .A(q[5]), .B(DB[656]), .Z(n33044) );
  IV U36953 ( .A(n33043), .Z(n37798) );
  XNOR U36954 ( .A(n33041), .B(n37800), .Z(n33043) );
  XNOR U36955 ( .A(q[4]), .B(DB[655]), .Z(n37800) );
  XNOR U36956 ( .A(q[3]), .B(DB[654]), .Z(n33041) );
  XOR U36957 ( .A(n37801), .B(n32810), .Z(n32661) );
  XOR U36958 ( .A(n37802), .B(n32786), .Z(n32810) );
  XOR U36959 ( .A(n37803), .B(n32778), .Z(n32786) );
  XOR U36960 ( .A(n37804), .B(n32767), .Z(n32778) );
  XNOR U36961 ( .A(q[30]), .B(DB[712]), .Z(n32767) );
  IV U36962 ( .A(n32766), .Z(n37804) );
  XNOR U36963 ( .A(n32764), .B(n37805), .Z(n32766) );
  XNOR U36964 ( .A(q[29]), .B(DB[711]), .Z(n37805) );
  XNOR U36965 ( .A(q[28]), .B(DB[710]), .Z(n32764) );
  IV U36966 ( .A(n32777), .Z(n37803) );
  XOR U36967 ( .A(n37806), .B(n37807), .Z(n32777) );
  XNOR U36968 ( .A(n32773), .B(n32775), .Z(n37807) );
  XNOR U36969 ( .A(q[24]), .B(DB[706]), .Z(n32775) );
  XNOR U36970 ( .A(q[27]), .B(DB[709]), .Z(n32773) );
  IV U36971 ( .A(n32772), .Z(n37806) );
  XNOR U36972 ( .A(n32770), .B(n37808), .Z(n32772) );
  XNOR U36973 ( .A(q[26]), .B(DB[708]), .Z(n37808) );
  XNOR U36974 ( .A(q[25]), .B(DB[707]), .Z(n32770) );
  IV U36975 ( .A(n32785), .Z(n37802) );
  XOR U36976 ( .A(n37809), .B(n37810), .Z(n32785) );
  XNOR U36977 ( .A(n32802), .B(n32783), .Z(n37810) );
  XNOR U36978 ( .A(q[16]), .B(DB[698]), .Z(n32783) );
  XOR U36979 ( .A(n37811), .B(n32791), .Z(n32802) );
  XNOR U36980 ( .A(q[23]), .B(DB[705]), .Z(n32791) );
  IV U36981 ( .A(n32790), .Z(n37811) );
  XNOR U36982 ( .A(n32788), .B(n37812), .Z(n32790) );
  XNOR U36983 ( .A(q[22]), .B(DB[704]), .Z(n37812) );
  XNOR U36984 ( .A(q[21]), .B(DB[703]), .Z(n32788) );
  IV U36985 ( .A(n32801), .Z(n37809) );
  XOR U36986 ( .A(n37813), .B(n37814), .Z(n32801) );
  XNOR U36987 ( .A(n32797), .B(n32799), .Z(n37814) );
  XNOR U36988 ( .A(q[17]), .B(DB[699]), .Z(n32799) );
  XNOR U36989 ( .A(q[20]), .B(DB[702]), .Z(n32797) );
  IV U36990 ( .A(n32796), .Z(n37813) );
  XNOR U36991 ( .A(n32794), .B(n37815), .Z(n32796) );
  XNOR U36992 ( .A(q[19]), .B(DB[701]), .Z(n37815) );
  XNOR U36993 ( .A(q[18]), .B(DB[700]), .Z(n32794) );
  IV U36994 ( .A(n32809), .Z(n37801) );
  XOR U36995 ( .A(n37816), .B(n37817), .Z(n32809) );
  XNOR U36996 ( .A(n32836), .B(n32807), .Z(n37817) );
  XNOR U36997 ( .A(q[0]), .B(DB[682]), .Z(n32807) );
  XOR U36998 ( .A(n37818), .B(n32828), .Z(n32836) );
  XOR U36999 ( .A(n37819), .B(n32816), .Z(n32828) );
  XNOR U37000 ( .A(q[15]), .B(DB[697]), .Z(n32816) );
  IV U37001 ( .A(n32815), .Z(n37819) );
  XNOR U37002 ( .A(n32813), .B(n37820), .Z(n32815) );
  XNOR U37003 ( .A(q[14]), .B(DB[696]), .Z(n37820) );
  XNOR U37004 ( .A(q[13]), .B(DB[695]), .Z(n32813) );
  IV U37005 ( .A(n32827), .Z(n37818) );
  XOR U37006 ( .A(n37821), .B(n37822), .Z(n32827) );
  XNOR U37007 ( .A(n32823), .B(n32825), .Z(n37822) );
  XNOR U37008 ( .A(q[9]), .B(DB[691]), .Z(n32825) );
  XNOR U37009 ( .A(q[12]), .B(DB[694]), .Z(n32823) );
  IV U37010 ( .A(n32822), .Z(n37821) );
  XNOR U37011 ( .A(n32820), .B(n37823), .Z(n32822) );
  XNOR U37012 ( .A(q[11]), .B(DB[693]), .Z(n37823) );
  XNOR U37013 ( .A(q[10]), .B(DB[692]), .Z(n32820) );
  IV U37014 ( .A(n32835), .Z(n37816) );
  XOR U37015 ( .A(n37824), .B(n37825), .Z(n32835) );
  XNOR U37016 ( .A(n32852), .B(n32833), .Z(n37825) );
  XNOR U37017 ( .A(q[1]), .B(DB[683]), .Z(n32833) );
  XOR U37018 ( .A(n37826), .B(n32841), .Z(n32852) );
  XNOR U37019 ( .A(q[8]), .B(DB[690]), .Z(n32841) );
  IV U37020 ( .A(n32840), .Z(n37826) );
  XNOR U37021 ( .A(n32838), .B(n37827), .Z(n32840) );
  XNOR U37022 ( .A(q[7]), .B(DB[689]), .Z(n37827) );
  XNOR U37023 ( .A(q[6]), .B(DB[688]), .Z(n32838) );
  IV U37024 ( .A(n32851), .Z(n37824) );
  XOR U37025 ( .A(n37828), .B(n37829), .Z(n32851) );
  XNOR U37026 ( .A(n32847), .B(n32849), .Z(n37829) );
  XNOR U37027 ( .A(q[2]), .B(DB[684]), .Z(n32849) );
  XNOR U37028 ( .A(q[5]), .B(DB[687]), .Z(n32847) );
  IV U37029 ( .A(n32846), .Z(n37828) );
  XNOR U37030 ( .A(n32844), .B(n37830), .Z(n32846) );
  XNOR U37031 ( .A(q[4]), .B(DB[686]), .Z(n37830) );
  XNOR U37032 ( .A(q[3]), .B(DB[685]), .Z(n32844) );
  XOR U37033 ( .A(n37831), .B(n32613), .Z(n32464) );
  XOR U37034 ( .A(n37832), .B(n32589), .Z(n32613) );
  XOR U37035 ( .A(n37833), .B(n32581), .Z(n32589) );
  XOR U37036 ( .A(n37834), .B(n32570), .Z(n32581) );
  XNOR U37037 ( .A(q[30]), .B(DB[743]), .Z(n32570) );
  IV U37038 ( .A(n32569), .Z(n37834) );
  XNOR U37039 ( .A(n32567), .B(n37835), .Z(n32569) );
  XNOR U37040 ( .A(q[29]), .B(DB[742]), .Z(n37835) );
  XNOR U37041 ( .A(q[28]), .B(DB[741]), .Z(n32567) );
  IV U37042 ( .A(n32580), .Z(n37833) );
  XOR U37043 ( .A(n37836), .B(n37837), .Z(n32580) );
  XNOR U37044 ( .A(n32576), .B(n32578), .Z(n37837) );
  XNOR U37045 ( .A(q[24]), .B(DB[737]), .Z(n32578) );
  XNOR U37046 ( .A(q[27]), .B(DB[740]), .Z(n32576) );
  IV U37047 ( .A(n32575), .Z(n37836) );
  XNOR U37048 ( .A(n32573), .B(n37838), .Z(n32575) );
  XNOR U37049 ( .A(q[26]), .B(DB[739]), .Z(n37838) );
  XNOR U37050 ( .A(q[25]), .B(DB[738]), .Z(n32573) );
  IV U37051 ( .A(n32588), .Z(n37832) );
  XOR U37052 ( .A(n37839), .B(n37840), .Z(n32588) );
  XNOR U37053 ( .A(n32605), .B(n32586), .Z(n37840) );
  XNOR U37054 ( .A(q[16]), .B(DB[729]), .Z(n32586) );
  XOR U37055 ( .A(n37841), .B(n32594), .Z(n32605) );
  XNOR U37056 ( .A(q[23]), .B(DB[736]), .Z(n32594) );
  IV U37057 ( .A(n32593), .Z(n37841) );
  XNOR U37058 ( .A(n32591), .B(n37842), .Z(n32593) );
  XNOR U37059 ( .A(q[22]), .B(DB[735]), .Z(n37842) );
  XNOR U37060 ( .A(q[21]), .B(DB[734]), .Z(n32591) );
  IV U37061 ( .A(n32604), .Z(n37839) );
  XOR U37062 ( .A(n37843), .B(n37844), .Z(n32604) );
  XNOR U37063 ( .A(n32600), .B(n32602), .Z(n37844) );
  XNOR U37064 ( .A(q[17]), .B(DB[730]), .Z(n32602) );
  XNOR U37065 ( .A(q[20]), .B(DB[733]), .Z(n32600) );
  IV U37066 ( .A(n32599), .Z(n37843) );
  XNOR U37067 ( .A(n32597), .B(n37845), .Z(n32599) );
  XNOR U37068 ( .A(q[19]), .B(DB[732]), .Z(n37845) );
  XNOR U37069 ( .A(q[18]), .B(DB[731]), .Z(n32597) );
  IV U37070 ( .A(n32612), .Z(n37831) );
  XOR U37071 ( .A(n37846), .B(n37847), .Z(n32612) );
  XNOR U37072 ( .A(n32639), .B(n32610), .Z(n37847) );
  XNOR U37073 ( .A(q[0]), .B(DB[713]), .Z(n32610) );
  XOR U37074 ( .A(n37848), .B(n32631), .Z(n32639) );
  XOR U37075 ( .A(n37849), .B(n32619), .Z(n32631) );
  XNOR U37076 ( .A(q[15]), .B(DB[728]), .Z(n32619) );
  IV U37077 ( .A(n32618), .Z(n37849) );
  XNOR U37078 ( .A(n32616), .B(n37850), .Z(n32618) );
  XNOR U37079 ( .A(q[14]), .B(DB[727]), .Z(n37850) );
  XNOR U37080 ( .A(q[13]), .B(DB[726]), .Z(n32616) );
  IV U37081 ( .A(n32630), .Z(n37848) );
  XOR U37082 ( .A(n37851), .B(n37852), .Z(n32630) );
  XNOR U37083 ( .A(n32626), .B(n32628), .Z(n37852) );
  XNOR U37084 ( .A(q[9]), .B(DB[722]), .Z(n32628) );
  XNOR U37085 ( .A(q[12]), .B(DB[725]), .Z(n32626) );
  IV U37086 ( .A(n32625), .Z(n37851) );
  XNOR U37087 ( .A(n32623), .B(n37853), .Z(n32625) );
  XNOR U37088 ( .A(q[11]), .B(DB[724]), .Z(n37853) );
  XNOR U37089 ( .A(q[10]), .B(DB[723]), .Z(n32623) );
  IV U37090 ( .A(n32638), .Z(n37846) );
  XOR U37091 ( .A(n37854), .B(n37855), .Z(n32638) );
  XNOR U37092 ( .A(n32655), .B(n32636), .Z(n37855) );
  XNOR U37093 ( .A(q[1]), .B(DB[714]), .Z(n32636) );
  XOR U37094 ( .A(n37856), .B(n32644), .Z(n32655) );
  XNOR U37095 ( .A(q[8]), .B(DB[721]), .Z(n32644) );
  IV U37096 ( .A(n32643), .Z(n37856) );
  XNOR U37097 ( .A(n32641), .B(n37857), .Z(n32643) );
  XNOR U37098 ( .A(q[7]), .B(DB[720]), .Z(n37857) );
  XNOR U37099 ( .A(q[6]), .B(DB[719]), .Z(n32641) );
  IV U37100 ( .A(n32654), .Z(n37854) );
  XOR U37101 ( .A(n37858), .B(n37859), .Z(n32654) );
  XNOR U37102 ( .A(n32650), .B(n32652), .Z(n37859) );
  XNOR U37103 ( .A(q[2]), .B(DB[715]), .Z(n32652) );
  XNOR U37104 ( .A(q[5]), .B(DB[718]), .Z(n32650) );
  IV U37105 ( .A(n32649), .Z(n37858) );
  XNOR U37106 ( .A(n32647), .B(n37860), .Z(n32649) );
  XNOR U37107 ( .A(q[4]), .B(DB[717]), .Z(n37860) );
  XNOR U37108 ( .A(q[3]), .B(DB[716]), .Z(n32647) );
  XOR U37109 ( .A(n37861), .B(n32416), .Z(n32267) );
  XOR U37110 ( .A(n37862), .B(n32392), .Z(n32416) );
  XOR U37111 ( .A(n37863), .B(n32384), .Z(n32392) );
  XOR U37112 ( .A(n37864), .B(n32373), .Z(n32384) );
  XNOR U37113 ( .A(q[30]), .B(DB[774]), .Z(n32373) );
  IV U37114 ( .A(n32372), .Z(n37864) );
  XNOR U37115 ( .A(n32370), .B(n37865), .Z(n32372) );
  XNOR U37116 ( .A(q[29]), .B(DB[773]), .Z(n37865) );
  XNOR U37117 ( .A(q[28]), .B(DB[772]), .Z(n32370) );
  IV U37118 ( .A(n32383), .Z(n37863) );
  XOR U37119 ( .A(n37866), .B(n37867), .Z(n32383) );
  XNOR U37120 ( .A(n32379), .B(n32381), .Z(n37867) );
  XNOR U37121 ( .A(q[24]), .B(DB[768]), .Z(n32381) );
  XNOR U37122 ( .A(q[27]), .B(DB[771]), .Z(n32379) );
  IV U37123 ( .A(n32378), .Z(n37866) );
  XNOR U37124 ( .A(n32376), .B(n37868), .Z(n32378) );
  XNOR U37125 ( .A(q[26]), .B(DB[770]), .Z(n37868) );
  XNOR U37126 ( .A(q[25]), .B(DB[769]), .Z(n32376) );
  IV U37127 ( .A(n32391), .Z(n37862) );
  XOR U37128 ( .A(n37869), .B(n37870), .Z(n32391) );
  XNOR U37129 ( .A(n32408), .B(n32389), .Z(n37870) );
  XNOR U37130 ( .A(q[16]), .B(DB[760]), .Z(n32389) );
  XOR U37131 ( .A(n37871), .B(n32397), .Z(n32408) );
  XNOR U37132 ( .A(q[23]), .B(DB[767]), .Z(n32397) );
  IV U37133 ( .A(n32396), .Z(n37871) );
  XNOR U37134 ( .A(n32394), .B(n37872), .Z(n32396) );
  XNOR U37135 ( .A(q[22]), .B(DB[766]), .Z(n37872) );
  XNOR U37136 ( .A(q[21]), .B(DB[765]), .Z(n32394) );
  IV U37137 ( .A(n32407), .Z(n37869) );
  XOR U37138 ( .A(n37873), .B(n37874), .Z(n32407) );
  XNOR U37139 ( .A(n32403), .B(n32405), .Z(n37874) );
  XNOR U37140 ( .A(q[17]), .B(DB[761]), .Z(n32405) );
  XNOR U37141 ( .A(q[20]), .B(DB[764]), .Z(n32403) );
  IV U37142 ( .A(n32402), .Z(n37873) );
  XNOR U37143 ( .A(n32400), .B(n37875), .Z(n32402) );
  XNOR U37144 ( .A(q[19]), .B(DB[763]), .Z(n37875) );
  XNOR U37145 ( .A(q[18]), .B(DB[762]), .Z(n32400) );
  IV U37146 ( .A(n32415), .Z(n37861) );
  XOR U37147 ( .A(n37876), .B(n37877), .Z(n32415) );
  XNOR U37148 ( .A(n32442), .B(n32413), .Z(n37877) );
  XNOR U37149 ( .A(q[0]), .B(DB[744]), .Z(n32413) );
  XOR U37150 ( .A(n37878), .B(n32434), .Z(n32442) );
  XOR U37151 ( .A(n37879), .B(n32422), .Z(n32434) );
  XNOR U37152 ( .A(q[15]), .B(DB[759]), .Z(n32422) );
  IV U37153 ( .A(n32421), .Z(n37879) );
  XNOR U37154 ( .A(n32419), .B(n37880), .Z(n32421) );
  XNOR U37155 ( .A(q[14]), .B(DB[758]), .Z(n37880) );
  XNOR U37156 ( .A(q[13]), .B(DB[757]), .Z(n32419) );
  IV U37157 ( .A(n32433), .Z(n37878) );
  XOR U37158 ( .A(n37881), .B(n37882), .Z(n32433) );
  XNOR U37159 ( .A(n32429), .B(n32431), .Z(n37882) );
  XNOR U37160 ( .A(q[9]), .B(DB[753]), .Z(n32431) );
  XNOR U37161 ( .A(q[12]), .B(DB[756]), .Z(n32429) );
  IV U37162 ( .A(n32428), .Z(n37881) );
  XNOR U37163 ( .A(n32426), .B(n37883), .Z(n32428) );
  XNOR U37164 ( .A(q[11]), .B(DB[755]), .Z(n37883) );
  XNOR U37165 ( .A(q[10]), .B(DB[754]), .Z(n32426) );
  IV U37166 ( .A(n32441), .Z(n37876) );
  XOR U37167 ( .A(n37884), .B(n37885), .Z(n32441) );
  XNOR U37168 ( .A(n32458), .B(n32439), .Z(n37885) );
  XNOR U37169 ( .A(q[1]), .B(DB[745]), .Z(n32439) );
  XOR U37170 ( .A(n37886), .B(n32447), .Z(n32458) );
  XNOR U37171 ( .A(q[8]), .B(DB[752]), .Z(n32447) );
  IV U37172 ( .A(n32446), .Z(n37886) );
  XNOR U37173 ( .A(n32444), .B(n37887), .Z(n32446) );
  XNOR U37174 ( .A(q[7]), .B(DB[751]), .Z(n37887) );
  XNOR U37175 ( .A(q[6]), .B(DB[750]), .Z(n32444) );
  IV U37176 ( .A(n32457), .Z(n37884) );
  XOR U37177 ( .A(n37888), .B(n37889), .Z(n32457) );
  XNOR U37178 ( .A(n32453), .B(n32455), .Z(n37889) );
  XNOR U37179 ( .A(q[2]), .B(DB[746]), .Z(n32455) );
  XNOR U37180 ( .A(q[5]), .B(DB[749]), .Z(n32453) );
  IV U37181 ( .A(n32452), .Z(n37888) );
  XNOR U37182 ( .A(n32450), .B(n37890), .Z(n32452) );
  XNOR U37183 ( .A(q[4]), .B(DB[748]), .Z(n37890) );
  XNOR U37184 ( .A(q[3]), .B(DB[747]), .Z(n32450) );
  XOR U37185 ( .A(n37891), .B(n32219), .Z(n32070) );
  XOR U37186 ( .A(n37892), .B(n32195), .Z(n32219) );
  XOR U37187 ( .A(n37893), .B(n32187), .Z(n32195) );
  XOR U37188 ( .A(n37894), .B(n32176), .Z(n32187) );
  XNOR U37189 ( .A(q[30]), .B(DB[805]), .Z(n32176) );
  IV U37190 ( .A(n32175), .Z(n37894) );
  XNOR U37191 ( .A(n32173), .B(n37895), .Z(n32175) );
  XNOR U37192 ( .A(q[29]), .B(DB[804]), .Z(n37895) );
  XNOR U37193 ( .A(q[28]), .B(DB[803]), .Z(n32173) );
  IV U37194 ( .A(n32186), .Z(n37893) );
  XOR U37195 ( .A(n37896), .B(n37897), .Z(n32186) );
  XNOR U37196 ( .A(n32182), .B(n32184), .Z(n37897) );
  XNOR U37197 ( .A(q[24]), .B(DB[799]), .Z(n32184) );
  XNOR U37198 ( .A(q[27]), .B(DB[802]), .Z(n32182) );
  IV U37199 ( .A(n32181), .Z(n37896) );
  XNOR U37200 ( .A(n32179), .B(n37898), .Z(n32181) );
  XNOR U37201 ( .A(q[26]), .B(DB[801]), .Z(n37898) );
  XNOR U37202 ( .A(q[25]), .B(DB[800]), .Z(n32179) );
  IV U37203 ( .A(n32194), .Z(n37892) );
  XOR U37204 ( .A(n37899), .B(n37900), .Z(n32194) );
  XNOR U37205 ( .A(n32211), .B(n32192), .Z(n37900) );
  XNOR U37206 ( .A(q[16]), .B(DB[791]), .Z(n32192) );
  XOR U37207 ( .A(n37901), .B(n32200), .Z(n32211) );
  XNOR U37208 ( .A(q[23]), .B(DB[798]), .Z(n32200) );
  IV U37209 ( .A(n32199), .Z(n37901) );
  XNOR U37210 ( .A(n32197), .B(n37902), .Z(n32199) );
  XNOR U37211 ( .A(q[22]), .B(DB[797]), .Z(n37902) );
  XNOR U37212 ( .A(q[21]), .B(DB[796]), .Z(n32197) );
  IV U37213 ( .A(n32210), .Z(n37899) );
  XOR U37214 ( .A(n37903), .B(n37904), .Z(n32210) );
  XNOR U37215 ( .A(n32206), .B(n32208), .Z(n37904) );
  XNOR U37216 ( .A(q[17]), .B(DB[792]), .Z(n32208) );
  XNOR U37217 ( .A(q[20]), .B(DB[795]), .Z(n32206) );
  IV U37218 ( .A(n32205), .Z(n37903) );
  XNOR U37219 ( .A(n32203), .B(n37905), .Z(n32205) );
  XNOR U37220 ( .A(q[19]), .B(DB[794]), .Z(n37905) );
  XNOR U37221 ( .A(q[18]), .B(DB[793]), .Z(n32203) );
  IV U37222 ( .A(n32218), .Z(n37891) );
  XOR U37223 ( .A(n37906), .B(n37907), .Z(n32218) );
  XNOR U37224 ( .A(n32245), .B(n32216), .Z(n37907) );
  XNOR U37225 ( .A(q[0]), .B(DB[775]), .Z(n32216) );
  XOR U37226 ( .A(n37908), .B(n32237), .Z(n32245) );
  XOR U37227 ( .A(n37909), .B(n32225), .Z(n32237) );
  XNOR U37228 ( .A(q[15]), .B(DB[790]), .Z(n32225) );
  IV U37229 ( .A(n32224), .Z(n37909) );
  XNOR U37230 ( .A(n32222), .B(n37910), .Z(n32224) );
  XNOR U37231 ( .A(q[14]), .B(DB[789]), .Z(n37910) );
  XNOR U37232 ( .A(q[13]), .B(DB[788]), .Z(n32222) );
  IV U37233 ( .A(n32236), .Z(n37908) );
  XOR U37234 ( .A(n37911), .B(n37912), .Z(n32236) );
  XNOR U37235 ( .A(n32232), .B(n32234), .Z(n37912) );
  XNOR U37236 ( .A(q[9]), .B(DB[784]), .Z(n32234) );
  XNOR U37237 ( .A(q[12]), .B(DB[787]), .Z(n32232) );
  IV U37238 ( .A(n32231), .Z(n37911) );
  XNOR U37239 ( .A(n32229), .B(n37913), .Z(n32231) );
  XNOR U37240 ( .A(q[11]), .B(DB[786]), .Z(n37913) );
  XNOR U37241 ( .A(q[10]), .B(DB[785]), .Z(n32229) );
  IV U37242 ( .A(n32244), .Z(n37906) );
  XOR U37243 ( .A(n37914), .B(n37915), .Z(n32244) );
  XNOR U37244 ( .A(n32261), .B(n32242), .Z(n37915) );
  XNOR U37245 ( .A(q[1]), .B(DB[776]), .Z(n32242) );
  XOR U37246 ( .A(n37916), .B(n32250), .Z(n32261) );
  XNOR U37247 ( .A(q[8]), .B(DB[783]), .Z(n32250) );
  IV U37248 ( .A(n32249), .Z(n37916) );
  XNOR U37249 ( .A(n32247), .B(n37917), .Z(n32249) );
  XNOR U37250 ( .A(q[7]), .B(DB[782]), .Z(n37917) );
  XNOR U37251 ( .A(q[6]), .B(DB[781]), .Z(n32247) );
  IV U37252 ( .A(n32260), .Z(n37914) );
  XOR U37253 ( .A(n37918), .B(n37919), .Z(n32260) );
  XNOR U37254 ( .A(n32256), .B(n32258), .Z(n37919) );
  XNOR U37255 ( .A(q[2]), .B(DB[777]), .Z(n32258) );
  XNOR U37256 ( .A(q[5]), .B(DB[780]), .Z(n32256) );
  IV U37257 ( .A(n32255), .Z(n37918) );
  XNOR U37258 ( .A(n32253), .B(n37920), .Z(n32255) );
  XNOR U37259 ( .A(q[4]), .B(DB[779]), .Z(n37920) );
  XNOR U37260 ( .A(q[3]), .B(DB[778]), .Z(n32253) );
  XOR U37261 ( .A(n37921), .B(n32022), .Z(n31873) );
  XOR U37262 ( .A(n37922), .B(n31998), .Z(n32022) );
  XOR U37263 ( .A(n37923), .B(n31990), .Z(n31998) );
  XOR U37264 ( .A(n37924), .B(n31979), .Z(n31990) );
  XNOR U37265 ( .A(q[30]), .B(DB[836]), .Z(n31979) );
  IV U37266 ( .A(n31978), .Z(n37924) );
  XNOR U37267 ( .A(n31976), .B(n37925), .Z(n31978) );
  XNOR U37268 ( .A(q[29]), .B(DB[835]), .Z(n37925) );
  XNOR U37269 ( .A(q[28]), .B(DB[834]), .Z(n31976) );
  IV U37270 ( .A(n31989), .Z(n37923) );
  XOR U37271 ( .A(n37926), .B(n37927), .Z(n31989) );
  XNOR U37272 ( .A(n31985), .B(n31987), .Z(n37927) );
  XNOR U37273 ( .A(q[24]), .B(DB[830]), .Z(n31987) );
  XNOR U37274 ( .A(q[27]), .B(DB[833]), .Z(n31985) );
  IV U37275 ( .A(n31984), .Z(n37926) );
  XNOR U37276 ( .A(n31982), .B(n37928), .Z(n31984) );
  XNOR U37277 ( .A(q[26]), .B(DB[832]), .Z(n37928) );
  XNOR U37278 ( .A(q[25]), .B(DB[831]), .Z(n31982) );
  IV U37279 ( .A(n31997), .Z(n37922) );
  XOR U37280 ( .A(n37929), .B(n37930), .Z(n31997) );
  XNOR U37281 ( .A(n32014), .B(n31995), .Z(n37930) );
  XNOR U37282 ( .A(q[16]), .B(DB[822]), .Z(n31995) );
  XOR U37283 ( .A(n37931), .B(n32003), .Z(n32014) );
  XNOR U37284 ( .A(q[23]), .B(DB[829]), .Z(n32003) );
  IV U37285 ( .A(n32002), .Z(n37931) );
  XNOR U37286 ( .A(n32000), .B(n37932), .Z(n32002) );
  XNOR U37287 ( .A(q[22]), .B(DB[828]), .Z(n37932) );
  XNOR U37288 ( .A(q[21]), .B(DB[827]), .Z(n32000) );
  IV U37289 ( .A(n32013), .Z(n37929) );
  XOR U37290 ( .A(n37933), .B(n37934), .Z(n32013) );
  XNOR U37291 ( .A(n32009), .B(n32011), .Z(n37934) );
  XNOR U37292 ( .A(q[17]), .B(DB[823]), .Z(n32011) );
  XNOR U37293 ( .A(q[20]), .B(DB[826]), .Z(n32009) );
  IV U37294 ( .A(n32008), .Z(n37933) );
  XNOR U37295 ( .A(n32006), .B(n37935), .Z(n32008) );
  XNOR U37296 ( .A(q[19]), .B(DB[825]), .Z(n37935) );
  XNOR U37297 ( .A(q[18]), .B(DB[824]), .Z(n32006) );
  IV U37298 ( .A(n32021), .Z(n37921) );
  XOR U37299 ( .A(n37936), .B(n37937), .Z(n32021) );
  XNOR U37300 ( .A(n32048), .B(n32019), .Z(n37937) );
  XNOR U37301 ( .A(q[0]), .B(DB[806]), .Z(n32019) );
  XOR U37302 ( .A(n37938), .B(n32040), .Z(n32048) );
  XOR U37303 ( .A(n37939), .B(n32028), .Z(n32040) );
  XNOR U37304 ( .A(q[15]), .B(DB[821]), .Z(n32028) );
  IV U37305 ( .A(n32027), .Z(n37939) );
  XNOR U37306 ( .A(n32025), .B(n37940), .Z(n32027) );
  XNOR U37307 ( .A(q[14]), .B(DB[820]), .Z(n37940) );
  XNOR U37308 ( .A(q[13]), .B(DB[819]), .Z(n32025) );
  IV U37309 ( .A(n32039), .Z(n37938) );
  XOR U37310 ( .A(n37941), .B(n37942), .Z(n32039) );
  XNOR U37311 ( .A(n32035), .B(n32037), .Z(n37942) );
  XNOR U37312 ( .A(q[9]), .B(DB[815]), .Z(n32037) );
  XNOR U37313 ( .A(q[12]), .B(DB[818]), .Z(n32035) );
  IV U37314 ( .A(n32034), .Z(n37941) );
  XNOR U37315 ( .A(n32032), .B(n37943), .Z(n32034) );
  XNOR U37316 ( .A(q[11]), .B(DB[817]), .Z(n37943) );
  XNOR U37317 ( .A(q[10]), .B(DB[816]), .Z(n32032) );
  IV U37318 ( .A(n32047), .Z(n37936) );
  XOR U37319 ( .A(n37944), .B(n37945), .Z(n32047) );
  XNOR U37320 ( .A(n32064), .B(n32045), .Z(n37945) );
  XNOR U37321 ( .A(q[1]), .B(DB[807]), .Z(n32045) );
  XOR U37322 ( .A(n37946), .B(n32053), .Z(n32064) );
  XNOR U37323 ( .A(q[8]), .B(DB[814]), .Z(n32053) );
  IV U37324 ( .A(n32052), .Z(n37946) );
  XNOR U37325 ( .A(n32050), .B(n37947), .Z(n32052) );
  XNOR U37326 ( .A(q[7]), .B(DB[813]), .Z(n37947) );
  XNOR U37327 ( .A(q[6]), .B(DB[812]), .Z(n32050) );
  IV U37328 ( .A(n32063), .Z(n37944) );
  XOR U37329 ( .A(n37948), .B(n37949), .Z(n32063) );
  XNOR U37330 ( .A(n32059), .B(n32061), .Z(n37949) );
  XNOR U37331 ( .A(q[2]), .B(DB[808]), .Z(n32061) );
  XNOR U37332 ( .A(q[5]), .B(DB[811]), .Z(n32059) );
  IV U37333 ( .A(n32058), .Z(n37948) );
  XNOR U37334 ( .A(n32056), .B(n37950), .Z(n32058) );
  XNOR U37335 ( .A(q[4]), .B(DB[810]), .Z(n37950) );
  XNOR U37336 ( .A(q[3]), .B(DB[809]), .Z(n32056) );
  XOR U37337 ( .A(n37951), .B(n31825), .Z(n31676) );
  XOR U37338 ( .A(n37952), .B(n31801), .Z(n31825) );
  XOR U37339 ( .A(n37953), .B(n31793), .Z(n31801) );
  XOR U37340 ( .A(n37954), .B(n31782), .Z(n31793) );
  XNOR U37341 ( .A(q[30]), .B(DB[867]), .Z(n31782) );
  IV U37342 ( .A(n31781), .Z(n37954) );
  XNOR U37343 ( .A(n31779), .B(n37955), .Z(n31781) );
  XNOR U37344 ( .A(q[29]), .B(DB[866]), .Z(n37955) );
  XNOR U37345 ( .A(q[28]), .B(DB[865]), .Z(n31779) );
  IV U37346 ( .A(n31792), .Z(n37953) );
  XOR U37347 ( .A(n37956), .B(n37957), .Z(n31792) );
  XNOR U37348 ( .A(n31788), .B(n31790), .Z(n37957) );
  XNOR U37349 ( .A(q[24]), .B(DB[861]), .Z(n31790) );
  XNOR U37350 ( .A(q[27]), .B(DB[864]), .Z(n31788) );
  IV U37351 ( .A(n31787), .Z(n37956) );
  XNOR U37352 ( .A(n31785), .B(n37958), .Z(n31787) );
  XNOR U37353 ( .A(q[26]), .B(DB[863]), .Z(n37958) );
  XNOR U37354 ( .A(q[25]), .B(DB[862]), .Z(n31785) );
  IV U37355 ( .A(n31800), .Z(n37952) );
  XOR U37356 ( .A(n37959), .B(n37960), .Z(n31800) );
  XNOR U37357 ( .A(n31817), .B(n31798), .Z(n37960) );
  XNOR U37358 ( .A(q[16]), .B(DB[853]), .Z(n31798) );
  XOR U37359 ( .A(n37961), .B(n31806), .Z(n31817) );
  XNOR U37360 ( .A(q[23]), .B(DB[860]), .Z(n31806) );
  IV U37361 ( .A(n31805), .Z(n37961) );
  XNOR U37362 ( .A(n31803), .B(n37962), .Z(n31805) );
  XNOR U37363 ( .A(q[22]), .B(DB[859]), .Z(n37962) );
  XNOR U37364 ( .A(q[21]), .B(DB[858]), .Z(n31803) );
  IV U37365 ( .A(n31816), .Z(n37959) );
  XOR U37366 ( .A(n37963), .B(n37964), .Z(n31816) );
  XNOR U37367 ( .A(n31812), .B(n31814), .Z(n37964) );
  XNOR U37368 ( .A(q[17]), .B(DB[854]), .Z(n31814) );
  XNOR U37369 ( .A(q[20]), .B(DB[857]), .Z(n31812) );
  IV U37370 ( .A(n31811), .Z(n37963) );
  XNOR U37371 ( .A(n31809), .B(n37965), .Z(n31811) );
  XNOR U37372 ( .A(q[19]), .B(DB[856]), .Z(n37965) );
  XNOR U37373 ( .A(q[18]), .B(DB[855]), .Z(n31809) );
  IV U37374 ( .A(n31824), .Z(n37951) );
  XOR U37375 ( .A(n37966), .B(n37967), .Z(n31824) );
  XNOR U37376 ( .A(n31851), .B(n31822), .Z(n37967) );
  XNOR U37377 ( .A(q[0]), .B(DB[837]), .Z(n31822) );
  XOR U37378 ( .A(n37968), .B(n31843), .Z(n31851) );
  XOR U37379 ( .A(n37969), .B(n31831), .Z(n31843) );
  XNOR U37380 ( .A(q[15]), .B(DB[852]), .Z(n31831) );
  IV U37381 ( .A(n31830), .Z(n37969) );
  XNOR U37382 ( .A(n31828), .B(n37970), .Z(n31830) );
  XNOR U37383 ( .A(q[14]), .B(DB[851]), .Z(n37970) );
  XNOR U37384 ( .A(q[13]), .B(DB[850]), .Z(n31828) );
  IV U37385 ( .A(n31842), .Z(n37968) );
  XOR U37386 ( .A(n37971), .B(n37972), .Z(n31842) );
  XNOR U37387 ( .A(n31838), .B(n31840), .Z(n37972) );
  XNOR U37388 ( .A(q[9]), .B(DB[846]), .Z(n31840) );
  XNOR U37389 ( .A(q[12]), .B(DB[849]), .Z(n31838) );
  IV U37390 ( .A(n31837), .Z(n37971) );
  XNOR U37391 ( .A(n31835), .B(n37973), .Z(n31837) );
  XNOR U37392 ( .A(q[11]), .B(DB[848]), .Z(n37973) );
  XNOR U37393 ( .A(q[10]), .B(DB[847]), .Z(n31835) );
  IV U37394 ( .A(n31850), .Z(n37966) );
  XOR U37395 ( .A(n37974), .B(n37975), .Z(n31850) );
  XNOR U37396 ( .A(n31867), .B(n31848), .Z(n37975) );
  XNOR U37397 ( .A(q[1]), .B(DB[838]), .Z(n31848) );
  XOR U37398 ( .A(n37976), .B(n31856), .Z(n31867) );
  XNOR U37399 ( .A(q[8]), .B(DB[845]), .Z(n31856) );
  IV U37400 ( .A(n31855), .Z(n37976) );
  XNOR U37401 ( .A(n31853), .B(n37977), .Z(n31855) );
  XNOR U37402 ( .A(q[7]), .B(DB[844]), .Z(n37977) );
  XNOR U37403 ( .A(q[6]), .B(DB[843]), .Z(n31853) );
  IV U37404 ( .A(n31866), .Z(n37974) );
  XOR U37405 ( .A(n37978), .B(n37979), .Z(n31866) );
  XNOR U37406 ( .A(n31862), .B(n31864), .Z(n37979) );
  XNOR U37407 ( .A(q[2]), .B(DB[839]), .Z(n31864) );
  XNOR U37408 ( .A(q[5]), .B(DB[842]), .Z(n31862) );
  IV U37409 ( .A(n31861), .Z(n37978) );
  XNOR U37410 ( .A(n31859), .B(n37980), .Z(n31861) );
  XNOR U37411 ( .A(q[4]), .B(DB[841]), .Z(n37980) );
  XNOR U37412 ( .A(q[3]), .B(DB[840]), .Z(n31859) );
  XOR U37413 ( .A(n37981), .B(n31628), .Z(n31479) );
  XOR U37414 ( .A(n37982), .B(n31604), .Z(n31628) );
  XOR U37415 ( .A(n37983), .B(n31596), .Z(n31604) );
  XOR U37416 ( .A(n37984), .B(n31585), .Z(n31596) );
  XNOR U37417 ( .A(q[30]), .B(DB[898]), .Z(n31585) );
  IV U37418 ( .A(n31584), .Z(n37984) );
  XNOR U37419 ( .A(n31582), .B(n37985), .Z(n31584) );
  XNOR U37420 ( .A(q[29]), .B(DB[897]), .Z(n37985) );
  XNOR U37421 ( .A(q[28]), .B(DB[896]), .Z(n31582) );
  IV U37422 ( .A(n31595), .Z(n37983) );
  XOR U37423 ( .A(n37986), .B(n37987), .Z(n31595) );
  XNOR U37424 ( .A(n31591), .B(n31593), .Z(n37987) );
  XNOR U37425 ( .A(q[24]), .B(DB[892]), .Z(n31593) );
  XNOR U37426 ( .A(q[27]), .B(DB[895]), .Z(n31591) );
  IV U37427 ( .A(n31590), .Z(n37986) );
  XNOR U37428 ( .A(n31588), .B(n37988), .Z(n31590) );
  XNOR U37429 ( .A(q[26]), .B(DB[894]), .Z(n37988) );
  XNOR U37430 ( .A(q[25]), .B(DB[893]), .Z(n31588) );
  IV U37431 ( .A(n31603), .Z(n37982) );
  XOR U37432 ( .A(n37989), .B(n37990), .Z(n31603) );
  XNOR U37433 ( .A(n31620), .B(n31601), .Z(n37990) );
  XNOR U37434 ( .A(q[16]), .B(DB[884]), .Z(n31601) );
  XOR U37435 ( .A(n37991), .B(n31609), .Z(n31620) );
  XNOR U37436 ( .A(q[23]), .B(DB[891]), .Z(n31609) );
  IV U37437 ( .A(n31608), .Z(n37991) );
  XNOR U37438 ( .A(n31606), .B(n37992), .Z(n31608) );
  XNOR U37439 ( .A(q[22]), .B(DB[890]), .Z(n37992) );
  XNOR U37440 ( .A(q[21]), .B(DB[889]), .Z(n31606) );
  IV U37441 ( .A(n31619), .Z(n37989) );
  XOR U37442 ( .A(n37993), .B(n37994), .Z(n31619) );
  XNOR U37443 ( .A(n31615), .B(n31617), .Z(n37994) );
  XNOR U37444 ( .A(q[17]), .B(DB[885]), .Z(n31617) );
  XNOR U37445 ( .A(q[20]), .B(DB[888]), .Z(n31615) );
  IV U37446 ( .A(n31614), .Z(n37993) );
  XNOR U37447 ( .A(n31612), .B(n37995), .Z(n31614) );
  XNOR U37448 ( .A(q[19]), .B(DB[887]), .Z(n37995) );
  XNOR U37449 ( .A(q[18]), .B(DB[886]), .Z(n31612) );
  IV U37450 ( .A(n31627), .Z(n37981) );
  XOR U37451 ( .A(n37996), .B(n37997), .Z(n31627) );
  XNOR U37452 ( .A(n31654), .B(n31625), .Z(n37997) );
  XNOR U37453 ( .A(q[0]), .B(DB[868]), .Z(n31625) );
  XOR U37454 ( .A(n37998), .B(n31646), .Z(n31654) );
  XOR U37455 ( .A(n37999), .B(n31634), .Z(n31646) );
  XNOR U37456 ( .A(q[15]), .B(DB[883]), .Z(n31634) );
  IV U37457 ( .A(n31633), .Z(n37999) );
  XNOR U37458 ( .A(n31631), .B(n38000), .Z(n31633) );
  XNOR U37459 ( .A(q[14]), .B(DB[882]), .Z(n38000) );
  XNOR U37460 ( .A(q[13]), .B(DB[881]), .Z(n31631) );
  IV U37461 ( .A(n31645), .Z(n37998) );
  XOR U37462 ( .A(n38001), .B(n38002), .Z(n31645) );
  XNOR U37463 ( .A(n31641), .B(n31643), .Z(n38002) );
  XNOR U37464 ( .A(q[9]), .B(DB[877]), .Z(n31643) );
  XNOR U37465 ( .A(q[12]), .B(DB[880]), .Z(n31641) );
  IV U37466 ( .A(n31640), .Z(n38001) );
  XNOR U37467 ( .A(n31638), .B(n38003), .Z(n31640) );
  XNOR U37468 ( .A(q[11]), .B(DB[879]), .Z(n38003) );
  XNOR U37469 ( .A(q[10]), .B(DB[878]), .Z(n31638) );
  IV U37470 ( .A(n31653), .Z(n37996) );
  XOR U37471 ( .A(n38004), .B(n38005), .Z(n31653) );
  XNOR U37472 ( .A(n31670), .B(n31651), .Z(n38005) );
  XNOR U37473 ( .A(q[1]), .B(DB[869]), .Z(n31651) );
  XOR U37474 ( .A(n38006), .B(n31659), .Z(n31670) );
  XNOR U37475 ( .A(q[8]), .B(DB[876]), .Z(n31659) );
  IV U37476 ( .A(n31658), .Z(n38006) );
  XNOR U37477 ( .A(n31656), .B(n38007), .Z(n31658) );
  XNOR U37478 ( .A(q[7]), .B(DB[875]), .Z(n38007) );
  XNOR U37479 ( .A(q[6]), .B(DB[874]), .Z(n31656) );
  IV U37480 ( .A(n31669), .Z(n38004) );
  XOR U37481 ( .A(n38008), .B(n38009), .Z(n31669) );
  XNOR U37482 ( .A(n31665), .B(n31667), .Z(n38009) );
  XNOR U37483 ( .A(q[2]), .B(DB[870]), .Z(n31667) );
  XNOR U37484 ( .A(q[5]), .B(DB[873]), .Z(n31665) );
  IV U37485 ( .A(n31664), .Z(n38008) );
  XNOR U37486 ( .A(n31662), .B(n38010), .Z(n31664) );
  XNOR U37487 ( .A(q[4]), .B(DB[872]), .Z(n38010) );
  XNOR U37488 ( .A(q[3]), .B(DB[871]), .Z(n31662) );
  XOR U37489 ( .A(n38011), .B(n31431), .Z(n31282) );
  XOR U37490 ( .A(n38012), .B(n31407), .Z(n31431) );
  XOR U37491 ( .A(n38013), .B(n31399), .Z(n31407) );
  XOR U37492 ( .A(n38014), .B(n31388), .Z(n31399) );
  XNOR U37493 ( .A(q[30]), .B(DB[929]), .Z(n31388) );
  IV U37494 ( .A(n31387), .Z(n38014) );
  XNOR U37495 ( .A(n31385), .B(n38015), .Z(n31387) );
  XNOR U37496 ( .A(q[29]), .B(DB[928]), .Z(n38015) );
  XNOR U37497 ( .A(q[28]), .B(DB[927]), .Z(n31385) );
  IV U37498 ( .A(n31398), .Z(n38013) );
  XOR U37499 ( .A(n38016), .B(n38017), .Z(n31398) );
  XNOR U37500 ( .A(n31394), .B(n31396), .Z(n38017) );
  XNOR U37501 ( .A(q[24]), .B(DB[923]), .Z(n31396) );
  XNOR U37502 ( .A(q[27]), .B(DB[926]), .Z(n31394) );
  IV U37503 ( .A(n31393), .Z(n38016) );
  XNOR U37504 ( .A(n31391), .B(n38018), .Z(n31393) );
  XNOR U37505 ( .A(q[26]), .B(DB[925]), .Z(n38018) );
  XNOR U37506 ( .A(q[25]), .B(DB[924]), .Z(n31391) );
  IV U37507 ( .A(n31406), .Z(n38012) );
  XOR U37508 ( .A(n38019), .B(n38020), .Z(n31406) );
  XNOR U37509 ( .A(n31423), .B(n31404), .Z(n38020) );
  XNOR U37510 ( .A(q[16]), .B(DB[915]), .Z(n31404) );
  XOR U37511 ( .A(n38021), .B(n31412), .Z(n31423) );
  XNOR U37512 ( .A(q[23]), .B(DB[922]), .Z(n31412) );
  IV U37513 ( .A(n31411), .Z(n38021) );
  XNOR U37514 ( .A(n31409), .B(n38022), .Z(n31411) );
  XNOR U37515 ( .A(q[22]), .B(DB[921]), .Z(n38022) );
  XNOR U37516 ( .A(q[21]), .B(DB[920]), .Z(n31409) );
  IV U37517 ( .A(n31422), .Z(n38019) );
  XOR U37518 ( .A(n38023), .B(n38024), .Z(n31422) );
  XNOR U37519 ( .A(n31418), .B(n31420), .Z(n38024) );
  XNOR U37520 ( .A(q[17]), .B(DB[916]), .Z(n31420) );
  XNOR U37521 ( .A(q[20]), .B(DB[919]), .Z(n31418) );
  IV U37522 ( .A(n31417), .Z(n38023) );
  XNOR U37523 ( .A(n31415), .B(n38025), .Z(n31417) );
  XNOR U37524 ( .A(q[19]), .B(DB[918]), .Z(n38025) );
  XNOR U37525 ( .A(q[18]), .B(DB[917]), .Z(n31415) );
  IV U37526 ( .A(n31430), .Z(n38011) );
  XOR U37527 ( .A(n38026), .B(n38027), .Z(n31430) );
  XNOR U37528 ( .A(n31457), .B(n31428), .Z(n38027) );
  XNOR U37529 ( .A(q[0]), .B(DB[899]), .Z(n31428) );
  XOR U37530 ( .A(n38028), .B(n31449), .Z(n31457) );
  XOR U37531 ( .A(n38029), .B(n31437), .Z(n31449) );
  XNOR U37532 ( .A(q[15]), .B(DB[914]), .Z(n31437) );
  IV U37533 ( .A(n31436), .Z(n38029) );
  XNOR U37534 ( .A(n31434), .B(n38030), .Z(n31436) );
  XNOR U37535 ( .A(q[14]), .B(DB[913]), .Z(n38030) );
  XNOR U37536 ( .A(q[13]), .B(DB[912]), .Z(n31434) );
  IV U37537 ( .A(n31448), .Z(n38028) );
  XOR U37538 ( .A(n38031), .B(n38032), .Z(n31448) );
  XNOR U37539 ( .A(n31444), .B(n31446), .Z(n38032) );
  XNOR U37540 ( .A(q[9]), .B(DB[908]), .Z(n31446) );
  XNOR U37541 ( .A(q[12]), .B(DB[911]), .Z(n31444) );
  IV U37542 ( .A(n31443), .Z(n38031) );
  XNOR U37543 ( .A(n31441), .B(n38033), .Z(n31443) );
  XNOR U37544 ( .A(q[11]), .B(DB[910]), .Z(n38033) );
  XNOR U37545 ( .A(q[10]), .B(DB[909]), .Z(n31441) );
  IV U37546 ( .A(n31456), .Z(n38026) );
  XOR U37547 ( .A(n38034), .B(n38035), .Z(n31456) );
  XNOR U37548 ( .A(n31473), .B(n31454), .Z(n38035) );
  XNOR U37549 ( .A(q[1]), .B(DB[900]), .Z(n31454) );
  XOR U37550 ( .A(n38036), .B(n31462), .Z(n31473) );
  XNOR U37551 ( .A(q[8]), .B(DB[907]), .Z(n31462) );
  IV U37552 ( .A(n31461), .Z(n38036) );
  XNOR U37553 ( .A(n31459), .B(n38037), .Z(n31461) );
  XNOR U37554 ( .A(q[7]), .B(DB[906]), .Z(n38037) );
  XNOR U37555 ( .A(q[6]), .B(DB[905]), .Z(n31459) );
  IV U37556 ( .A(n31472), .Z(n38034) );
  XOR U37557 ( .A(n38038), .B(n38039), .Z(n31472) );
  XNOR U37558 ( .A(n31468), .B(n31470), .Z(n38039) );
  XNOR U37559 ( .A(q[2]), .B(DB[901]), .Z(n31470) );
  XNOR U37560 ( .A(q[5]), .B(DB[904]), .Z(n31468) );
  IV U37561 ( .A(n31467), .Z(n38038) );
  XNOR U37562 ( .A(n31465), .B(n38040), .Z(n31467) );
  XNOR U37563 ( .A(q[4]), .B(DB[903]), .Z(n38040) );
  XNOR U37564 ( .A(q[3]), .B(DB[902]), .Z(n31465) );
  XOR U37565 ( .A(n38041), .B(n31234), .Z(n31085) );
  XOR U37566 ( .A(n38042), .B(n31210), .Z(n31234) );
  XOR U37567 ( .A(n38043), .B(n31202), .Z(n31210) );
  XOR U37568 ( .A(n38044), .B(n31191), .Z(n31202) );
  XNOR U37569 ( .A(q[30]), .B(DB[960]), .Z(n31191) );
  IV U37570 ( .A(n31190), .Z(n38044) );
  XNOR U37571 ( .A(n31188), .B(n38045), .Z(n31190) );
  XNOR U37572 ( .A(q[29]), .B(DB[959]), .Z(n38045) );
  XNOR U37573 ( .A(q[28]), .B(DB[958]), .Z(n31188) );
  IV U37574 ( .A(n31201), .Z(n38043) );
  XOR U37575 ( .A(n38046), .B(n38047), .Z(n31201) );
  XNOR U37576 ( .A(n31197), .B(n31199), .Z(n38047) );
  XNOR U37577 ( .A(q[24]), .B(DB[954]), .Z(n31199) );
  XNOR U37578 ( .A(q[27]), .B(DB[957]), .Z(n31197) );
  IV U37579 ( .A(n31196), .Z(n38046) );
  XNOR U37580 ( .A(n31194), .B(n38048), .Z(n31196) );
  XNOR U37581 ( .A(q[26]), .B(DB[956]), .Z(n38048) );
  XNOR U37582 ( .A(q[25]), .B(DB[955]), .Z(n31194) );
  IV U37583 ( .A(n31209), .Z(n38042) );
  XOR U37584 ( .A(n38049), .B(n38050), .Z(n31209) );
  XNOR U37585 ( .A(n31226), .B(n31207), .Z(n38050) );
  XNOR U37586 ( .A(q[16]), .B(DB[946]), .Z(n31207) );
  XOR U37587 ( .A(n38051), .B(n31215), .Z(n31226) );
  XNOR U37588 ( .A(q[23]), .B(DB[953]), .Z(n31215) );
  IV U37589 ( .A(n31214), .Z(n38051) );
  XNOR U37590 ( .A(n31212), .B(n38052), .Z(n31214) );
  XNOR U37591 ( .A(q[22]), .B(DB[952]), .Z(n38052) );
  XNOR U37592 ( .A(q[21]), .B(DB[951]), .Z(n31212) );
  IV U37593 ( .A(n31225), .Z(n38049) );
  XOR U37594 ( .A(n38053), .B(n38054), .Z(n31225) );
  XNOR U37595 ( .A(n31221), .B(n31223), .Z(n38054) );
  XNOR U37596 ( .A(q[17]), .B(DB[947]), .Z(n31223) );
  XNOR U37597 ( .A(q[20]), .B(DB[950]), .Z(n31221) );
  IV U37598 ( .A(n31220), .Z(n38053) );
  XNOR U37599 ( .A(n31218), .B(n38055), .Z(n31220) );
  XNOR U37600 ( .A(q[19]), .B(DB[949]), .Z(n38055) );
  XNOR U37601 ( .A(q[18]), .B(DB[948]), .Z(n31218) );
  IV U37602 ( .A(n31233), .Z(n38041) );
  XOR U37603 ( .A(n38056), .B(n38057), .Z(n31233) );
  XNOR U37604 ( .A(n31260), .B(n31231), .Z(n38057) );
  XNOR U37605 ( .A(q[0]), .B(DB[930]), .Z(n31231) );
  XOR U37606 ( .A(n38058), .B(n31252), .Z(n31260) );
  XOR U37607 ( .A(n38059), .B(n31240), .Z(n31252) );
  XNOR U37608 ( .A(q[15]), .B(DB[945]), .Z(n31240) );
  IV U37609 ( .A(n31239), .Z(n38059) );
  XNOR U37610 ( .A(n31237), .B(n38060), .Z(n31239) );
  XNOR U37611 ( .A(q[14]), .B(DB[944]), .Z(n38060) );
  XNOR U37612 ( .A(q[13]), .B(DB[943]), .Z(n31237) );
  IV U37613 ( .A(n31251), .Z(n38058) );
  XOR U37614 ( .A(n38061), .B(n38062), .Z(n31251) );
  XNOR U37615 ( .A(n31247), .B(n31249), .Z(n38062) );
  XNOR U37616 ( .A(q[9]), .B(DB[939]), .Z(n31249) );
  XNOR U37617 ( .A(q[12]), .B(DB[942]), .Z(n31247) );
  IV U37618 ( .A(n31246), .Z(n38061) );
  XNOR U37619 ( .A(n31244), .B(n38063), .Z(n31246) );
  XNOR U37620 ( .A(q[11]), .B(DB[941]), .Z(n38063) );
  XNOR U37621 ( .A(q[10]), .B(DB[940]), .Z(n31244) );
  IV U37622 ( .A(n31259), .Z(n38056) );
  XOR U37623 ( .A(n38064), .B(n38065), .Z(n31259) );
  XNOR U37624 ( .A(n31276), .B(n31257), .Z(n38065) );
  XNOR U37625 ( .A(q[1]), .B(DB[931]), .Z(n31257) );
  XOR U37626 ( .A(n38066), .B(n31265), .Z(n31276) );
  XNOR U37627 ( .A(q[8]), .B(DB[938]), .Z(n31265) );
  IV U37628 ( .A(n31264), .Z(n38066) );
  XNOR U37629 ( .A(n31262), .B(n38067), .Z(n31264) );
  XNOR U37630 ( .A(q[7]), .B(DB[937]), .Z(n38067) );
  XNOR U37631 ( .A(q[6]), .B(DB[936]), .Z(n31262) );
  IV U37632 ( .A(n31275), .Z(n38064) );
  XOR U37633 ( .A(n38068), .B(n38069), .Z(n31275) );
  XNOR U37634 ( .A(n31271), .B(n31273), .Z(n38069) );
  XNOR U37635 ( .A(q[2]), .B(DB[932]), .Z(n31273) );
  XNOR U37636 ( .A(q[5]), .B(DB[935]), .Z(n31271) );
  IV U37637 ( .A(n31270), .Z(n38068) );
  XNOR U37638 ( .A(n31268), .B(n38070), .Z(n31270) );
  XNOR U37639 ( .A(q[4]), .B(DB[934]), .Z(n38070) );
  XNOR U37640 ( .A(q[3]), .B(DB[933]), .Z(n31268) );
  XOR U37641 ( .A(n38071), .B(n31037), .Z(n30888) );
  XOR U37642 ( .A(n38072), .B(n31013), .Z(n31037) );
  XOR U37643 ( .A(n38073), .B(n31005), .Z(n31013) );
  XOR U37644 ( .A(n38074), .B(n30994), .Z(n31005) );
  XNOR U37645 ( .A(q[30]), .B(DB[991]), .Z(n30994) );
  IV U37646 ( .A(n30993), .Z(n38074) );
  XNOR U37647 ( .A(n30991), .B(n38075), .Z(n30993) );
  XNOR U37648 ( .A(q[29]), .B(DB[990]), .Z(n38075) );
  XNOR U37649 ( .A(q[28]), .B(DB[989]), .Z(n30991) );
  IV U37650 ( .A(n31004), .Z(n38073) );
  XOR U37651 ( .A(n38076), .B(n38077), .Z(n31004) );
  XNOR U37652 ( .A(n31000), .B(n31002), .Z(n38077) );
  XNOR U37653 ( .A(q[24]), .B(DB[985]), .Z(n31002) );
  XNOR U37654 ( .A(q[27]), .B(DB[988]), .Z(n31000) );
  IV U37655 ( .A(n30999), .Z(n38076) );
  XNOR U37656 ( .A(n30997), .B(n38078), .Z(n30999) );
  XNOR U37657 ( .A(q[26]), .B(DB[987]), .Z(n38078) );
  XNOR U37658 ( .A(q[25]), .B(DB[986]), .Z(n30997) );
  IV U37659 ( .A(n31012), .Z(n38072) );
  XOR U37660 ( .A(n38079), .B(n38080), .Z(n31012) );
  XNOR U37661 ( .A(n31029), .B(n31010), .Z(n38080) );
  XNOR U37662 ( .A(q[16]), .B(DB[977]), .Z(n31010) );
  XOR U37663 ( .A(n38081), .B(n31018), .Z(n31029) );
  XNOR U37664 ( .A(q[23]), .B(DB[984]), .Z(n31018) );
  IV U37665 ( .A(n31017), .Z(n38081) );
  XNOR U37666 ( .A(n31015), .B(n38082), .Z(n31017) );
  XNOR U37667 ( .A(q[22]), .B(DB[983]), .Z(n38082) );
  XNOR U37668 ( .A(q[21]), .B(DB[982]), .Z(n31015) );
  IV U37669 ( .A(n31028), .Z(n38079) );
  XOR U37670 ( .A(n38083), .B(n38084), .Z(n31028) );
  XNOR U37671 ( .A(n31024), .B(n31026), .Z(n38084) );
  XNOR U37672 ( .A(q[17]), .B(DB[978]), .Z(n31026) );
  XNOR U37673 ( .A(q[20]), .B(DB[981]), .Z(n31024) );
  IV U37674 ( .A(n31023), .Z(n38083) );
  XNOR U37675 ( .A(n31021), .B(n38085), .Z(n31023) );
  XNOR U37676 ( .A(q[19]), .B(DB[980]), .Z(n38085) );
  XNOR U37677 ( .A(q[18]), .B(DB[979]), .Z(n31021) );
  IV U37678 ( .A(n31036), .Z(n38071) );
  XOR U37679 ( .A(n38086), .B(n38087), .Z(n31036) );
  XNOR U37680 ( .A(n31063), .B(n31034), .Z(n38087) );
  XNOR U37681 ( .A(q[0]), .B(DB[961]), .Z(n31034) );
  XOR U37682 ( .A(n38088), .B(n31055), .Z(n31063) );
  XOR U37683 ( .A(n38089), .B(n31043), .Z(n31055) );
  XNOR U37684 ( .A(q[15]), .B(DB[976]), .Z(n31043) );
  IV U37685 ( .A(n31042), .Z(n38089) );
  XNOR U37686 ( .A(n31040), .B(n38090), .Z(n31042) );
  XNOR U37687 ( .A(q[14]), .B(DB[975]), .Z(n38090) );
  XNOR U37688 ( .A(q[13]), .B(DB[974]), .Z(n31040) );
  IV U37689 ( .A(n31054), .Z(n38088) );
  XOR U37690 ( .A(n38091), .B(n38092), .Z(n31054) );
  XNOR U37691 ( .A(n31050), .B(n31052), .Z(n38092) );
  XNOR U37692 ( .A(q[9]), .B(DB[970]), .Z(n31052) );
  XNOR U37693 ( .A(q[12]), .B(DB[973]), .Z(n31050) );
  IV U37694 ( .A(n31049), .Z(n38091) );
  XNOR U37695 ( .A(n31047), .B(n38093), .Z(n31049) );
  XNOR U37696 ( .A(q[11]), .B(DB[972]), .Z(n38093) );
  XNOR U37697 ( .A(q[10]), .B(DB[971]), .Z(n31047) );
  IV U37698 ( .A(n31062), .Z(n38086) );
  XOR U37699 ( .A(n38094), .B(n38095), .Z(n31062) );
  XNOR U37700 ( .A(n31079), .B(n31060), .Z(n38095) );
  XNOR U37701 ( .A(q[1]), .B(DB[962]), .Z(n31060) );
  XOR U37702 ( .A(n38096), .B(n31068), .Z(n31079) );
  XNOR U37703 ( .A(q[8]), .B(DB[969]), .Z(n31068) );
  IV U37704 ( .A(n31067), .Z(n38096) );
  XNOR U37705 ( .A(n31065), .B(n38097), .Z(n31067) );
  XNOR U37706 ( .A(q[7]), .B(DB[968]), .Z(n38097) );
  XNOR U37707 ( .A(q[6]), .B(DB[967]), .Z(n31065) );
  IV U37708 ( .A(n31078), .Z(n38094) );
  XOR U37709 ( .A(n38098), .B(n38099), .Z(n31078) );
  XNOR U37710 ( .A(n31074), .B(n31076), .Z(n38099) );
  XNOR U37711 ( .A(q[2]), .B(DB[963]), .Z(n31076) );
  XNOR U37712 ( .A(q[5]), .B(DB[966]), .Z(n31074) );
  IV U37713 ( .A(n31073), .Z(n38098) );
  XNOR U37714 ( .A(n31071), .B(n38100), .Z(n31073) );
  XNOR U37715 ( .A(q[4]), .B(DB[965]), .Z(n38100) );
  XNOR U37716 ( .A(q[3]), .B(DB[964]), .Z(n31071) );
  XOR U37717 ( .A(n38101), .B(n30840), .Z(n30691) );
  XOR U37718 ( .A(n38102), .B(n30816), .Z(n30840) );
  XOR U37719 ( .A(n38103), .B(n30808), .Z(n30816) );
  XOR U37720 ( .A(n38104), .B(n30797), .Z(n30808) );
  XNOR U37721 ( .A(q[30]), .B(DB[1022]), .Z(n30797) );
  IV U37722 ( .A(n30796), .Z(n38104) );
  XNOR U37723 ( .A(n30794), .B(n38105), .Z(n30796) );
  XNOR U37724 ( .A(q[29]), .B(DB[1021]), .Z(n38105) );
  XNOR U37725 ( .A(q[28]), .B(DB[1020]), .Z(n30794) );
  IV U37726 ( .A(n30807), .Z(n38103) );
  XOR U37727 ( .A(n38106), .B(n38107), .Z(n30807) );
  XNOR U37728 ( .A(n30803), .B(n30805), .Z(n38107) );
  XNOR U37729 ( .A(q[24]), .B(DB[1016]), .Z(n30805) );
  XNOR U37730 ( .A(q[27]), .B(DB[1019]), .Z(n30803) );
  IV U37731 ( .A(n30802), .Z(n38106) );
  XNOR U37732 ( .A(n30800), .B(n38108), .Z(n30802) );
  XNOR U37733 ( .A(q[26]), .B(DB[1018]), .Z(n38108) );
  XNOR U37734 ( .A(q[25]), .B(DB[1017]), .Z(n30800) );
  IV U37735 ( .A(n30815), .Z(n38102) );
  XOR U37736 ( .A(n38109), .B(n38110), .Z(n30815) );
  XNOR U37737 ( .A(n30832), .B(n30813), .Z(n38110) );
  XNOR U37738 ( .A(q[16]), .B(DB[1008]), .Z(n30813) );
  XOR U37739 ( .A(n38111), .B(n30821), .Z(n30832) );
  XNOR U37740 ( .A(q[23]), .B(DB[1015]), .Z(n30821) );
  IV U37741 ( .A(n30820), .Z(n38111) );
  XNOR U37742 ( .A(n30818), .B(n38112), .Z(n30820) );
  XNOR U37743 ( .A(q[22]), .B(DB[1014]), .Z(n38112) );
  XNOR U37744 ( .A(q[21]), .B(DB[1013]), .Z(n30818) );
  IV U37745 ( .A(n30831), .Z(n38109) );
  XOR U37746 ( .A(n38113), .B(n38114), .Z(n30831) );
  XNOR U37747 ( .A(n30827), .B(n30829), .Z(n38114) );
  XNOR U37748 ( .A(q[17]), .B(DB[1009]), .Z(n30829) );
  XNOR U37749 ( .A(q[20]), .B(DB[1012]), .Z(n30827) );
  IV U37750 ( .A(n30826), .Z(n38113) );
  XNOR U37751 ( .A(n30824), .B(n38115), .Z(n30826) );
  XNOR U37752 ( .A(q[19]), .B(DB[1011]), .Z(n38115) );
  XNOR U37753 ( .A(q[18]), .B(DB[1010]), .Z(n30824) );
  IV U37754 ( .A(n30839), .Z(n38101) );
  XOR U37755 ( .A(n38116), .B(n38117), .Z(n30839) );
  XNOR U37756 ( .A(n30866), .B(n30837), .Z(n38117) );
  XNOR U37757 ( .A(q[0]), .B(DB[992]), .Z(n30837) );
  XOR U37758 ( .A(n38118), .B(n30858), .Z(n30866) );
  XOR U37759 ( .A(n38119), .B(n30846), .Z(n30858) );
  XNOR U37760 ( .A(q[15]), .B(DB[1007]), .Z(n30846) );
  IV U37761 ( .A(n30845), .Z(n38119) );
  XNOR U37762 ( .A(n30843), .B(n38120), .Z(n30845) );
  XNOR U37763 ( .A(q[14]), .B(DB[1006]), .Z(n38120) );
  XNOR U37764 ( .A(q[13]), .B(DB[1005]), .Z(n30843) );
  IV U37765 ( .A(n30857), .Z(n38118) );
  XOR U37766 ( .A(n38121), .B(n38122), .Z(n30857) );
  XNOR U37767 ( .A(n30853), .B(n30855), .Z(n38122) );
  XNOR U37768 ( .A(q[9]), .B(DB[1001]), .Z(n30855) );
  XNOR U37769 ( .A(q[12]), .B(DB[1004]), .Z(n30853) );
  IV U37770 ( .A(n30852), .Z(n38121) );
  XNOR U37771 ( .A(n30850), .B(n38123), .Z(n30852) );
  XNOR U37772 ( .A(q[11]), .B(DB[1003]), .Z(n38123) );
  XNOR U37773 ( .A(q[10]), .B(DB[1002]), .Z(n30850) );
  IV U37774 ( .A(n30865), .Z(n38116) );
  XOR U37775 ( .A(n38124), .B(n38125), .Z(n30865) );
  XNOR U37776 ( .A(n30882), .B(n30863), .Z(n38125) );
  XNOR U37777 ( .A(q[1]), .B(DB[993]), .Z(n30863) );
  XOR U37778 ( .A(n38126), .B(n30871), .Z(n30882) );
  XNOR U37779 ( .A(q[8]), .B(DB[1000]), .Z(n30871) );
  IV U37780 ( .A(n30870), .Z(n38126) );
  XNOR U37781 ( .A(n30868), .B(n38127), .Z(n30870) );
  XNOR U37782 ( .A(q[7]), .B(DB[999]), .Z(n38127) );
  XNOR U37783 ( .A(q[6]), .B(DB[998]), .Z(n30868) );
  IV U37784 ( .A(n30881), .Z(n38124) );
  XOR U37785 ( .A(n38128), .B(n38129), .Z(n30881) );
  XNOR U37786 ( .A(n30877), .B(n30879), .Z(n38129) );
  XNOR U37787 ( .A(q[2]), .B(DB[994]), .Z(n30879) );
  XNOR U37788 ( .A(q[5]), .B(DB[997]), .Z(n30877) );
  IV U37789 ( .A(n30876), .Z(n38128) );
  XNOR U37790 ( .A(n30874), .B(n38130), .Z(n30876) );
  XNOR U37791 ( .A(q[4]), .B(DB[996]), .Z(n38130) );
  XNOR U37792 ( .A(q[3]), .B(DB[995]), .Z(n30874) );
  XOR U37793 ( .A(n38131), .B(n30643), .Z(n30494) );
  XOR U37794 ( .A(n38132), .B(n30619), .Z(n30643) );
  XOR U37795 ( .A(n38133), .B(n30611), .Z(n30619) );
  XOR U37796 ( .A(n38134), .B(n30600), .Z(n30611) );
  XNOR U37797 ( .A(q[30]), .B(DB[1053]), .Z(n30600) );
  IV U37798 ( .A(n30599), .Z(n38134) );
  XNOR U37799 ( .A(n30597), .B(n38135), .Z(n30599) );
  XNOR U37800 ( .A(q[29]), .B(DB[1052]), .Z(n38135) );
  XNOR U37801 ( .A(q[28]), .B(DB[1051]), .Z(n30597) );
  IV U37802 ( .A(n30610), .Z(n38133) );
  XOR U37803 ( .A(n38136), .B(n38137), .Z(n30610) );
  XNOR U37804 ( .A(n30606), .B(n30608), .Z(n38137) );
  XNOR U37805 ( .A(q[24]), .B(DB[1047]), .Z(n30608) );
  XNOR U37806 ( .A(q[27]), .B(DB[1050]), .Z(n30606) );
  IV U37807 ( .A(n30605), .Z(n38136) );
  XNOR U37808 ( .A(n30603), .B(n38138), .Z(n30605) );
  XNOR U37809 ( .A(q[26]), .B(DB[1049]), .Z(n38138) );
  XNOR U37810 ( .A(q[25]), .B(DB[1048]), .Z(n30603) );
  IV U37811 ( .A(n30618), .Z(n38132) );
  XOR U37812 ( .A(n38139), .B(n38140), .Z(n30618) );
  XNOR U37813 ( .A(n30635), .B(n30616), .Z(n38140) );
  XNOR U37814 ( .A(q[16]), .B(DB[1039]), .Z(n30616) );
  XOR U37815 ( .A(n38141), .B(n30624), .Z(n30635) );
  XNOR U37816 ( .A(q[23]), .B(DB[1046]), .Z(n30624) );
  IV U37817 ( .A(n30623), .Z(n38141) );
  XNOR U37818 ( .A(n30621), .B(n38142), .Z(n30623) );
  XNOR U37819 ( .A(q[22]), .B(DB[1045]), .Z(n38142) );
  XNOR U37820 ( .A(q[21]), .B(DB[1044]), .Z(n30621) );
  IV U37821 ( .A(n30634), .Z(n38139) );
  XOR U37822 ( .A(n38143), .B(n38144), .Z(n30634) );
  XNOR U37823 ( .A(n30630), .B(n30632), .Z(n38144) );
  XNOR U37824 ( .A(q[17]), .B(DB[1040]), .Z(n30632) );
  XNOR U37825 ( .A(q[20]), .B(DB[1043]), .Z(n30630) );
  IV U37826 ( .A(n30629), .Z(n38143) );
  XNOR U37827 ( .A(n30627), .B(n38145), .Z(n30629) );
  XNOR U37828 ( .A(q[19]), .B(DB[1042]), .Z(n38145) );
  XNOR U37829 ( .A(q[18]), .B(DB[1041]), .Z(n30627) );
  IV U37830 ( .A(n30642), .Z(n38131) );
  XOR U37831 ( .A(n38146), .B(n38147), .Z(n30642) );
  XNOR U37832 ( .A(n30669), .B(n30640), .Z(n38147) );
  XNOR U37833 ( .A(q[0]), .B(DB[1023]), .Z(n30640) );
  XOR U37834 ( .A(n38148), .B(n30661), .Z(n30669) );
  XOR U37835 ( .A(n38149), .B(n30649), .Z(n30661) );
  XNOR U37836 ( .A(q[15]), .B(DB[1038]), .Z(n30649) );
  IV U37837 ( .A(n30648), .Z(n38149) );
  XNOR U37838 ( .A(n30646), .B(n38150), .Z(n30648) );
  XNOR U37839 ( .A(q[14]), .B(DB[1037]), .Z(n38150) );
  XNOR U37840 ( .A(q[13]), .B(DB[1036]), .Z(n30646) );
  IV U37841 ( .A(n30660), .Z(n38148) );
  XOR U37842 ( .A(n38151), .B(n38152), .Z(n30660) );
  XNOR U37843 ( .A(n30656), .B(n30658), .Z(n38152) );
  XNOR U37844 ( .A(q[9]), .B(DB[1032]), .Z(n30658) );
  XNOR U37845 ( .A(q[12]), .B(DB[1035]), .Z(n30656) );
  IV U37846 ( .A(n30655), .Z(n38151) );
  XNOR U37847 ( .A(n30653), .B(n38153), .Z(n30655) );
  XNOR U37848 ( .A(q[11]), .B(DB[1034]), .Z(n38153) );
  XNOR U37849 ( .A(q[10]), .B(DB[1033]), .Z(n30653) );
  IV U37850 ( .A(n30668), .Z(n38146) );
  XOR U37851 ( .A(n38154), .B(n38155), .Z(n30668) );
  XNOR U37852 ( .A(n30685), .B(n30666), .Z(n38155) );
  XNOR U37853 ( .A(q[1]), .B(DB[1024]), .Z(n30666) );
  XOR U37854 ( .A(n38156), .B(n30674), .Z(n30685) );
  XNOR U37855 ( .A(q[8]), .B(DB[1031]), .Z(n30674) );
  IV U37856 ( .A(n30673), .Z(n38156) );
  XNOR U37857 ( .A(n30671), .B(n38157), .Z(n30673) );
  XNOR U37858 ( .A(q[7]), .B(DB[1030]), .Z(n38157) );
  XNOR U37859 ( .A(q[6]), .B(DB[1029]), .Z(n30671) );
  IV U37860 ( .A(n30684), .Z(n38154) );
  XOR U37861 ( .A(n38158), .B(n38159), .Z(n30684) );
  XNOR U37862 ( .A(n30680), .B(n30682), .Z(n38159) );
  XNOR U37863 ( .A(q[2]), .B(DB[1025]), .Z(n30682) );
  XNOR U37864 ( .A(q[5]), .B(DB[1028]), .Z(n30680) );
  IV U37865 ( .A(n30679), .Z(n38158) );
  XNOR U37866 ( .A(n30677), .B(n38160), .Z(n30679) );
  XNOR U37867 ( .A(q[4]), .B(DB[1027]), .Z(n38160) );
  XNOR U37868 ( .A(q[3]), .B(DB[1026]), .Z(n30677) );
  XOR U37869 ( .A(n38161), .B(n30446), .Z(n30297) );
  XOR U37870 ( .A(n38162), .B(n30422), .Z(n30446) );
  XOR U37871 ( .A(n38163), .B(n30414), .Z(n30422) );
  XOR U37872 ( .A(n38164), .B(n30403), .Z(n30414) );
  XNOR U37873 ( .A(q[30]), .B(DB[1084]), .Z(n30403) );
  IV U37874 ( .A(n30402), .Z(n38164) );
  XNOR U37875 ( .A(n30400), .B(n38165), .Z(n30402) );
  XNOR U37876 ( .A(q[29]), .B(DB[1083]), .Z(n38165) );
  XNOR U37877 ( .A(q[28]), .B(DB[1082]), .Z(n30400) );
  IV U37878 ( .A(n30413), .Z(n38163) );
  XOR U37879 ( .A(n38166), .B(n38167), .Z(n30413) );
  XNOR U37880 ( .A(n30409), .B(n30411), .Z(n38167) );
  XNOR U37881 ( .A(q[24]), .B(DB[1078]), .Z(n30411) );
  XNOR U37882 ( .A(q[27]), .B(DB[1081]), .Z(n30409) );
  IV U37883 ( .A(n30408), .Z(n38166) );
  XNOR U37884 ( .A(n30406), .B(n38168), .Z(n30408) );
  XNOR U37885 ( .A(q[26]), .B(DB[1080]), .Z(n38168) );
  XNOR U37886 ( .A(q[25]), .B(DB[1079]), .Z(n30406) );
  IV U37887 ( .A(n30421), .Z(n38162) );
  XOR U37888 ( .A(n38169), .B(n38170), .Z(n30421) );
  XNOR U37889 ( .A(n30438), .B(n30419), .Z(n38170) );
  XNOR U37890 ( .A(q[16]), .B(DB[1070]), .Z(n30419) );
  XOR U37891 ( .A(n38171), .B(n30427), .Z(n30438) );
  XNOR U37892 ( .A(q[23]), .B(DB[1077]), .Z(n30427) );
  IV U37893 ( .A(n30426), .Z(n38171) );
  XNOR U37894 ( .A(n30424), .B(n38172), .Z(n30426) );
  XNOR U37895 ( .A(q[22]), .B(DB[1076]), .Z(n38172) );
  XNOR U37896 ( .A(q[21]), .B(DB[1075]), .Z(n30424) );
  IV U37897 ( .A(n30437), .Z(n38169) );
  XOR U37898 ( .A(n38173), .B(n38174), .Z(n30437) );
  XNOR U37899 ( .A(n30433), .B(n30435), .Z(n38174) );
  XNOR U37900 ( .A(q[17]), .B(DB[1071]), .Z(n30435) );
  XNOR U37901 ( .A(q[20]), .B(DB[1074]), .Z(n30433) );
  IV U37902 ( .A(n30432), .Z(n38173) );
  XNOR U37903 ( .A(n30430), .B(n38175), .Z(n30432) );
  XNOR U37904 ( .A(q[19]), .B(DB[1073]), .Z(n38175) );
  XNOR U37905 ( .A(q[18]), .B(DB[1072]), .Z(n30430) );
  IV U37906 ( .A(n30445), .Z(n38161) );
  XOR U37907 ( .A(n38176), .B(n38177), .Z(n30445) );
  XNOR U37908 ( .A(n30472), .B(n30443), .Z(n38177) );
  XNOR U37909 ( .A(q[0]), .B(DB[1054]), .Z(n30443) );
  XOR U37910 ( .A(n38178), .B(n30464), .Z(n30472) );
  XOR U37911 ( .A(n38179), .B(n30452), .Z(n30464) );
  XNOR U37912 ( .A(q[15]), .B(DB[1069]), .Z(n30452) );
  IV U37913 ( .A(n30451), .Z(n38179) );
  XNOR U37914 ( .A(n30449), .B(n38180), .Z(n30451) );
  XNOR U37915 ( .A(q[14]), .B(DB[1068]), .Z(n38180) );
  XNOR U37916 ( .A(q[13]), .B(DB[1067]), .Z(n30449) );
  IV U37917 ( .A(n30463), .Z(n38178) );
  XOR U37918 ( .A(n38181), .B(n38182), .Z(n30463) );
  XNOR U37919 ( .A(n30459), .B(n30461), .Z(n38182) );
  XNOR U37920 ( .A(q[9]), .B(DB[1063]), .Z(n30461) );
  XNOR U37921 ( .A(q[12]), .B(DB[1066]), .Z(n30459) );
  IV U37922 ( .A(n30458), .Z(n38181) );
  XNOR U37923 ( .A(n30456), .B(n38183), .Z(n30458) );
  XNOR U37924 ( .A(q[11]), .B(DB[1065]), .Z(n38183) );
  XNOR U37925 ( .A(q[10]), .B(DB[1064]), .Z(n30456) );
  IV U37926 ( .A(n30471), .Z(n38176) );
  XOR U37927 ( .A(n38184), .B(n38185), .Z(n30471) );
  XNOR U37928 ( .A(n30488), .B(n30469), .Z(n38185) );
  XNOR U37929 ( .A(q[1]), .B(DB[1055]), .Z(n30469) );
  XOR U37930 ( .A(n38186), .B(n30477), .Z(n30488) );
  XNOR U37931 ( .A(q[8]), .B(DB[1062]), .Z(n30477) );
  IV U37932 ( .A(n30476), .Z(n38186) );
  XNOR U37933 ( .A(n30474), .B(n38187), .Z(n30476) );
  XNOR U37934 ( .A(q[7]), .B(DB[1061]), .Z(n38187) );
  XNOR U37935 ( .A(q[6]), .B(DB[1060]), .Z(n30474) );
  IV U37936 ( .A(n30487), .Z(n38184) );
  XOR U37937 ( .A(n38188), .B(n38189), .Z(n30487) );
  XNOR U37938 ( .A(n30483), .B(n30485), .Z(n38189) );
  XNOR U37939 ( .A(q[2]), .B(DB[1056]), .Z(n30485) );
  XNOR U37940 ( .A(q[5]), .B(DB[1059]), .Z(n30483) );
  IV U37941 ( .A(n30482), .Z(n38188) );
  XNOR U37942 ( .A(n30480), .B(n38190), .Z(n30482) );
  XNOR U37943 ( .A(q[4]), .B(DB[1058]), .Z(n38190) );
  XNOR U37944 ( .A(q[3]), .B(DB[1057]), .Z(n30480) );
  XOR U37945 ( .A(n38191), .B(n30249), .Z(n30100) );
  XOR U37946 ( .A(n38192), .B(n30225), .Z(n30249) );
  XOR U37947 ( .A(n38193), .B(n30217), .Z(n30225) );
  XOR U37948 ( .A(n38194), .B(n30206), .Z(n30217) );
  XNOR U37949 ( .A(q[30]), .B(DB[1115]), .Z(n30206) );
  IV U37950 ( .A(n30205), .Z(n38194) );
  XNOR U37951 ( .A(n30203), .B(n38195), .Z(n30205) );
  XNOR U37952 ( .A(q[29]), .B(DB[1114]), .Z(n38195) );
  XNOR U37953 ( .A(q[28]), .B(DB[1113]), .Z(n30203) );
  IV U37954 ( .A(n30216), .Z(n38193) );
  XOR U37955 ( .A(n38196), .B(n38197), .Z(n30216) );
  XNOR U37956 ( .A(n30212), .B(n30214), .Z(n38197) );
  XNOR U37957 ( .A(q[24]), .B(DB[1109]), .Z(n30214) );
  XNOR U37958 ( .A(q[27]), .B(DB[1112]), .Z(n30212) );
  IV U37959 ( .A(n30211), .Z(n38196) );
  XNOR U37960 ( .A(n30209), .B(n38198), .Z(n30211) );
  XNOR U37961 ( .A(q[26]), .B(DB[1111]), .Z(n38198) );
  XNOR U37962 ( .A(q[25]), .B(DB[1110]), .Z(n30209) );
  IV U37963 ( .A(n30224), .Z(n38192) );
  XOR U37964 ( .A(n38199), .B(n38200), .Z(n30224) );
  XNOR U37965 ( .A(n30241), .B(n30222), .Z(n38200) );
  XNOR U37966 ( .A(q[16]), .B(DB[1101]), .Z(n30222) );
  XOR U37967 ( .A(n38201), .B(n30230), .Z(n30241) );
  XNOR U37968 ( .A(q[23]), .B(DB[1108]), .Z(n30230) );
  IV U37969 ( .A(n30229), .Z(n38201) );
  XNOR U37970 ( .A(n30227), .B(n38202), .Z(n30229) );
  XNOR U37971 ( .A(q[22]), .B(DB[1107]), .Z(n38202) );
  XNOR U37972 ( .A(q[21]), .B(DB[1106]), .Z(n30227) );
  IV U37973 ( .A(n30240), .Z(n38199) );
  XOR U37974 ( .A(n38203), .B(n38204), .Z(n30240) );
  XNOR U37975 ( .A(n30236), .B(n30238), .Z(n38204) );
  XNOR U37976 ( .A(q[17]), .B(DB[1102]), .Z(n30238) );
  XNOR U37977 ( .A(q[20]), .B(DB[1105]), .Z(n30236) );
  IV U37978 ( .A(n30235), .Z(n38203) );
  XNOR U37979 ( .A(n30233), .B(n38205), .Z(n30235) );
  XNOR U37980 ( .A(q[19]), .B(DB[1104]), .Z(n38205) );
  XNOR U37981 ( .A(q[18]), .B(DB[1103]), .Z(n30233) );
  IV U37982 ( .A(n30248), .Z(n38191) );
  XOR U37983 ( .A(n38206), .B(n38207), .Z(n30248) );
  XNOR U37984 ( .A(n30275), .B(n30246), .Z(n38207) );
  XNOR U37985 ( .A(q[0]), .B(DB[1085]), .Z(n30246) );
  XOR U37986 ( .A(n38208), .B(n30267), .Z(n30275) );
  XOR U37987 ( .A(n38209), .B(n30255), .Z(n30267) );
  XNOR U37988 ( .A(q[15]), .B(DB[1100]), .Z(n30255) );
  IV U37989 ( .A(n30254), .Z(n38209) );
  XNOR U37990 ( .A(n30252), .B(n38210), .Z(n30254) );
  XNOR U37991 ( .A(q[14]), .B(DB[1099]), .Z(n38210) );
  XNOR U37992 ( .A(q[13]), .B(DB[1098]), .Z(n30252) );
  IV U37993 ( .A(n30266), .Z(n38208) );
  XOR U37994 ( .A(n38211), .B(n38212), .Z(n30266) );
  XNOR U37995 ( .A(n30262), .B(n30264), .Z(n38212) );
  XNOR U37996 ( .A(q[9]), .B(DB[1094]), .Z(n30264) );
  XNOR U37997 ( .A(q[12]), .B(DB[1097]), .Z(n30262) );
  IV U37998 ( .A(n30261), .Z(n38211) );
  XNOR U37999 ( .A(n30259), .B(n38213), .Z(n30261) );
  XNOR U38000 ( .A(q[11]), .B(DB[1096]), .Z(n38213) );
  XNOR U38001 ( .A(q[10]), .B(DB[1095]), .Z(n30259) );
  IV U38002 ( .A(n30274), .Z(n38206) );
  XOR U38003 ( .A(n38214), .B(n38215), .Z(n30274) );
  XNOR U38004 ( .A(n30291), .B(n30272), .Z(n38215) );
  XNOR U38005 ( .A(q[1]), .B(DB[1086]), .Z(n30272) );
  XOR U38006 ( .A(n38216), .B(n30280), .Z(n30291) );
  XNOR U38007 ( .A(q[8]), .B(DB[1093]), .Z(n30280) );
  IV U38008 ( .A(n30279), .Z(n38216) );
  XNOR U38009 ( .A(n30277), .B(n38217), .Z(n30279) );
  XNOR U38010 ( .A(q[7]), .B(DB[1092]), .Z(n38217) );
  XNOR U38011 ( .A(q[6]), .B(DB[1091]), .Z(n30277) );
  IV U38012 ( .A(n30290), .Z(n38214) );
  XOR U38013 ( .A(n38218), .B(n38219), .Z(n30290) );
  XNOR U38014 ( .A(n30286), .B(n30288), .Z(n38219) );
  XNOR U38015 ( .A(q[2]), .B(DB[1087]), .Z(n30288) );
  XNOR U38016 ( .A(q[5]), .B(DB[1090]), .Z(n30286) );
  IV U38017 ( .A(n30285), .Z(n38218) );
  XNOR U38018 ( .A(n30283), .B(n38220), .Z(n30285) );
  XNOR U38019 ( .A(q[4]), .B(DB[1089]), .Z(n38220) );
  XNOR U38020 ( .A(q[3]), .B(DB[1088]), .Z(n30283) );
  XOR U38021 ( .A(n38221), .B(n30052), .Z(n29903) );
  XOR U38022 ( .A(n38222), .B(n30028), .Z(n30052) );
  XOR U38023 ( .A(n38223), .B(n30020), .Z(n30028) );
  XOR U38024 ( .A(n38224), .B(n30009), .Z(n30020) );
  XNOR U38025 ( .A(q[30]), .B(DB[1146]), .Z(n30009) );
  IV U38026 ( .A(n30008), .Z(n38224) );
  XNOR U38027 ( .A(n30006), .B(n38225), .Z(n30008) );
  XNOR U38028 ( .A(q[29]), .B(DB[1145]), .Z(n38225) );
  XNOR U38029 ( .A(q[28]), .B(DB[1144]), .Z(n30006) );
  IV U38030 ( .A(n30019), .Z(n38223) );
  XOR U38031 ( .A(n38226), .B(n38227), .Z(n30019) );
  XNOR U38032 ( .A(n30015), .B(n30017), .Z(n38227) );
  XNOR U38033 ( .A(q[24]), .B(DB[1140]), .Z(n30017) );
  XNOR U38034 ( .A(q[27]), .B(DB[1143]), .Z(n30015) );
  IV U38035 ( .A(n30014), .Z(n38226) );
  XNOR U38036 ( .A(n30012), .B(n38228), .Z(n30014) );
  XNOR U38037 ( .A(q[26]), .B(DB[1142]), .Z(n38228) );
  XNOR U38038 ( .A(q[25]), .B(DB[1141]), .Z(n30012) );
  IV U38039 ( .A(n30027), .Z(n38222) );
  XOR U38040 ( .A(n38229), .B(n38230), .Z(n30027) );
  XNOR U38041 ( .A(n30044), .B(n30025), .Z(n38230) );
  XNOR U38042 ( .A(q[16]), .B(DB[1132]), .Z(n30025) );
  XOR U38043 ( .A(n38231), .B(n30033), .Z(n30044) );
  XNOR U38044 ( .A(q[23]), .B(DB[1139]), .Z(n30033) );
  IV U38045 ( .A(n30032), .Z(n38231) );
  XNOR U38046 ( .A(n30030), .B(n38232), .Z(n30032) );
  XNOR U38047 ( .A(q[22]), .B(DB[1138]), .Z(n38232) );
  XNOR U38048 ( .A(q[21]), .B(DB[1137]), .Z(n30030) );
  IV U38049 ( .A(n30043), .Z(n38229) );
  XOR U38050 ( .A(n38233), .B(n38234), .Z(n30043) );
  XNOR U38051 ( .A(n30039), .B(n30041), .Z(n38234) );
  XNOR U38052 ( .A(q[17]), .B(DB[1133]), .Z(n30041) );
  XNOR U38053 ( .A(q[20]), .B(DB[1136]), .Z(n30039) );
  IV U38054 ( .A(n30038), .Z(n38233) );
  XNOR U38055 ( .A(n30036), .B(n38235), .Z(n30038) );
  XNOR U38056 ( .A(q[19]), .B(DB[1135]), .Z(n38235) );
  XNOR U38057 ( .A(q[18]), .B(DB[1134]), .Z(n30036) );
  IV U38058 ( .A(n30051), .Z(n38221) );
  XOR U38059 ( .A(n38236), .B(n38237), .Z(n30051) );
  XNOR U38060 ( .A(n30078), .B(n30049), .Z(n38237) );
  XNOR U38061 ( .A(q[0]), .B(DB[1116]), .Z(n30049) );
  XOR U38062 ( .A(n38238), .B(n30070), .Z(n30078) );
  XOR U38063 ( .A(n38239), .B(n30058), .Z(n30070) );
  XNOR U38064 ( .A(q[15]), .B(DB[1131]), .Z(n30058) );
  IV U38065 ( .A(n30057), .Z(n38239) );
  XNOR U38066 ( .A(n30055), .B(n38240), .Z(n30057) );
  XNOR U38067 ( .A(q[14]), .B(DB[1130]), .Z(n38240) );
  XNOR U38068 ( .A(q[13]), .B(DB[1129]), .Z(n30055) );
  IV U38069 ( .A(n30069), .Z(n38238) );
  XOR U38070 ( .A(n38241), .B(n38242), .Z(n30069) );
  XNOR U38071 ( .A(n30065), .B(n30067), .Z(n38242) );
  XNOR U38072 ( .A(q[9]), .B(DB[1125]), .Z(n30067) );
  XNOR U38073 ( .A(q[12]), .B(DB[1128]), .Z(n30065) );
  IV U38074 ( .A(n30064), .Z(n38241) );
  XNOR U38075 ( .A(n30062), .B(n38243), .Z(n30064) );
  XNOR U38076 ( .A(q[11]), .B(DB[1127]), .Z(n38243) );
  XNOR U38077 ( .A(q[10]), .B(DB[1126]), .Z(n30062) );
  IV U38078 ( .A(n30077), .Z(n38236) );
  XOR U38079 ( .A(n38244), .B(n38245), .Z(n30077) );
  XNOR U38080 ( .A(n30094), .B(n30075), .Z(n38245) );
  XNOR U38081 ( .A(q[1]), .B(DB[1117]), .Z(n30075) );
  XOR U38082 ( .A(n38246), .B(n30083), .Z(n30094) );
  XNOR U38083 ( .A(q[8]), .B(DB[1124]), .Z(n30083) );
  IV U38084 ( .A(n30082), .Z(n38246) );
  XNOR U38085 ( .A(n30080), .B(n38247), .Z(n30082) );
  XNOR U38086 ( .A(q[7]), .B(DB[1123]), .Z(n38247) );
  XNOR U38087 ( .A(q[6]), .B(DB[1122]), .Z(n30080) );
  IV U38088 ( .A(n30093), .Z(n38244) );
  XOR U38089 ( .A(n38248), .B(n38249), .Z(n30093) );
  XNOR U38090 ( .A(n30089), .B(n30091), .Z(n38249) );
  XNOR U38091 ( .A(q[2]), .B(DB[1118]), .Z(n30091) );
  XNOR U38092 ( .A(q[5]), .B(DB[1121]), .Z(n30089) );
  IV U38093 ( .A(n30088), .Z(n38248) );
  XNOR U38094 ( .A(n30086), .B(n38250), .Z(n30088) );
  XNOR U38095 ( .A(q[4]), .B(DB[1120]), .Z(n38250) );
  XNOR U38096 ( .A(q[3]), .B(DB[1119]), .Z(n30086) );
  XOR U38097 ( .A(n38251), .B(n29855), .Z(n29706) );
  XOR U38098 ( .A(n38252), .B(n29831), .Z(n29855) );
  XOR U38099 ( .A(n38253), .B(n29823), .Z(n29831) );
  XOR U38100 ( .A(n38254), .B(n29812), .Z(n29823) );
  XNOR U38101 ( .A(q[30]), .B(DB[1177]), .Z(n29812) );
  IV U38102 ( .A(n29811), .Z(n38254) );
  XNOR U38103 ( .A(n29809), .B(n38255), .Z(n29811) );
  XNOR U38104 ( .A(q[29]), .B(DB[1176]), .Z(n38255) );
  XNOR U38105 ( .A(q[28]), .B(DB[1175]), .Z(n29809) );
  IV U38106 ( .A(n29822), .Z(n38253) );
  XOR U38107 ( .A(n38256), .B(n38257), .Z(n29822) );
  XNOR U38108 ( .A(n29818), .B(n29820), .Z(n38257) );
  XNOR U38109 ( .A(q[24]), .B(DB[1171]), .Z(n29820) );
  XNOR U38110 ( .A(q[27]), .B(DB[1174]), .Z(n29818) );
  IV U38111 ( .A(n29817), .Z(n38256) );
  XNOR U38112 ( .A(n29815), .B(n38258), .Z(n29817) );
  XNOR U38113 ( .A(q[26]), .B(DB[1173]), .Z(n38258) );
  XNOR U38114 ( .A(q[25]), .B(DB[1172]), .Z(n29815) );
  IV U38115 ( .A(n29830), .Z(n38252) );
  XOR U38116 ( .A(n38259), .B(n38260), .Z(n29830) );
  XNOR U38117 ( .A(n29847), .B(n29828), .Z(n38260) );
  XNOR U38118 ( .A(q[16]), .B(DB[1163]), .Z(n29828) );
  XOR U38119 ( .A(n38261), .B(n29836), .Z(n29847) );
  XNOR U38120 ( .A(q[23]), .B(DB[1170]), .Z(n29836) );
  IV U38121 ( .A(n29835), .Z(n38261) );
  XNOR U38122 ( .A(n29833), .B(n38262), .Z(n29835) );
  XNOR U38123 ( .A(q[22]), .B(DB[1169]), .Z(n38262) );
  XNOR U38124 ( .A(q[21]), .B(DB[1168]), .Z(n29833) );
  IV U38125 ( .A(n29846), .Z(n38259) );
  XOR U38126 ( .A(n38263), .B(n38264), .Z(n29846) );
  XNOR U38127 ( .A(n29842), .B(n29844), .Z(n38264) );
  XNOR U38128 ( .A(q[17]), .B(DB[1164]), .Z(n29844) );
  XNOR U38129 ( .A(q[20]), .B(DB[1167]), .Z(n29842) );
  IV U38130 ( .A(n29841), .Z(n38263) );
  XNOR U38131 ( .A(n29839), .B(n38265), .Z(n29841) );
  XNOR U38132 ( .A(q[19]), .B(DB[1166]), .Z(n38265) );
  XNOR U38133 ( .A(q[18]), .B(DB[1165]), .Z(n29839) );
  IV U38134 ( .A(n29854), .Z(n38251) );
  XOR U38135 ( .A(n38266), .B(n38267), .Z(n29854) );
  XNOR U38136 ( .A(n29881), .B(n29852), .Z(n38267) );
  XNOR U38137 ( .A(q[0]), .B(DB[1147]), .Z(n29852) );
  XOR U38138 ( .A(n38268), .B(n29873), .Z(n29881) );
  XOR U38139 ( .A(n38269), .B(n29861), .Z(n29873) );
  XNOR U38140 ( .A(q[15]), .B(DB[1162]), .Z(n29861) );
  IV U38141 ( .A(n29860), .Z(n38269) );
  XNOR U38142 ( .A(n29858), .B(n38270), .Z(n29860) );
  XNOR U38143 ( .A(q[14]), .B(DB[1161]), .Z(n38270) );
  XNOR U38144 ( .A(q[13]), .B(DB[1160]), .Z(n29858) );
  IV U38145 ( .A(n29872), .Z(n38268) );
  XOR U38146 ( .A(n38271), .B(n38272), .Z(n29872) );
  XNOR U38147 ( .A(n29868), .B(n29870), .Z(n38272) );
  XNOR U38148 ( .A(q[9]), .B(DB[1156]), .Z(n29870) );
  XNOR U38149 ( .A(q[12]), .B(DB[1159]), .Z(n29868) );
  IV U38150 ( .A(n29867), .Z(n38271) );
  XNOR U38151 ( .A(n29865), .B(n38273), .Z(n29867) );
  XNOR U38152 ( .A(q[11]), .B(DB[1158]), .Z(n38273) );
  XNOR U38153 ( .A(q[10]), .B(DB[1157]), .Z(n29865) );
  IV U38154 ( .A(n29880), .Z(n38266) );
  XOR U38155 ( .A(n38274), .B(n38275), .Z(n29880) );
  XNOR U38156 ( .A(n29897), .B(n29878), .Z(n38275) );
  XNOR U38157 ( .A(q[1]), .B(DB[1148]), .Z(n29878) );
  XOR U38158 ( .A(n38276), .B(n29886), .Z(n29897) );
  XNOR U38159 ( .A(q[8]), .B(DB[1155]), .Z(n29886) );
  IV U38160 ( .A(n29885), .Z(n38276) );
  XNOR U38161 ( .A(n29883), .B(n38277), .Z(n29885) );
  XNOR U38162 ( .A(q[7]), .B(DB[1154]), .Z(n38277) );
  XNOR U38163 ( .A(q[6]), .B(DB[1153]), .Z(n29883) );
  IV U38164 ( .A(n29896), .Z(n38274) );
  XOR U38165 ( .A(n38278), .B(n38279), .Z(n29896) );
  XNOR U38166 ( .A(n29892), .B(n29894), .Z(n38279) );
  XNOR U38167 ( .A(q[2]), .B(DB[1149]), .Z(n29894) );
  XNOR U38168 ( .A(q[5]), .B(DB[1152]), .Z(n29892) );
  IV U38169 ( .A(n29891), .Z(n38278) );
  XNOR U38170 ( .A(n29889), .B(n38280), .Z(n29891) );
  XNOR U38171 ( .A(q[4]), .B(DB[1151]), .Z(n38280) );
  XNOR U38172 ( .A(q[3]), .B(DB[1150]), .Z(n29889) );
  XOR U38173 ( .A(n38281), .B(n29658), .Z(n29509) );
  XOR U38174 ( .A(n38282), .B(n29634), .Z(n29658) );
  XOR U38175 ( .A(n38283), .B(n29626), .Z(n29634) );
  XOR U38176 ( .A(n38284), .B(n29615), .Z(n29626) );
  XNOR U38177 ( .A(q[30]), .B(DB[1208]), .Z(n29615) );
  IV U38178 ( .A(n29614), .Z(n38284) );
  XNOR U38179 ( .A(n29612), .B(n38285), .Z(n29614) );
  XNOR U38180 ( .A(q[29]), .B(DB[1207]), .Z(n38285) );
  XNOR U38181 ( .A(q[28]), .B(DB[1206]), .Z(n29612) );
  IV U38182 ( .A(n29625), .Z(n38283) );
  XOR U38183 ( .A(n38286), .B(n38287), .Z(n29625) );
  XNOR U38184 ( .A(n29621), .B(n29623), .Z(n38287) );
  XNOR U38185 ( .A(q[24]), .B(DB[1202]), .Z(n29623) );
  XNOR U38186 ( .A(q[27]), .B(DB[1205]), .Z(n29621) );
  IV U38187 ( .A(n29620), .Z(n38286) );
  XNOR U38188 ( .A(n29618), .B(n38288), .Z(n29620) );
  XNOR U38189 ( .A(q[26]), .B(DB[1204]), .Z(n38288) );
  XNOR U38190 ( .A(q[25]), .B(DB[1203]), .Z(n29618) );
  IV U38191 ( .A(n29633), .Z(n38282) );
  XOR U38192 ( .A(n38289), .B(n38290), .Z(n29633) );
  XNOR U38193 ( .A(n29650), .B(n29631), .Z(n38290) );
  XNOR U38194 ( .A(q[16]), .B(DB[1194]), .Z(n29631) );
  XOR U38195 ( .A(n38291), .B(n29639), .Z(n29650) );
  XNOR U38196 ( .A(q[23]), .B(DB[1201]), .Z(n29639) );
  IV U38197 ( .A(n29638), .Z(n38291) );
  XNOR U38198 ( .A(n29636), .B(n38292), .Z(n29638) );
  XNOR U38199 ( .A(q[22]), .B(DB[1200]), .Z(n38292) );
  XNOR U38200 ( .A(q[21]), .B(DB[1199]), .Z(n29636) );
  IV U38201 ( .A(n29649), .Z(n38289) );
  XOR U38202 ( .A(n38293), .B(n38294), .Z(n29649) );
  XNOR U38203 ( .A(n29645), .B(n29647), .Z(n38294) );
  XNOR U38204 ( .A(q[17]), .B(DB[1195]), .Z(n29647) );
  XNOR U38205 ( .A(q[20]), .B(DB[1198]), .Z(n29645) );
  IV U38206 ( .A(n29644), .Z(n38293) );
  XNOR U38207 ( .A(n29642), .B(n38295), .Z(n29644) );
  XNOR U38208 ( .A(q[19]), .B(DB[1197]), .Z(n38295) );
  XNOR U38209 ( .A(q[18]), .B(DB[1196]), .Z(n29642) );
  IV U38210 ( .A(n29657), .Z(n38281) );
  XOR U38211 ( .A(n38296), .B(n38297), .Z(n29657) );
  XNOR U38212 ( .A(n29684), .B(n29655), .Z(n38297) );
  XNOR U38213 ( .A(q[0]), .B(DB[1178]), .Z(n29655) );
  XOR U38214 ( .A(n38298), .B(n29676), .Z(n29684) );
  XOR U38215 ( .A(n38299), .B(n29664), .Z(n29676) );
  XNOR U38216 ( .A(q[15]), .B(DB[1193]), .Z(n29664) );
  IV U38217 ( .A(n29663), .Z(n38299) );
  XNOR U38218 ( .A(n29661), .B(n38300), .Z(n29663) );
  XNOR U38219 ( .A(q[14]), .B(DB[1192]), .Z(n38300) );
  XNOR U38220 ( .A(q[13]), .B(DB[1191]), .Z(n29661) );
  IV U38221 ( .A(n29675), .Z(n38298) );
  XOR U38222 ( .A(n38301), .B(n38302), .Z(n29675) );
  XNOR U38223 ( .A(n29671), .B(n29673), .Z(n38302) );
  XNOR U38224 ( .A(q[9]), .B(DB[1187]), .Z(n29673) );
  XNOR U38225 ( .A(q[12]), .B(DB[1190]), .Z(n29671) );
  IV U38226 ( .A(n29670), .Z(n38301) );
  XNOR U38227 ( .A(n29668), .B(n38303), .Z(n29670) );
  XNOR U38228 ( .A(q[11]), .B(DB[1189]), .Z(n38303) );
  XNOR U38229 ( .A(q[10]), .B(DB[1188]), .Z(n29668) );
  IV U38230 ( .A(n29683), .Z(n38296) );
  XOR U38231 ( .A(n38304), .B(n38305), .Z(n29683) );
  XNOR U38232 ( .A(n29700), .B(n29681), .Z(n38305) );
  XNOR U38233 ( .A(q[1]), .B(DB[1179]), .Z(n29681) );
  XOR U38234 ( .A(n38306), .B(n29689), .Z(n29700) );
  XNOR U38235 ( .A(q[8]), .B(DB[1186]), .Z(n29689) );
  IV U38236 ( .A(n29688), .Z(n38306) );
  XNOR U38237 ( .A(n29686), .B(n38307), .Z(n29688) );
  XNOR U38238 ( .A(q[7]), .B(DB[1185]), .Z(n38307) );
  XNOR U38239 ( .A(q[6]), .B(DB[1184]), .Z(n29686) );
  IV U38240 ( .A(n29699), .Z(n38304) );
  XOR U38241 ( .A(n38308), .B(n38309), .Z(n29699) );
  XNOR U38242 ( .A(n29695), .B(n29697), .Z(n38309) );
  XNOR U38243 ( .A(q[2]), .B(DB[1180]), .Z(n29697) );
  XNOR U38244 ( .A(q[5]), .B(DB[1183]), .Z(n29695) );
  IV U38245 ( .A(n29694), .Z(n38308) );
  XNOR U38246 ( .A(n29692), .B(n38310), .Z(n29694) );
  XNOR U38247 ( .A(q[4]), .B(DB[1182]), .Z(n38310) );
  XNOR U38248 ( .A(q[3]), .B(DB[1181]), .Z(n29692) );
  XOR U38249 ( .A(n38311), .B(n29461), .Z(n29312) );
  XOR U38250 ( .A(n38312), .B(n29437), .Z(n29461) );
  XOR U38251 ( .A(n38313), .B(n29429), .Z(n29437) );
  XOR U38252 ( .A(n38314), .B(n29418), .Z(n29429) );
  XNOR U38253 ( .A(q[30]), .B(DB[1239]), .Z(n29418) );
  IV U38254 ( .A(n29417), .Z(n38314) );
  XNOR U38255 ( .A(n29415), .B(n38315), .Z(n29417) );
  XNOR U38256 ( .A(q[29]), .B(DB[1238]), .Z(n38315) );
  XNOR U38257 ( .A(q[28]), .B(DB[1237]), .Z(n29415) );
  IV U38258 ( .A(n29428), .Z(n38313) );
  XOR U38259 ( .A(n38316), .B(n38317), .Z(n29428) );
  XNOR U38260 ( .A(n29424), .B(n29426), .Z(n38317) );
  XNOR U38261 ( .A(q[24]), .B(DB[1233]), .Z(n29426) );
  XNOR U38262 ( .A(q[27]), .B(DB[1236]), .Z(n29424) );
  IV U38263 ( .A(n29423), .Z(n38316) );
  XNOR U38264 ( .A(n29421), .B(n38318), .Z(n29423) );
  XNOR U38265 ( .A(q[26]), .B(DB[1235]), .Z(n38318) );
  XNOR U38266 ( .A(q[25]), .B(DB[1234]), .Z(n29421) );
  IV U38267 ( .A(n29436), .Z(n38312) );
  XOR U38268 ( .A(n38319), .B(n38320), .Z(n29436) );
  XNOR U38269 ( .A(n29453), .B(n29434), .Z(n38320) );
  XNOR U38270 ( .A(q[16]), .B(DB[1225]), .Z(n29434) );
  XOR U38271 ( .A(n38321), .B(n29442), .Z(n29453) );
  XNOR U38272 ( .A(q[23]), .B(DB[1232]), .Z(n29442) );
  IV U38273 ( .A(n29441), .Z(n38321) );
  XNOR U38274 ( .A(n29439), .B(n38322), .Z(n29441) );
  XNOR U38275 ( .A(q[22]), .B(DB[1231]), .Z(n38322) );
  XNOR U38276 ( .A(q[21]), .B(DB[1230]), .Z(n29439) );
  IV U38277 ( .A(n29452), .Z(n38319) );
  XOR U38278 ( .A(n38323), .B(n38324), .Z(n29452) );
  XNOR U38279 ( .A(n29448), .B(n29450), .Z(n38324) );
  XNOR U38280 ( .A(q[17]), .B(DB[1226]), .Z(n29450) );
  XNOR U38281 ( .A(q[20]), .B(DB[1229]), .Z(n29448) );
  IV U38282 ( .A(n29447), .Z(n38323) );
  XNOR U38283 ( .A(n29445), .B(n38325), .Z(n29447) );
  XNOR U38284 ( .A(q[19]), .B(DB[1228]), .Z(n38325) );
  XNOR U38285 ( .A(q[18]), .B(DB[1227]), .Z(n29445) );
  IV U38286 ( .A(n29460), .Z(n38311) );
  XOR U38287 ( .A(n38326), .B(n38327), .Z(n29460) );
  XNOR U38288 ( .A(n29487), .B(n29458), .Z(n38327) );
  XNOR U38289 ( .A(q[0]), .B(DB[1209]), .Z(n29458) );
  XOR U38290 ( .A(n38328), .B(n29479), .Z(n29487) );
  XOR U38291 ( .A(n38329), .B(n29467), .Z(n29479) );
  XNOR U38292 ( .A(q[15]), .B(DB[1224]), .Z(n29467) );
  IV U38293 ( .A(n29466), .Z(n38329) );
  XNOR U38294 ( .A(n29464), .B(n38330), .Z(n29466) );
  XNOR U38295 ( .A(q[14]), .B(DB[1223]), .Z(n38330) );
  XNOR U38296 ( .A(q[13]), .B(DB[1222]), .Z(n29464) );
  IV U38297 ( .A(n29478), .Z(n38328) );
  XOR U38298 ( .A(n38331), .B(n38332), .Z(n29478) );
  XNOR U38299 ( .A(n29474), .B(n29476), .Z(n38332) );
  XNOR U38300 ( .A(q[9]), .B(DB[1218]), .Z(n29476) );
  XNOR U38301 ( .A(q[12]), .B(DB[1221]), .Z(n29474) );
  IV U38302 ( .A(n29473), .Z(n38331) );
  XNOR U38303 ( .A(n29471), .B(n38333), .Z(n29473) );
  XNOR U38304 ( .A(q[11]), .B(DB[1220]), .Z(n38333) );
  XNOR U38305 ( .A(q[10]), .B(DB[1219]), .Z(n29471) );
  IV U38306 ( .A(n29486), .Z(n38326) );
  XOR U38307 ( .A(n38334), .B(n38335), .Z(n29486) );
  XNOR U38308 ( .A(n29503), .B(n29484), .Z(n38335) );
  XNOR U38309 ( .A(q[1]), .B(DB[1210]), .Z(n29484) );
  XOR U38310 ( .A(n38336), .B(n29492), .Z(n29503) );
  XNOR U38311 ( .A(q[8]), .B(DB[1217]), .Z(n29492) );
  IV U38312 ( .A(n29491), .Z(n38336) );
  XNOR U38313 ( .A(n29489), .B(n38337), .Z(n29491) );
  XNOR U38314 ( .A(q[7]), .B(DB[1216]), .Z(n38337) );
  XNOR U38315 ( .A(q[6]), .B(DB[1215]), .Z(n29489) );
  IV U38316 ( .A(n29502), .Z(n38334) );
  XOR U38317 ( .A(n38338), .B(n38339), .Z(n29502) );
  XNOR U38318 ( .A(n29498), .B(n29500), .Z(n38339) );
  XNOR U38319 ( .A(q[2]), .B(DB[1211]), .Z(n29500) );
  XNOR U38320 ( .A(q[5]), .B(DB[1214]), .Z(n29498) );
  IV U38321 ( .A(n29497), .Z(n38338) );
  XNOR U38322 ( .A(n29495), .B(n38340), .Z(n29497) );
  XNOR U38323 ( .A(q[4]), .B(DB[1213]), .Z(n38340) );
  XNOR U38324 ( .A(q[3]), .B(DB[1212]), .Z(n29495) );
  XOR U38325 ( .A(n38341), .B(n29264), .Z(n29115) );
  XOR U38326 ( .A(n38342), .B(n29240), .Z(n29264) );
  XOR U38327 ( .A(n38343), .B(n29232), .Z(n29240) );
  XOR U38328 ( .A(n38344), .B(n29221), .Z(n29232) );
  XNOR U38329 ( .A(q[30]), .B(DB[1270]), .Z(n29221) );
  IV U38330 ( .A(n29220), .Z(n38344) );
  XNOR U38331 ( .A(n29218), .B(n38345), .Z(n29220) );
  XNOR U38332 ( .A(q[29]), .B(DB[1269]), .Z(n38345) );
  XNOR U38333 ( .A(q[28]), .B(DB[1268]), .Z(n29218) );
  IV U38334 ( .A(n29231), .Z(n38343) );
  XOR U38335 ( .A(n38346), .B(n38347), .Z(n29231) );
  XNOR U38336 ( .A(n29227), .B(n29229), .Z(n38347) );
  XNOR U38337 ( .A(q[24]), .B(DB[1264]), .Z(n29229) );
  XNOR U38338 ( .A(q[27]), .B(DB[1267]), .Z(n29227) );
  IV U38339 ( .A(n29226), .Z(n38346) );
  XNOR U38340 ( .A(n29224), .B(n38348), .Z(n29226) );
  XNOR U38341 ( .A(q[26]), .B(DB[1266]), .Z(n38348) );
  XNOR U38342 ( .A(q[25]), .B(DB[1265]), .Z(n29224) );
  IV U38343 ( .A(n29239), .Z(n38342) );
  XOR U38344 ( .A(n38349), .B(n38350), .Z(n29239) );
  XNOR U38345 ( .A(n29256), .B(n29237), .Z(n38350) );
  XNOR U38346 ( .A(q[16]), .B(DB[1256]), .Z(n29237) );
  XOR U38347 ( .A(n38351), .B(n29245), .Z(n29256) );
  XNOR U38348 ( .A(q[23]), .B(DB[1263]), .Z(n29245) );
  IV U38349 ( .A(n29244), .Z(n38351) );
  XNOR U38350 ( .A(n29242), .B(n38352), .Z(n29244) );
  XNOR U38351 ( .A(q[22]), .B(DB[1262]), .Z(n38352) );
  XNOR U38352 ( .A(q[21]), .B(DB[1261]), .Z(n29242) );
  IV U38353 ( .A(n29255), .Z(n38349) );
  XOR U38354 ( .A(n38353), .B(n38354), .Z(n29255) );
  XNOR U38355 ( .A(n29251), .B(n29253), .Z(n38354) );
  XNOR U38356 ( .A(q[17]), .B(DB[1257]), .Z(n29253) );
  XNOR U38357 ( .A(q[20]), .B(DB[1260]), .Z(n29251) );
  IV U38358 ( .A(n29250), .Z(n38353) );
  XNOR U38359 ( .A(n29248), .B(n38355), .Z(n29250) );
  XNOR U38360 ( .A(q[19]), .B(DB[1259]), .Z(n38355) );
  XNOR U38361 ( .A(q[18]), .B(DB[1258]), .Z(n29248) );
  IV U38362 ( .A(n29263), .Z(n38341) );
  XOR U38363 ( .A(n38356), .B(n38357), .Z(n29263) );
  XNOR U38364 ( .A(n29290), .B(n29261), .Z(n38357) );
  XNOR U38365 ( .A(q[0]), .B(DB[1240]), .Z(n29261) );
  XOR U38366 ( .A(n38358), .B(n29282), .Z(n29290) );
  XOR U38367 ( .A(n38359), .B(n29270), .Z(n29282) );
  XNOR U38368 ( .A(q[15]), .B(DB[1255]), .Z(n29270) );
  IV U38369 ( .A(n29269), .Z(n38359) );
  XNOR U38370 ( .A(n29267), .B(n38360), .Z(n29269) );
  XNOR U38371 ( .A(q[14]), .B(DB[1254]), .Z(n38360) );
  XNOR U38372 ( .A(q[13]), .B(DB[1253]), .Z(n29267) );
  IV U38373 ( .A(n29281), .Z(n38358) );
  XOR U38374 ( .A(n38361), .B(n38362), .Z(n29281) );
  XNOR U38375 ( .A(n29277), .B(n29279), .Z(n38362) );
  XNOR U38376 ( .A(q[9]), .B(DB[1249]), .Z(n29279) );
  XNOR U38377 ( .A(q[12]), .B(DB[1252]), .Z(n29277) );
  IV U38378 ( .A(n29276), .Z(n38361) );
  XNOR U38379 ( .A(n29274), .B(n38363), .Z(n29276) );
  XNOR U38380 ( .A(q[11]), .B(DB[1251]), .Z(n38363) );
  XNOR U38381 ( .A(q[10]), .B(DB[1250]), .Z(n29274) );
  IV U38382 ( .A(n29289), .Z(n38356) );
  XOR U38383 ( .A(n38364), .B(n38365), .Z(n29289) );
  XNOR U38384 ( .A(n29306), .B(n29287), .Z(n38365) );
  XNOR U38385 ( .A(q[1]), .B(DB[1241]), .Z(n29287) );
  XOR U38386 ( .A(n38366), .B(n29295), .Z(n29306) );
  XNOR U38387 ( .A(q[8]), .B(DB[1248]), .Z(n29295) );
  IV U38388 ( .A(n29294), .Z(n38366) );
  XNOR U38389 ( .A(n29292), .B(n38367), .Z(n29294) );
  XNOR U38390 ( .A(q[7]), .B(DB[1247]), .Z(n38367) );
  XNOR U38391 ( .A(q[6]), .B(DB[1246]), .Z(n29292) );
  IV U38392 ( .A(n29305), .Z(n38364) );
  XOR U38393 ( .A(n38368), .B(n38369), .Z(n29305) );
  XNOR U38394 ( .A(n29301), .B(n29303), .Z(n38369) );
  XNOR U38395 ( .A(q[2]), .B(DB[1242]), .Z(n29303) );
  XNOR U38396 ( .A(q[5]), .B(DB[1245]), .Z(n29301) );
  IV U38397 ( .A(n29300), .Z(n38368) );
  XNOR U38398 ( .A(n29298), .B(n38370), .Z(n29300) );
  XNOR U38399 ( .A(q[4]), .B(DB[1244]), .Z(n38370) );
  XNOR U38400 ( .A(q[3]), .B(DB[1243]), .Z(n29298) );
  XOR U38401 ( .A(n38371), .B(n29067), .Z(n28918) );
  XOR U38402 ( .A(n38372), .B(n29043), .Z(n29067) );
  XOR U38403 ( .A(n38373), .B(n29035), .Z(n29043) );
  XOR U38404 ( .A(n38374), .B(n29024), .Z(n29035) );
  XNOR U38405 ( .A(q[30]), .B(DB[1301]), .Z(n29024) );
  IV U38406 ( .A(n29023), .Z(n38374) );
  XNOR U38407 ( .A(n29021), .B(n38375), .Z(n29023) );
  XNOR U38408 ( .A(q[29]), .B(DB[1300]), .Z(n38375) );
  XNOR U38409 ( .A(q[28]), .B(DB[1299]), .Z(n29021) );
  IV U38410 ( .A(n29034), .Z(n38373) );
  XOR U38411 ( .A(n38376), .B(n38377), .Z(n29034) );
  XNOR U38412 ( .A(n29030), .B(n29032), .Z(n38377) );
  XNOR U38413 ( .A(q[24]), .B(DB[1295]), .Z(n29032) );
  XNOR U38414 ( .A(q[27]), .B(DB[1298]), .Z(n29030) );
  IV U38415 ( .A(n29029), .Z(n38376) );
  XNOR U38416 ( .A(n29027), .B(n38378), .Z(n29029) );
  XNOR U38417 ( .A(q[26]), .B(DB[1297]), .Z(n38378) );
  XNOR U38418 ( .A(q[25]), .B(DB[1296]), .Z(n29027) );
  IV U38419 ( .A(n29042), .Z(n38372) );
  XOR U38420 ( .A(n38379), .B(n38380), .Z(n29042) );
  XNOR U38421 ( .A(n29059), .B(n29040), .Z(n38380) );
  XNOR U38422 ( .A(q[16]), .B(DB[1287]), .Z(n29040) );
  XOR U38423 ( .A(n38381), .B(n29048), .Z(n29059) );
  XNOR U38424 ( .A(q[23]), .B(DB[1294]), .Z(n29048) );
  IV U38425 ( .A(n29047), .Z(n38381) );
  XNOR U38426 ( .A(n29045), .B(n38382), .Z(n29047) );
  XNOR U38427 ( .A(q[22]), .B(DB[1293]), .Z(n38382) );
  XNOR U38428 ( .A(q[21]), .B(DB[1292]), .Z(n29045) );
  IV U38429 ( .A(n29058), .Z(n38379) );
  XOR U38430 ( .A(n38383), .B(n38384), .Z(n29058) );
  XNOR U38431 ( .A(n29054), .B(n29056), .Z(n38384) );
  XNOR U38432 ( .A(q[17]), .B(DB[1288]), .Z(n29056) );
  XNOR U38433 ( .A(q[20]), .B(DB[1291]), .Z(n29054) );
  IV U38434 ( .A(n29053), .Z(n38383) );
  XNOR U38435 ( .A(n29051), .B(n38385), .Z(n29053) );
  XNOR U38436 ( .A(q[19]), .B(DB[1290]), .Z(n38385) );
  XNOR U38437 ( .A(q[18]), .B(DB[1289]), .Z(n29051) );
  IV U38438 ( .A(n29066), .Z(n38371) );
  XOR U38439 ( .A(n38386), .B(n38387), .Z(n29066) );
  XNOR U38440 ( .A(n29093), .B(n29064), .Z(n38387) );
  XNOR U38441 ( .A(q[0]), .B(DB[1271]), .Z(n29064) );
  XOR U38442 ( .A(n38388), .B(n29085), .Z(n29093) );
  XOR U38443 ( .A(n38389), .B(n29073), .Z(n29085) );
  XNOR U38444 ( .A(q[15]), .B(DB[1286]), .Z(n29073) );
  IV U38445 ( .A(n29072), .Z(n38389) );
  XNOR U38446 ( .A(n29070), .B(n38390), .Z(n29072) );
  XNOR U38447 ( .A(q[14]), .B(DB[1285]), .Z(n38390) );
  XNOR U38448 ( .A(q[13]), .B(DB[1284]), .Z(n29070) );
  IV U38449 ( .A(n29084), .Z(n38388) );
  XOR U38450 ( .A(n38391), .B(n38392), .Z(n29084) );
  XNOR U38451 ( .A(n29080), .B(n29082), .Z(n38392) );
  XNOR U38452 ( .A(q[9]), .B(DB[1280]), .Z(n29082) );
  XNOR U38453 ( .A(q[12]), .B(DB[1283]), .Z(n29080) );
  IV U38454 ( .A(n29079), .Z(n38391) );
  XNOR U38455 ( .A(n29077), .B(n38393), .Z(n29079) );
  XNOR U38456 ( .A(q[11]), .B(DB[1282]), .Z(n38393) );
  XNOR U38457 ( .A(q[10]), .B(DB[1281]), .Z(n29077) );
  IV U38458 ( .A(n29092), .Z(n38386) );
  XOR U38459 ( .A(n38394), .B(n38395), .Z(n29092) );
  XNOR U38460 ( .A(n29109), .B(n29090), .Z(n38395) );
  XNOR U38461 ( .A(q[1]), .B(DB[1272]), .Z(n29090) );
  XOR U38462 ( .A(n38396), .B(n29098), .Z(n29109) );
  XNOR U38463 ( .A(q[8]), .B(DB[1279]), .Z(n29098) );
  IV U38464 ( .A(n29097), .Z(n38396) );
  XNOR U38465 ( .A(n29095), .B(n38397), .Z(n29097) );
  XNOR U38466 ( .A(q[7]), .B(DB[1278]), .Z(n38397) );
  XNOR U38467 ( .A(q[6]), .B(DB[1277]), .Z(n29095) );
  IV U38468 ( .A(n29108), .Z(n38394) );
  XOR U38469 ( .A(n38398), .B(n38399), .Z(n29108) );
  XNOR U38470 ( .A(n29104), .B(n29106), .Z(n38399) );
  XNOR U38471 ( .A(q[2]), .B(DB[1273]), .Z(n29106) );
  XNOR U38472 ( .A(q[5]), .B(DB[1276]), .Z(n29104) );
  IV U38473 ( .A(n29103), .Z(n38398) );
  XNOR U38474 ( .A(n29101), .B(n38400), .Z(n29103) );
  XNOR U38475 ( .A(q[4]), .B(DB[1275]), .Z(n38400) );
  XNOR U38476 ( .A(q[3]), .B(DB[1274]), .Z(n29101) );
  XOR U38477 ( .A(n38401), .B(n28870), .Z(n28721) );
  XOR U38478 ( .A(n38402), .B(n28846), .Z(n28870) );
  XOR U38479 ( .A(n38403), .B(n28838), .Z(n28846) );
  XOR U38480 ( .A(n38404), .B(n28827), .Z(n28838) );
  XNOR U38481 ( .A(q[30]), .B(DB[1332]), .Z(n28827) );
  IV U38482 ( .A(n28826), .Z(n38404) );
  XNOR U38483 ( .A(n28824), .B(n38405), .Z(n28826) );
  XNOR U38484 ( .A(q[29]), .B(DB[1331]), .Z(n38405) );
  XNOR U38485 ( .A(q[28]), .B(DB[1330]), .Z(n28824) );
  IV U38486 ( .A(n28837), .Z(n38403) );
  XOR U38487 ( .A(n38406), .B(n38407), .Z(n28837) );
  XNOR U38488 ( .A(n28833), .B(n28835), .Z(n38407) );
  XNOR U38489 ( .A(q[24]), .B(DB[1326]), .Z(n28835) );
  XNOR U38490 ( .A(q[27]), .B(DB[1329]), .Z(n28833) );
  IV U38491 ( .A(n28832), .Z(n38406) );
  XNOR U38492 ( .A(n28830), .B(n38408), .Z(n28832) );
  XNOR U38493 ( .A(q[26]), .B(DB[1328]), .Z(n38408) );
  XNOR U38494 ( .A(q[25]), .B(DB[1327]), .Z(n28830) );
  IV U38495 ( .A(n28845), .Z(n38402) );
  XOR U38496 ( .A(n38409), .B(n38410), .Z(n28845) );
  XNOR U38497 ( .A(n28862), .B(n28843), .Z(n38410) );
  XNOR U38498 ( .A(q[16]), .B(DB[1318]), .Z(n28843) );
  XOR U38499 ( .A(n38411), .B(n28851), .Z(n28862) );
  XNOR U38500 ( .A(q[23]), .B(DB[1325]), .Z(n28851) );
  IV U38501 ( .A(n28850), .Z(n38411) );
  XNOR U38502 ( .A(n28848), .B(n38412), .Z(n28850) );
  XNOR U38503 ( .A(q[22]), .B(DB[1324]), .Z(n38412) );
  XNOR U38504 ( .A(q[21]), .B(DB[1323]), .Z(n28848) );
  IV U38505 ( .A(n28861), .Z(n38409) );
  XOR U38506 ( .A(n38413), .B(n38414), .Z(n28861) );
  XNOR U38507 ( .A(n28857), .B(n28859), .Z(n38414) );
  XNOR U38508 ( .A(q[17]), .B(DB[1319]), .Z(n28859) );
  XNOR U38509 ( .A(q[20]), .B(DB[1322]), .Z(n28857) );
  IV U38510 ( .A(n28856), .Z(n38413) );
  XNOR U38511 ( .A(n28854), .B(n38415), .Z(n28856) );
  XNOR U38512 ( .A(q[19]), .B(DB[1321]), .Z(n38415) );
  XNOR U38513 ( .A(q[18]), .B(DB[1320]), .Z(n28854) );
  IV U38514 ( .A(n28869), .Z(n38401) );
  XOR U38515 ( .A(n38416), .B(n38417), .Z(n28869) );
  XNOR U38516 ( .A(n28896), .B(n28867), .Z(n38417) );
  XNOR U38517 ( .A(q[0]), .B(DB[1302]), .Z(n28867) );
  XOR U38518 ( .A(n38418), .B(n28888), .Z(n28896) );
  XOR U38519 ( .A(n38419), .B(n28876), .Z(n28888) );
  XNOR U38520 ( .A(q[15]), .B(DB[1317]), .Z(n28876) );
  IV U38521 ( .A(n28875), .Z(n38419) );
  XNOR U38522 ( .A(n28873), .B(n38420), .Z(n28875) );
  XNOR U38523 ( .A(q[14]), .B(DB[1316]), .Z(n38420) );
  XNOR U38524 ( .A(q[13]), .B(DB[1315]), .Z(n28873) );
  IV U38525 ( .A(n28887), .Z(n38418) );
  XOR U38526 ( .A(n38421), .B(n38422), .Z(n28887) );
  XNOR U38527 ( .A(n28883), .B(n28885), .Z(n38422) );
  XNOR U38528 ( .A(q[9]), .B(DB[1311]), .Z(n28885) );
  XNOR U38529 ( .A(q[12]), .B(DB[1314]), .Z(n28883) );
  IV U38530 ( .A(n28882), .Z(n38421) );
  XNOR U38531 ( .A(n28880), .B(n38423), .Z(n28882) );
  XNOR U38532 ( .A(q[11]), .B(DB[1313]), .Z(n38423) );
  XNOR U38533 ( .A(q[10]), .B(DB[1312]), .Z(n28880) );
  IV U38534 ( .A(n28895), .Z(n38416) );
  XOR U38535 ( .A(n38424), .B(n38425), .Z(n28895) );
  XNOR U38536 ( .A(n28912), .B(n28893), .Z(n38425) );
  XNOR U38537 ( .A(q[1]), .B(DB[1303]), .Z(n28893) );
  XOR U38538 ( .A(n38426), .B(n28901), .Z(n28912) );
  XNOR U38539 ( .A(q[8]), .B(DB[1310]), .Z(n28901) );
  IV U38540 ( .A(n28900), .Z(n38426) );
  XNOR U38541 ( .A(n28898), .B(n38427), .Z(n28900) );
  XNOR U38542 ( .A(q[7]), .B(DB[1309]), .Z(n38427) );
  XNOR U38543 ( .A(q[6]), .B(DB[1308]), .Z(n28898) );
  IV U38544 ( .A(n28911), .Z(n38424) );
  XOR U38545 ( .A(n38428), .B(n38429), .Z(n28911) );
  XNOR U38546 ( .A(n28907), .B(n28909), .Z(n38429) );
  XNOR U38547 ( .A(q[2]), .B(DB[1304]), .Z(n28909) );
  XNOR U38548 ( .A(q[5]), .B(DB[1307]), .Z(n28907) );
  IV U38549 ( .A(n28906), .Z(n38428) );
  XNOR U38550 ( .A(n28904), .B(n38430), .Z(n28906) );
  XNOR U38551 ( .A(q[4]), .B(DB[1306]), .Z(n38430) );
  XNOR U38552 ( .A(q[3]), .B(DB[1305]), .Z(n28904) );
  XOR U38553 ( .A(n38431), .B(n28673), .Z(n28524) );
  XOR U38554 ( .A(n38432), .B(n28649), .Z(n28673) );
  XOR U38555 ( .A(n38433), .B(n28641), .Z(n28649) );
  XOR U38556 ( .A(n38434), .B(n28630), .Z(n28641) );
  XNOR U38557 ( .A(q[30]), .B(DB[1363]), .Z(n28630) );
  IV U38558 ( .A(n28629), .Z(n38434) );
  XNOR U38559 ( .A(n28627), .B(n38435), .Z(n28629) );
  XNOR U38560 ( .A(q[29]), .B(DB[1362]), .Z(n38435) );
  XNOR U38561 ( .A(q[28]), .B(DB[1361]), .Z(n28627) );
  IV U38562 ( .A(n28640), .Z(n38433) );
  XOR U38563 ( .A(n38436), .B(n38437), .Z(n28640) );
  XNOR U38564 ( .A(n28636), .B(n28638), .Z(n38437) );
  XNOR U38565 ( .A(q[24]), .B(DB[1357]), .Z(n28638) );
  XNOR U38566 ( .A(q[27]), .B(DB[1360]), .Z(n28636) );
  IV U38567 ( .A(n28635), .Z(n38436) );
  XNOR U38568 ( .A(n28633), .B(n38438), .Z(n28635) );
  XNOR U38569 ( .A(q[26]), .B(DB[1359]), .Z(n38438) );
  XNOR U38570 ( .A(q[25]), .B(DB[1358]), .Z(n28633) );
  IV U38571 ( .A(n28648), .Z(n38432) );
  XOR U38572 ( .A(n38439), .B(n38440), .Z(n28648) );
  XNOR U38573 ( .A(n28665), .B(n28646), .Z(n38440) );
  XNOR U38574 ( .A(q[16]), .B(DB[1349]), .Z(n28646) );
  XOR U38575 ( .A(n38441), .B(n28654), .Z(n28665) );
  XNOR U38576 ( .A(q[23]), .B(DB[1356]), .Z(n28654) );
  IV U38577 ( .A(n28653), .Z(n38441) );
  XNOR U38578 ( .A(n28651), .B(n38442), .Z(n28653) );
  XNOR U38579 ( .A(q[22]), .B(DB[1355]), .Z(n38442) );
  XNOR U38580 ( .A(q[21]), .B(DB[1354]), .Z(n28651) );
  IV U38581 ( .A(n28664), .Z(n38439) );
  XOR U38582 ( .A(n38443), .B(n38444), .Z(n28664) );
  XNOR U38583 ( .A(n28660), .B(n28662), .Z(n38444) );
  XNOR U38584 ( .A(q[17]), .B(DB[1350]), .Z(n28662) );
  XNOR U38585 ( .A(q[20]), .B(DB[1353]), .Z(n28660) );
  IV U38586 ( .A(n28659), .Z(n38443) );
  XNOR U38587 ( .A(n28657), .B(n38445), .Z(n28659) );
  XNOR U38588 ( .A(q[19]), .B(DB[1352]), .Z(n38445) );
  XNOR U38589 ( .A(q[18]), .B(DB[1351]), .Z(n28657) );
  IV U38590 ( .A(n28672), .Z(n38431) );
  XOR U38591 ( .A(n38446), .B(n38447), .Z(n28672) );
  XNOR U38592 ( .A(n28699), .B(n28670), .Z(n38447) );
  XNOR U38593 ( .A(q[0]), .B(DB[1333]), .Z(n28670) );
  XOR U38594 ( .A(n38448), .B(n28691), .Z(n28699) );
  XOR U38595 ( .A(n38449), .B(n28679), .Z(n28691) );
  XNOR U38596 ( .A(q[15]), .B(DB[1348]), .Z(n28679) );
  IV U38597 ( .A(n28678), .Z(n38449) );
  XNOR U38598 ( .A(n28676), .B(n38450), .Z(n28678) );
  XNOR U38599 ( .A(q[14]), .B(DB[1347]), .Z(n38450) );
  XNOR U38600 ( .A(q[13]), .B(DB[1346]), .Z(n28676) );
  IV U38601 ( .A(n28690), .Z(n38448) );
  XOR U38602 ( .A(n38451), .B(n38452), .Z(n28690) );
  XNOR U38603 ( .A(n28686), .B(n28688), .Z(n38452) );
  XNOR U38604 ( .A(q[9]), .B(DB[1342]), .Z(n28688) );
  XNOR U38605 ( .A(q[12]), .B(DB[1345]), .Z(n28686) );
  IV U38606 ( .A(n28685), .Z(n38451) );
  XNOR U38607 ( .A(n28683), .B(n38453), .Z(n28685) );
  XNOR U38608 ( .A(q[11]), .B(DB[1344]), .Z(n38453) );
  XNOR U38609 ( .A(q[10]), .B(DB[1343]), .Z(n28683) );
  IV U38610 ( .A(n28698), .Z(n38446) );
  XOR U38611 ( .A(n38454), .B(n38455), .Z(n28698) );
  XNOR U38612 ( .A(n28715), .B(n28696), .Z(n38455) );
  XNOR U38613 ( .A(q[1]), .B(DB[1334]), .Z(n28696) );
  XOR U38614 ( .A(n38456), .B(n28704), .Z(n28715) );
  XNOR U38615 ( .A(q[8]), .B(DB[1341]), .Z(n28704) );
  IV U38616 ( .A(n28703), .Z(n38456) );
  XNOR U38617 ( .A(n28701), .B(n38457), .Z(n28703) );
  XNOR U38618 ( .A(q[7]), .B(DB[1340]), .Z(n38457) );
  XNOR U38619 ( .A(q[6]), .B(DB[1339]), .Z(n28701) );
  IV U38620 ( .A(n28714), .Z(n38454) );
  XOR U38621 ( .A(n38458), .B(n38459), .Z(n28714) );
  XNOR U38622 ( .A(n28710), .B(n28712), .Z(n38459) );
  XNOR U38623 ( .A(q[2]), .B(DB[1335]), .Z(n28712) );
  XNOR U38624 ( .A(q[5]), .B(DB[1338]), .Z(n28710) );
  IV U38625 ( .A(n28709), .Z(n38458) );
  XNOR U38626 ( .A(n28707), .B(n38460), .Z(n28709) );
  XNOR U38627 ( .A(q[4]), .B(DB[1337]), .Z(n38460) );
  XNOR U38628 ( .A(q[3]), .B(DB[1336]), .Z(n28707) );
  XOR U38629 ( .A(n38461), .B(n28476), .Z(n28327) );
  XOR U38630 ( .A(n38462), .B(n28452), .Z(n28476) );
  XOR U38631 ( .A(n38463), .B(n28444), .Z(n28452) );
  XOR U38632 ( .A(n38464), .B(n28433), .Z(n28444) );
  XNOR U38633 ( .A(q[30]), .B(DB[1394]), .Z(n28433) );
  IV U38634 ( .A(n28432), .Z(n38464) );
  XNOR U38635 ( .A(n28430), .B(n38465), .Z(n28432) );
  XNOR U38636 ( .A(q[29]), .B(DB[1393]), .Z(n38465) );
  XNOR U38637 ( .A(q[28]), .B(DB[1392]), .Z(n28430) );
  IV U38638 ( .A(n28443), .Z(n38463) );
  XOR U38639 ( .A(n38466), .B(n38467), .Z(n28443) );
  XNOR U38640 ( .A(n28439), .B(n28441), .Z(n38467) );
  XNOR U38641 ( .A(q[24]), .B(DB[1388]), .Z(n28441) );
  XNOR U38642 ( .A(q[27]), .B(DB[1391]), .Z(n28439) );
  IV U38643 ( .A(n28438), .Z(n38466) );
  XNOR U38644 ( .A(n28436), .B(n38468), .Z(n28438) );
  XNOR U38645 ( .A(q[26]), .B(DB[1390]), .Z(n38468) );
  XNOR U38646 ( .A(q[25]), .B(DB[1389]), .Z(n28436) );
  IV U38647 ( .A(n28451), .Z(n38462) );
  XOR U38648 ( .A(n38469), .B(n38470), .Z(n28451) );
  XNOR U38649 ( .A(n28468), .B(n28449), .Z(n38470) );
  XNOR U38650 ( .A(q[16]), .B(DB[1380]), .Z(n28449) );
  XOR U38651 ( .A(n38471), .B(n28457), .Z(n28468) );
  XNOR U38652 ( .A(q[23]), .B(DB[1387]), .Z(n28457) );
  IV U38653 ( .A(n28456), .Z(n38471) );
  XNOR U38654 ( .A(n28454), .B(n38472), .Z(n28456) );
  XNOR U38655 ( .A(q[22]), .B(DB[1386]), .Z(n38472) );
  XNOR U38656 ( .A(q[21]), .B(DB[1385]), .Z(n28454) );
  IV U38657 ( .A(n28467), .Z(n38469) );
  XOR U38658 ( .A(n38473), .B(n38474), .Z(n28467) );
  XNOR U38659 ( .A(n28463), .B(n28465), .Z(n38474) );
  XNOR U38660 ( .A(q[17]), .B(DB[1381]), .Z(n28465) );
  XNOR U38661 ( .A(q[20]), .B(DB[1384]), .Z(n28463) );
  IV U38662 ( .A(n28462), .Z(n38473) );
  XNOR U38663 ( .A(n28460), .B(n38475), .Z(n28462) );
  XNOR U38664 ( .A(q[19]), .B(DB[1383]), .Z(n38475) );
  XNOR U38665 ( .A(q[18]), .B(DB[1382]), .Z(n28460) );
  IV U38666 ( .A(n28475), .Z(n38461) );
  XOR U38667 ( .A(n38476), .B(n38477), .Z(n28475) );
  XNOR U38668 ( .A(n28502), .B(n28473), .Z(n38477) );
  XNOR U38669 ( .A(q[0]), .B(DB[1364]), .Z(n28473) );
  XOR U38670 ( .A(n38478), .B(n28494), .Z(n28502) );
  XOR U38671 ( .A(n38479), .B(n28482), .Z(n28494) );
  XNOR U38672 ( .A(q[15]), .B(DB[1379]), .Z(n28482) );
  IV U38673 ( .A(n28481), .Z(n38479) );
  XNOR U38674 ( .A(n28479), .B(n38480), .Z(n28481) );
  XNOR U38675 ( .A(q[14]), .B(DB[1378]), .Z(n38480) );
  XNOR U38676 ( .A(q[13]), .B(DB[1377]), .Z(n28479) );
  IV U38677 ( .A(n28493), .Z(n38478) );
  XOR U38678 ( .A(n38481), .B(n38482), .Z(n28493) );
  XNOR U38679 ( .A(n28489), .B(n28491), .Z(n38482) );
  XNOR U38680 ( .A(q[9]), .B(DB[1373]), .Z(n28491) );
  XNOR U38681 ( .A(q[12]), .B(DB[1376]), .Z(n28489) );
  IV U38682 ( .A(n28488), .Z(n38481) );
  XNOR U38683 ( .A(n28486), .B(n38483), .Z(n28488) );
  XNOR U38684 ( .A(q[11]), .B(DB[1375]), .Z(n38483) );
  XNOR U38685 ( .A(q[10]), .B(DB[1374]), .Z(n28486) );
  IV U38686 ( .A(n28501), .Z(n38476) );
  XOR U38687 ( .A(n38484), .B(n38485), .Z(n28501) );
  XNOR U38688 ( .A(n28518), .B(n28499), .Z(n38485) );
  XNOR U38689 ( .A(q[1]), .B(DB[1365]), .Z(n28499) );
  XOR U38690 ( .A(n38486), .B(n28507), .Z(n28518) );
  XNOR U38691 ( .A(q[8]), .B(DB[1372]), .Z(n28507) );
  IV U38692 ( .A(n28506), .Z(n38486) );
  XNOR U38693 ( .A(n28504), .B(n38487), .Z(n28506) );
  XNOR U38694 ( .A(q[7]), .B(DB[1371]), .Z(n38487) );
  XNOR U38695 ( .A(q[6]), .B(DB[1370]), .Z(n28504) );
  IV U38696 ( .A(n28517), .Z(n38484) );
  XOR U38697 ( .A(n38488), .B(n38489), .Z(n28517) );
  XNOR U38698 ( .A(n28513), .B(n28515), .Z(n38489) );
  XNOR U38699 ( .A(q[2]), .B(DB[1366]), .Z(n28515) );
  XNOR U38700 ( .A(q[5]), .B(DB[1369]), .Z(n28513) );
  IV U38701 ( .A(n28512), .Z(n38488) );
  XNOR U38702 ( .A(n28510), .B(n38490), .Z(n28512) );
  XNOR U38703 ( .A(q[4]), .B(DB[1368]), .Z(n38490) );
  XNOR U38704 ( .A(q[3]), .B(DB[1367]), .Z(n28510) );
  XOR U38705 ( .A(n38491), .B(n28279), .Z(n28130) );
  XOR U38706 ( .A(n38492), .B(n28255), .Z(n28279) );
  XOR U38707 ( .A(n38493), .B(n28247), .Z(n28255) );
  XOR U38708 ( .A(n38494), .B(n28236), .Z(n28247) );
  XNOR U38709 ( .A(q[30]), .B(DB[1425]), .Z(n28236) );
  IV U38710 ( .A(n28235), .Z(n38494) );
  XNOR U38711 ( .A(n28233), .B(n38495), .Z(n28235) );
  XNOR U38712 ( .A(q[29]), .B(DB[1424]), .Z(n38495) );
  XNOR U38713 ( .A(q[28]), .B(DB[1423]), .Z(n28233) );
  IV U38714 ( .A(n28246), .Z(n38493) );
  XOR U38715 ( .A(n38496), .B(n38497), .Z(n28246) );
  XNOR U38716 ( .A(n28242), .B(n28244), .Z(n38497) );
  XNOR U38717 ( .A(q[24]), .B(DB[1419]), .Z(n28244) );
  XNOR U38718 ( .A(q[27]), .B(DB[1422]), .Z(n28242) );
  IV U38719 ( .A(n28241), .Z(n38496) );
  XNOR U38720 ( .A(n28239), .B(n38498), .Z(n28241) );
  XNOR U38721 ( .A(q[26]), .B(DB[1421]), .Z(n38498) );
  XNOR U38722 ( .A(q[25]), .B(DB[1420]), .Z(n28239) );
  IV U38723 ( .A(n28254), .Z(n38492) );
  XOR U38724 ( .A(n38499), .B(n38500), .Z(n28254) );
  XNOR U38725 ( .A(n28271), .B(n28252), .Z(n38500) );
  XNOR U38726 ( .A(q[16]), .B(DB[1411]), .Z(n28252) );
  XOR U38727 ( .A(n38501), .B(n28260), .Z(n28271) );
  XNOR U38728 ( .A(q[23]), .B(DB[1418]), .Z(n28260) );
  IV U38729 ( .A(n28259), .Z(n38501) );
  XNOR U38730 ( .A(n28257), .B(n38502), .Z(n28259) );
  XNOR U38731 ( .A(q[22]), .B(DB[1417]), .Z(n38502) );
  XNOR U38732 ( .A(q[21]), .B(DB[1416]), .Z(n28257) );
  IV U38733 ( .A(n28270), .Z(n38499) );
  XOR U38734 ( .A(n38503), .B(n38504), .Z(n28270) );
  XNOR U38735 ( .A(n28266), .B(n28268), .Z(n38504) );
  XNOR U38736 ( .A(q[17]), .B(DB[1412]), .Z(n28268) );
  XNOR U38737 ( .A(q[20]), .B(DB[1415]), .Z(n28266) );
  IV U38738 ( .A(n28265), .Z(n38503) );
  XNOR U38739 ( .A(n28263), .B(n38505), .Z(n28265) );
  XNOR U38740 ( .A(q[19]), .B(DB[1414]), .Z(n38505) );
  XNOR U38741 ( .A(q[18]), .B(DB[1413]), .Z(n28263) );
  IV U38742 ( .A(n28278), .Z(n38491) );
  XOR U38743 ( .A(n38506), .B(n38507), .Z(n28278) );
  XNOR U38744 ( .A(n28305), .B(n28276), .Z(n38507) );
  XNOR U38745 ( .A(q[0]), .B(DB[1395]), .Z(n28276) );
  XOR U38746 ( .A(n38508), .B(n28297), .Z(n28305) );
  XOR U38747 ( .A(n38509), .B(n28285), .Z(n28297) );
  XNOR U38748 ( .A(q[15]), .B(DB[1410]), .Z(n28285) );
  IV U38749 ( .A(n28284), .Z(n38509) );
  XNOR U38750 ( .A(n28282), .B(n38510), .Z(n28284) );
  XNOR U38751 ( .A(q[14]), .B(DB[1409]), .Z(n38510) );
  XNOR U38752 ( .A(q[13]), .B(DB[1408]), .Z(n28282) );
  IV U38753 ( .A(n28296), .Z(n38508) );
  XOR U38754 ( .A(n38511), .B(n38512), .Z(n28296) );
  XNOR U38755 ( .A(n28292), .B(n28294), .Z(n38512) );
  XNOR U38756 ( .A(q[9]), .B(DB[1404]), .Z(n28294) );
  XNOR U38757 ( .A(q[12]), .B(DB[1407]), .Z(n28292) );
  IV U38758 ( .A(n28291), .Z(n38511) );
  XNOR U38759 ( .A(n28289), .B(n38513), .Z(n28291) );
  XNOR U38760 ( .A(q[11]), .B(DB[1406]), .Z(n38513) );
  XNOR U38761 ( .A(q[10]), .B(DB[1405]), .Z(n28289) );
  IV U38762 ( .A(n28304), .Z(n38506) );
  XOR U38763 ( .A(n38514), .B(n38515), .Z(n28304) );
  XNOR U38764 ( .A(n28321), .B(n28302), .Z(n38515) );
  XNOR U38765 ( .A(q[1]), .B(DB[1396]), .Z(n28302) );
  XOR U38766 ( .A(n38516), .B(n28310), .Z(n28321) );
  XNOR U38767 ( .A(q[8]), .B(DB[1403]), .Z(n28310) );
  IV U38768 ( .A(n28309), .Z(n38516) );
  XNOR U38769 ( .A(n28307), .B(n38517), .Z(n28309) );
  XNOR U38770 ( .A(q[7]), .B(DB[1402]), .Z(n38517) );
  XNOR U38771 ( .A(q[6]), .B(DB[1401]), .Z(n28307) );
  IV U38772 ( .A(n28320), .Z(n38514) );
  XOR U38773 ( .A(n38518), .B(n38519), .Z(n28320) );
  XNOR U38774 ( .A(n28316), .B(n28318), .Z(n38519) );
  XNOR U38775 ( .A(q[2]), .B(DB[1397]), .Z(n28318) );
  XNOR U38776 ( .A(q[5]), .B(DB[1400]), .Z(n28316) );
  IV U38777 ( .A(n28315), .Z(n38518) );
  XNOR U38778 ( .A(n28313), .B(n38520), .Z(n28315) );
  XNOR U38779 ( .A(q[4]), .B(DB[1399]), .Z(n38520) );
  XNOR U38780 ( .A(q[3]), .B(DB[1398]), .Z(n28313) );
  XOR U38781 ( .A(n38521), .B(n28082), .Z(n27933) );
  XOR U38782 ( .A(n38522), .B(n28058), .Z(n28082) );
  XOR U38783 ( .A(n38523), .B(n28050), .Z(n28058) );
  XOR U38784 ( .A(n38524), .B(n28039), .Z(n28050) );
  XNOR U38785 ( .A(q[30]), .B(DB[1456]), .Z(n28039) );
  IV U38786 ( .A(n28038), .Z(n38524) );
  XNOR U38787 ( .A(n28036), .B(n38525), .Z(n28038) );
  XNOR U38788 ( .A(q[29]), .B(DB[1455]), .Z(n38525) );
  XNOR U38789 ( .A(q[28]), .B(DB[1454]), .Z(n28036) );
  IV U38790 ( .A(n28049), .Z(n38523) );
  XOR U38791 ( .A(n38526), .B(n38527), .Z(n28049) );
  XNOR U38792 ( .A(n28045), .B(n28047), .Z(n38527) );
  XNOR U38793 ( .A(q[24]), .B(DB[1450]), .Z(n28047) );
  XNOR U38794 ( .A(q[27]), .B(DB[1453]), .Z(n28045) );
  IV U38795 ( .A(n28044), .Z(n38526) );
  XNOR U38796 ( .A(n28042), .B(n38528), .Z(n28044) );
  XNOR U38797 ( .A(q[26]), .B(DB[1452]), .Z(n38528) );
  XNOR U38798 ( .A(q[25]), .B(DB[1451]), .Z(n28042) );
  IV U38799 ( .A(n28057), .Z(n38522) );
  XOR U38800 ( .A(n38529), .B(n38530), .Z(n28057) );
  XNOR U38801 ( .A(n28074), .B(n28055), .Z(n38530) );
  XNOR U38802 ( .A(q[16]), .B(DB[1442]), .Z(n28055) );
  XOR U38803 ( .A(n38531), .B(n28063), .Z(n28074) );
  XNOR U38804 ( .A(q[23]), .B(DB[1449]), .Z(n28063) );
  IV U38805 ( .A(n28062), .Z(n38531) );
  XNOR U38806 ( .A(n28060), .B(n38532), .Z(n28062) );
  XNOR U38807 ( .A(q[22]), .B(DB[1448]), .Z(n38532) );
  XNOR U38808 ( .A(q[21]), .B(DB[1447]), .Z(n28060) );
  IV U38809 ( .A(n28073), .Z(n38529) );
  XOR U38810 ( .A(n38533), .B(n38534), .Z(n28073) );
  XNOR U38811 ( .A(n28069), .B(n28071), .Z(n38534) );
  XNOR U38812 ( .A(q[17]), .B(DB[1443]), .Z(n28071) );
  XNOR U38813 ( .A(q[20]), .B(DB[1446]), .Z(n28069) );
  IV U38814 ( .A(n28068), .Z(n38533) );
  XNOR U38815 ( .A(n28066), .B(n38535), .Z(n28068) );
  XNOR U38816 ( .A(q[19]), .B(DB[1445]), .Z(n38535) );
  XNOR U38817 ( .A(q[18]), .B(DB[1444]), .Z(n28066) );
  IV U38818 ( .A(n28081), .Z(n38521) );
  XOR U38819 ( .A(n38536), .B(n38537), .Z(n28081) );
  XNOR U38820 ( .A(n28108), .B(n28079), .Z(n38537) );
  XNOR U38821 ( .A(q[0]), .B(DB[1426]), .Z(n28079) );
  XOR U38822 ( .A(n38538), .B(n28100), .Z(n28108) );
  XOR U38823 ( .A(n38539), .B(n28088), .Z(n28100) );
  XNOR U38824 ( .A(q[15]), .B(DB[1441]), .Z(n28088) );
  IV U38825 ( .A(n28087), .Z(n38539) );
  XNOR U38826 ( .A(n28085), .B(n38540), .Z(n28087) );
  XNOR U38827 ( .A(q[14]), .B(DB[1440]), .Z(n38540) );
  XNOR U38828 ( .A(q[13]), .B(DB[1439]), .Z(n28085) );
  IV U38829 ( .A(n28099), .Z(n38538) );
  XOR U38830 ( .A(n38541), .B(n38542), .Z(n28099) );
  XNOR U38831 ( .A(n28095), .B(n28097), .Z(n38542) );
  XNOR U38832 ( .A(q[9]), .B(DB[1435]), .Z(n28097) );
  XNOR U38833 ( .A(q[12]), .B(DB[1438]), .Z(n28095) );
  IV U38834 ( .A(n28094), .Z(n38541) );
  XNOR U38835 ( .A(n28092), .B(n38543), .Z(n28094) );
  XNOR U38836 ( .A(q[11]), .B(DB[1437]), .Z(n38543) );
  XNOR U38837 ( .A(q[10]), .B(DB[1436]), .Z(n28092) );
  IV U38838 ( .A(n28107), .Z(n38536) );
  XOR U38839 ( .A(n38544), .B(n38545), .Z(n28107) );
  XNOR U38840 ( .A(n28124), .B(n28105), .Z(n38545) );
  XNOR U38841 ( .A(q[1]), .B(DB[1427]), .Z(n28105) );
  XOR U38842 ( .A(n38546), .B(n28113), .Z(n28124) );
  XNOR U38843 ( .A(q[8]), .B(DB[1434]), .Z(n28113) );
  IV U38844 ( .A(n28112), .Z(n38546) );
  XNOR U38845 ( .A(n28110), .B(n38547), .Z(n28112) );
  XNOR U38846 ( .A(q[7]), .B(DB[1433]), .Z(n38547) );
  XNOR U38847 ( .A(q[6]), .B(DB[1432]), .Z(n28110) );
  IV U38848 ( .A(n28123), .Z(n38544) );
  XOR U38849 ( .A(n38548), .B(n38549), .Z(n28123) );
  XNOR U38850 ( .A(n28119), .B(n28121), .Z(n38549) );
  XNOR U38851 ( .A(q[2]), .B(DB[1428]), .Z(n28121) );
  XNOR U38852 ( .A(q[5]), .B(DB[1431]), .Z(n28119) );
  IV U38853 ( .A(n28118), .Z(n38548) );
  XNOR U38854 ( .A(n28116), .B(n38550), .Z(n28118) );
  XNOR U38855 ( .A(q[4]), .B(DB[1430]), .Z(n38550) );
  XNOR U38856 ( .A(q[3]), .B(DB[1429]), .Z(n28116) );
  XOR U38857 ( .A(n38551), .B(n27885), .Z(n27736) );
  XOR U38858 ( .A(n38552), .B(n27861), .Z(n27885) );
  XOR U38859 ( .A(n38553), .B(n27853), .Z(n27861) );
  XOR U38860 ( .A(n38554), .B(n27842), .Z(n27853) );
  XNOR U38861 ( .A(q[30]), .B(DB[1487]), .Z(n27842) );
  IV U38862 ( .A(n27841), .Z(n38554) );
  XNOR U38863 ( .A(n27839), .B(n38555), .Z(n27841) );
  XNOR U38864 ( .A(q[29]), .B(DB[1486]), .Z(n38555) );
  XNOR U38865 ( .A(q[28]), .B(DB[1485]), .Z(n27839) );
  IV U38866 ( .A(n27852), .Z(n38553) );
  XOR U38867 ( .A(n38556), .B(n38557), .Z(n27852) );
  XNOR U38868 ( .A(n27848), .B(n27850), .Z(n38557) );
  XNOR U38869 ( .A(q[24]), .B(DB[1481]), .Z(n27850) );
  XNOR U38870 ( .A(q[27]), .B(DB[1484]), .Z(n27848) );
  IV U38871 ( .A(n27847), .Z(n38556) );
  XNOR U38872 ( .A(n27845), .B(n38558), .Z(n27847) );
  XNOR U38873 ( .A(q[26]), .B(DB[1483]), .Z(n38558) );
  XNOR U38874 ( .A(q[25]), .B(DB[1482]), .Z(n27845) );
  IV U38875 ( .A(n27860), .Z(n38552) );
  XOR U38876 ( .A(n38559), .B(n38560), .Z(n27860) );
  XNOR U38877 ( .A(n27877), .B(n27858), .Z(n38560) );
  XNOR U38878 ( .A(q[16]), .B(DB[1473]), .Z(n27858) );
  XOR U38879 ( .A(n38561), .B(n27866), .Z(n27877) );
  XNOR U38880 ( .A(q[23]), .B(DB[1480]), .Z(n27866) );
  IV U38881 ( .A(n27865), .Z(n38561) );
  XNOR U38882 ( .A(n27863), .B(n38562), .Z(n27865) );
  XNOR U38883 ( .A(q[22]), .B(DB[1479]), .Z(n38562) );
  XNOR U38884 ( .A(q[21]), .B(DB[1478]), .Z(n27863) );
  IV U38885 ( .A(n27876), .Z(n38559) );
  XOR U38886 ( .A(n38563), .B(n38564), .Z(n27876) );
  XNOR U38887 ( .A(n27872), .B(n27874), .Z(n38564) );
  XNOR U38888 ( .A(q[17]), .B(DB[1474]), .Z(n27874) );
  XNOR U38889 ( .A(q[20]), .B(DB[1477]), .Z(n27872) );
  IV U38890 ( .A(n27871), .Z(n38563) );
  XNOR U38891 ( .A(n27869), .B(n38565), .Z(n27871) );
  XNOR U38892 ( .A(q[19]), .B(DB[1476]), .Z(n38565) );
  XNOR U38893 ( .A(q[18]), .B(DB[1475]), .Z(n27869) );
  IV U38894 ( .A(n27884), .Z(n38551) );
  XOR U38895 ( .A(n38566), .B(n38567), .Z(n27884) );
  XNOR U38896 ( .A(n27911), .B(n27882), .Z(n38567) );
  XNOR U38897 ( .A(q[0]), .B(DB[1457]), .Z(n27882) );
  XOR U38898 ( .A(n38568), .B(n27903), .Z(n27911) );
  XOR U38899 ( .A(n38569), .B(n27891), .Z(n27903) );
  XNOR U38900 ( .A(q[15]), .B(DB[1472]), .Z(n27891) );
  IV U38901 ( .A(n27890), .Z(n38569) );
  XNOR U38902 ( .A(n27888), .B(n38570), .Z(n27890) );
  XNOR U38903 ( .A(q[14]), .B(DB[1471]), .Z(n38570) );
  XNOR U38904 ( .A(q[13]), .B(DB[1470]), .Z(n27888) );
  IV U38905 ( .A(n27902), .Z(n38568) );
  XOR U38906 ( .A(n38571), .B(n38572), .Z(n27902) );
  XNOR U38907 ( .A(n27898), .B(n27900), .Z(n38572) );
  XNOR U38908 ( .A(q[9]), .B(DB[1466]), .Z(n27900) );
  XNOR U38909 ( .A(q[12]), .B(DB[1469]), .Z(n27898) );
  IV U38910 ( .A(n27897), .Z(n38571) );
  XNOR U38911 ( .A(n27895), .B(n38573), .Z(n27897) );
  XNOR U38912 ( .A(q[11]), .B(DB[1468]), .Z(n38573) );
  XNOR U38913 ( .A(q[10]), .B(DB[1467]), .Z(n27895) );
  IV U38914 ( .A(n27910), .Z(n38566) );
  XOR U38915 ( .A(n38574), .B(n38575), .Z(n27910) );
  XNOR U38916 ( .A(n27927), .B(n27908), .Z(n38575) );
  XNOR U38917 ( .A(q[1]), .B(DB[1458]), .Z(n27908) );
  XOR U38918 ( .A(n38576), .B(n27916), .Z(n27927) );
  XNOR U38919 ( .A(q[8]), .B(DB[1465]), .Z(n27916) );
  IV U38920 ( .A(n27915), .Z(n38576) );
  XNOR U38921 ( .A(n27913), .B(n38577), .Z(n27915) );
  XNOR U38922 ( .A(q[7]), .B(DB[1464]), .Z(n38577) );
  XNOR U38923 ( .A(q[6]), .B(DB[1463]), .Z(n27913) );
  IV U38924 ( .A(n27926), .Z(n38574) );
  XOR U38925 ( .A(n38578), .B(n38579), .Z(n27926) );
  XNOR U38926 ( .A(n27922), .B(n27924), .Z(n38579) );
  XNOR U38927 ( .A(q[2]), .B(DB[1459]), .Z(n27924) );
  XNOR U38928 ( .A(q[5]), .B(DB[1462]), .Z(n27922) );
  IV U38929 ( .A(n27921), .Z(n38578) );
  XNOR U38930 ( .A(n27919), .B(n38580), .Z(n27921) );
  XNOR U38931 ( .A(q[4]), .B(DB[1461]), .Z(n38580) );
  XNOR U38932 ( .A(q[3]), .B(DB[1460]), .Z(n27919) );
  XOR U38933 ( .A(n38581), .B(n27688), .Z(n27539) );
  XOR U38934 ( .A(n38582), .B(n27664), .Z(n27688) );
  XOR U38935 ( .A(n38583), .B(n27656), .Z(n27664) );
  XOR U38936 ( .A(n38584), .B(n27645), .Z(n27656) );
  XNOR U38937 ( .A(q[30]), .B(DB[1518]), .Z(n27645) );
  IV U38938 ( .A(n27644), .Z(n38584) );
  XNOR U38939 ( .A(n27642), .B(n38585), .Z(n27644) );
  XNOR U38940 ( .A(q[29]), .B(DB[1517]), .Z(n38585) );
  XNOR U38941 ( .A(q[28]), .B(DB[1516]), .Z(n27642) );
  IV U38942 ( .A(n27655), .Z(n38583) );
  XOR U38943 ( .A(n38586), .B(n38587), .Z(n27655) );
  XNOR U38944 ( .A(n27651), .B(n27653), .Z(n38587) );
  XNOR U38945 ( .A(q[24]), .B(DB[1512]), .Z(n27653) );
  XNOR U38946 ( .A(q[27]), .B(DB[1515]), .Z(n27651) );
  IV U38947 ( .A(n27650), .Z(n38586) );
  XNOR U38948 ( .A(n27648), .B(n38588), .Z(n27650) );
  XNOR U38949 ( .A(q[26]), .B(DB[1514]), .Z(n38588) );
  XNOR U38950 ( .A(q[25]), .B(DB[1513]), .Z(n27648) );
  IV U38951 ( .A(n27663), .Z(n38582) );
  XOR U38952 ( .A(n38589), .B(n38590), .Z(n27663) );
  XNOR U38953 ( .A(n27680), .B(n27661), .Z(n38590) );
  XNOR U38954 ( .A(q[16]), .B(DB[1504]), .Z(n27661) );
  XOR U38955 ( .A(n38591), .B(n27669), .Z(n27680) );
  XNOR U38956 ( .A(q[23]), .B(DB[1511]), .Z(n27669) );
  IV U38957 ( .A(n27668), .Z(n38591) );
  XNOR U38958 ( .A(n27666), .B(n38592), .Z(n27668) );
  XNOR U38959 ( .A(q[22]), .B(DB[1510]), .Z(n38592) );
  XNOR U38960 ( .A(q[21]), .B(DB[1509]), .Z(n27666) );
  IV U38961 ( .A(n27679), .Z(n38589) );
  XOR U38962 ( .A(n38593), .B(n38594), .Z(n27679) );
  XNOR U38963 ( .A(n27675), .B(n27677), .Z(n38594) );
  XNOR U38964 ( .A(q[17]), .B(DB[1505]), .Z(n27677) );
  XNOR U38965 ( .A(q[20]), .B(DB[1508]), .Z(n27675) );
  IV U38966 ( .A(n27674), .Z(n38593) );
  XNOR U38967 ( .A(n27672), .B(n38595), .Z(n27674) );
  XNOR U38968 ( .A(q[19]), .B(DB[1507]), .Z(n38595) );
  XNOR U38969 ( .A(q[18]), .B(DB[1506]), .Z(n27672) );
  IV U38970 ( .A(n27687), .Z(n38581) );
  XOR U38971 ( .A(n38596), .B(n38597), .Z(n27687) );
  XNOR U38972 ( .A(n27714), .B(n27685), .Z(n38597) );
  XNOR U38973 ( .A(q[0]), .B(DB[1488]), .Z(n27685) );
  XOR U38974 ( .A(n38598), .B(n27706), .Z(n27714) );
  XOR U38975 ( .A(n38599), .B(n27694), .Z(n27706) );
  XNOR U38976 ( .A(q[15]), .B(DB[1503]), .Z(n27694) );
  IV U38977 ( .A(n27693), .Z(n38599) );
  XNOR U38978 ( .A(n27691), .B(n38600), .Z(n27693) );
  XNOR U38979 ( .A(q[14]), .B(DB[1502]), .Z(n38600) );
  XNOR U38980 ( .A(q[13]), .B(DB[1501]), .Z(n27691) );
  IV U38981 ( .A(n27705), .Z(n38598) );
  XOR U38982 ( .A(n38601), .B(n38602), .Z(n27705) );
  XNOR U38983 ( .A(n27701), .B(n27703), .Z(n38602) );
  XNOR U38984 ( .A(q[9]), .B(DB[1497]), .Z(n27703) );
  XNOR U38985 ( .A(q[12]), .B(DB[1500]), .Z(n27701) );
  IV U38986 ( .A(n27700), .Z(n38601) );
  XNOR U38987 ( .A(n27698), .B(n38603), .Z(n27700) );
  XNOR U38988 ( .A(q[11]), .B(DB[1499]), .Z(n38603) );
  XNOR U38989 ( .A(q[10]), .B(DB[1498]), .Z(n27698) );
  IV U38990 ( .A(n27713), .Z(n38596) );
  XOR U38991 ( .A(n38604), .B(n38605), .Z(n27713) );
  XNOR U38992 ( .A(n27730), .B(n27711), .Z(n38605) );
  XNOR U38993 ( .A(q[1]), .B(DB[1489]), .Z(n27711) );
  XOR U38994 ( .A(n38606), .B(n27719), .Z(n27730) );
  XNOR U38995 ( .A(q[8]), .B(DB[1496]), .Z(n27719) );
  IV U38996 ( .A(n27718), .Z(n38606) );
  XNOR U38997 ( .A(n27716), .B(n38607), .Z(n27718) );
  XNOR U38998 ( .A(q[7]), .B(DB[1495]), .Z(n38607) );
  XNOR U38999 ( .A(q[6]), .B(DB[1494]), .Z(n27716) );
  IV U39000 ( .A(n27729), .Z(n38604) );
  XOR U39001 ( .A(n38608), .B(n38609), .Z(n27729) );
  XNOR U39002 ( .A(n27725), .B(n27727), .Z(n38609) );
  XNOR U39003 ( .A(q[2]), .B(DB[1490]), .Z(n27727) );
  XNOR U39004 ( .A(q[5]), .B(DB[1493]), .Z(n27725) );
  IV U39005 ( .A(n27724), .Z(n38608) );
  XNOR U39006 ( .A(n27722), .B(n38610), .Z(n27724) );
  XNOR U39007 ( .A(q[4]), .B(DB[1492]), .Z(n38610) );
  XNOR U39008 ( .A(q[3]), .B(DB[1491]), .Z(n27722) );
  XOR U39009 ( .A(n38611), .B(n27491), .Z(n27342) );
  XOR U39010 ( .A(n38612), .B(n27467), .Z(n27491) );
  XOR U39011 ( .A(n38613), .B(n27459), .Z(n27467) );
  XOR U39012 ( .A(n38614), .B(n27448), .Z(n27459) );
  XNOR U39013 ( .A(q[30]), .B(DB[1549]), .Z(n27448) );
  IV U39014 ( .A(n27447), .Z(n38614) );
  XNOR U39015 ( .A(n27445), .B(n38615), .Z(n27447) );
  XNOR U39016 ( .A(q[29]), .B(DB[1548]), .Z(n38615) );
  XNOR U39017 ( .A(q[28]), .B(DB[1547]), .Z(n27445) );
  IV U39018 ( .A(n27458), .Z(n38613) );
  XOR U39019 ( .A(n38616), .B(n38617), .Z(n27458) );
  XNOR U39020 ( .A(n27454), .B(n27456), .Z(n38617) );
  XNOR U39021 ( .A(q[24]), .B(DB[1543]), .Z(n27456) );
  XNOR U39022 ( .A(q[27]), .B(DB[1546]), .Z(n27454) );
  IV U39023 ( .A(n27453), .Z(n38616) );
  XNOR U39024 ( .A(n27451), .B(n38618), .Z(n27453) );
  XNOR U39025 ( .A(q[26]), .B(DB[1545]), .Z(n38618) );
  XNOR U39026 ( .A(q[25]), .B(DB[1544]), .Z(n27451) );
  IV U39027 ( .A(n27466), .Z(n38612) );
  XOR U39028 ( .A(n38619), .B(n38620), .Z(n27466) );
  XNOR U39029 ( .A(n27483), .B(n27464), .Z(n38620) );
  XNOR U39030 ( .A(q[16]), .B(DB[1535]), .Z(n27464) );
  XOR U39031 ( .A(n38621), .B(n27472), .Z(n27483) );
  XNOR U39032 ( .A(q[23]), .B(DB[1542]), .Z(n27472) );
  IV U39033 ( .A(n27471), .Z(n38621) );
  XNOR U39034 ( .A(n27469), .B(n38622), .Z(n27471) );
  XNOR U39035 ( .A(q[22]), .B(DB[1541]), .Z(n38622) );
  XNOR U39036 ( .A(q[21]), .B(DB[1540]), .Z(n27469) );
  IV U39037 ( .A(n27482), .Z(n38619) );
  XOR U39038 ( .A(n38623), .B(n38624), .Z(n27482) );
  XNOR U39039 ( .A(n27478), .B(n27480), .Z(n38624) );
  XNOR U39040 ( .A(q[17]), .B(DB[1536]), .Z(n27480) );
  XNOR U39041 ( .A(q[20]), .B(DB[1539]), .Z(n27478) );
  IV U39042 ( .A(n27477), .Z(n38623) );
  XNOR U39043 ( .A(n27475), .B(n38625), .Z(n27477) );
  XNOR U39044 ( .A(q[19]), .B(DB[1538]), .Z(n38625) );
  XNOR U39045 ( .A(q[18]), .B(DB[1537]), .Z(n27475) );
  IV U39046 ( .A(n27490), .Z(n38611) );
  XOR U39047 ( .A(n38626), .B(n38627), .Z(n27490) );
  XNOR U39048 ( .A(n27517), .B(n27488), .Z(n38627) );
  XNOR U39049 ( .A(q[0]), .B(DB[1519]), .Z(n27488) );
  XOR U39050 ( .A(n38628), .B(n27509), .Z(n27517) );
  XOR U39051 ( .A(n38629), .B(n27497), .Z(n27509) );
  XNOR U39052 ( .A(q[15]), .B(DB[1534]), .Z(n27497) );
  IV U39053 ( .A(n27496), .Z(n38629) );
  XNOR U39054 ( .A(n27494), .B(n38630), .Z(n27496) );
  XNOR U39055 ( .A(q[14]), .B(DB[1533]), .Z(n38630) );
  XNOR U39056 ( .A(q[13]), .B(DB[1532]), .Z(n27494) );
  IV U39057 ( .A(n27508), .Z(n38628) );
  XOR U39058 ( .A(n38631), .B(n38632), .Z(n27508) );
  XNOR U39059 ( .A(n27504), .B(n27506), .Z(n38632) );
  XNOR U39060 ( .A(q[9]), .B(DB[1528]), .Z(n27506) );
  XNOR U39061 ( .A(q[12]), .B(DB[1531]), .Z(n27504) );
  IV U39062 ( .A(n27503), .Z(n38631) );
  XNOR U39063 ( .A(n27501), .B(n38633), .Z(n27503) );
  XNOR U39064 ( .A(q[11]), .B(DB[1530]), .Z(n38633) );
  XNOR U39065 ( .A(q[10]), .B(DB[1529]), .Z(n27501) );
  IV U39066 ( .A(n27516), .Z(n38626) );
  XOR U39067 ( .A(n38634), .B(n38635), .Z(n27516) );
  XNOR U39068 ( .A(n27533), .B(n27514), .Z(n38635) );
  XNOR U39069 ( .A(q[1]), .B(DB[1520]), .Z(n27514) );
  XOR U39070 ( .A(n38636), .B(n27522), .Z(n27533) );
  XNOR U39071 ( .A(q[8]), .B(DB[1527]), .Z(n27522) );
  IV U39072 ( .A(n27521), .Z(n38636) );
  XNOR U39073 ( .A(n27519), .B(n38637), .Z(n27521) );
  XNOR U39074 ( .A(q[7]), .B(DB[1526]), .Z(n38637) );
  XNOR U39075 ( .A(q[6]), .B(DB[1525]), .Z(n27519) );
  IV U39076 ( .A(n27532), .Z(n38634) );
  XOR U39077 ( .A(n38638), .B(n38639), .Z(n27532) );
  XNOR U39078 ( .A(n27528), .B(n27530), .Z(n38639) );
  XNOR U39079 ( .A(q[2]), .B(DB[1521]), .Z(n27530) );
  XNOR U39080 ( .A(q[5]), .B(DB[1524]), .Z(n27528) );
  IV U39081 ( .A(n27527), .Z(n38638) );
  XNOR U39082 ( .A(n27525), .B(n38640), .Z(n27527) );
  XNOR U39083 ( .A(q[4]), .B(DB[1523]), .Z(n38640) );
  XNOR U39084 ( .A(q[3]), .B(DB[1522]), .Z(n27525) );
  XOR U39085 ( .A(n38641), .B(n27294), .Z(n27145) );
  XOR U39086 ( .A(n38642), .B(n27270), .Z(n27294) );
  XOR U39087 ( .A(n38643), .B(n27262), .Z(n27270) );
  XOR U39088 ( .A(n38644), .B(n27251), .Z(n27262) );
  XNOR U39089 ( .A(q[30]), .B(DB[1580]), .Z(n27251) );
  IV U39090 ( .A(n27250), .Z(n38644) );
  XNOR U39091 ( .A(n27248), .B(n38645), .Z(n27250) );
  XNOR U39092 ( .A(q[29]), .B(DB[1579]), .Z(n38645) );
  XNOR U39093 ( .A(q[28]), .B(DB[1578]), .Z(n27248) );
  IV U39094 ( .A(n27261), .Z(n38643) );
  XOR U39095 ( .A(n38646), .B(n38647), .Z(n27261) );
  XNOR U39096 ( .A(n27257), .B(n27259), .Z(n38647) );
  XNOR U39097 ( .A(q[24]), .B(DB[1574]), .Z(n27259) );
  XNOR U39098 ( .A(q[27]), .B(DB[1577]), .Z(n27257) );
  IV U39099 ( .A(n27256), .Z(n38646) );
  XNOR U39100 ( .A(n27254), .B(n38648), .Z(n27256) );
  XNOR U39101 ( .A(q[26]), .B(DB[1576]), .Z(n38648) );
  XNOR U39102 ( .A(q[25]), .B(DB[1575]), .Z(n27254) );
  IV U39103 ( .A(n27269), .Z(n38642) );
  XOR U39104 ( .A(n38649), .B(n38650), .Z(n27269) );
  XNOR U39105 ( .A(n27286), .B(n27267), .Z(n38650) );
  XNOR U39106 ( .A(q[16]), .B(DB[1566]), .Z(n27267) );
  XOR U39107 ( .A(n38651), .B(n27275), .Z(n27286) );
  XNOR U39108 ( .A(q[23]), .B(DB[1573]), .Z(n27275) );
  IV U39109 ( .A(n27274), .Z(n38651) );
  XNOR U39110 ( .A(n27272), .B(n38652), .Z(n27274) );
  XNOR U39111 ( .A(q[22]), .B(DB[1572]), .Z(n38652) );
  XNOR U39112 ( .A(q[21]), .B(DB[1571]), .Z(n27272) );
  IV U39113 ( .A(n27285), .Z(n38649) );
  XOR U39114 ( .A(n38653), .B(n38654), .Z(n27285) );
  XNOR U39115 ( .A(n27281), .B(n27283), .Z(n38654) );
  XNOR U39116 ( .A(q[17]), .B(DB[1567]), .Z(n27283) );
  XNOR U39117 ( .A(q[20]), .B(DB[1570]), .Z(n27281) );
  IV U39118 ( .A(n27280), .Z(n38653) );
  XNOR U39119 ( .A(n27278), .B(n38655), .Z(n27280) );
  XNOR U39120 ( .A(q[19]), .B(DB[1569]), .Z(n38655) );
  XNOR U39121 ( .A(q[18]), .B(DB[1568]), .Z(n27278) );
  IV U39122 ( .A(n27293), .Z(n38641) );
  XOR U39123 ( .A(n38656), .B(n38657), .Z(n27293) );
  XNOR U39124 ( .A(n27320), .B(n27291), .Z(n38657) );
  XNOR U39125 ( .A(q[0]), .B(DB[1550]), .Z(n27291) );
  XOR U39126 ( .A(n38658), .B(n27312), .Z(n27320) );
  XOR U39127 ( .A(n38659), .B(n27300), .Z(n27312) );
  XNOR U39128 ( .A(q[15]), .B(DB[1565]), .Z(n27300) );
  IV U39129 ( .A(n27299), .Z(n38659) );
  XNOR U39130 ( .A(n27297), .B(n38660), .Z(n27299) );
  XNOR U39131 ( .A(q[14]), .B(DB[1564]), .Z(n38660) );
  XNOR U39132 ( .A(q[13]), .B(DB[1563]), .Z(n27297) );
  IV U39133 ( .A(n27311), .Z(n38658) );
  XOR U39134 ( .A(n38661), .B(n38662), .Z(n27311) );
  XNOR U39135 ( .A(n27307), .B(n27309), .Z(n38662) );
  XNOR U39136 ( .A(q[9]), .B(DB[1559]), .Z(n27309) );
  XNOR U39137 ( .A(q[12]), .B(DB[1562]), .Z(n27307) );
  IV U39138 ( .A(n27306), .Z(n38661) );
  XNOR U39139 ( .A(n27304), .B(n38663), .Z(n27306) );
  XNOR U39140 ( .A(q[11]), .B(DB[1561]), .Z(n38663) );
  XNOR U39141 ( .A(q[10]), .B(DB[1560]), .Z(n27304) );
  IV U39142 ( .A(n27319), .Z(n38656) );
  XOR U39143 ( .A(n38664), .B(n38665), .Z(n27319) );
  XNOR U39144 ( .A(n27336), .B(n27317), .Z(n38665) );
  XNOR U39145 ( .A(q[1]), .B(DB[1551]), .Z(n27317) );
  XOR U39146 ( .A(n38666), .B(n27325), .Z(n27336) );
  XNOR U39147 ( .A(q[8]), .B(DB[1558]), .Z(n27325) );
  IV U39148 ( .A(n27324), .Z(n38666) );
  XNOR U39149 ( .A(n27322), .B(n38667), .Z(n27324) );
  XNOR U39150 ( .A(q[7]), .B(DB[1557]), .Z(n38667) );
  XNOR U39151 ( .A(q[6]), .B(DB[1556]), .Z(n27322) );
  IV U39152 ( .A(n27335), .Z(n38664) );
  XOR U39153 ( .A(n38668), .B(n38669), .Z(n27335) );
  XNOR U39154 ( .A(n27331), .B(n27333), .Z(n38669) );
  XNOR U39155 ( .A(q[2]), .B(DB[1552]), .Z(n27333) );
  XNOR U39156 ( .A(q[5]), .B(DB[1555]), .Z(n27331) );
  IV U39157 ( .A(n27330), .Z(n38668) );
  XNOR U39158 ( .A(n27328), .B(n38670), .Z(n27330) );
  XNOR U39159 ( .A(q[4]), .B(DB[1554]), .Z(n38670) );
  XNOR U39160 ( .A(q[3]), .B(DB[1553]), .Z(n27328) );
  XOR U39161 ( .A(n38671), .B(n27097), .Z(n26948) );
  XOR U39162 ( .A(n38672), .B(n27073), .Z(n27097) );
  XOR U39163 ( .A(n38673), .B(n27065), .Z(n27073) );
  XOR U39164 ( .A(n38674), .B(n27054), .Z(n27065) );
  XNOR U39165 ( .A(q[30]), .B(DB[1611]), .Z(n27054) );
  IV U39166 ( .A(n27053), .Z(n38674) );
  XNOR U39167 ( .A(n27051), .B(n38675), .Z(n27053) );
  XNOR U39168 ( .A(q[29]), .B(DB[1610]), .Z(n38675) );
  XNOR U39169 ( .A(q[28]), .B(DB[1609]), .Z(n27051) );
  IV U39170 ( .A(n27064), .Z(n38673) );
  XOR U39171 ( .A(n38676), .B(n38677), .Z(n27064) );
  XNOR U39172 ( .A(n27060), .B(n27062), .Z(n38677) );
  XNOR U39173 ( .A(q[24]), .B(DB[1605]), .Z(n27062) );
  XNOR U39174 ( .A(q[27]), .B(DB[1608]), .Z(n27060) );
  IV U39175 ( .A(n27059), .Z(n38676) );
  XNOR U39176 ( .A(n27057), .B(n38678), .Z(n27059) );
  XNOR U39177 ( .A(q[26]), .B(DB[1607]), .Z(n38678) );
  XNOR U39178 ( .A(q[25]), .B(DB[1606]), .Z(n27057) );
  IV U39179 ( .A(n27072), .Z(n38672) );
  XOR U39180 ( .A(n38679), .B(n38680), .Z(n27072) );
  XNOR U39181 ( .A(n27089), .B(n27070), .Z(n38680) );
  XNOR U39182 ( .A(q[16]), .B(DB[1597]), .Z(n27070) );
  XOR U39183 ( .A(n38681), .B(n27078), .Z(n27089) );
  XNOR U39184 ( .A(q[23]), .B(DB[1604]), .Z(n27078) );
  IV U39185 ( .A(n27077), .Z(n38681) );
  XNOR U39186 ( .A(n27075), .B(n38682), .Z(n27077) );
  XNOR U39187 ( .A(q[22]), .B(DB[1603]), .Z(n38682) );
  XNOR U39188 ( .A(q[21]), .B(DB[1602]), .Z(n27075) );
  IV U39189 ( .A(n27088), .Z(n38679) );
  XOR U39190 ( .A(n38683), .B(n38684), .Z(n27088) );
  XNOR U39191 ( .A(n27084), .B(n27086), .Z(n38684) );
  XNOR U39192 ( .A(q[17]), .B(DB[1598]), .Z(n27086) );
  XNOR U39193 ( .A(q[20]), .B(DB[1601]), .Z(n27084) );
  IV U39194 ( .A(n27083), .Z(n38683) );
  XNOR U39195 ( .A(n27081), .B(n38685), .Z(n27083) );
  XNOR U39196 ( .A(q[19]), .B(DB[1600]), .Z(n38685) );
  XNOR U39197 ( .A(q[18]), .B(DB[1599]), .Z(n27081) );
  IV U39198 ( .A(n27096), .Z(n38671) );
  XOR U39199 ( .A(n38686), .B(n38687), .Z(n27096) );
  XNOR U39200 ( .A(n27123), .B(n27094), .Z(n38687) );
  XNOR U39201 ( .A(q[0]), .B(DB[1581]), .Z(n27094) );
  XOR U39202 ( .A(n38688), .B(n27115), .Z(n27123) );
  XOR U39203 ( .A(n38689), .B(n27103), .Z(n27115) );
  XNOR U39204 ( .A(q[15]), .B(DB[1596]), .Z(n27103) );
  IV U39205 ( .A(n27102), .Z(n38689) );
  XNOR U39206 ( .A(n27100), .B(n38690), .Z(n27102) );
  XNOR U39207 ( .A(q[14]), .B(DB[1595]), .Z(n38690) );
  XNOR U39208 ( .A(q[13]), .B(DB[1594]), .Z(n27100) );
  IV U39209 ( .A(n27114), .Z(n38688) );
  XOR U39210 ( .A(n38691), .B(n38692), .Z(n27114) );
  XNOR U39211 ( .A(n27110), .B(n27112), .Z(n38692) );
  XNOR U39212 ( .A(q[9]), .B(DB[1590]), .Z(n27112) );
  XNOR U39213 ( .A(q[12]), .B(DB[1593]), .Z(n27110) );
  IV U39214 ( .A(n27109), .Z(n38691) );
  XNOR U39215 ( .A(n27107), .B(n38693), .Z(n27109) );
  XNOR U39216 ( .A(q[11]), .B(DB[1592]), .Z(n38693) );
  XNOR U39217 ( .A(q[10]), .B(DB[1591]), .Z(n27107) );
  IV U39218 ( .A(n27122), .Z(n38686) );
  XOR U39219 ( .A(n38694), .B(n38695), .Z(n27122) );
  XNOR U39220 ( .A(n27139), .B(n27120), .Z(n38695) );
  XNOR U39221 ( .A(q[1]), .B(DB[1582]), .Z(n27120) );
  XOR U39222 ( .A(n38696), .B(n27128), .Z(n27139) );
  XNOR U39223 ( .A(q[8]), .B(DB[1589]), .Z(n27128) );
  IV U39224 ( .A(n27127), .Z(n38696) );
  XNOR U39225 ( .A(n27125), .B(n38697), .Z(n27127) );
  XNOR U39226 ( .A(q[7]), .B(DB[1588]), .Z(n38697) );
  XNOR U39227 ( .A(q[6]), .B(DB[1587]), .Z(n27125) );
  IV U39228 ( .A(n27138), .Z(n38694) );
  XOR U39229 ( .A(n38698), .B(n38699), .Z(n27138) );
  XNOR U39230 ( .A(n27134), .B(n27136), .Z(n38699) );
  XNOR U39231 ( .A(q[2]), .B(DB[1583]), .Z(n27136) );
  XNOR U39232 ( .A(q[5]), .B(DB[1586]), .Z(n27134) );
  IV U39233 ( .A(n27133), .Z(n38698) );
  XNOR U39234 ( .A(n27131), .B(n38700), .Z(n27133) );
  XNOR U39235 ( .A(q[4]), .B(DB[1585]), .Z(n38700) );
  XNOR U39236 ( .A(q[3]), .B(DB[1584]), .Z(n27131) );
  XOR U39237 ( .A(n38701), .B(n26900), .Z(n26751) );
  XOR U39238 ( .A(n38702), .B(n26876), .Z(n26900) );
  XOR U39239 ( .A(n38703), .B(n26868), .Z(n26876) );
  XOR U39240 ( .A(n38704), .B(n26857), .Z(n26868) );
  XNOR U39241 ( .A(q[30]), .B(DB[1642]), .Z(n26857) );
  IV U39242 ( .A(n26856), .Z(n38704) );
  XNOR U39243 ( .A(n26854), .B(n38705), .Z(n26856) );
  XNOR U39244 ( .A(q[29]), .B(DB[1641]), .Z(n38705) );
  XNOR U39245 ( .A(q[28]), .B(DB[1640]), .Z(n26854) );
  IV U39246 ( .A(n26867), .Z(n38703) );
  XOR U39247 ( .A(n38706), .B(n38707), .Z(n26867) );
  XNOR U39248 ( .A(n26863), .B(n26865), .Z(n38707) );
  XNOR U39249 ( .A(q[24]), .B(DB[1636]), .Z(n26865) );
  XNOR U39250 ( .A(q[27]), .B(DB[1639]), .Z(n26863) );
  IV U39251 ( .A(n26862), .Z(n38706) );
  XNOR U39252 ( .A(n26860), .B(n38708), .Z(n26862) );
  XNOR U39253 ( .A(q[26]), .B(DB[1638]), .Z(n38708) );
  XNOR U39254 ( .A(q[25]), .B(DB[1637]), .Z(n26860) );
  IV U39255 ( .A(n26875), .Z(n38702) );
  XOR U39256 ( .A(n38709), .B(n38710), .Z(n26875) );
  XNOR U39257 ( .A(n26892), .B(n26873), .Z(n38710) );
  XNOR U39258 ( .A(q[16]), .B(DB[1628]), .Z(n26873) );
  XOR U39259 ( .A(n38711), .B(n26881), .Z(n26892) );
  XNOR U39260 ( .A(q[23]), .B(DB[1635]), .Z(n26881) );
  IV U39261 ( .A(n26880), .Z(n38711) );
  XNOR U39262 ( .A(n26878), .B(n38712), .Z(n26880) );
  XNOR U39263 ( .A(q[22]), .B(DB[1634]), .Z(n38712) );
  XNOR U39264 ( .A(q[21]), .B(DB[1633]), .Z(n26878) );
  IV U39265 ( .A(n26891), .Z(n38709) );
  XOR U39266 ( .A(n38713), .B(n38714), .Z(n26891) );
  XNOR U39267 ( .A(n26887), .B(n26889), .Z(n38714) );
  XNOR U39268 ( .A(q[17]), .B(DB[1629]), .Z(n26889) );
  XNOR U39269 ( .A(q[20]), .B(DB[1632]), .Z(n26887) );
  IV U39270 ( .A(n26886), .Z(n38713) );
  XNOR U39271 ( .A(n26884), .B(n38715), .Z(n26886) );
  XNOR U39272 ( .A(q[19]), .B(DB[1631]), .Z(n38715) );
  XNOR U39273 ( .A(q[18]), .B(DB[1630]), .Z(n26884) );
  IV U39274 ( .A(n26899), .Z(n38701) );
  XOR U39275 ( .A(n38716), .B(n38717), .Z(n26899) );
  XNOR U39276 ( .A(n26926), .B(n26897), .Z(n38717) );
  XNOR U39277 ( .A(q[0]), .B(DB[1612]), .Z(n26897) );
  XOR U39278 ( .A(n38718), .B(n26918), .Z(n26926) );
  XOR U39279 ( .A(n38719), .B(n26906), .Z(n26918) );
  XNOR U39280 ( .A(q[15]), .B(DB[1627]), .Z(n26906) );
  IV U39281 ( .A(n26905), .Z(n38719) );
  XNOR U39282 ( .A(n26903), .B(n38720), .Z(n26905) );
  XNOR U39283 ( .A(q[14]), .B(DB[1626]), .Z(n38720) );
  XNOR U39284 ( .A(q[13]), .B(DB[1625]), .Z(n26903) );
  IV U39285 ( .A(n26917), .Z(n38718) );
  XOR U39286 ( .A(n38721), .B(n38722), .Z(n26917) );
  XNOR U39287 ( .A(n26913), .B(n26915), .Z(n38722) );
  XNOR U39288 ( .A(q[9]), .B(DB[1621]), .Z(n26915) );
  XNOR U39289 ( .A(q[12]), .B(DB[1624]), .Z(n26913) );
  IV U39290 ( .A(n26912), .Z(n38721) );
  XNOR U39291 ( .A(n26910), .B(n38723), .Z(n26912) );
  XNOR U39292 ( .A(q[11]), .B(DB[1623]), .Z(n38723) );
  XNOR U39293 ( .A(q[10]), .B(DB[1622]), .Z(n26910) );
  IV U39294 ( .A(n26925), .Z(n38716) );
  XOR U39295 ( .A(n38724), .B(n38725), .Z(n26925) );
  XNOR U39296 ( .A(n26942), .B(n26923), .Z(n38725) );
  XNOR U39297 ( .A(q[1]), .B(DB[1613]), .Z(n26923) );
  XOR U39298 ( .A(n38726), .B(n26931), .Z(n26942) );
  XNOR U39299 ( .A(q[8]), .B(DB[1620]), .Z(n26931) );
  IV U39300 ( .A(n26930), .Z(n38726) );
  XNOR U39301 ( .A(n26928), .B(n38727), .Z(n26930) );
  XNOR U39302 ( .A(q[7]), .B(DB[1619]), .Z(n38727) );
  XNOR U39303 ( .A(q[6]), .B(DB[1618]), .Z(n26928) );
  IV U39304 ( .A(n26941), .Z(n38724) );
  XOR U39305 ( .A(n38728), .B(n38729), .Z(n26941) );
  XNOR U39306 ( .A(n26937), .B(n26939), .Z(n38729) );
  XNOR U39307 ( .A(q[2]), .B(DB[1614]), .Z(n26939) );
  XNOR U39308 ( .A(q[5]), .B(DB[1617]), .Z(n26937) );
  IV U39309 ( .A(n26936), .Z(n38728) );
  XNOR U39310 ( .A(n26934), .B(n38730), .Z(n26936) );
  XNOR U39311 ( .A(q[4]), .B(DB[1616]), .Z(n38730) );
  XNOR U39312 ( .A(q[3]), .B(DB[1615]), .Z(n26934) );
  XOR U39313 ( .A(n38731), .B(n26703), .Z(n26554) );
  XOR U39314 ( .A(n38732), .B(n26679), .Z(n26703) );
  XOR U39315 ( .A(n38733), .B(n26671), .Z(n26679) );
  XOR U39316 ( .A(n38734), .B(n26660), .Z(n26671) );
  XNOR U39317 ( .A(q[30]), .B(DB[1673]), .Z(n26660) );
  IV U39318 ( .A(n26659), .Z(n38734) );
  XNOR U39319 ( .A(n26657), .B(n38735), .Z(n26659) );
  XNOR U39320 ( .A(q[29]), .B(DB[1672]), .Z(n38735) );
  XNOR U39321 ( .A(q[28]), .B(DB[1671]), .Z(n26657) );
  IV U39322 ( .A(n26670), .Z(n38733) );
  XOR U39323 ( .A(n38736), .B(n38737), .Z(n26670) );
  XNOR U39324 ( .A(n26666), .B(n26668), .Z(n38737) );
  XNOR U39325 ( .A(q[24]), .B(DB[1667]), .Z(n26668) );
  XNOR U39326 ( .A(q[27]), .B(DB[1670]), .Z(n26666) );
  IV U39327 ( .A(n26665), .Z(n38736) );
  XNOR U39328 ( .A(n26663), .B(n38738), .Z(n26665) );
  XNOR U39329 ( .A(q[26]), .B(DB[1669]), .Z(n38738) );
  XNOR U39330 ( .A(q[25]), .B(DB[1668]), .Z(n26663) );
  IV U39331 ( .A(n26678), .Z(n38732) );
  XOR U39332 ( .A(n38739), .B(n38740), .Z(n26678) );
  XNOR U39333 ( .A(n26695), .B(n26676), .Z(n38740) );
  XNOR U39334 ( .A(q[16]), .B(DB[1659]), .Z(n26676) );
  XOR U39335 ( .A(n38741), .B(n26684), .Z(n26695) );
  XNOR U39336 ( .A(q[23]), .B(DB[1666]), .Z(n26684) );
  IV U39337 ( .A(n26683), .Z(n38741) );
  XNOR U39338 ( .A(n26681), .B(n38742), .Z(n26683) );
  XNOR U39339 ( .A(q[22]), .B(DB[1665]), .Z(n38742) );
  XNOR U39340 ( .A(q[21]), .B(DB[1664]), .Z(n26681) );
  IV U39341 ( .A(n26694), .Z(n38739) );
  XOR U39342 ( .A(n38743), .B(n38744), .Z(n26694) );
  XNOR U39343 ( .A(n26690), .B(n26692), .Z(n38744) );
  XNOR U39344 ( .A(q[17]), .B(DB[1660]), .Z(n26692) );
  XNOR U39345 ( .A(q[20]), .B(DB[1663]), .Z(n26690) );
  IV U39346 ( .A(n26689), .Z(n38743) );
  XNOR U39347 ( .A(n26687), .B(n38745), .Z(n26689) );
  XNOR U39348 ( .A(q[19]), .B(DB[1662]), .Z(n38745) );
  XNOR U39349 ( .A(q[18]), .B(DB[1661]), .Z(n26687) );
  IV U39350 ( .A(n26702), .Z(n38731) );
  XOR U39351 ( .A(n38746), .B(n38747), .Z(n26702) );
  XNOR U39352 ( .A(n26729), .B(n26700), .Z(n38747) );
  XNOR U39353 ( .A(q[0]), .B(DB[1643]), .Z(n26700) );
  XOR U39354 ( .A(n38748), .B(n26721), .Z(n26729) );
  XOR U39355 ( .A(n38749), .B(n26709), .Z(n26721) );
  XNOR U39356 ( .A(q[15]), .B(DB[1658]), .Z(n26709) );
  IV U39357 ( .A(n26708), .Z(n38749) );
  XNOR U39358 ( .A(n26706), .B(n38750), .Z(n26708) );
  XNOR U39359 ( .A(q[14]), .B(DB[1657]), .Z(n38750) );
  XNOR U39360 ( .A(q[13]), .B(DB[1656]), .Z(n26706) );
  IV U39361 ( .A(n26720), .Z(n38748) );
  XOR U39362 ( .A(n38751), .B(n38752), .Z(n26720) );
  XNOR U39363 ( .A(n26716), .B(n26718), .Z(n38752) );
  XNOR U39364 ( .A(q[9]), .B(DB[1652]), .Z(n26718) );
  XNOR U39365 ( .A(q[12]), .B(DB[1655]), .Z(n26716) );
  IV U39366 ( .A(n26715), .Z(n38751) );
  XNOR U39367 ( .A(n26713), .B(n38753), .Z(n26715) );
  XNOR U39368 ( .A(q[11]), .B(DB[1654]), .Z(n38753) );
  XNOR U39369 ( .A(q[10]), .B(DB[1653]), .Z(n26713) );
  IV U39370 ( .A(n26728), .Z(n38746) );
  XOR U39371 ( .A(n38754), .B(n38755), .Z(n26728) );
  XNOR U39372 ( .A(n26745), .B(n26726), .Z(n38755) );
  XNOR U39373 ( .A(q[1]), .B(DB[1644]), .Z(n26726) );
  XOR U39374 ( .A(n38756), .B(n26734), .Z(n26745) );
  XNOR U39375 ( .A(q[8]), .B(DB[1651]), .Z(n26734) );
  IV U39376 ( .A(n26733), .Z(n38756) );
  XNOR U39377 ( .A(n26731), .B(n38757), .Z(n26733) );
  XNOR U39378 ( .A(q[7]), .B(DB[1650]), .Z(n38757) );
  XNOR U39379 ( .A(q[6]), .B(DB[1649]), .Z(n26731) );
  IV U39380 ( .A(n26744), .Z(n38754) );
  XOR U39381 ( .A(n38758), .B(n38759), .Z(n26744) );
  XNOR U39382 ( .A(n26740), .B(n26742), .Z(n38759) );
  XNOR U39383 ( .A(q[2]), .B(DB[1645]), .Z(n26742) );
  XNOR U39384 ( .A(q[5]), .B(DB[1648]), .Z(n26740) );
  IV U39385 ( .A(n26739), .Z(n38758) );
  XNOR U39386 ( .A(n26737), .B(n38760), .Z(n26739) );
  XNOR U39387 ( .A(q[4]), .B(DB[1647]), .Z(n38760) );
  XNOR U39388 ( .A(q[3]), .B(DB[1646]), .Z(n26737) );
  XOR U39389 ( .A(n38761), .B(n26506), .Z(n26357) );
  XOR U39390 ( .A(n38762), .B(n26482), .Z(n26506) );
  XOR U39391 ( .A(n38763), .B(n26474), .Z(n26482) );
  XOR U39392 ( .A(n38764), .B(n26463), .Z(n26474) );
  XNOR U39393 ( .A(q[30]), .B(DB[1704]), .Z(n26463) );
  IV U39394 ( .A(n26462), .Z(n38764) );
  XNOR U39395 ( .A(n26460), .B(n38765), .Z(n26462) );
  XNOR U39396 ( .A(q[29]), .B(DB[1703]), .Z(n38765) );
  XNOR U39397 ( .A(q[28]), .B(DB[1702]), .Z(n26460) );
  IV U39398 ( .A(n26473), .Z(n38763) );
  XOR U39399 ( .A(n38766), .B(n38767), .Z(n26473) );
  XNOR U39400 ( .A(n26469), .B(n26471), .Z(n38767) );
  XNOR U39401 ( .A(q[24]), .B(DB[1698]), .Z(n26471) );
  XNOR U39402 ( .A(q[27]), .B(DB[1701]), .Z(n26469) );
  IV U39403 ( .A(n26468), .Z(n38766) );
  XNOR U39404 ( .A(n26466), .B(n38768), .Z(n26468) );
  XNOR U39405 ( .A(q[26]), .B(DB[1700]), .Z(n38768) );
  XNOR U39406 ( .A(q[25]), .B(DB[1699]), .Z(n26466) );
  IV U39407 ( .A(n26481), .Z(n38762) );
  XOR U39408 ( .A(n38769), .B(n38770), .Z(n26481) );
  XNOR U39409 ( .A(n26498), .B(n26479), .Z(n38770) );
  XNOR U39410 ( .A(q[16]), .B(DB[1690]), .Z(n26479) );
  XOR U39411 ( .A(n38771), .B(n26487), .Z(n26498) );
  XNOR U39412 ( .A(q[23]), .B(DB[1697]), .Z(n26487) );
  IV U39413 ( .A(n26486), .Z(n38771) );
  XNOR U39414 ( .A(n26484), .B(n38772), .Z(n26486) );
  XNOR U39415 ( .A(q[22]), .B(DB[1696]), .Z(n38772) );
  XNOR U39416 ( .A(q[21]), .B(DB[1695]), .Z(n26484) );
  IV U39417 ( .A(n26497), .Z(n38769) );
  XOR U39418 ( .A(n38773), .B(n38774), .Z(n26497) );
  XNOR U39419 ( .A(n26493), .B(n26495), .Z(n38774) );
  XNOR U39420 ( .A(q[17]), .B(DB[1691]), .Z(n26495) );
  XNOR U39421 ( .A(q[20]), .B(DB[1694]), .Z(n26493) );
  IV U39422 ( .A(n26492), .Z(n38773) );
  XNOR U39423 ( .A(n26490), .B(n38775), .Z(n26492) );
  XNOR U39424 ( .A(q[19]), .B(DB[1693]), .Z(n38775) );
  XNOR U39425 ( .A(q[18]), .B(DB[1692]), .Z(n26490) );
  IV U39426 ( .A(n26505), .Z(n38761) );
  XOR U39427 ( .A(n38776), .B(n38777), .Z(n26505) );
  XNOR U39428 ( .A(n26532), .B(n26503), .Z(n38777) );
  XNOR U39429 ( .A(q[0]), .B(DB[1674]), .Z(n26503) );
  XOR U39430 ( .A(n38778), .B(n26524), .Z(n26532) );
  XOR U39431 ( .A(n38779), .B(n26512), .Z(n26524) );
  XNOR U39432 ( .A(q[15]), .B(DB[1689]), .Z(n26512) );
  IV U39433 ( .A(n26511), .Z(n38779) );
  XNOR U39434 ( .A(n26509), .B(n38780), .Z(n26511) );
  XNOR U39435 ( .A(q[14]), .B(DB[1688]), .Z(n38780) );
  XNOR U39436 ( .A(q[13]), .B(DB[1687]), .Z(n26509) );
  IV U39437 ( .A(n26523), .Z(n38778) );
  XOR U39438 ( .A(n38781), .B(n38782), .Z(n26523) );
  XNOR U39439 ( .A(n26519), .B(n26521), .Z(n38782) );
  XNOR U39440 ( .A(q[9]), .B(DB[1683]), .Z(n26521) );
  XNOR U39441 ( .A(q[12]), .B(DB[1686]), .Z(n26519) );
  IV U39442 ( .A(n26518), .Z(n38781) );
  XNOR U39443 ( .A(n26516), .B(n38783), .Z(n26518) );
  XNOR U39444 ( .A(q[11]), .B(DB[1685]), .Z(n38783) );
  XNOR U39445 ( .A(q[10]), .B(DB[1684]), .Z(n26516) );
  IV U39446 ( .A(n26531), .Z(n38776) );
  XOR U39447 ( .A(n38784), .B(n38785), .Z(n26531) );
  XNOR U39448 ( .A(n26548), .B(n26529), .Z(n38785) );
  XNOR U39449 ( .A(q[1]), .B(DB[1675]), .Z(n26529) );
  XOR U39450 ( .A(n38786), .B(n26537), .Z(n26548) );
  XNOR U39451 ( .A(q[8]), .B(DB[1682]), .Z(n26537) );
  IV U39452 ( .A(n26536), .Z(n38786) );
  XNOR U39453 ( .A(n26534), .B(n38787), .Z(n26536) );
  XNOR U39454 ( .A(q[7]), .B(DB[1681]), .Z(n38787) );
  XNOR U39455 ( .A(q[6]), .B(DB[1680]), .Z(n26534) );
  IV U39456 ( .A(n26547), .Z(n38784) );
  XOR U39457 ( .A(n38788), .B(n38789), .Z(n26547) );
  XNOR U39458 ( .A(n26543), .B(n26545), .Z(n38789) );
  XNOR U39459 ( .A(q[2]), .B(DB[1676]), .Z(n26545) );
  XNOR U39460 ( .A(q[5]), .B(DB[1679]), .Z(n26543) );
  IV U39461 ( .A(n26542), .Z(n38788) );
  XNOR U39462 ( .A(n26540), .B(n38790), .Z(n26542) );
  XNOR U39463 ( .A(q[4]), .B(DB[1678]), .Z(n38790) );
  XNOR U39464 ( .A(q[3]), .B(DB[1677]), .Z(n26540) );
  XOR U39465 ( .A(n38791), .B(n26309), .Z(n26160) );
  XOR U39466 ( .A(n38792), .B(n26285), .Z(n26309) );
  XOR U39467 ( .A(n38793), .B(n26277), .Z(n26285) );
  XOR U39468 ( .A(n38794), .B(n26266), .Z(n26277) );
  XNOR U39469 ( .A(q[30]), .B(DB[1735]), .Z(n26266) );
  IV U39470 ( .A(n26265), .Z(n38794) );
  XNOR U39471 ( .A(n26263), .B(n38795), .Z(n26265) );
  XNOR U39472 ( .A(q[29]), .B(DB[1734]), .Z(n38795) );
  XNOR U39473 ( .A(q[28]), .B(DB[1733]), .Z(n26263) );
  IV U39474 ( .A(n26276), .Z(n38793) );
  XOR U39475 ( .A(n38796), .B(n38797), .Z(n26276) );
  XNOR U39476 ( .A(n26272), .B(n26274), .Z(n38797) );
  XNOR U39477 ( .A(q[24]), .B(DB[1729]), .Z(n26274) );
  XNOR U39478 ( .A(q[27]), .B(DB[1732]), .Z(n26272) );
  IV U39479 ( .A(n26271), .Z(n38796) );
  XNOR U39480 ( .A(n26269), .B(n38798), .Z(n26271) );
  XNOR U39481 ( .A(q[26]), .B(DB[1731]), .Z(n38798) );
  XNOR U39482 ( .A(q[25]), .B(DB[1730]), .Z(n26269) );
  IV U39483 ( .A(n26284), .Z(n38792) );
  XOR U39484 ( .A(n38799), .B(n38800), .Z(n26284) );
  XNOR U39485 ( .A(n26301), .B(n26282), .Z(n38800) );
  XNOR U39486 ( .A(q[16]), .B(DB[1721]), .Z(n26282) );
  XOR U39487 ( .A(n38801), .B(n26290), .Z(n26301) );
  XNOR U39488 ( .A(q[23]), .B(DB[1728]), .Z(n26290) );
  IV U39489 ( .A(n26289), .Z(n38801) );
  XNOR U39490 ( .A(n26287), .B(n38802), .Z(n26289) );
  XNOR U39491 ( .A(q[22]), .B(DB[1727]), .Z(n38802) );
  XNOR U39492 ( .A(q[21]), .B(DB[1726]), .Z(n26287) );
  IV U39493 ( .A(n26300), .Z(n38799) );
  XOR U39494 ( .A(n38803), .B(n38804), .Z(n26300) );
  XNOR U39495 ( .A(n26296), .B(n26298), .Z(n38804) );
  XNOR U39496 ( .A(q[17]), .B(DB[1722]), .Z(n26298) );
  XNOR U39497 ( .A(q[20]), .B(DB[1725]), .Z(n26296) );
  IV U39498 ( .A(n26295), .Z(n38803) );
  XNOR U39499 ( .A(n26293), .B(n38805), .Z(n26295) );
  XNOR U39500 ( .A(q[19]), .B(DB[1724]), .Z(n38805) );
  XNOR U39501 ( .A(q[18]), .B(DB[1723]), .Z(n26293) );
  IV U39502 ( .A(n26308), .Z(n38791) );
  XOR U39503 ( .A(n38806), .B(n38807), .Z(n26308) );
  XNOR U39504 ( .A(n26335), .B(n26306), .Z(n38807) );
  XNOR U39505 ( .A(q[0]), .B(DB[1705]), .Z(n26306) );
  XOR U39506 ( .A(n38808), .B(n26327), .Z(n26335) );
  XOR U39507 ( .A(n38809), .B(n26315), .Z(n26327) );
  XNOR U39508 ( .A(q[15]), .B(DB[1720]), .Z(n26315) );
  IV U39509 ( .A(n26314), .Z(n38809) );
  XNOR U39510 ( .A(n26312), .B(n38810), .Z(n26314) );
  XNOR U39511 ( .A(q[14]), .B(DB[1719]), .Z(n38810) );
  XNOR U39512 ( .A(q[13]), .B(DB[1718]), .Z(n26312) );
  IV U39513 ( .A(n26326), .Z(n38808) );
  XOR U39514 ( .A(n38811), .B(n38812), .Z(n26326) );
  XNOR U39515 ( .A(n26322), .B(n26324), .Z(n38812) );
  XNOR U39516 ( .A(q[9]), .B(DB[1714]), .Z(n26324) );
  XNOR U39517 ( .A(q[12]), .B(DB[1717]), .Z(n26322) );
  IV U39518 ( .A(n26321), .Z(n38811) );
  XNOR U39519 ( .A(n26319), .B(n38813), .Z(n26321) );
  XNOR U39520 ( .A(q[11]), .B(DB[1716]), .Z(n38813) );
  XNOR U39521 ( .A(q[10]), .B(DB[1715]), .Z(n26319) );
  IV U39522 ( .A(n26334), .Z(n38806) );
  XOR U39523 ( .A(n38814), .B(n38815), .Z(n26334) );
  XNOR U39524 ( .A(n26351), .B(n26332), .Z(n38815) );
  XNOR U39525 ( .A(q[1]), .B(DB[1706]), .Z(n26332) );
  XOR U39526 ( .A(n38816), .B(n26340), .Z(n26351) );
  XNOR U39527 ( .A(q[8]), .B(DB[1713]), .Z(n26340) );
  IV U39528 ( .A(n26339), .Z(n38816) );
  XNOR U39529 ( .A(n26337), .B(n38817), .Z(n26339) );
  XNOR U39530 ( .A(q[7]), .B(DB[1712]), .Z(n38817) );
  XNOR U39531 ( .A(q[6]), .B(DB[1711]), .Z(n26337) );
  IV U39532 ( .A(n26350), .Z(n38814) );
  XOR U39533 ( .A(n38818), .B(n38819), .Z(n26350) );
  XNOR U39534 ( .A(n26346), .B(n26348), .Z(n38819) );
  XNOR U39535 ( .A(q[2]), .B(DB[1707]), .Z(n26348) );
  XNOR U39536 ( .A(q[5]), .B(DB[1710]), .Z(n26346) );
  IV U39537 ( .A(n26345), .Z(n38818) );
  XNOR U39538 ( .A(n26343), .B(n38820), .Z(n26345) );
  XNOR U39539 ( .A(q[4]), .B(DB[1709]), .Z(n38820) );
  XNOR U39540 ( .A(q[3]), .B(DB[1708]), .Z(n26343) );
  XOR U39541 ( .A(n38821), .B(n26112), .Z(n25963) );
  XOR U39542 ( .A(n38822), .B(n26088), .Z(n26112) );
  XOR U39543 ( .A(n38823), .B(n26080), .Z(n26088) );
  XOR U39544 ( .A(n38824), .B(n26069), .Z(n26080) );
  XNOR U39545 ( .A(q[30]), .B(DB[1766]), .Z(n26069) );
  IV U39546 ( .A(n26068), .Z(n38824) );
  XNOR U39547 ( .A(n26066), .B(n38825), .Z(n26068) );
  XNOR U39548 ( .A(q[29]), .B(DB[1765]), .Z(n38825) );
  XNOR U39549 ( .A(q[28]), .B(DB[1764]), .Z(n26066) );
  IV U39550 ( .A(n26079), .Z(n38823) );
  XOR U39551 ( .A(n38826), .B(n38827), .Z(n26079) );
  XNOR U39552 ( .A(n26075), .B(n26077), .Z(n38827) );
  XNOR U39553 ( .A(q[24]), .B(DB[1760]), .Z(n26077) );
  XNOR U39554 ( .A(q[27]), .B(DB[1763]), .Z(n26075) );
  IV U39555 ( .A(n26074), .Z(n38826) );
  XNOR U39556 ( .A(n26072), .B(n38828), .Z(n26074) );
  XNOR U39557 ( .A(q[26]), .B(DB[1762]), .Z(n38828) );
  XNOR U39558 ( .A(q[25]), .B(DB[1761]), .Z(n26072) );
  IV U39559 ( .A(n26087), .Z(n38822) );
  XOR U39560 ( .A(n38829), .B(n38830), .Z(n26087) );
  XNOR U39561 ( .A(n26104), .B(n26085), .Z(n38830) );
  XNOR U39562 ( .A(q[16]), .B(DB[1752]), .Z(n26085) );
  XOR U39563 ( .A(n38831), .B(n26093), .Z(n26104) );
  XNOR U39564 ( .A(q[23]), .B(DB[1759]), .Z(n26093) );
  IV U39565 ( .A(n26092), .Z(n38831) );
  XNOR U39566 ( .A(n26090), .B(n38832), .Z(n26092) );
  XNOR U39567 ( .A(q[22]), .B(DB[1758]), .Z(n38832) );
  XNOR U39568 ( .A(q[21]), .B(DB[1757]), .Z(n26090) );
  IV U39569 ( .A(n26103), .Z(n38829) );
  XOR U39570 ( .A(n38833), .B(n38834), .Z(n26103) );
  XNOR U39571 ( .A(n26099), .B(n26101), .Z(n38834) );
  XNOR U39572 ( .A(q[17]), .B(DB[1753]), .Z(n26101) );
  XNOR U39573 ( .A(q[20]), .B(DB[1756]), .Z(n26099) );
  IV U39574 ( .A(n26098), .Z(n38833) );
  XNOR U39575 ( .A(n26096), .B(n38835), .Z(n26098) );
  XNOR U39576 ( .A(q[19]), .B(DB[1755]), .Z(n38835) );
  XNOR U39577 ( .A(q[18]), .B(DB[1754]), .Z(n26096) );
  IV U39578 ( .A(n26111), .Z(n38821) );
  XOR U39579 ( .A(n38836), .B(n38837), .Z(n26111) );
  XNOR U39580 ( .A(n26138), .B(n26109), .Z(n38837) );
  XNOR U39581 ( .A(q[0]), .B(DB[1736]), .Z(n26109) );
  XOR U39582 ( .A(n38838), .B(n26130), .Z(n26138) );
  XOR U39583 ( .A(n38839), .B(n26118), .Z(n26130) );
  XNOR U39584 ( .A(q[15]), .B(DB[1751]), .Z(n26118) );
  IV U39585 ( .A(n26117), .Z(n38839) );
  XNOR U39586 ( .A(n26115), .B(n38840), .Z(n26117) );
  XNOR U39587 ( .A(q[14]), .B(DB[1750]), .Z(n38840) );
  XNOR U39588 ( .A(q[13]), .B(DB[1749]), .Z(n26115) );
  IV U39589 ( .A(n26129), .Z(n38838) );
  XOR U39590 ( .A(n38841), .B(n38842), .Z(n26129) );
  XNOR U39591 ( .A(n26125), .B(n26127), .Z(n38842) );
  XNOR U39592 ( .A(q[9]), .B(DB[1745]), .Z(n26127) );
  XNOR U39593 ( .A(q[12]), .B(DB[1748]), .Z(n26125) );
  IV U39594 ( .A(n26124), .Z(n38841) );
  XNOR U39595 ( .A(n26122), .B(n38843), .Z(n26124) );
  XNOR U39596 ( .A(q[11]), .B(DB[1747]), .Z(n38843) );
  XNOR U39597 ( .A(q[10]), .B(DB[1746]), .Z(n26122) );
  IV U39598 ( .A(n26137), .Z(n38836) );
  XOR U39599 ( .A(n38844), .B(n38845), .Z(n26137) );
  XNOR U39600 ( .A(n26154), .B(n26135), .Z(n38845) );
  XNOR U39601 ( .A(q[1]), .B(DB[1737]), .Z(n26135) );
  XOR U39602 ( .A(n38846), .B(n26143), .Z(n26154) );
  XNOR U39603 ( .A(q[8]), .B(DB[1744]), .Z(n26143) );
  IV U39604 ( .A(n26142), .Z(n38846) );
  XNOR U39605 ( .A(n26140), .B(n38847), .Z(n26142) );
  XNOR U39606 ( .A(q[7]), .B(DB[1743]), .Z(n38847) );
  XNOR U39607 ( .A(q[6]), .B(DB[1742]), .Z(n26140) );
  IV U39608 ( .A(n26153), .Z(n38844) );
  XOR U39609 ( .A(n38848), .B(n38849), .Z(n26153) );
  XNOR U39610 ( .A(n26149), .B(n26151), .Z(n38849) );
  XNOR U39611 ( .A(q[2]), .B(DB[1738]), .Z(n26151) );
  XNOR U39612 ( .A(q[5]), .B(DB[1741]), .Z(n26149) );
  IV U39613 ( .A(n26148), .Z(n38848) );
  XNOR U39614 ( .A(n26146), .B(n38850), .Z(n26148) );
  XNOR U39615 ( .A(q[4]), .B(DB[1740]), .Z(n38850) );
  XNOR U39616 ( .A(q[3]), .B(DB[1739]), .Z(n26146) );
  XOR U39617 ( .A(n38851), .B(n25915), .Z(n25766) );
  XOR U39618 ( .A(n38852), .B(n25891), .Z(n25915) );
  XOR U39619 ( .A(n38853), .B(n25883), .Z(n25891) );
  XOR U39620 ( .A(n38854), .B(n25872), .Z(n25883) );
  XNOR U39621 ( .A(q[30]), .B(DB[1797]), .Z(n25872) );
  IV U39622 ( .A(n25871), .Z(n38854) );
  XNOR U39623 ( .A(n25869), .B(n38855), .Z(n25871) );
  XNOR U39624 ( .A(q[29]), .B(DB[1796]), .Z(n38855) );
  XNOR U39625 ( .A(q[28]), .B(DB[1795]), .Z(n25869) );
  IV U39626 ( .A(n25882), .Z(n38853) );
  XOR U39627 ( .A(n38856), .B(n38857), .Z(n25882) );
  XNOR U39628 ( .A(n25878), .B(n25880), .Z(n38857) );
  XNOR U39629 ( .A(q[24]), .B(DB[1791]), .Z(n25880) );
  XNOR U39630 ( .A(q[27]), .B(DB[1794]), .Z(n25878) );
  IV U39631 ( .A(n25877), .Z(n38856) );
  XNOR U39632 ( .A(n25875), .B(n38858), .Z(n25877) );
  XNOR U39633 ( .A(q[26]), .B(DB[1793]), .Z(n38858) );
  XNOR U39634 ( .A(q[25]), .B(DB[1792]), .Z(n25875) );
  IV U39635 ( .A(n25890), .Z(n38852) );
  XOR U39636 ( .A(n38859), .B(n38860), .Z(n25890) );
  XNOR U39637 ( .A(n25907), .B(n25888), .Z(n38860) );
  XNOR U39638 ( .A(q[16]), .B(DB[1783]), .Z(n25888) );
  XOR U39639 ( .A(n38861), .B(n25896), .Z(n25907) );
  XNOR U39640 ( .A(q[23]), .B(DB[1790]), .Z(n25896) );
  IV U39641 ( .A(n25895), .Z(n38861) );
  XNOR U39642 ( .A(n25893), .B(n38862), .Z(n25895) );
  XNOR U39643 ( .A(q[22]), .B(DB[1789]), .Z(n38862) );
  XNOR U39644 ( .A(q[21]), .B(DB[1788]), .Z(n25893) );
  IV U39645 ( .A(n25906), .Z(n38859) );
  XOR U39646 ( .A(n38863), .B(n38864), .Z(n25906) );
  XNOR U39647 ( .A(n25902), .B(n25904), .Z(n38864) );
  XNOR U39648 ( .A(q[17]), .B(DB[1784]), .Z(n25904) );
  XNOR U39649 ( .A(q[20]), .B(DB[1787]), .Z(n25902) );
  IV U39650 ( .A(n25901), .Z(n38863) );
  XNOR U39651 ( .A(n25899), .B(n38865), .Z(n25901) );
  XNOR U39652 ( .A(q[19]), .B(DB[1786]), .Z(n38865) );
  XNOR U39653 ( .A(q[18]), .B(DB[1785]), .Z(n25899) );
  IV U39654 ( .A(n25914), .Z(n38851) );
  XOR U39655 ( .A(n38866), .B(n38867), .Z(n25914) );
  XNOR U39656 ( .A(n25941), .B(n25912), .Z(n38867) );
  XNOR U39657 ( .A(q[0]), .B(DB[1767]), .Z(n25912) );
  XOR U39658 ( .A(n38868), .B(n25933), .Z(n25941) );
  XOR U39659 ( .A(n38869), .B(n25921), .Z(n25933) );
  XNOR U39660 ( .A(q[15]), .B(DB[1782]), .Z(n25921) );
  IV U39661 ( .A(n25920), .Z(n38869) );
  XNOR U39662 ( .A(n25918), .B(n38870), .Z(n25920) );
  XNOR U39663 ( .A(q[14]), .B(DB[1781]), .Z(n38870) );
  XNOR U39664 ( .A(q[13]), .B(DB[1780]), .Z(n25918) );
  IV U39665 ( .A(n25932), .Z(n38868) );
  XOR U39666 ( .A(n38871), .B(n38872), .Z(n25932) );
  XNOR U39667 ( .A(n25928), .B(n25930), .Z(n38872) );
  XNOR U39668 ( .A(q[9]), .B(DB[1776]), .Z(n25930) );
  XNOR U39669 ( .A(q[12]), .B(DB[1779]), .Z(n25928) );
  IV U39670 ( .A(n25927), .Z(n38871) );
  XNOR U39671 ( .A(n25925), .B(n38873), .Z(n25927) );
  XNOR U39672 ( .A(q[11]), .B(DB[1778]), .Z(n38873) );
  XNOR U39673 ( .A(q[10]), .B(DB[1777]), .Z(n25925) );
  IV U39674 ( .A(n25940), .Z(n38866) );
  XOR U39675 ( .A(n38874), .B(n38875), .Z(n25940) );
  XNOR U39676 ( .A(n25957), .B(n25938), .Z(n38875) );
  XNOR U39677 ( .A(q[1]), .B(DB[1768]), .Z(n25938) );
  XOR U39678 ( .A(n38876), .B(n25946), .Z(n25957) );
  XNOR U39679 ( .A(q[8]), .B(DB[1775]), .Z(n25946) );
  IV U39680 ( .A(n25945), .Z(n38876) );
  XNOR U39681 ( .A(n25943), .B(n38877), .Z(n25945) );
  XNOR U39682 ( .A(q[7]), .B(DB[1774]), .Z(n38877) );
  XNOR U39683 ( .A(q[6]), .B(DB[1773]), .Z(n25943) );
  IV U39684 ( .A(n25956), .Z(n38874) );
  XOR U39685 ( .A(n38878), .B(n38879), .Z(n25956) );
  XNOR U39686 ( .A(n25952), .B(n25954), .Z(n38879) );
  XNOR U39687 ( .A(q[2]), .B(DB[1769]), .Z(n25954) );
  XNOR U39688 ( .A(q[5]), .B(DB[1772]), .Z(n25952) );
  IV U39689 ( .A(n25951), .Z(n38878) );
  XNOR U39690 ( .A(n25949), .B(n38880), .Z(n25951) );
  XNOR U39691 ( .A(q[4]), .B(DB[1771]), .Z(n38880) );
  XNOR U39692 ( .A(q[3]), .B(DB[1770]), .Z(n25949) );
  XOR U39693 ( .A(n38881), .B(n25718), .Z(n25569) );
  XOR U39694 ( .A(n38882), .B(n25694), .Z(n25718) );
  XOR U39695 ( .A(n38883), .B(n25686), .Z(n25694) );
  XOR U39696 ( .A(n38884), .B(n25675), .Z(n25686) );
  XNOR U39697 ( .A(q[30]), .B(DB[1828]), .Z(n25675) );
  IV U39698 ( .A(n25674), .Z(n38884) );
  XNOR U39699 ( .A(n25672), .B(n38885), .Z(n25674) );
  XNOR U39700 ( .A(q[29]), .B(DB[1827]), .Z(n38885) );
  XNOR U39701 ( .A(q[28]), .B(DB[1826]), .Z(n25672) );
  IV U39702 ( .A(n25685), .Z(n38883) );
  XOR U39703 ( .A(n38886), .B(n38887), .Z(n25685) );
  XNOR U39704 ( .A(n25681), .B(n25683), .Z(n38887) );
  XNOR U39705 ( .A(q[24]), .B(DB[1822]), .Z(n25683) );
  XNOR U39706 ( .A(q[27]), .B(DB[1825]), .Z(n25681) );
  IV U39707 ( .A(n25680), .Z(n38886) );
  XNOR U39708 ( .A(n25678), .B(n38888), .Z(n25680) );
  XNOR U39709 ( .A(q[26]), .B(DB[1824]), .Z(n38888) );
  XNOR U39710 ( .A(q[25]), .B(DB[1823]), .Z(n25678) );
  IV U39711 ( .A(n25693), .Z(n38882) );
  XOR U39712 ( .A(n38889), .B(n38890), .Z(n25693) );
  XNOR U39713 ( .A(n25710), .B(n25691), .Z(n38890) );
  XNOR U39714 ( .A(q[16]), .B(DB[1814]), .Z(n25691) );
  XOR U39715 ( .A(n38891), .B(n25699), .Z(n25710) );
  XNOR U39716 ( .A(q[23]), .B(DB[1821]), .Z(n25699) );
  IV U39717 ( .A(n25698), .Z(n38891) );
  XNOR U39718 ( .A(n25696), .B(n38892), .Z(n25698) );
  XNOR U39719 ( .A(q[22]), .B(DB[1820]), .Z(n38892) );
  XNOR U39720 ( .A(q[21]), .B(DB[1819]), .Z(n25696) );
  IV U39721 ( .A(n25709), .Z(n38889) );
  XOR U39722 ( .A(n38893), .B(n38894), .Z(n25709) );
  XNOR U39723 ( .A(n25705), .B(n25707), .Z(n38894) );
  XNOR U39724 ( .A(q[17]), .B(DB[1815]), .Z(n25707) );
  XNOR U39725 ( .A(q[20]), .B(DB[1818]), .Z(n25705) );
  IV U39726 ( .A(n25704), .Z(n38893) );
  XNOR U39727 ( .A(n25702), .B(n38895), .Z(n25704) );
  XNOR U39728 ( .A(q[19]), .B(DB[1817]), .Z(n38895) );
  XNOR U39729 ( .A(q[18]), .B(DB[1816]), .Z(n25702) );
  IV U39730 ( .A(n25717), .Z(n38881) );
  XOR U39731 ( .A(n38896), .B(n38897), .Z(n25717) );
  XNOR U39732 ( .A(n25744), .B(n25715), .Z(n38897) );
  XNOR U39733 ( .A(q[0]), .B(DB[1798]), .Z(n25715) );
  XOR U39734 ( .A(n38898), .B(n25736), .Z(n25744) );
  XOR U39735 ( .A(n38899), .B(n25724), .Z(n25736) );
  XNOR U39736 ( .A(q[15]), .B(DB[1813]), .Z(n25724) );
  IV U39737 ( .A(n25723), .Z(n38899) );
  XNOR U39738 ( .A(n25721), .B(n38900), .Z(n25723) );
  XNOR U39739 ( .A(q[14]), .B(DB[1812]), .Z(n38900) );
  XNOR U39740 ( .A(q[13]), .B(DB[1811]), .Z(n25721) );
  IV U39741 ( .A(n25735), .Z(n38898) );
  XOR U39742 ( .A(n38901), .B(n38902), .Z(n25735) );
  XNOR U39743 ( .A(n25731), .B(n25733), .Z(n38902) );
  XNOR U39744 ( .A(q[9]), .B(DB[1807]), .Z(n25733) );
  XNOR U39745 ( .A(q[12]), .B(DB[1810]), .Z(n25731) );
  IV U39746 ( .A(n25730), .Z(n38901) );
  XNOR U39747 ( .A(n25728), .B(n38903), .Z(n25730) );
  XNOR U39748 ( .A(q[11]), .B(DB[1809]), .Z(n38903) );
  XNOR U39749 ( .A(q[10]), .B(DB[1808]), .Z(n25728) );
  IV U39750 ( .A(n25743), .Z(n38896) );
  XOR U39751 ( .A(n38904), .B(n38905), .Z(n25743) );
  XNOR U39752 ( .A(n25760), .B(n25741), .Z(n38905) );
  XNOR U39753 ( .A(q[1]), .B(DB[1799]), .Z(n25741) );
  XOR U39754 ( .A(n38906), .B(n25749), .Z(n25760) );
  XNOR U39755 ( .A(q[8]), .B(DB[1806]), .Z(n25749) );
  IV U39756 ( .A(n25748), .Z(n38906) );
  XNOR U39757 ( .A(n25746), .B(n38907), .Z(n25748) );
  XNOR U39758 ( .A(q[7]), .B(DB[1805]), .Z(n38907) );
  XNOR U39759 ( .A(q[6]), .B(DB[1804]), .Z(n25746) );
  IV U39760 ( .A(n25759), .Z(n38904) );
  XOR U39761 ( .A(n38908), .B(n38909), .Z(n25759) );
  XNOR U39762 ( .A(n25755), .B(n25757), .Z(n38909) );
  XNOR U39763 ( .A(q[2]), .B(DB[1800]), .Z(n25757) );
  XNOR U39764 ( .A(q[5]), .B(DB[1803]), .Z(n25755) );
  IV U39765 ( .A(n25754), .Z(n38908) );
  XNOR U39766 ( .A(n25752), .B(n38910), .Z(n25754) );
  XNOR U39767 ( .A(q[4]), .B(DB[1802]), .Z(n38910) );
  XNOR U39768 ( .A(q[3]), .B(DB[1801]), .Z(n25752) );
  XOR U39769 ( .A(n38911), .B(n25521), .Z(n25372) );
  XOR U39770 ( .A(n38912), .B(n25497), .Z(n25521) );
  XOR U39771 ( .A(n38913), .B(n25489), .Z(n25497) );
  XOR U39772 ( .A(n38914), .B(n25478), .Z(n25489) );
  XNOR U39773 ( .A(q[30]), .B(DB[1859]), .Z(n25478) );
  IV U39774 ( .A(n25477), .Z(n38914) );
  XNOR U39775 ( .A(n25475), .B(n38915), .Z(n25477) );
  XNOR U39776 ( .A(q[29]), .B(DB[1858]), .Z(n38915) );
  XNOR U39777 ( .A(q[28]), .B(DB[1857]), .Z(n25475) );
  IV U39778 ( .A(n25488), .Z(n38913) );
  XOR U39779 ( .A(n38916), .B(n38917), .Z(n25488) );
  XNOR U39780 ( .A(n25484), .B(n25486), .Z(n38917) );
  XNOR U39781 ( .A(q[24]), .B(DB[1853]), .Z(n25486) );
  XNOR U39782 ( .A(q[27]), .B(DB[1856]), .Z(n25484) );
  IV U39783 ( .A(n25483), .Z(n38916) );
  XNOR U39784 ( .A(n25481), .B(n38918), .Z(n25483) );
  XNOR U39785 ( .A(q[26]), .B(DB[1855]), .Z(n38918) );
  XNOR U39786 ( .A(q[25]), .B(DB[1854]), .Z(n25481) );
  IV U39787 ( .A(n25496), .Z(n38912) );
  XOR U39788 ( .A(n38919), .B(n38920), .Z(n25496) );
  XNOR U39789 ( .A(n25513), .B(n25494), .Z(n38920) );
  XNOR U39790 ( .A(q[16]), .B(DB[1845]), .Z(n25494) );
  XOR U39791 ( .A(n38921), .B(n25502), .Z(n25513) );
  XNOR U39792 ( .A(q[23]), .B(DB[1852]), .Z(n25502) );
  IV U39793 ( .A(n25501), .Z(n38921) );
  XNOR U39794 ( .A(n25499), .B(n38922), .Z(n25501) );
  XNOR U39795 ( .A(q[22]), .B(DB[1851]), .Z(n38922) );
  XNOR U39796 ( .A(q[21]), .B(DB[1850]), .Z(n25499) );
  IV U39797 ( .A(n25512), .Z(n38919) );
  XOR U39798 ( .A(n38923), .B(n38924), .Z(n25512) );
  XNOR U39799 ( .A(n25508), .B(n25510), .Z(n38924) );
  XNOR U39800 ( .A(q[17]), .B(DB[1846]), .Z(n25510) );
  XNOR U39801 ( .A(q[20]), .B(DB[1849]), .Z(n25508) );
  IV U39802 ( .A(n25507), .Z(n38923) );
  XNOR U39803 ( .A(n25505), .B(n38925), .Z(n25507) );
  XNOR U39804 ( .A(q[19]), .B(DB[1848]), .Z(n38925) );
  XNOR U39805 ( .A(q[18]), .B(DB[1847]), .Z(n25505) );
  IV U39806 ( .A(n25520), .Z(n38911) );
  XOR U39807 ( .A(n38926), .B(n38927), .Z(n25520) );
  XNOR U39808 ( .A(n25547), .B(n25518), .Z(n38927) );
  XNOR U39809 ( .A(q[0]), .B(DB[1829]), .Z(n25518) );
  XOR U39810 ( .A(n38928), .B(n25539), .Z(n25547) );
  XOR U39811 ( .A(n38929), .B(n25527), .Z(n25539) );
  XNOR U39812 ( .A(q[15]), .B(DB[1844]), .Z(n25527) );
  IV U39813 ( .A(n25526), .Z(n38929) );
  XNOR U39814 ( .A(n25524), .B(n38930), .Z(n25526) );
  XNOR U39815 ( .A(q[14]), .B(DB[1843]), .Z(n38930) );
  XNOR U39816 ( .A(q[13]), .B(DB[1842]), .Z(n25524) );
  IV U39817 ( .A(n25538), .Z(n38928) );
  XOR U39818 ( .A(n38931), .B(n38932), .Z(n25538) );
  XNOR U39819 ( .A(n25534), .B(n25536), .Z(n38932) );
  XNOR U39820 ( .A(q[9]), .B(DB[1838]), .Z(n25536) );
  XNOR U39821 ( .A(q[12]), .B(DB[1841]), .Z(n25534) );
  IV U39822 ( .A(n25533), .Z(n38931) );
  XNOR U39823 ( .A(n25531), .B(n38933), .Z(n25533) );
  XNOR U39824 ( .A(q[11]), .B(DB[1840]), .Z(n38933) );
  XNOR U39825 ( .A(q[10]), .B(DB[1839]), .Z(n25531) );
  IV U39826 ( .A(n25546), .Z(n38926) );
  XOR U39827 ( .A(n38934), .B(n38935), .Z(n25546) );
  XNOR U39828 ( .A(n25563), .B(n25544), .Z(n38935) );
  XNOR U39829 ( .A(q[1]), .B(DB[1830]), .Z(n25544) );
  XOR U39830 ( .A(n38936), .B(n25552), .Z(n25563) );
  XNOR U39831 ( .A(q[8]), .B(DB[1837]), .Z(n25552) );
  IV U39832 ( .A(n25551), .Z(n38936) );
  XNOR U39833 ( .A(n25549), .B(n38937), .Z(n25551) );
  XNOR U39834 ( .A(q[7]), .B(DB[1836]), .Z(n38937) );
  XNOR U39835 ( .A(q[6]), .B(DB[1835]), .Z(n25549) );
  IV U39836 ( .A(n25562), .Z(n38934) );
  XOR U39837 ( .A(n38938), .B(n38939), .Z(n25562) );
  XNOR U39838 ( .A(n25558), .B(n25560), .Z(n38939) );
  XNOR U39839 ( .A(q[2]), .B(DB[1831]), .Z(n25560) );
  XNOR U39840 ( .A(q[5]), .B(DB[1834]), .Z(n25558) );
  IV U39841 ( .A(n25557), .Z(n38938) );
  XNOR U39842 ( .A(n25555), .B(n38940), .Z(n25557) );
  XNOR U39843 ( .A(q[4]), .B(DB[1833]), .Z(n38940) );
  XNOR U39844 ( .A(q[3]), .B(DB[1832]), .Z(n25555) );
  XOR U39845 ( .A(n38941), .B(n25324), .Z(n25175) );
  XOR U39846 ( .A(n38942), .B(n25300), .Z(n25324) );
  XOR U39847 ( .A(n38943), .B(n25292), .Z(n25300) );
  XOR U39848 ( .A(n38944), .B(n25281), .Z(n25292) );
  XNOR U39849 ( .A(q[30]), .B(DB[1890]), .Z(n25281) );
  IV U39850 ( .A(n25280), .Z(n38944) );
  XNOR U39851 ( .A(n25278), .B(n38945), .Z(n25280) );
  XNOR U39852 ( .A(q[29]), .B(DB[1889]), .Z(n38945) );
  XNOR U39853 ( .A(q[28]), .B(DB[1888]), .Z(n25278) );
  IV U39854 ( .A(n25291), .Z(n38943) );
  XOR U39855 ( .A(n38946), .B(n38947), .Z(n25291) );
  XNOR U39856 ( .A(n25287), .B(n25289), .Z(n38947) );
  XNOR U39857 ( .A(q[24]), .B(DB[1884]), .Z(n25289) );
  XNOR U39858 ( .A(q[27]), .B(DB[1887]), .Z(n25287) );
  IV U39859 ( .A(n25286), .Z(n38946) );
  XNOR U39860 ( .A(n25284), .B(n38948), .Z(n25286) );
  XNOR U39861 ( .A(q[26]), .B(DB[1886]), .Z(n38948) );
  XNOR U39862 ( .A(q[25]), .B(DB[1885]), .Z(n25284) );
  IV U39863 ( .A(n25299), .Z(n38942) );
  XOR U39864 ( .A(n38949), .B(n38950), .Z(n25299) );
  XNOR U39865 ( .A(n25316), .B(n25297), .Z(n38950) );
  XNOR U39866 ( .A(q[16]), .B(DB[1876]), .Z(n25297) );
  XOR U39867 ( .A(n38951), .B(n25305), .Z(n25316) );
  XNOR U39868 ( .A(q[23]), .B(DB[1883]), .Z(n25305) );
  IV U39869 ( .A(n25304), .Z(n38951) );
  XNOR U39870 ( .A(n25302), .B(n38952), .Z(n25304) );
  XNOR U39871 ( .A(q[22]), .B(DB[1882]), .Z(n38952) );
  XNOR U39872 ( .A(q[21]), .B(DB[1881]), .Z(n25302) );
  IV U39873 ( .A(n25315), .Z(n38949) );
  XOR U39874 ( .A(n38953), .B(n38954), .Z(n25315) );
  XNOR U39875 ( .A(n25311), .B(n25313), .Z(n38954) );
  XNOR U39876 ( .A(q[17]), .B(DB[1877]), .Z(n25313) );
  XNOR U39877 ( .A(q[20]), .B(DB[1880]), .Z(n25311) );
  IV U39878 ( .A(n25310), .Z(n38953) );
  XNOR U39879 ( .A(n25308), .B(n38955), .Z(n25310) );
  XNOR U39880 ( .A(q[19]), .B(DB[1879]), .Z(n38955) );
  XNOR U39881 ( .A(q[18]), .B(DB[1878]), .Z(n25308) );
  IV U39882 ( .A(n25323), .Z(n38941) );
  XOR U39883 ( .A(n38956), .B(n38957), .Z(n25323) );
  XNOR U39884 ( .A(n25350), .B(n25321), .Z(n38957) );
  XNOR U39885 ( .A(q[0]), .B(DB[1860]), .Z(n25321) );
  XOR U39886 ( .A(n38958), .B(n25342), .Z(n25350) );
  XOR U39887 ( .A(n38959), .B(n25330), .Z(n25342) );
  XNOR U39888 ( .A(q[15]), .B(DB[1875]), .Z(n25330) );
  IV U39889 ( .A(n25329), .Z(n38959) );
  XNOR U39890 ( .A(n25327), .B(n38960), .Z(n25329) );
  XNOR U39891 ( .A(q[14]), .B(DB[1874]), .Z(n38960) );
  XNOR U39892 ( .A(q[13]), .B(DB[1873]), .Z(n25327) );
  IV U39893 ( .A(n25341), .Z(n38958) );
  XOR U39894 ( .A(n38961), .B(n38962), .Z(n25341) );
  XNOR U39895 ( .A(n25337), .B(n25339), .Z(n38962) );
  XNOR U39896 ( .A(q[9]), .B(DB[1869]), .Z(n25339) );
  XNOR U39897 ( .A(q[12]), .B(DB[1872]), .Z(n25337) );
  IV U39898 ( .A(n25336), .Z(n38961) );
  XNOR U39899 ( .A(n25334), .B(n38963), .Z(n25336) );
  XNOR U39900 ( .A(q[11]), .B(DB[1871]), .Z(n38963) );
  XNOR U39901 ( .A(q[10]), .B(DB[1870]), .Z(n25334) );
  IV U39902 ( .A(n25349), .Z(n38956) );
  XOR U39903 ( .A(n38964), .B(n38965), .Z(n25349) );
  XNOR U39904 ( .A(n25366), .B(n25347), .Z(n38965) );
  XNOR U39905 ( .A(q[1]), .B(DB[1861]), .Z(n25347) );
  XOR U39906 ( .A(n38966), .B(n25355), .Z(n25366) );
  XNOR U39907 ( .A(q[8]), .B(DB[1868]), .Z(n25355) );
  IV U39908 ( .A(n25354), .Z(n38966) );
  XNOR U39909 ( .A(n25352), .B(n38967), .Z(n25354) );
  XNOR U39910 ( .A(q[7]), .B(DB[1867]), .Z(n38967) );
  XNOR U39911 ( .A(q[6]), .B(DB[1866]), .Z(n25352) );
  IV U39912 ( .A(n25365), .Z(n38964) );
  XOR U39913 ( .A(n38968), .B(n38969), .Z(n25365) );
  XNOR U39914 ( .A(n25361), .B(n25363), .Z(n38969) );
  XNOR U39915 ( .A(q[2]), .B(DB[1862]), .Z(n25363) );
  XNOR U39916 ( .A(q[5]), .B(DB[1865]), .Z(n25361) );
  IV U39917 ( .A(n25360), .Z(n38968) );
  XNOR U39918 ( .A(n25358), .B(n38970), .Z(n25360) );
  XNOR U39919 ( .A(q[4]), .B(DB[1864]), .Z(n38970) );
  XNOR U39920 ( .A(q[3]), .B(DB[1863]), .Z(n25358) );
  XOR U39921 ( .A(n38971), .B(n25127), .Z(n24978) );
  XOR U39922 ( .A(n38972), .B(n25103), .Z(n25127) );
  XOR U39923 ( .A(n38973), .B(n25095), .Z(n25103) );
  XOR U39924 ( .A(n38974), .B(n25084), .Z(n25095) );
  XNOR U39925 ( .A(q[30]), .B(DB[1921]), .Z(n25084) );
  IV U39926 ( .A(n25083), .Z(n38974) );
  XNOR U39927 ( .A(n25081), .B(n38975), .Z(n25083) );
  XNOR U39928 ( .A(q[29]), .B(DB[1920]), .Z(n38975) );
  XNOR U39929 ( .A(q[28]), .B(DB[1919]), .Z(n25081) );
  IV U39930 ( .A(n25094), .Z(n38973) );
  XOR U39931 ( .A(n38976), .B(n38977), .Z(n25094) );
  XNOR U39932 ( .A(n25090), .B(n25092), .Z(n38977) );
  XNOR U39933 ( .A(q[24]), .B(DB[1915]), .Z(n25092) );
  XNOR U39934 ( .A(q[27]), .B(DB[1918]), .Z(n25090) );
  IV U39935 ( .A(n25089), .Z(n38976) );
  XNOR U39936 ( .A(n25087), .B(n38978), .Z(n25089) );
  XNOR U39937 ( .A(q[26]), .B(DB[1917]), .Z(n38978) );
  XNOR U39938 ( .A(q[25]), .B(DB[1916]), .Z(n25087) );
  IV U39939 ( .A(n25102), .Z(n38972) );
  XOR U39940 ( .A(n38979), .B(n38980), .Z(n25102) );
  XNOR U39941 ( .A(n25119), .B(n25100), .Z(n38980) );
  XNOR U39942 ( .A(q[16]), .B(DB[1907]), .Z(n25100) );
  XOR U39943 ( .A(n38981), .B(n25108), .Z(n25119) );
  XNOR U39944 ( .A(q[23]), .B(DB[1914]), .Z(n25108) );
  IV U39945 ( .A(n25107), .Z(n38981) );
  XNOR U39946 ( .A(n25105), .B(n38982), .Z(n25107) );
  XNOR U39947 ( .A(q[22]), .B(DB[1913]), .Z(n38982) );
  XNOR U39948 ( .A(q[21]), .B(DB[1912]), .Z(n25105) );
  IV U39949 ( .A(n25118), .Z(n38979) );
  XOR U39950 ( .A(n38983), .B(n38984), .Z(n25118) );
  XNOR U39951 ( .A(n25114), .B(n25116), .Z(n38984) );
  XNOR U39952 ( .A(q[17]), .B(DB[1908]), .Z(n25116) );
  XNOR U39953 ( .A(q[20]), .B(DB[1911]), .Z(n25114) );
  IV U39954 ( .A(n25113), .Z(n38983) );
  XNOR U39955 ( .A(n25111), .B(n38985), .Z(n25113) );
  XNOR U39956 ( .A(q[19]), .B(DB[1910]), .Z(n38985) );
  XNOR U39957 ( .A(q[18]), .B(DB[1909]), .Z(n25111) );
  IV U39958 ( .A(n25126), .Z(n38971) );
  XOR U39959 ( .A(n38986), .B(n38987), .Z(n25126) );
  XNOR U39960 ( .A(n25153), .B(n25124), .Z(n38987) );
  XNOR U39961 ( .A(q[0]), .B(DB[1891]), .Z(n25124) );
  XOR U39962 ( .A(n38988), .B(n25145), .Z(n25153) );
  XOR U39963 ( .A(n38989), .B(n25133), .Z(n25145) );
  XNOR U39964 ( .A(q[15]), .B(DB[1906]), .Z(n25133) );
  IV U39965 ( .A(n25132), .Z(n38989) );
  XNOR U39966 ( .A(n25130), .B(n38990), .Z(n25132) );
  XNOR U39967 ( .A(q[14]), .B(DB[1905]), .Z(n38990) );
  XNOR U39968 ( .A(q[13]), .B(DB[1904]), .Z(n25130) );
  IV U39969 ( .A(n25144), .Z(n38988) );
  XOR U39970 ( .A(n38991), .B(n38992), .Z(n25144) );
  XNOR U39971 ( .A(n25140), .B(n25142), .Z(n38992) );
  XNOR U39972 ( .A(q[9]), .B(DB[1900]), .Z(n25142) );
  XNOR U39973 ( .A(q[12]), .B(DB[1903]), .Z(n25140) );
  IV U39974 ( .A(n25139), .Z(n38991) );
  XNOR U39975 ( .A(n25137), .B(n38993), .Z(n25139) );
  XNOR U39976 ( .A(q[11]), .B(DB[1902]), .Z(n38993) );
  XNOR U39977 ( .A(q[10]), .B(DB[1901]), .Z(n25137) );
  IV U39978 ( .A(n25152), .Z(n38986) );
  XOR U39979 ( .A(n38994), .B(n38995), .Z(n25152) );
  XNOR U39980 ( .A(n25169), .B(n25150), .Z(n38995) );
  XNOR U39981 ( .A(q[1]), .B(DB[1892]), .Z(n25150) );
  XOR U39982 ( .A(n38996), .B(n25158), .Z(n25169) );
  XNOR U39983 ( .A(q[8]), .B(DB[1899]), .Z(n25158) );
  IV U39984 ( .A(n25157), .Z(n38996) );
  XNOR U39985 ( .A(n25155), .B(n38997), .Z(n25157) );
  XNOR U39986 ( .A(q[7]), .B(DB[1898]), .Z(n38997) );
  XNOR U39987 ( .A(q[6]), .B(DB[1897]), .Z(n25155) );
  IV U39988 ( .A(n25168), .Z(n38994) );
  XOR U39989 ( .A(n38998), .B(n38999), .Z(n25168) );
  XNOR U39990 ( .A(n25164), .B(n25166), .Z(n38999) );
  XNOR U39991 ( .A(q[2]), .B(DB[1893]), .Z(n25166) );
  XNOR U39992 ( .A(q[5]), .B(DB[1896]), .Z(n25164) );
  IV U39993 ( .A(n25163), .Z(n38998) );
  XNOR U39994 ( .A(n25161), .B(n39000), .Z(n25163) );
  XNOR U39995 ( .A(q[4]), .B(DB[1895]), .Z(n39000) );
  XNOR U39996 ( .A(q[3]), .B(DB[1894]), .Z(n25161) );
  XOR U39997 ( .A(n39001), .B(n24930), .Z(n24781) );
  XOR U39998 ( .A(n39002), .B(n24906), .Z(n24930) );
  XOR U39999 ( .A(n39003), .B(n24898), .Z(n24906) );
  XOR U40000 ( .A(n39004), .B(n24887), .Z(n24898) );
  XNOR U40001 ( .A(q[30]), .B(DB[1952]), .Z(n24887) );
  IV U40002 ( .A(n24886), .Z(n39004) );
  XNOR U40003 ( .A(n24884), .B(n39005), .Z(n24886) );
  XNOR U40004 ( .A(q[29]), .B(DB[1951]), .Z(n39005) );
  XNOR U40005 ( .A(q[28]), .B(DB[1950]), .Z(n24884) );
  IV U40006 ( .A(n24897), .Z(n39003) );
  XOR U40007 ( .A(n39006), .B(n39007), .Z(n24897) );
  XNOR U40008 ( .A(n24893), .B(n24895), .Z(n39007) );
  XNOR U40009 ( .A(q[24]), .B(DB[1946]), .Z(n24895) );
  XNOR U40010 ( .A(q[27]), .B(DB[1949]), .Z(n24893) );
  IV U40011 ( .A(n24892), .Z(n39006) );
  XNOR U40012 ( .A(n24890), .B(n39008), .Z(n24892) );
  XNOR U40013 ( .A(q[26]), .B(DB[1948]), .Z(n39008) );
  XNOR U40014 ( .A(q[25]), .B(DB[1947]), .Z(n24890) );
  IV U40015 ( .A(n24905), .Z(n39002) );
  XOR U40016 ( .A(n39009), .B(n39010), .Z(n24905) );
  XNOR U40017 ( .A(n24922), .B(n24903), .Z(n39010) );
  XNOR U40018 ( .A(q[16]), .B(DB[1938]), .Z(n24903) );
  XOR U40019 ( .A(n39011), .B(n24911), .Z(n24922) );
  XNOR U40020 ( .A(q[23]), .B(DB[1945]), .Z(n24911) );
  IV U40021 ( .A(n24910), .Z(n39011) );
  XNOR U40022 ( .A(n24908), .B(n39012), .Z(n24910) );
  XNOR U40023 ( .A(q[22]), .B(DB[1944]), .Z(n39012) );
  XNOR U40024 ( .A(q[21]), .B(DB[1943]), .Z(n24908) );
  IV U40025 ( .A(n24921), .Z(n39009) );
  XOR U40026 ( .A(n39013), .B(n39014), .Z(n24921) );
  XNOR U40027 ( .A(n24917), .B(n24919), .Z(n39014) );
  XNOR U40028 ( .A(q[17]), .B(DB[1939]), .Z(n24919) );
  XNOR U40029 ( .A(q[20]), .B(DB[1942]), .Z(n24917) );
  IV U40030 ( .A(n24916), .Z(n39013) );
  XNOR U40031 ( .A(n24914), .B(n39015), .Z(n24916) );
  XNOR U40032 ( .A(q[19]), .B(DB[1941]), .Z(n39015) );
  XNOR U40033 ( .A(q[18]), .B(DB[1940]), .Z(n24914) );
  IV U40034 ( .A(n24929), .Z(n39001) );
  XOR U40035 ( .A(n39016), .B(n39017), .Z(n24929) );
  XNOR U40036 ( .A(n24956), .B(n24927), .Z(n39017) );
  XNOR U40037 ( .A(q[0]), .B(DB[1922]), .Z(n24927) );
  XOR U40038 ( .A(n39018), .B(n24948), .Z(n24956) );
  XOR U40039 ( .A(n39019), .B(n24936), .Z(n24948) );
  XNOR U40040 ( .A(q[15]), .B(DB[1937]), .Z(n24936) );
  IV U40041 ( .A(n24935), .Z(n39019) );
  XNOR U40042 ( .A(n24933), .B(n39020), .Z(n24935) );
  XNOR U40043 ( .A(q[14]), .B(DB[1936]), .Z(n39020) );
  XNOR U40044 ( .A(q[13]), .B(DB[1935]), .Z(n24933) );
  IV U40045 ( .A(n24947), .Z(n39018) );
  XOR U40046 ( .A(n39021), .B(n39022), .Z(n24947) );
  XNOR U40047 ( .A(n24943), .B(n24945), .Z(n39022) );
  XNOR U40048 ( .A(q[9]), .B(DB[1931]), .Z(n24945) );
  XNOR U40049 ( .A(q[12]), .B(DB[1934]), .Z(n24943) );
  IV U40050 ( .A(n24942), .Z(n39021) );
  XNOR U40051 ( .A(n24940), .B(n39023), .Z(n24942) );
  XNOR U40052 ( .A(q[11]), .B(DB[1933]), .Z(n39023) );
  XNOR U40053 ( .A(q[10]), .B(DB[1932]), .Z(n24940) );
  IV U40054 ( .A(n24955), .Z(n39016) );
  XOR U40055 ( .A(n39024), .B(n39025), .Z(n24955) );
  XNOR U40056 ( .A(n24972), .B(n24953), .Z(n39025) );
  XNOR U40057 ( .A(q[1]), .B(DB[1923]), .Z(n24953) );
  XOR U40058 ( .A(n39026), .B(n24961), .Z(n24972) );
  XNOR U40059 ( .A(q[8]), .B(DB[1930]), .Z(n24961) );
  IV U40060 ( .A(n24960), .Z(n39026) );
  XNOR U40061 ( .A(n24958), .B(n39027), .Z(n24960) );
  XNOR U40062 ( .A(q[7]), .B(DB[1929]), .Z(n39027) );
  XNOR U40063 ( .A(q[6]), .B(DB[1928]), .Z(n24958) );
  IV U40064 ( .A(n24971), .Z(n39024) );
  XOR U40065 ( .A(n39028), .B(n39029), .Z(n24971) );
  XNOR U40066 ( .A(n24967), .B(n24969), .Z(n39029) );
  XNOR U40067 ( .A(q[2]), .B(DB[1924]), .Z(n24969) );
  XNOR U40068 ( .A(q[5]), .B(DB[1927]), .Z(n24967) );
  IV U40069 ( .A(n24966), .Z(n39028) );
  XNOR U40070 ( .A(n24964), .B(n39030), .Z(n24966) );
  XNOR U40071 ( .A(q[4]), .B(DB[1926]), .Z(n39030) );
  XNOR U40072 ( .A(q[3]), .B(DB[1925]), .Z(n24964) );
  XOR U40073 ( .A(n39031), .B(n24733), .Z(n24584) );
  XOR U40074 ( .A(n39032), .B(n24709), .Z(n24733) );
  XOR U40075 ( .A(n39033), .B(n24701), .Z(n24709) );
  XOR U40076 ( .A(n39034), .B(n24690), .Z(n24701) );
  XNOR U40077 ( .A(q[30]), .B(DB[1983]), .Z(n24690) );
  IV U40078 ( .A(n24689), .Z(n39034) );
  XNOR U40079 ( .A(n24687), .B(n39035), .Z(n24689) );
  XNOR U40080 ( .A(q[29]), .B(DB[1982]), .Z(n39035) );
  XNOR U40081 ( .A(q[28]), .B(DB[1981]), .Z(n24687) );
  IV U40082 ( .A(n24700), .Z(n39033) );
  XOR U40083 ( .A(n39036), .B(n39037), .Z(n24700) );
  XNOR U40084 ( .A(n24696), .B(n24698), .Z(n39037) );
  XNOR U40085 ( .A(q[24]), .B(DB[1977]), .Z(n24698) );
  XNOR U40086 ( .A(q[27]), .B(DB[1980]), .Z(n24696) );
  IV U40087 ( .A(n24695), .Z(n39036) );
  XNOR U40088 ( .A(n24693), .B(n39038), .Z(n24695) );
  XNOR U40089 ( .A(q[26]), .B(DB[1979]), .Z(n39038) );
  XNOR U40090 ( .A(q[25]), .B(DB[1978]), .Z(n24693) );
  IV U40091 ( .A(n24708), .Z(n39032) );
  XOR U40092 ( .A(n39039), .B(n39040), .Z(n24708) );
  XNOR U40093 ( .A(n24725), .B(n24706), .Z(n39040) );
  XNOR U40094 ( .A(q[16]), .B(DB[1969]), .Z(n24706) );
  XOR U40095 ( .A(n39041), .B(n24714), .Z(n24725) );
  XNOR U40096 ( .A(q[23]), .B(DB[1976]), .Z(n24714) );
  IV U40097 ( .A(n24713), .Z(n39041) );
  XNOR U40098 ( .A(n24711), .B(n39042), .Z(n24713) );
  XNOR U40099 ( .A(q[22]), .B(DB[1975]), .Z(n39042) );
  XNOR U40100 ( .A(q[21]), .B(DB[1974]), .Z(n24711) );
  IV U40101 ( .A(n24724), .Z(n39039) );
  XOR U40102 ( .A(n39043), .B(n39044), .Z(n24724) );
  XNOR U40103 ( .A(n24720), .B(n24722), .Z(n39044) );
  XNOR U40104 ( .A(q[17]), .B(DB[1970]), .Z(n24722) );
  XNOR U40105 ( .A(q[20]), .B(DB[1973]), .Z(n24720) );
  IV U40106 ( .A(n24719), .Z(n39043) );
  XNOR U40107 ( .A(n24717), .B(n39045), .Z(n24719) );
  XNOR U40108 ( .A(q[19]), .B(DB[1972]), .Z(n39045) );
  XNOR U40109 ( .A(q[18]), .B(DB[1971]), .Z(n24717) );
  IV U40110 ( .A(n24732), .Z(n39031) );
  XOR U40111 ( .A(n39046), .B(n39047), .Z(n24732) );
  XNOR U40112 ( .A(n24759), .B(n24730), .Z(n39047) );
  XNOR U40113 ( .A(q[0]), .B(DB[1953]), .Z(n24730) );
  XOR U40114 ( .A(n39048), .B(n24751), .Z(n24759) );
  XOR U40115 ( .A(n39049), .B(n24739), .Z(n24751) );
  XNOR U40116 ( .A(q[15]), .B(DB[1968]), .Z(n24739) );
  IV U40117 ( .A(n24738), .Z(n39049) );
  XNOR U40118 ( .A(n24736), .B(n39050), .Z(n24738) );
  XNOR U40119 ( .A(q[14]), .B(DB[1967]), .Z(n39050) );
  XNOR U40120 ( .A(q[13]), .B(DB[1966]), .Z(n24736) );
  IV U40121 ( .A(n24750), .Z(n39048) );
  XOR U40122 ( .A(n39051), .B(n39052), .Z(n24750) );
  XNOR U40123 ( .A(n24746), .B(n24748), .Z(n39052) );
  XNOR U40124 ( .A(q[9]), .B(DB[1962]), .Z(n24748) );
  XNOR U40125 ( .A(q[12]), .B(DB[1965]), .Z(n24746) );
  IV U40126 ( .A(n24745), .Z(n39051) );
  XNOR U40127 ( .A(n24743), .B(n39053), .Z(n24745) );
  XNOR U40128 ( .A(q[11]), .B(DB[1964]), .Z(n39053) );
  XNOR U40129 ( .A(q[10]), .B(DB[1963]), .Z(n24743) );
  IV U40130 ( .A(n24758), .Z(n39046) );
  XOR U40131 ( .A(n39054), .B(n39055), .Z(n24758) );
  XNOR U40132 ( .A(n24775), .B(n24756), .Z(n39055) );
  XNOR U40133 ( .A(q[1]), .B(DB[1954]), .Z(n24756) );
  XOR U40134 ( .A(n39056), .B(n24764), .Z(n24775) );
  XNOR U40135 ( .A(q[8]), .B(DB[1961]), .Z(n24764) );
  IV U40136 ( .A(n24763), .Z(n39056) );
  XNOR U40137 ( .A(n24761), .B(n39057), .Z(n24763) );
  XNOR U40138 ( .A(q[7]), .B(DB[1960]), .Z(n39057) );
  XNOR U40139 ( .A(q[6]), .B(DB[1959]), .Z(n24761) );
  IV U40140 ( .A(n24774), .Z(n39054) );
  XOR U40141 ( .A(n39058), .B(n39059), .Z(n24774) );
  XNOR U40142 ( .A(n24770), .B(n24772), .Z(n39059) );
  XNOR U40143 ( .A(q[2]), .B(DB[1955]), .Z(n24772) );
  XNOR U40144 ( .A(q[5]), .B(DB[1958]), .Z(n24770) );
  IV U40145 ( .A(n24769), .Z(n39058) );
  XNOR U40146 ( .A(n24767), .B(n39060), .Z(n24769) );
  XNOR U40147 ( .A(q[4]), .B(DB[1957]), .Z(n39060) );
  XNOR U40148 ( .A(q[3]), .B(DB[1956]), .Z(n24767) );
  XOR U40149 ( .A(n39061), .B(n24536), .Z(n24387) );
  XOR U40150 ( .A(n39062), .B(n24512), .Z(n24536) );
  XOR U40151 ( .A(n39063), .B(n24504), .Z(n24512) );
  XOR U40152 ( .A(n39064), .B(n24493), .Z(n24504) );
  XNOR U40153 ( .A(q[30]), .B(DB[2014]), .Z(n24493) );
  IV U40154 ( .A(n24492), .Z(n39064) );
  XNOR U40155 ( .A(n24490), .B(n39065), .Z(n24492) );
  XNOR U40156 ( .A(q[29]), .B(DB[2013]), .Z(n39065) );
  XNOR U40157 ( .A(q[28]), .B(DB[2012]), .Z(n24490) );
  IV U40158 ( .A(n24503), .Z(n39063) );
  XOR U40159 ( .A(n39066), .B(n39067), .Z(n24503) );
  XNOR U40160 ( .A(n24499), .B(n24501), .Z(n39067) );
  XNOR U40161 ( .A(q[24]), .B(DB[2008]), .Z(n24501) );
  XNOR U40162 ( .A(q[27]), .B(DB[2011]), .Z(n24499) );
  IV U40163 ( .A(n24498), .Z(n39066) );
  XNOR U40164 ( .A(n24496), .B(n39068), .Z(n24498) );
  XNOR U40165 ( .A(q[26]), .B(DB[2010]), .Z(n39068) );
  XNOR U40166 ( .A(q[25]), .B(DB[2009]), .Z(n24496) );
  IV U40167 ( .A(n24511), .Z(n39062) );
  XOR U40168 ( .A(n39069), .B(n39070), .Z(n24511) );
  XNOR U40169 ( .A(n24528), .B(n24509), .Z(n39070) );
  XNOR U40170 ( .A(q[16]), .B(DB[2000]), .Z(n24509) );
  XOR U40171 ( .A(n39071), .B(n24517), .Z(n24528) );
  XNOR U40172 ( .A(q[23]), .B(DB[2007]), .Z(n24517) );
  IV U40173 ( .A(n24516), .Z(n39071) );
  XNOR U40174 ( .A(n24514), .B(n39072), .Z(n24516) );
  XNOR U40175 ( .A(q[22]), .B(DB[2006]), .Z(n39072) );
  XNOR U40176 ( .A(q[21]), .B(DB[2005]), .Z(n24514) );
  IV U40177 ( .A(n24527), .Z(n39069) );
  XOR U40178 ( .A(n39073), .B(n39074), .Z(n24527) );
  XNOR U40179 ( .A(n24523), .B(n24525), .Z(n39074) );
  XNOR U40180 ( .A(q[17]), .B(DB[2001]), .Z(n24525) );
  XNOR U40181 ( .A(q[20]), .B(DB[2004]), .Z(n24523) );
  IV U40182 ( .A(n24522), .Z(n39073) );
  XNOR U40183 ( .A(n24520), .B(n39075), .Z(n24522) );
  XNOR U40184 ( .A(q[19]), .B(DB[2003]), .Z(n39075) );
  XNOR U40185 ( .A(q[18]), .B(DB[2002]), .Z(n24520) );
  IV U40186 ( .A(n24535), .Z(n39061) );
  XOR U40187 ( .A(n39076), .B(n39077), .Z(n24535) );
  XNOR U40188 ( .A(n24562), .B(n24533), .Z(n39077) );
  XNOR U40189 ( .A(q[0]), .B(DB[1984]), .Z(n24533) );
  XOR U40190 ( .A(n39078), .B(n24554), .Z(n24562) );
  XOR U40191 ( .A(n39079), .B(n24542), .Z(n24554) );
  XNOR U40192 ( .A(q[15]), .B(DB[1999]), .Z(n24542) );
  IV U40193 ( .A(n24541), .Z(n39079) );
  XNOR U40194 ( .A(n24539), .B(n39080), .Z(n24541) );
  XNOR U40195 ( .A(q[14]), .B(DB[1998]), .Z(n39080) );
  XNOR U40196 ( .A(q[13]), .B(DB[1997]), .Z(n24539) );
  IV U40197 ( .A(n24553), .Z(n39078) );
  XOR U40198 ( .A(n39081), .B(n39082), .Z(n24553) );
  XNOR U40199 ( .A(n24549), .B(n24551), .Z(n39082) );
  XNOR U40200 ( .A(q[9]), .B(DB[1993]), .Z(n24551) );
  XNOR U40201 ( .A(q[12]), .B(DB[1996]), .Z(n24549) );
  IV U40202 ( .A(n24548), .Z(n39081) );
  XNOR U40203 ( .A(n24546), .B(n39083), .Z(n24548) );
  XNOR U40204 ( .A(q[11]), .B(DB[1995]), .Z(n39083) );
  XNOR U40205 ( .A(q[10]), .B(DB[1994]), .Z(n24546) );
  IV U40206 ( .A(n24561), .Z(n39076) );
  XOR U40207 ( .A(n39084), .B(n39085), .Z(n24561) );
  XNOR U40208 ( .A(n24578), .B(n24559), .Z(n39085) );
  XNOR U40209 ( .A(q[1]), .B(DB[1985]), .Z(n24559) );
  XOR U40210 ( .A(n39086), .B(n24567), .Z(n24578) );
  XNOR U40211 ( .A(q[8]), .B(DB[1992]), .Z(n24567) );
  IV U40212 ( .A(n24566), .Z(n39086) );
  XNOR U40213 ( .A(n24564), .B(n39087), .Z(n24566) );
  XNOR U40214 ( .A(q[7]), .B(DB[1991]), .Z(n39087) );
  XNOR U40215 ( .A(q[6]), .B(DB[1990]), .Z(n24564) );
  IV U40216 ( .A(n24577), .Z(n39084) );
  XOR U40217 ( .A(n39088), .B(n39089), .Z(n24577) );
  XNOR U40218 ( .A(n24573), .B(n24575), .Z(n39089) );
  XNOR U40219 ( .A(q[2]), .B(DB[1986]), .Z(n24575) );
  XNOR U40220 ( .A(q[5]), .B(DB[1989]), .Z(n24573) );
  IV U40221 ( .A(n24572), .Z(n39088) );
  XNOR U40222 ( .A(n24570), .B(n39090), .Z(n24572) );
  XNOR U40223 ( .A(q[4]), .B(DB[1988]), .Z(n39090) );
  XNOR U40224 ( .A(q[3]), .B(DB[1987]), .Z(n24570) );
  XOR U40225 ( .A(n39091), .B(n24339), .Z(n24190) );
  XOR U40226 ( .A(n39092), .B(n24315), .Z(n24339) );
  XOR U40227 ( .A(n39093), .B(n24307), .Z(n24315) );
  XOR U40228 ( .A(n39094), .B(n24296), .Z(n24307) );
  XNOR U40229 ( .A(q[30]), .B(DB[2045]), .Z(n24296) );
  IV U40230 ( .A(n24295), .Z(n39094) );
  XNOR U40231 ( .A(n24293), .B(n39095), .Z(n24295) );
  XNOR U40232 ( .A(q[29]), .B(DB[2044]), .Z(n39095) );
  XNOR U40233 ( .A(q[28]), .B(DB[2043]), .Z(n24293) );
  IV U40234 ( .A(n24306), .Z(n39093) );
  XOR U40235 ( .A(n39096), .B(n39097), .Z(n24306) );
  XNOR U40236 ( .A(n24302), .B(n24304), .Z(n39097) );
  XNOR U40237 ( .A(q[24]), .B(DB[2039]), .Z(n24304) );
  XNOR U40238 ( .A(q[27]), .B(DB[2042]), .Z(n24302) );
  IV U40239 ( .A(n24301), .Z(n39096) );
  XNOR U40240 ( .A(n24299), .B(n39098), .Z(n24301) );
  XNOR U40241 ( .A(q[26]), .B(DB[2041]), .Z(n39098) );
  XNOR U40242 ( .A(q[25]), .B(DB[2040]), .Z(n24299) );
  IV U40243 ( .A(n24314), .Z(n39092) );
  XOR U40244 ( .A(n39099), .B(n39100), .Z(n24314) );
  XNOR U40245 ( .A(n24331), .B(n24312), .Z(n39100) );
  XNOR U40246 ( .A(q[16]), .B(DB[2031]), .Z(n24312) );
  XOR U40247 ( .A(n39101), .B(n24320), .Z(n24331) );
  XNOR U40248 ( .A(q[23]), .B(DB[2038]), .Z(n24320) );
  IV U40249 ( .A(n24319), .Z(n39101) );
  XNOR U40250 ( .A(n24317), .B(n39102), .Z(n24319) );
  XNOR U40251 ( .A(q[22]), .B(DB[2037]), .Z(n39102) );
  XNOR U40252 ( .A(q[21]), .B(DB[2036]), .Z(n24317) );
  IV U40253 ( .A(n24330), .Z(n39099) );
  XOR U40254 ( .A(n39103), .B(n39104), .Z(n24330) );
  XNOR U40255 ( .A(n24326), .B(n24328), .Z(n39104) );
  XNOR U40256 ( .A(q[17]), .B(DB[2032]), .Z(n24328) );
  XNOR U40257 ( .A(q[20]), .B(DB[2035]), .Z(n24326) );
  IV U40258 ( .A(n24325), .Z(n39103) );
  XNOR U40259 ( .A(n24323), .B(n39105), .Z(n24325) );
  XNOR U40260 ( .A(q[19]), .B(DB[2034]), .Z(n39105) );
  XNOR U40261 ( .A(q[18]), .B(DB[2033]), .Z(n24323) );
  IV U40262 ( .A(n24338), .Z(n39091) );
  XOR U40263 ( .A(n39106), .B(n39107), .Z(n24338) );
  XNOR U40264 ( .A(n24365), .B(n24336), .Z(n39107) );
  XNOR U40265 ( .A(q[0]), .B(DB[2015]), .Z(n24336) );
  XOR U40266 ( .A(n39108), .B(n24357), .Z(n24365) );
  XOR U40267 ( .A(n39109), .B(n24345), .Z(n24357) );
  XNOR U40268 ( .A(q[15]), .B(DB[2030]), .Z(n24345) );
  IV U40269 ( .A(n24344), .Z(n39109) );
  XNOR U40270 ( .A(n24342), .B(n39110), .Z(n24344) );
  XNOR U40271 ( .A(q[14]), .B(DB[2029]), .Z(n39110) );
  XNOR U40272 ( .A(q[13]), .B(DB[2028]), .Z(n24342) );
  IV U40273 ( .A(n24356), .Z(n39108) );
  XOR U40274 ( .A(n39111), .B(n39112), .Z(n24356) );
  XNOR U40275 ( .A(n24352), .B(n24354), .Z(n39112) );
  XNOR U40276 ( .A(q[9]), .B(DB[2024]), .Z(n24354) );
  XNOR U40277 ( .A(q[12]), .B(DB[2027]), .Z(n24352) );
  IV U40278 ( .A(n24351), .Z(n39111) );
  XNOR U40279 ( .A(n24349), .B(n39113), .Z(n24351) );
  XNOR U40280 ( .A(q[11]), .B(DB[2026]), .Z(n39113) );
  XNOR U40281 ( .A(q[10]), .B(DB[2025]), .Z(n24349) );
  IV U40282 ( .A(n24364), .Z(n39106) );
  XOR U40283 ( .A(n39114), .B(n39115), .Z(n24364) );
  XNOR U40284 ( .A(n24381), .B(n24362), .Z(n39115) );
  XNOR U40285 ( .A(q[1]), .B(DB[2016]), .Z(n24362) );
  XOR U40286 ( .A(n39116), .B(n24370), .Z(n24381) );
  XNOR U40287 ( .A(q[8]), .B(DB[2023]), .Z(n24370) );
  IV U40288 ( .A(n24369), .Z(n39116) );
  XNOR U40289 ( .A(n24367), .B(n39117), .Z(n24369) );
  XNOR U40290 ( .A(q[7]), .B(DB[2022]), .Z(n39117) );
  XNOR U40291 ( .A(q[6]), .B(DB[2021]), .Z(n24367) );
  IV U40292 ( .A(n24380), .Z(n39114) );
  XOR U40293 ( .A(n39118), .B(n39119), .Z(n24380) );
  XNOR U40294 ( .A(n24376), .B(n24378), .Z(n39119) );
  XNOR U40295 ( .A(q[2]), .B(DB[2017]), .Z(n24378) );
  XNOR U40296 ( .A(q[5]), .B(DB[2020]), .Z(n24376) );
  IV U40297 ( .A(n24375), .Z(n39118) );
  XNOR U40298 ( .A(n24373), .B(n39120), .Z(n24375) );
  XNOR U40299 ( .A(q[4]), .B(DB[2019]), .Z(n39120) );
  XNOR U40300 ( .A(q[3]), .B(DB[2018]), .Z(n24373) );
  XOR U40301 ( .A(n39121), .B(n24142), .Z(n23993) );
  XOR U40302 ( .A(n39122), .B(n24118), .Z(n24142) );
  XOR U40303 ( .A(n39123), .B(n24110), .Z(n24118) );
  XOR U40304 ( .A(n39124), .B(n24099), .Z(n24110) );
  XNOR U40305 ( .A(q[30]), .B(DB[2076]), .Z(n24099) );
  IV U40306 ( .A(n24098), .Z(n39124) );
  XNOR U40307 ( .A(n24096), .B(n39125), .Z(n24098) );
  XNOR U40308 ( .A(q[29]), .B(DB[2075]), .Z(n39125) );
  XNOR U40309 ( .A(q[28]), .B(DB[2074]), .Z(n24096) );
  IV U40310 ( .A(n24109), .Z(n39123) );
  XOR U40311 ( .A(n39126), .B(n39127), .Z(n24109) );
  XNOR U40312 ( .A(n24105), .B(n24107), .Z(n39127) );
  XNOR U40313 ( .A(q[24]), .B(DB[2070]), .Z(n24107) );
  XNOR U40314 ( .A(q[27]), .B(DB[2073]), .Z(n24105) );
  IV U40315 ( .A(n24104), .Z(n39126) );
  XNOR U40316 ( .A(n24102), .B(n39128), .Z(n24104) );
  XNOR U40317 ( .A(q[26]), .B(DB[2072]), .Z(n39128) );
  XNOR U40318 ( .A(q[25]), .B(DB[2071]), .Z(n24102) );
  IV U40319 ( .A(n24117), .Z(n39122) );
  XOR U40320 ( .A(n39129), .B(n39130), .Z(n24117) );
  XNOR U40321 ( .A(n24134), .B(n24115), .Z(n39130) );
  XNOR U40322 ( .A(q[16]), .B(DB[2062]), .Z(n24115) );
  XOR U40323 ( .A(n39131), .B(n24123), .Z(n24134) );
  XNOR U40324 ( .A(q[23]), .B(DB[2069]), .Z(n24123) );
  IV U40325 ( .A(n24122), .Z(n39131) );
  XNOR U40326 ( .A(n24120), .B(n39132), .Z(n24122) );
  XNOR U40327 ( .A(q[22]), .B(DB[2068]), .Z(n39132) );
  XNOR U40328 ( .A(q[21]), .B(DB[2067]), .Z(n24120) );
  IV U40329 ( .A(n24133), .Z(n39129) );
  XOR U40330 ( .A(n39133), .B(n39134), .Z(n24133) );
  XNOR U40331 ( .A(n24129), .B(n24131), .Z(n39134) );
  XNOR U40332 ( .A(q[17]), .B(DB[2063]), .Z(n24131) );
  XNOR U40333 ( .A(q[20]), .B(DB[2066]), .Z(n24129) );
  IV U40334 ( .A(n24128), .Z(n39133) );
  XNOR U40335 ( .A(n24126), .B(n39135), .Z(n24128) );
  XNOR U40336 ( .A(q[19]), .B(DB[2065]), .Z(n39135) );
  XNOR U40337 ( .A(q[18]), .B(DB[2064]), .Z(n24126) );
  IV U40338 ( .A(n24141), .Z(n39121) );
  XOR U40339 ( .A(n39136), .B(n39137), .Z(n24141) );
  XNOR U40340 ( .A(n24168), .B(n24139), .Z(n39137) );
  XNOR U40341 ( .A(q[0]), .B(DB[2046]), .Z(n24139) );
  XOR U40342 ( .A(n39138), .B(n24160), .Z(n24168) );
  XOR U40343 ( .A(n39139), .B(n24148), .Z(n24160) );
  XNOR U40344 ( .A(q[15]), .B(DB[2061]), .Z(n24148) );
  IV U40345 ( .A(n24147), .Z(n39139) );
  XNOR U40346 ( .A(n24145), .B(n39140), .Z(n24147) );
  XNOR U40347 ( .A(q[14]), .B(DB[2060]), .Z(n39140) );
  XNOR U40348 ( .A(q[13]), .B(DB[2059]), .Z(n24145) );
  IV U40349 ( .A(n24159), .Z(n39138) );
  XOR U40350 ( .A(n39141), .B(n39142), .Z(n24159) );
  XNOR U40351 ( .A(n24155), .B(n24157), .Z(n39142) );
  XNOR U40352 ( .A(q[9]), .B(DB[2055]), .Z(n24157) );
  XNOR U40353 ( .A(q[12]), .B(DB[2058]), .Z(n24155) );
  IV U40354 ( .A(n24154), .Z(n39141) );
  XNOR U40355 ( .A(n24152), .B(n39143), .Z(n24154) );
  XNOR U40356 ( .A(q[11]), .B(DB[2057]), .Z(n39143) );
  XNOR U40357 ( .A(q[10]), .B(DB[2056]), .Z(n24152) );
  IV U40358 ( .A(n24167), .Z(n39136) );
  XOR U40359 ( .A(n39144), .B(n39145), .Z(n24167) );
  XNOR U40360 ( .A(n24184), .B(n24165), .Z(n39145) );
  XNOR U40361 ( .A(q[1]), .B(DB[2047]), .Z(n24165) );
  XOR U40362 ( .A(n39146), .B(n24173), .Z(n24184) );
  XNOR U40363 ( .A(q[8]), .B(DB[2054]), .Z(n24173) );
  IV U40364 ( .A(n24172), .Z(n39146) );
  XNOR U40365 ( .A(n24170), .B(n39147), .Z(n24172) );
  XNOR U40366 ( .A(q[7]), .B(DB[2053]), .Z(n39147) );
  XNOR U40367 ( .A(q[6]), .B(DB[2052]), .Z(n24170) );
  IV U40368 ( .A(n24183), .Z(n39144) );
  XOR U40369 ( .A(n39148), .B(n39149), .Z(n24183) );
  XNOR U40370 ( .A(n24179), .B(n24181), .Z(n39149) );
  XNOR U40371 ( .A(q[2]), .B(DB[2048]), .Z(n24181) );
  XNOR U40372 ( .A(q[5]), .B(DB[2051]), .Z(n24179) );
  IV U40373 ( .A(n24178), .Z(n39148) );
  XNOR U40374 ( .A(n24176), .B(n39150), .Z(n24178) );
  XNOR U40375 ( .A(q[4]), .B(DB[2050]), .Z(n39150) );
  XNOR U40376 ( .A(q[3]), .B(DB[2049]), .Z(n24176) );
  XOR U40377 ( .A(n39151), .B(n23945), .Z(n23796) );
  XOR U40378 ( .A(n39152), .B(n23921), .Z(n23945) );
  XOR U40379 ( .A(n39153), .B(n23913), .Z(n23921) );
  XOR U40380 ( .A(n39154), .B(n23902), .Z(n23913) );
  XNOR U40381 ( .A(q[30]), .B(DB[2107]), .Z(n23902) );
  IV U40382 ( .A(n23901), .Z(n39154) );
  XNOR U40383 ( .A(n23899), .B(n39155), .Z(n23901) );
  XNOR U40384 ( .A(q[29]), .B(DB[2106]), .Z(n39155) );
  XNOR U40385 ( .A(q[28]), .B(DB[2105]), .Z(n23899) );
  IV U40386 ( .A(n23912), .Z(n39153) );
  XOR U40387 ( .A(n39156), .B(n39157), .Z(n23912) );
  XNOR U40388 ( .A(n23908), .B(n23910), .Z(n39157) );
  XNOR U40389 ( .A(q[24]), .B(DB[2101]), .Z(n23910) );
  XNOR U40390 ( .A(q[27]), .B(DB[2104]), .Z(n23908) );
  IV U40391 ( .A(n23907), .Z(n39156) );
  XNOR U40392 ( .A(n23905), .B(n39158), .Z(n23907) );
  XNOR U40393 ( .A(q[26]), .B(DB[2103]), .Z(n39158) );
  XNOR U40394 ( .A(q[25]), .B(DB[2102]), .Z(n23905) );
  IV U40395 ( .A(n23920), .Z(n39152) );
  XOR U40396 ( .A(n39159), .B(n39160), .Z(n23920) );
  XNOR U40397 ( .A(n23937), .B(n23918), .Z(n39160) );
  XNOR U40398 ( .A(q[16]), .B(DB[2093]), .Z(n23918) );
  XOR U40399 ( .A(n39161), .B(n23926), .Z(n23937) );
  XNOR U40400 ( .A(q[23]), .B(DB[2100]), .Z(n23926) );
  IV U40401 ( .A(n23925), .Z(n39161) );
  XNOR U40402 ( .A(n23923), .B(n39162), .Z(n23925) );
  XNOR U40403 ( .A(q[22]), .B(DB[2099]), .Z(n39162) );
  XNOR U40404 ( .A(q[21]), .B(DB[2098]), .Z(n23923) );
  IV U40405 ( .A(n23936), .Z(n39159) );
  XOR U40406 ( .A(n39163), .B(n39164), .Z(n23936) );
  XNOR U40407 ( .A(n23932), .B(n23934), .Z(n39164) );
  XNOR U40408 ( .A(q[17]), .B(DB[2094]), .Z(n23934) );
  XNOR U40409 ( .A(q[20]), .B(DB[2097]), .Z(n23932) );
  IV U40410 ( .A(n23931), .Z(n39163) );
  XNOR U40411 ( .A(n23929), .B(n39165), .Z(n23931) );
  XNOR U40412 ( .A(q[19]), .B(DB[2096]), .Z(n39165) );
  XNOR U40413 ( .A(q[18]), .B(DB[2095]), .Z(n23929) );
  IV U40414 ( .A(n23944), .Z(n39151) );
  XOR U40415 ( .A(n39166), .B(n39167), .Z(n23944) );
  XNOR U40416 ( .A(n23971), .B(n23942), .Z(n39167) );
  XNOR U40417 ( .A(q[0]), .B(DB[2077]), .Z(n23942) );
  XOR U40418 ( .A(n39168), .B(n23963), .Z(n23971) );
  XOR U40419 ( .A(n39169), .B(n23951), .Z(n23963) );
  XNOR U40420 ( .A(q[15]), .B(DB[2092]), .Z(n23951) );
  IV U40421 ( .A(n23950), .Z(n39169) );
  XNOR U40422 ( .A(n23948), .B(n39170), .Z(n23950) );
  XNOR U40423 ( .A(q[14]), .B(DB[2091]), .Z(n39170) );
  XNOR U40424 ( .A(q[13]), .B(DB[2090]), .Z(n23948) );
  IV U40425 ( .A(n23962), .Z(n39168) );
  XOR U40426 ( .A(n39171), .B(n39172), .Z(n23962) );
  XNOR U40427 ( .A(n23958), .B(n23960), .Z(n39172) );
  XNOR U40428 ( .A(q[9]), .B(DB[2086]), .Z(n23960) );
  XNOR U40429 ( .A(q[12]), .B(DB[2089]), .Z(n23958) );
  IV U40430 ( .A(n23957), .Z(n39171) );
  XNOR U40431 ( .A(n23955), .B(n39173), .Z(n23957) );
  XNOR U40432 ( .A(q[11]), .B(DB[2088]), .Z(n39173) );
  XNOR U40433 ( .A(q[10]), .B(DB[2087]), .Z(n23955) );
  IV U40434 ( .A(n23970), .Z(n39166) );
  XOR U40435 ( .A(n39174), .B(n39175), .Z(n23970) );
  XNOR U40436 ( .A(n23987), .B(n23968), .Z(n39175) );
  XNOR U40437 ( .A(q[1]), .B(DB[2078]), .Z(n23968) );
  XOR U40438 ( .A(n39176), .B(n23976), .Z(n23987) );
  XNOR U40439 ( .A(q[8]), .B(DB[2085]), .Z(n23976) );
  IV U40440 ( .A(n23975), .Z(n39176) );
  XNOR U40441 ( .A(n23973), .B(n39177), .Z(n23975) );
  XNOR U40442 ( .A(q[7]), .B(DB[2084]), .Z(n39177) );
  XNOR U40443 ( .A(q[6]), .B(DB[2083]), .Z(n23973) );
  IV U40444 ( .A(n23986), .Z(n39174) );
  XOR U40445 ( .A(n39178), .B(n39179), .Z(n23986) );
  XNOR U40446 ( .A(n23982), .B(n23984), .Z(n39179) );
  XNOR U40447 ( .A(q[2]), .B(DB[2079]), .Z(n23984) );
  XNOR U40448 ( .A(q[5]), .B(DB[2082]), .Z(n23982) );
  IV U40449 ( .A(n23981), .Z(n39178) );
  XNOR U40450 ( .A(n23979), .B(n39180), .Z(n23981) );
  XNOR U40451 ( .A(q[4]), .B(DB[2081]), .Z(n39180) );
  XNOR U40452 ( .A(q[3]), .B(DB[2080]), .Z(n23979) );
  XOR U40453 ( .A(n39181), .B(n23748), .Z(n23599) );
  XOR U40454 ( .A(n39182), .B(n23724), .Z(n23748) );
  XOR U40455 ( .A(n39183), .B(n23716), .Z(n23724) );
  XOR U40456 ( .A(n39184), .B(n23705), .Z(n23716) );
  XNOR U40457 ( .A(q[30]), .B(DB[2138]), .Z(n23705) );
  IV U40458 ( .A(n23704), .Z(n39184) );
  XNOR U40459 ( .A(n23702), .B(n39185), .Z(n23704) );
  XNOR U40460 ( .A(q[29]), .B(DB[2137]), .Z(n39185) );
  XNOR U40461 ( .A(q[28]), .B(DB[2136]), .Z(n23702) );
  IV U40462 ( .A(n23715), .Z(n39183) );
  XOR U40463 ( .A(n39186), .B(n39187), .Z(n23715) );
  XNOR U40464 ( .A(n23711), .B(n23713), .Z(n39187) );
  XNOR U40465 ( .A(q[24]), .B(DB[2132]), .Z(n23713) );
  XNOR U40466 ( .A(q[27]), .B(DB[2135]), .Z(n23711) );
  IV U40467 ( .A(n23710), .Z(n39186) );
  XNOR U40468 ( .A(n23708), .B(n39188), .Z(n23710) );
  XNOR U40469 ( .A(q[26]), .B(DB[2134]), .Z(n39188) );
  XNOR U40470 ( .A(q[25]), .B(DB[2133]), .Z(n23708) );
  IV U40471 ( .A(n23723), .Z(n39182) );
  XOR U40472 ( .A(n39189), .B(n39190), .Z(n23723) );
  XNOR U40473 ( .A(n23740), .B(n23721), .Z(n39190) );
  XNOR U40474 ( .A(q[16]), .B(DB[2124]), .Z(n23721) );
  XOR U40475 ( .A(n39191), .B(n23729), .Z(n23740) );
  XNOR U40476 ( .A(q[23]), .B(DB[2131]), .Z(n23729) );
  IV U40477 ( .A(n23728), .Z(n39191) );
  XNOR U40478 ( .A(n23726), .B(n39192), .Z(n23728) );
  XNOR U40479 ( .A(q[22]), .B(DB[2130]), .Z(n39192) );
  XNOR U40480 ( .A(q[21]), .B(DB[2129]), .Z(n23726) );
  IV U40481 ( .A(n23739), .Z(n39189) );
  XOR U40482 ( .A(n39193), .B(n39194), .Z(n23739) );
  XNOR U40483 ( .A(n23735), .B(n23737), .Z(n39194) );
  XNOR U40484 ( .A(q[17]), .B(DB[2125]), .Z(n23737) );
  XNOR U40485 ( .A(q[20]), .B(DB[2128]), .Z(n23735) );
  IV U40486 ( .A(n23734), .Z(n39193) );
  XNOR U40487 ( .A(n23732), .B(n39195), .Z(n23734) );
  XNOR U40488 ( .A(q[19]), .B(DB[2127]), .Z(n39195) );
  XNOR U40489 ( .A(q[18]), .B(DB[2126]), .Z(n23732) );
  IV U40490 ( .A(n23747), .Z(n39181) );
  XOR U40491 ( .A(n39196), .B(n39197), .Z(n23747) );
  XNOR U40492 ( .A(n23774), .B(n23745), .Z(n39197) );
  XNOR U40493 ( .A(q[0]), .B(DB[2108]), .Z(n23745) );
  XOR U40494 ( .A(n39198), .B(n23766), .Z(n23774) );
  XOR U40495 ( .A(n39199), .B(n23754), .Z(n23766) );
  XNOR U40496 ( .A(q[15]), .B(DB[2123]), .Z(n23754) );
  IV U40497 ( .A(n23753), .Z(n39199) );
  XNOR U40498 ( .A(n23751), .B(n39200), .Z(n23753) );
  XNOR U40499 ( .A(q[14]), .B(DB[2122]), .Z(n39200) );
  XNOR U40500 ( .A(q[13]), .B(DB[2121]), .Z(n23751) );
  IV U40501 ( .A(n23765), .Z(n39198) );
  XOR U40502 ( .A(n39201), .B(n39202), .Z(n23765) );
  XNOR U40503 ( .A(n23761), .B(n23763), .Z(n39202) );
  XNOR U40504 ( .A(q[9]), .B(DB[2117]), .Z(n23763) );
  XNOR U40505 ( .A(q[12]), .B(DB[2120]), .Z(n23761) );
  IV U40506 ( .A(n23760), .Z(n39201) );
  XNOR U40507 ( .A(n23758), .B(n39203), .Z(n23760) );
  XNOR U40508 ( .A(q[11]), .B(DB[2119]), .Z(n39203) );
  XNOR U40509 ( .A(q[10]), .B(DB[2118]), .Z(n23758) );
  IV U40510 ( .A(n23773), .Z(n39196) );
  XOR U40511 ( .A(n39204), .B(n39205), .Z(n23773) );
  XNOR U40512 ( .A(n23790), .B(n23771), .Z(n39205) );
  XNOR U40513 ( .A(q[1]), .B(DB[2109]), .Z(n23771) );
  XOR U40514 ( .A(n39206), .B(n23779), .Z(n23790) );
  XNOR U40515 ( .A(q[8]), .B(DB[2116]), .Z(n23779) );
  IV U40516 ( .A(n23778), .Z(n39206) );
  XNOR U40517 ( .A(n23776), .B(n39207), .Z(n23778) );
  XNOR U40518 ( .A(q[7]), .B(DB[2115]), .Z(n39207) );
  XNOR U40519 ( .A(q[6]), .B(DB[2114]), .Z(n23776) );
  IV U40520 ( .A(n23789), .Z(n39204) );
  XOR U40521 ( .A(n39208), .B(n39209), .Z(n23789) );
  XNOR U40522 ( .A(n23785), .B(n23787), .Z(n39209) );
  XNOR U40523 ( .A(q[2]), .B(DB[2110]), .Z(n23787) );
  XNOR U40524 ( .A(q[5]), .B(DB[2113]), .Z(n23785) );
  IV U40525 ( .A(n23784), .Z(n39208) );
  XNOR U40526 ( .A(n23782), .B(n39210), .Z(n23784) );
  XNOR U40527 ( .A(q[4]), .B(DB[2112]), .Z(n39210) );
  XNOR U40528 ( .A(q[3]), .B(DB[2111]), .Z(n23782) );
  XOR U40529 ( .A(n39211), .B(n23551), .Z(n23402) );
  XOR U40530 ( .A(n39212), .B(n23527), .Z(n23551) );
  XOR U40531 ( .A(n39213), .B(n23519), .Z(n23527) );
  XOR U40532 ( .A(n39214), .B(n23508), .Z(n23519) );
  XNOR U40533 ( .A(q[30]), .B(DB[2169]), .Z(n23508) );
  IV U40534 ( .A(n23507), .Z(n39214) );
  XNOR U40535 ( .A(n23505), .B(n39215), .Z(n23507) );
  XNOR U40536 ( .A(q[29]), .B(DB[2168]), .Z(n39215) );
  XNOR U40537 ( .A(q[28]), .B(DB[2167]), .Z(n23505) );
  IV U40538 ( .A(n23518), .Z(n39213) );
  XOR U40539 ( .A(n39216), .B(n39217), .Z(n23518) );
  XNOR U40540 ( .A(n23514), .B(n23516), .Z(n39217) );
  XNOR U40541 ( .A(q[24]), .B(DB[2163]), .Z(n23516) );
  XNOR U40542 ( .A(q[27]), .B(DB[2166]), .Z(n23514) );
  IV U40543 ( .A(n23513), .Z(n39216) );
  XNOR U40544 ( .A(n23511), .B(n39218), .Z(n23513) );
  XNOR U40545 ( .A(q[26]), .B(DB[2165]), .Z(n39218) );
  XNOR U40546 ( .A(q[25]), .B(DB[2164]), .Z(n23511) );
  IV U40547 ( .A(n23526), .Z(n39212) );
  XOR U40548 ( .A(n39219), .B(n39220), .Z(n23526) );
  XNOR U40549 ( .A(n23543), .B(n23524), .Z(n39220) );
  XNOR U40550 ( .A(q[16]), .B(DB[2155]), .Z(n23524) );
  XOR U40551 ( .A(n39221), .B(n23532), .Z(n23543) );
  XNOR U40552 ( .A(q[23]), .B(DB[2162]), .Z(n23532) );
  IV U40553 ( .A(n23531), .Z(n39221) );
  XNOR U40554 ( .A(n23529), .B(n39222), .Z(n23531) );
  XNOR U40555 ( .A(q[22]), .B(DB[2161]), .Z(n39222) );
  XNOR U40556 ( .A(q[21]), .B(DB[2160]), .Z(n23529) );
  IV U40557 ( .A(n23542), .Z(n39219) );
  XOR U40558 ( .A(n39223), .B(n39224), .Z(n23542) );
  XNOR U40559 ( .A(n23538), .B(n23540), .Z(n39224) );
  XNOR U40560 ( .A(q[17]), .B(DB[2156]), .Z(n23540) );
  XNOR U40561 ( .A(q[20]), .B(DB[2159]), .Z(n23538) );
  IV U40562 ( .A(n23537), .Z(n39223) );
  XNOR U40563 ( .A(n23535), .B(n39225), .Z(n23537) );
  XNOR U40564 ( .A(q[19]), .B(DB[2158]), .Z(n39225) );
  XNOR U40565 ( .A(q[18]), .B(DB[2157]), .Z(n23535) );
  IV U40566 ( .A(n23550), .Z(n39211) );
  XOR U40567 ( .A(n39226), .B(n39227), .Z(n23550) );
  XNOR U40568 ( .A(n23577), .B(n23548), .Z(n39227) );
  XNOR U40569 ( .A(q[0]), .B(DB[2139]), .Z(n23548) );
  XOR U40570 ( .A(n39228), .B(n23569), .Z(n23577) );
  XOR U40571 ( .A(n39229), .B(n23557), .Z(n23569) );
  XNOR U40572 ( .A(q[15]), .B(DB[2154]), .Z(n23557) );
  IV U40573 ( .A(n23556), .Z(n39229) );
  XNOR U40574 ( .A(n23554), .B(n39230), .Z(n23556) );
  XNOR U40575 ( .A(q[14]), .B(DB[2153]), .Z(n39230) );
  XNOR U40576 ( .A(q[13]), .B(DB[2152]), .Z(n23554) );
  IV U40577 ( .A(n23568), .Z(n39228) );
  XOR U40578 ( .A(n39231), .B(n39232), .Z(n23568) );
  XNOR U40579 ( .A(n23564), .B(n23566), .Z(n39232) );
  XNOR U40580 ( .A(q[9]), .B(DB[2148]), .Z(n23566) );
  XNOR U40581 ( .A(q[12]), .B(DB[2151]), .Z(n23564) );
  IV U40582 ( .A(n23563), .Z(n39231) );
  XNOR U40583 ( .A(n23561), .B(n39233), .Z(n23563) );
  XNOR U40584 ( .A(q[11]), .B(DB[2150]), .Z(n39233) );
  XNOR U40585 ( .A(q[10]), .B(DB[2149]), .Z(n23561) );
  IV U40586 ( .A(n23576), .Z(n39226) );
  XOR U40587 ( .A(n39234), .B(n39235), .Z(n23576) );
  XNOR U40588 ( .A(n23593), .B(n23574), .Z(n39235) );
  XNOR U40589 ( .A(q[1]), .B(DB[2140]), .Z(n23574) );
  XOR U40590 ( .A(n39236), .B(n23582), .Z(n23593) );
  XNOR U40591 ( .A(q[8]), .B(DB[2147]), .Z(n23582) );
  IV U40592 ( .A(n23581), .Z(n39236) );
  XNOR U40593 ( .A(n23579), .B(n39237), .Z(n23581) );
  XNOR U40594 ( .A(q[7]), .B(DB[2146]), .Z(n39237) );
  XNOR U40595 ( .A(q[6]), .B(DB[2145]), .Z(n23579) );
  IV U40596 ( .A(n23592), .Z(n39234) );
  XOR U40597 ( .A(n39238), .B(n39239), .Z(n23592) );
  XNOR U40598 ( .A(n23588), .B(n23590), .Z(n39239) );
  XNOR U40599 ( .A(q[2]), .B(DB[2141]), .Z(n23590) );
  XNOR U40600 ( .A(q[5]), .B(DB[2144]), .Z(n23588) );
  IV U40601 ( .A(n23587), .Z(n39238) );
  XNOR U40602 ( .A(n23585), .B(n39240), .Z(n23587) );
  XNOR U40603 ( .A(q[4]), .B(DB[2143]), .Z(n39240) );
  XNOR U40604 ( .A(q[3]), .B(DB[2142]), .Z(n23585) );
  XOR U40605 ( .A(n39241), .B(n23354), .Z(n23205) );
  XOR U40606 ( .A(n39242), .B(n23330), .Z(n23354) );
  XOR U40607 ( .A(n39243), .B(n23322), .Z(n23330) );
  XOR U40608 ( .A(n39244), .B(n23311), .Z(n23322) );
  XNOR U40609 ( .A(q[30]), .B(DB[2200]), .Z(n23311) );
  IV U40610 ( .A(n23310), .Z(n39244) );
  XNOR U40611 ( .A(n23308), .B(n39245), .Z(n23310) );
  XNOR U40612 ( .A(q[29]), .B(DB[2199]), .Z(n39245) );
  XNOR U40613 ( .A(q[28]), .B(DB[2198]), .Z(n23308) );
  IV U40614 ( .A(n23321), .Z(n39243) );
  XOR U40615 ( .A(n39246), .B(n39247), .Z(n23321) );
  XNOR U40616 ( .A(n23317), .B(n23319), .Z(n39247) );
  XNOR U40617 ( .A(q[24]), .B(DB[2194]), .Z(n23319) );
  XNOR U40618 ( .A(q[27]), .B(DB[2197]), .Z(n23317) );
  IV U40619 ( .A(n23316), .Z(n39246) );
  XNOR U40620 ( .A(n23314), .B(n39248), .Z(n23316) );
  XNOR U40621 ( .A(q[26]), .B(DB[2196]), .Z(n39248) );
  XNOR U40622 ( .A(q[25]), .B(DB[2195]), .Z(n23314) );
  IV U40623 ( .A(n23329), .Z(n39242) );
  XOR U40624 ( .A(n39249), .B(n39250), .Z(n23329) );
  XNOR U40625 ( .A(n23346), .B(n23327), .Z(n39250) );
  XNOR U40626 ( .A(q[16]), .B(DB[2186]), .Z(n23327) );
  XOR U40627 ( .A(n39251), .B(n23335), .Z(n23346) );
  XNOR U40628 ( .A(q[23]), .B(DB[2193]), .Z(n23335) );
  IV U40629 ( .A(n23334), .Z(n39251) );
  XNOR U40630 ( .A(n23332), .B(n39252), .Z(n23334) );
  XNOR U40631 ( .A(q[22]), .B(DB[2192]), .Z(n39252) );
  XNOR U40632 ( .A(q[21]), .B(DB[2191]), .Z(n23332) );
  IV U40633 ( .A(n23345), .Z(n39249) );
  XOR U40634 ( .A(n39253), .B(n39254), .Z(n23345) );
  XNOR U40635 ( .A(n23341), .B(n23343), .Z(n39254) );
  XNOR U40636 ( .A(q[17]), .B(DB[2187]), .Z(n23343) );
  XNOR U40637 ( .A(q[20]), .B(DB[2190]), .Z(n23341) );
  IV U40638 ( .A(n23340), .Z(n39253) );
  XNOR U40639 ( .A(n23338), .B(n39255), .Z(n23340) );
  XNOR U40640 ( .A(q[19]), .B(DB[2189]), .Z(n39255) );
  XNOR U40641 ( .A(q[18]), .B(DB[2188]), .Z(n23338) );
  IV U40642 ( .A(n23353), .Z(n39241) );
  XOR U40643 ( .A(n39256), .B(n39257), .Z(n23353) );
  XNOR U40644 ( .A(n23380), .B(n23351), .Z(n39257) );
  XNOR U40645 ( .A(q[0]), .B(DB[2170]), .Z(n23351) );
  XOR U40646 ( .A(n39258), .B(n23372), .Z(n23380) );
  XOR U40647 ( .A(n39259), .B(n23360), .Z(n23372) );
  XNOR U40648 ( .A(q[15]), .B(DB[2185]), .Z(n23360) );
  IV U40649 ( .A(n23359), .Z(n39259) );
  XNOR U40650 ( .A(n23357), .B(n39260), .Z(n23359) );
  XNOR U40651 ( .A(q[14]), .B(DB[2184]), .Z(n39260) );
  XNOR U40652 ( .A(q[13]), .B(DB[2183]), .Z(n23357) );
  IV U40653 ( .A(n23371), .Z(n39258) );
  XOR U40654 ( .A(n39261), .B(n39262), .Z(n23371) );
  XNOR U40655 ( .A(n23367), .B(n23369), .Z(n39262) );
  XNOR U40656 ( .A(q[9]), .B(DB[2179]), .Z(n23369) );
  XNOR U40657 ( .A(q[12]), .B(DB[2182]), .Z(n23367) );
  IV U40658 ( .A(n23366), .Z(n39261) );
  XNOR U40659 ( .A(n23364), .B(n39263), .Z(n23366) );
  XNOR U40660 ( .A(q[11]), .B(DB[2181]), .Z(n39263) );
  XNOR U40661 ( .A(q[10]), .B(DB[2180]), .Z(n23364) );
  IV U40662 ( .A(n23379), .Z(n39256) );
  XOR U40663 ( .A(n39264), .B(n39265), .Z(n23379) );
  XNOR U40664 ( .A(n23396), .B(n23377), .Z(n39265) );
  XNOR U40665 ( .A(q[1]), .B(DB[2171]), .Z(n23377) );
  XOR U40666 ( .A(n39266), .B(n23385), .Z(n23396) );
  XNOR U40667 ( .A(q[8]), .B(DB[2178]), .Z(n23385) );
  IV U40668 ( .A(n23384), .Z(n39266) );
  XNOR U40669 ( .A(n23382), .B(n39267), .Z(n23384) );
  XNOR U40670 ( .A(q[7]), .B(DB[2177]), .Z(n39267) );
  XNOR U40671 ( .A(q[6]), .B(DB[2176]), .Z(n23382) );
  IV U40672 ( .A(n23395), .Z(n39264) );
  XOR U40673 ( .A(n39268), .B(n39269), .Z(n23395) );
  XNOR U40674 ( .A(n23391), .B(n23393), .Z(n39269) );
  XNOR U40675 ( .A(q[2]), .B(DB[2172]), .Z(n23393) );
  XNOR U40676 ( .A(q[5]), .B(DB[2175]), .Z(n23391) );
  IV U40677 ( .A(n23390), .Z(n39268) );
  XNOR U40678 ( .A(n23388), .B(n39270), .Z(n23390) );
  XNOR U40679 ( .A(q[4]), .B(DB[2174]), .Z(n39270) );
  XNOR U40680 ( .A(q[3]), .B(DB[2173]), .Z(n23388) );
  XOR U40681 ( .A(n39271), .B(n23157), .Z(n23008) );
  XOR U40682 ( .A(n39272), .B(n23133), .Z(n23157) );
  XOR U40683 ( .A(n39273), .B(n23125), .Z(n23133) );
  XOR U40684 ( .A(n39274), .B(n23114), .Z(n23125) );
  XNOR U40685 ( .A(q[30]), .B(DB[2231]), .Z(n23114) );
  IV U40686 ( .A(n23113), .Z(n39274) );
  XNOR U40687 ( .A(n23111), .B(n39275), .Z(n23113) );
  XNOR U40688 ( .A(q[29]), .B(DB[2230]), .Z(n39275) );
  XNOR U40689 ( .A(q[28]), .B(DB[2229]), .Z(n23111) );
  IV U40690 ( .A(n23124), .Z(n39273) );
  XOR U40691 ( .A(n39276), .B(n39277), .Z(n23124) );
  XNOR U40692 ( .A(n23120), .B(n23122), .Z(n39277) );
  XNOR U40693 ( .A(q[24]), .B(DB[2225]), .Z(n23122) );
  XNOR U40694 ( .A(q[27]), .B(DB[2228]), .Z(n23120) );
  IV U40695 ( .A(n23119), .Z(n39276) );
  XNOR U40696 ( .A(n23117), .B(n39278), .Z(n23119) );
  XNOR U40697 ( .A(q[26]), .B(DB[2227]), .Z(n39278) );
  XNOR U40698 ( .A(q[25]), .B(DB[2226]), .Z(n23117) );
  IV U40699 ( .A(n23132), .Z(n39272) );
  XOR U40700 ( .A(n39279), .B(n39280), .Z(n23132) );
  XNOR U40701 ( .A(n23149), .B(n23130), .Z(n39280) );
  XNOR U40702 ( .A(q[16]), .B(DB[2217]), .Z(n23130) );
  XOR U40703 ( .A(n39281), .B(n23138), .Z(n23149) );
  XNOR U40704 ( .A(q[23]), .B(DB[2224]), .Z(n23138) );
  IV U40705 ( .A(n23137), .Z(n39281) );
  XNOR U40706 ( .A(n23135), .B(n39282), .Z(n23137) );
  XNOR U40707 ( .A(q[22]), .B(DB[2223]), .Z(n39282) );
  XNOR U40708 ( .A(q[21]), .B(DB[2222]), .Z(n23135) );
  IV U40709 ( .A(n23148), .Z(n39279) );
  XOR U40710 ( .A(n39283), .B(n39284), .Z(n23148) );
  XNOR U40711 ( .A(n23144), .B(n23146), .Z(n39284) );
  XNOR U40712 ( .A(q[17]), .B(DB[2218]), .Z(n23146) );
  XNOR U40713 ( .A(q[20]), .B(DB[2221]), .Z(n23144) );
  IV U40714 ( .A(n23143), .Z(n39283) );
  XNOR U40715 ( .A(n23141), .B(n39285), .Z(n23143) );
  XNOR U40716 ( .A(q[19]), .B(DB[2220]), .Z(n39285) );
  XNOR U40717 ( .A(q[18]), .B(DB[2219]), .Z(n23141) );
  IV U40718 ( .A(n23156), .Z(n39271) );
  XOR U40719 ( .A(n39286), .B(n39287), .Z(n23156) );
  XNOR U40720 ( .A(n23183), .B(n23154), .Z(n39287) );
  XNOR U40721 ( .A(q[0]), .B(DB[2201]), .Z(n23154) );
  XOR U40722 ( .A(n39288), .B(n23175), .Z(n23183) );
  XOR U40723 ( .A(n39289), .B(n23163), .Z(n23175) );
  XNOR U40724 ( .A(q[15]), .B(DB[2216]), .Z(n23163) );
  IV U40725 ( .A(n23162), .Z(n39289) );
  XNOR U40726 ( .A(n23160), .B(n39290), .Z(n23162) );
  XNOR U40727 ( .A(q[14]), .B(DB[2215]), .Z(n39290) );
  XNOR U40728 ( .A(q[13]), .B(DB[2214]), .Z(n23160) );
  IV U40729 ( .A(n23174), .Z(n39288) );
  XOR U40730 ( .A(n39291), .B(n39292), .Z(n23174) );
  XNOR U40731 ( .A(n23170), .B(n23172), .Z(n39292) );
  XNOR U40732 ( .A(q[9]), .B(DB[2210]), .Z(n23172) );
  XNOR U40733 ( .A(q[12]), .B(DB[2213]), .Z(n23170) );
  IV U40734 ( .A(n23169), .Z(n39291) );
  XNOR U40735 ( .A(n23167), .B(n39293), .Z(n23169) );
  XNOR U40736 ( .A(q[11]), .B(DB[2212]), .Z(n39293) );
  XNOR U40737 ( .A(q[10]), .B(DB[2211]), .Z(n23167) );
  IV U40738 ( .A(n23182), .Z(n39286) );
  XOR U40739 ( .A(n39294), .B(n39295), .Z(n23182) );
  XNOR U40740 ( .A(n23199), .B(n23180), .Z(n39295) );
  XNOR U40741 ( .A(q[1]), .B(DB[2202]), .Z(n23180) );
  XOR U40742 ( .A(n39296), .B(n23188), .Z(n23199) );
  XNOR U40743 ( .A(q[8]), .B(DB[2209]), .Z(n23188) );
  IV U40744 ( .A(n23187), .Z(n39296) );
  XNOR U40745 ( .A(n23185), .B(n39297), .Z(n23187) );
  XNOR U40746 ( .A(q[7]), .B(DB[2208]), .Z(n39297) );
  XNOR U40747 ( .A(q[6]), .B(DB[2207]), .Z(n23185) );
  IV U40748 ( .A(n23198), .Z(n39294) );
  XOR U40749 ( .A(n39298), .B(n39299), .Z(n23198) );
  XNOR U40750 ( .A(n23194), .B(n23196), .Z(n39299) );
  XNOR U40751 ( .A(q[2]), .B(DB[2203]), .Z(n23196) );
  XNOR U40752 ( .A(q[5]), .B(DB[2206]), .Z(n23194) );
  IV U40753 ( .A(n23193), .Z(n39298) );
  XNOR U40754 ( .A(n23191), .B(n39300), .Z(n23193) );
  XNOR U40755 ( .A(q[4]), .B(DB[2205]), .Z(n39300) );
  XNOR U40756 ( .A(q[3]), .B(DB[2204]), .Z(n23191) );
  XOR U40757 ( .A(n39301), .B(n22960), .Z(n22811) );
  XOR U40758 ( .A(n39302), .B(n22936), .Z(n22960) );
  XOR U40759 ( .A(n39303), .B(n22928), .Z(n22936) );
  XOR U40760 ( .A(n39304), .B(n22917), .Z(n22928) );
  XNOR U40761 ( .A(q[30]), .B(DB[2262]), .Z(n22917) );
  IV U40762 ( .A(n22916), .Z(n39304) );
  XNOR U40763 ( .A(n22914), .B(n39305), .Z(n22916) );
  XNOR U40764 ( .A(q[29]), .B(DB[2261]), .Z(n39305) );
  XNOR U40765 ( .A(q[28]), .B(DB[2260]), .Z(n22914) );
  IV U40766 ( .A(n22927), .Z(n39303) );
  XOR U40767 ( .A(n39306), .B(n39307), .Z(n22927) );
  XNOR U40768 ( .A(n22923), .B(n22925), .Z(n39307) );
  XNOR U40769 ( .A(q[24]), .B(DB[2256]), .Z(n22925) );
  XNOR U40770 ( .A(q[27]), .B(DB[2259]), .Z(n22923) );
  IV U40771 ( .A(n22922), .Z(n39306) );
  XNOR U40772 ( .A(n22920), .B(n39308), .Z(n22922) );
  XNOR U40773 ( .A(q[26]), .B(DB[2258]), .Z(n39308) );
  XNOR U40774 ( .A(q[25]), .B(DB[2257]), .Z(n22920) );
  IV U40775 ( .A(n22935), .Z(n39302) );
  XOR U40776 ( .A(n39309), .B(n39310), .Z(n22935) );
  XNOR U40777 ( .A(n22952), .B(n22933), .Z(n39310) );
  XNOR U40778 ( .A(q[16]), .B(DB[2248]), .Z(n22933) );
  XOR U40779 ( .A(n39311), .B(n22941), .Z(n22952) );
  XNOR U40780 ( .A(q[23]), .B(DB[2255]), .Z(n22941) );
  IV U40781 ( .A(n22940), .Z(n39311) );
  XNOR U40782 ( .A(n22938), .B(n39312), .Z(n22940) );
  XNOR U40783 ( .A(q[22]), .B(DB[2254]), .Z(n39312) );
  XNOR U40784 ( .A(q[21]), .B(DB[2253]), .Z(n22938) );
  IV U40785 ( .A(n22951), .Z(n39309) );
  XOR U40786 ( .A(n39313), .B(n39314), .Z(n22951) );
  XNOR U40787 ( .A(n22947), .B(n22949), .Z(n39314) );
  XNOR U40788 ( .A(q[17]), .B(DB[2249]), .Z(n22949) );
  XNOR U40789 ( .A(q[20]), .B(DB[2252]), .Z(n22947) );
  IV U40790 ( .A(n22946), .Z(n39313) );
  XNOR U40791 ( .A(n22944), .B(n39315), .Z(n22946) );
  XNOR U40792 ( .A(q[19]), .B(DB[2251]), .Z(n39315) );
  XNOR U40793 ( .A(q[18]), .B(DB[2250]), .Z(n22944) );
  IV U40794 ( .A(n22959), .Z(n39301) );
  XOR U40795 ( .A(n39316), .B(n39317), .Z(n22959) );
  XNOR U40796 ( .A(n22986), .B(n22957), .Z(n39317) );
  XNOR U40797 ( .A(q[0]), .B(DB[2232]), .Z(n22957) );
  XOR U40798 ( .A(n39318), .B(n22978), .Z(n22986) );
  XOR U40799 ( .A(n39319), .B(n22966), .Z(n22978) );
  XNOR U40800 ( .A(q[15]), .B(DB[2247]), .Z(n22966) );
  IV U40801 ( .A(n22965), .Z(n39319) );
  XNOR U40802 ( .A(n22963), .B(n39320), .Z(n22965) );
  XNOR U40803 ( .A(q[14]), .B(DB[2246]), .Z(n39320) );
  XNOR U40804 ( .A(q[13]), .B(DB[2245]), .Z(n22963) );
  IV U40805 ( .A(n22977), .Z(n39318) );
  XOR U40806 ( .A(n39321), .B(n39322), .Z(n22977) );
  XNOR U40807 ( .A(n22973), .B(n22975), .Z(n39322) );
  XNOR U40808 ( .A(q[9]), .B(DB[2241]), .Z(n22975) );
  XNOR U40809 ( .A(q[12]), .B(DB[2244]), .Z(n22973) );
  IV U40810 ( .A(n22972), .Z(n39321) );
  XNOR U40811 ( .A(n22970), .B(n39323), .Z(n22972) );
  XNOR U40812 ( .A(q[11]), .B(DB[2243]), .Z(n39323) );
  XNOR U40813 ( .A(q[10]), .B(DB[2242]), .Z(n22970) );
  IV U40814 ( .A(n22985), .Z(n39316) );
  XOR U40815 ( .A(n39324), .B(n39325), .Z(n22985) );
  XNOR U40816 ( .A(n23002), .B(n22983), .Z(n39325) );
  XNOR U40817 ( .A(q[1]), .B(DB[2233]), .Z(n22983) );
  XOR U40818 ( .A(n39326), .B(n22991), .Z(n23002) );
  XNOR U40819 ( .A(q[8]), .B(DB[2240]), .Z(n22991) );
  IV U40820 ( .A(n22990), .Z(n39326) );
  XNOR U40821 ( .A(n22988), .B(n39327), .Z(n22990) );
  XNOR U40822 ( .A(q[7]), .B(DB[2239]), .Z(n39327) );
  XNOR U40823 ( .A(q[6]), .B(DB[2238]), .Z(n22988) );
  IV U40824 ( .A(n23001), .Z(n39324) );
  XOR U40825 ( .A(n39328), .B(n39329), .Z(n23001) );
  XNOR U40826 ( .A(n22997), .B(n22999), .Z(n39329) );
  XNOR U40827 ( .A(q[2]), .B(DB[2234]), .Z(n22999) );
  XNOR U40828 ( .A(q[5]), .B(DB[2237]), .Z(n22997) );
  IV U40829 ( .A(n22996), .Z(n39328) );
  XNOR U40830 ( .A(n22994), .B(n39330), .Z(n22996) );
  XNOR U40831 ( .A(q[4]), .B(DB[2236]), .Z(n39330) );
  XNOR U40832 ( .A(q[3]), .B(DB[2235]), .Z(n22994) );
  XOR U40833 ( .A(n39331), .B(n22763), .Z(n22614) );
  XOR U40834 ( .A(n39332), .B(n22739), .Z(n22763) );
  XOR U40835 ( .A(n39333), .B(n22731), .Z(n22739) );
  XOR U40836 ( .A(n39334), .B(n22720), .Z(n22731) );
  XNOR U40837 ( .A(q[30]), .B(DB[2293]), .Z(n22720) );
  IV U40838 ( .A(n22719), .Z(n39334) );
  XNOR U40839 ( .A(n22717), .B(n39335), .Z(n22719) );
  XNOR U40840 ( .A(q[29]), .B(DB[2292]), .Z(n39335) );
  XNOR U40841 ( .A(q[28]), .B(DB[2291]), .Z(n22717) );
  IV U40842 ( .A(n22730), .Z(n39333) );
  XOR U40843 ( .A(n39336), .B(n39337), .Z(n22730) );
  XNOR U40844 ( .A(n22726), .B(n22728), .Z(n39337) );
  XNOR U40845 ( .A(q[24]), .B(DB[2287]), .Z(n22728) );
  XNOR U40846 ( .A(q[27]), .B(DB[2290]), .Z(n22726) );
  IV U40847 ( .A(n22725), .Z(n39336) );
  XNOR U40848 ( .A(n22723), .B(n39338), .Z(n22725) );
  XNOR U40849 ( .A(q[26]), .B(DB[2289]), .Z(n39338) );
  XNOR U40850 ( .A(q[25]), .B(DB[2288]), .Z(n22723) );
  IV U40851 ( .A(n22738), .Z(n39332) );
  XOR U40852 ( .A(n39339), .B(n39340), .Z(n22738) );
  XNOR U40853 ( .A(n22755), .B(n22736), .Z(n39340) );
  XNOR U40854 ( .A(q[16]), .B(DB[2279]), .Z(n22736) );
  XOR U40855 ( .A(n39341), .B(n22744), .Z(n22755) );
  XNOR U40856 ( .A(q[23]), .B(DB[2286]), .Z(n22744) );
  IV U40857 ( .A(n22743), .Z(n39341) );
  XNOR U40858 ( .A(n22741), .B(n39342), .Z(n22743) );
  XNOR U40859 ( .A(q[22]), .B(DB[2285]), .Z(n39342) );
  XNOR U40860 ( .A(q[21]), .B(DB[2284]), .Z(n22741) );
  IV U40861 ( .A(n22754), .Z(n39339) );
  XOR U40862 ( .A(n39343), .B(n39344), .Z(n22754) );
  XNOR U40863 ( .A(n22750), .B(n22752), .Z(n39344) );
  XNOR U40864 ( .A(q[17]), .B(DB[2280]), .Z(n22752) );
  XNOR U40865 ( .A(q[20]), .B(DB[2283]), .Z(n22750) );
  IV U40866 ( .A(n22749), .Z(n39343) );
  XNOR U40867 ( .A(n22747), .B(n39345), .Z(n22749) );
  XNOR U40868 ( .A(q[19]), .B(DB[2282]), .Z(n39345) );
  XNOR U40869 ( .A(q[18]), .B(DB[2281]), .Z(n22747) );
  IV U40870 ( .A(n22762), .Z(n39331) );
  XOR U40871 ( .A(n39346), .B(n39347), .Z(n22762) );
  XNOR U40872 ( .A(n22789), .B(n22760), .Z(n39347) );
  XNOR U40873 ( .A(q[0]), .B(DB[2263]), .Z(n22760) );
  XOR U40874 ( .A(n39348), .B(n22781), .Z(n22789) );
  XOR U40875 ( .A(n39349), .B(n22769), .Z(n22781) );
  XNOR U40876 ( .A(q[15]), .B(DB[2278]), .Z(n22769) );
  IV U40877 ( .A(n22768), .Z(n39349) );
  XNOR U40878 ( .A(n22766), .B(n39350), .Z(n22768) );
  XNOR U40879 ( .A(q[14]), .B(DB[2277]), .Z(n39350) );
  XNOR U40880 ( .A(q[13]), .B(DB[2276]), .Z(n22766) );
  IV U40881 ( .A(n22780), .Z(n39348) );
  XOR U40882 ( .A(n39351), .B(n39352), .Z(n22780) );
  XNOR U40883 ( .A(n22776), .B(n22778), .Z(n39352) );
  XNOR U40884 ( .A(q[9]), .B(DB[2272]), .Z(n22778) );
  XNOR U40885 ( .A(q[12]), .B(DB[2275]), .Z(n22776) );
  IV U40886 ( .A(n22775), .Z(n39351) );
  XNOR U40887 ( .A(n22773), .B(n39353), .Z(n22775) );
  XNOR U40888 ( .A(q[11]), .B(DB[2274]), .Z(n39353) );
  XNOR U40889 ( .A(q[10]), .B(DB[2273]), .Z(n22773) );
  IV U40890 ( .A(n22788), .Z(n39346) );
  XOR U40891 ( .A(n39354), .B(n39355), .Z(n22788) );
  XNOR U40892 ( .A(n22805), .B(n22786), .Z(n39355) );
  XNOR U40893 ( .A(q[1]), .B(DB[2264]), .Z(n22786) );
  XOR U40894 ( .A(n39356), .B(n22794), .Z(n22805) );
  XNOR U40895 ( .A(q[8]), .B(DB[2271]), .Z(n22794) );
  IV U40896 ( .A(n22793), .Z(n39356) );
  XNOR U40897 ( .A(n22791), .B(n39357), .Z(n22793) );
  XNOR U40898 ( .A(q[7]), .B(DB[2270]), .Z(n39357) );
  XNOR U40899 ( .A(q[6]), .B(DB[2269]), .Z(n22791) );
  IV U40900 ( .A(n22804), .Z(n39354) );
  XOR U40901 ( .A(n39358), .B(n39359), .Z(n22804) );
  XNOR U40902 ( .A(n22800), .B(n22802), .Z(n39359) );
  XNOR U40903 ( .A(q[2]), .B(DB[2265]), .Z(n22802) );
  XNOR U40904 ( .A(q[5]), .B(DB[2268]), .Z(n22800) );
  IV U40905 ( .A(n22799), .Z(n39358) );
  XNOR U40906 ( .A(n22797), .B(n39360), .Z(n22799) );
  XNOR U40907 ( .A(q[4]), .B(DB[2267]), .Z(n39360) );
  XNOR U40908 ( .A(q[3]), .B(DB[2266]), .Z(n22797) );
  XOR U40909 ( .A(n39361), .B(n22566), .Z(n22417) );
  XOR U40910 ( .A(n39362), .B(n22542), .Z(n22566) );
  XOR U40911 ( .A(n39363), .B(n22534), .Z(n22542) );
  XOR U40912 ( .A(n39364), .B(n22523), .Z(n22534) );
  XNOR U40913 ( .A(q[30]), .B(DB[2324]), .Z(n22523) );
  IV U40914 ( .A(n22522), .Z(n39364) );
  XNOR U40915 ( .A(n22520), .B(n39365), .Z(n22522) );
  XNOR U40916 ( .A(q[29]), .B(DB[2323]), .Z(n39365) );
  XNOR U40917 ( .A(q[28]), .B(DB[2322]), .Z(n22520) );
  IV U40918 ( .A(n22533), .Z(n39363) );
  XOR U40919 ( .A(n39366), .B(n39367), .Z(n22533) );
  XNOR U40920 ( .A(n22529), .B(n22531), .Z(n39367) );
  XNOR U40921 ( .A(q[24]), .B(DB[2318]), .Z(n22531) );
  XNOR U40922 ( .A(q[27]), .B(DB[2321]), .Z(n22529) );
  IV U40923 ( .A(n22528), .Z(n39366) );
  XNOR U40924 ( .A(n22526), .B(n39368), .Z(n22528) );
  XNOR U40925 ( .A(q[26]), .B(DB[2320]), .Z(n39368) );
  XNOR U40926 ( .A(q[25]), .B(DB[2319]), .Z(n22526) );
  IV U40927 ( .A(n22541), .Z(n39362) );
  XOR U40928 ( .A(n39369), .B(n39370), .Z(n22541) );
  XNOR U40929 ( .A(n22558), .B(n22539), .Z(n39370) );
  XNOR U40930 ( .A(q[16]), .B(DB[2310]), .Z(n22539) );
  XOR U40931 ( .A(n39371), .B(n22547), .Z(n22558) );
  XNOR U40932 ( .A(q[23]), .B(DB[2317]), .Z(n22547) );
  IV U40933 ( .A(n22546), .Z(n39371) );
  XNOR U40934 ( .A(n22544), .B(n39372), .Z(n22546) );
  XNOR U40935 ( .A(q[22]), .B(DB[2316]), .Z(n39372) );
  XNOR U40936 ( .A(q[21]), .B(DB[2315]), .Z(n22544) );
  IV U40937 ( .A(n22557), .Z(n39369) );
  XOR U40938 ( .A(n39373), .B(n39374), .Z(n22557) );
  XNOR U40939 ( .A(n22553), .B(n22555), .Z(n39374) );
  XNOR U40940 ( .A(q[17]), .B(DB[2311]), .Z(n22555) );
  XNOR U40941 ( .A(q[20]), .B(DB[2314]), .Z(n22553) );
  IV U40942 ( .A(n22552), .Z(n39373) );
  XNOR U40943 ( .A(n22550), .B(n39375), .Z(n22552) );
  XNOR U40944 ( .A(q[19]), .B(DB[2313]), .Z(n39375) );
  XNOR U40945 ( .A(q[18]), .B(DB[2312]), .Z(n22550) );
  IV U40946 ( .A(n22565), .Z(n39361) );
  XOR U40947 ( .A(n39376), .B(n39377), .Z(n22565) );
  XNOR U40948 ( .A(n22592), .B(n22563), .Z(n39377) );
  XNOR U40949 ( .A(q[0]), .B(DB[2294]), .Z(n22563) );
  XOR U40950 ( .A(n39378), .B(n22584), .Z(n22592) );
  XOR U40951 ( .A(n39379), .B(n22572), .Z(n22584) );
  XNOR U40952 ( .A(q[15]), .B(DB[2309]), .Z(n22572) );
  IV U40953 ( .A(n22571), .Z(n39379) );
  XNOR U40954 ( .A(n22569), .B(n39380), .Z(n22571) );
  XNOR U40955 ( .A(q[14]), .B(DB[2308]), .Z(n39380) );
  XNOR U40956 ( .A(q[13]), .B(DB[2307]), .Z(n22569) );
  IV U40957 ( .A(n22583), .Z(n39378) );
  XOR U40958 ( .A(n39381), .B(n39382), .Z(n22583) );
  XNOR U40959 ( .A(n22579), .B(n22581), .Z(n39382) );
  XNOR U40960 ( .A(q[9]), .B(DB[2303]), .Z(n22581) );
  XNOR U40961 ( .A(q[12]), .B(DB[2306]), .Z(n22579) );
  IV U40962 ( .A(n22578), .Z(n39381) );
  XNOR U40963 ( .A(n22576), .B(n39383), .Z(n22578) );
  XNOR U40964 ( .A(q[11]), .B(DB[2305]), .Z(n39383) );
  XNOR U40965 ( .A(q[10]), .B(DB[2304]), .Z(n22576) );
  IV U40966 ( .A(n22591), .Z(n39376) );
  XOR U40967 ( .A(n39384), .B(n39385), .Z(n22591) );
  XNOR U40968 ( .A(n22608), .B(n22589), .Z(n39385) );
  XNOR U40969 ( .A(q[1]), .B(DB[2295]), .Z(n22589) );
  XOR U40970 ( .A(n39386), .B(n22597), .Z(n22608) );
  XNOR U40971 ( .A(q[8]), .B(DB[2302]), .Z(n22597) );
  IV U40972 ( .A(n22596), .Z(n39386) );
  XNOR U40973 ( .A(n22594), .B(n39387), .Z(n22596) );
  XNOR U40974 ( .A(q[7]), .B(DB[2301]), .Z(n39387) );
  XNOR U40975 ( .A(q[6]), .B(DB[2300]), .Z(n22594) );
  IV U40976 ( .A(n22607), .Z(n39384) );
  XOR U40977 ( .A(n39388), .B(n39389), .Z(n22607) );
  XNOR U40978 ( .A(n22603), .B(n22605), .Z(n39389) );
  XNOR U40979 ( .A(q[2]), .B(DB[2296]), .Z(n22605) );
  XNOR U40980 ( .A(q[5]), .B(DB[2299]), .Z(n22603) );
  IV U40981 ( .A(n22602), .Z(n39388) );
  XNOR U40982 ( .A(n22600), .B(n39390), .Z(n22602) );
  XNOR U40983 ( .A(q[4]), .B(DB[2298]), .Z(n39390) );
  XNOR U40984 ( .A(q[3]), .B(DB[2297]), .Z(n22600) );
  XOR U40985 ( .A(n39391), .B(n22369), .Z(n22220) );
  XOR U40986 ( .A(n39392), .B(n22345), .Z(n22369) );
  XOR U40987 ( .A(n39393), .B(n22337), .Z(n22345) );
  XOR U40988 ( .A(n39394), .B(n22326), .Z(n22337) );
  XNOR U40989 ( .A(q[30]), .B(DB[2355]), .Z(n22326) );
  IV U40990 ( .A(n22325), .Z(n39394) );
  XNOR U40991 ( .A(n22323), .B(n39395), .Z(n22325) );
  XNOR U40992 ( .A(q[29]), .B(DB[2354]), .Z(n39395) );
  XNOR U40993 ( .A(q[28]), .B(DB[2353]), .Z(n22323) );
  IV U40994 ( .A(n22336), .Z(n39393) );
  XOR U40995 ( .A(n39396), .B(n39397), .Z(n22336) );
  XNOR U40996 ( .A(n22332), .B(n22334), .Z(n39397) );
  XNOR U40997 ( .A(q[24]), .B(DB[2349]), .Z(n22334) );
  XNOR U40998 ( .A(q[27]), .B(DB[2352]), .Z(n22332) );
  IV U40999 ( .A(n22331), .Z(n39396) );
  XNOR U41000 ( .A(n22329), .B(n39398), .Z(n22331) );
  XNOR U41001 ( .A(q[26]), .B(DB[2351]), .Z(n39398) );
  XNOR U41002 ( .A(q[25]), .B(DB[2350]), .Z(n22329) );
  IV U41003 ( .A(n22344), .Z(n39392) );
  XOR U41004 ( .A(n39399), .B(n39400), .Z(n22344) );
  XNOR U41005 ( .A(n22361), .B(n22342), .Z(n39400) );
  XNOR U41006 ( .A(q[16]), .B(DB[2341]), .Z(n22342) );
  XOR U41007 ( .A(n39401), .B(n22350), .Z(n22361) );
  XNOR U41008 ( .A(q[23]), .B(DB[2348]), .Z(n22350) );
  IV U41009 ( .A(n22349), .Z(n39401) );
  XNOR U41010 ( .A(n22347), .B(n39402), .Z(n22349) );
  XNOR U41011 ( .A(q[22]), .B(DB[2347]), .Z(n39402) );
  XNOR U41012 ( .A(q[21]), .B(DB[2346]), .Z(n22347) );
  IV U41013 ( .A(n22360), .Z(n39399) );
  XOR U41014 ( .A(n39403), .B(n39404), .Z(n22360) );
  XNOR U41015 ( .A(n22356), .B(n22358), .Z(n39404) );
  XNOR U41016 ( .A(q[17]), .B(DB[2342]), .Z(n22358) );
  XNOR U41017 ( .A(q[20]), .B(DB[2345]), .Z(n22356) );
  IV U41018 ( .A(n22355), .Z(n39403) );
  XNOR U41019 ( .A(n22353), .B(n39405), .Z(n22355) );
  XNOR U41020 ( .A(q[19]), .B(DB[2344]), .Z(n39405) );
  XNOR U41021 ( .A(q[18]), .B(DB[2343]), .Z(n22353) );
  IV U41022 ( .A(n22368), .Z(n39391) );
  XOR U41023 ( .A(n39406), .B(n39407), .Z(n22368) );
  XNOR U41024 ( .A(n22395), .B(n22366), .Z(n39407) );
  XNOR U41025 ( .A(q[0]), .B(DB[2325]), .Z(n22366) );
  XOR U41026 ( .A(n39408), .B(n22387), .Z(n22395) );
  XOR U41027 ( .A(n39409), .B(n22375), .Z(n22387) );
  XNOR U41028 ( .A(q[15]), .B(DB[2340]), .Z(n22375) );
  IV U41029 ( .A(n22374), .Z(n39409) );
  XNOR U41030 ( .A(n22372), .B(n39410), .Z(n22374) );
  XNOR U41031 ( .A(q[14]), .B(DB[2339]), .Z(n39410) );
  XNOR U41032 ( .A(q[13]), .B(DB[2338]), .Z(n22372) );
  IV U41033 ( .A(n22386), .Z(n39408) );
  XOR U41034 ( .A(n39411), .B(n39412), .Z(n22386) );
  XNOR U41035 ( .A(n22382), .B(n22384), .Z(n39412) );
  XNOR U41036 ( .A(q[9]), .B(DB[2334]), .Z(n22384) );
  XNOR U41037 ( .A(q[12]), .B(DB[2337]), .Z(n22382) );
  IV U41038 ( .A(n22381), .Z(n39411) );
  XNOR U41039 ( .A(n22379), .B(n39413), .Z(n22381) );
  XNOR U41040 ( .A(q[11]), .B(DB[2336]), .Z(n39413) );
  XNOR U41041 ( .A(q[10]), .B(DB[2335]), .Z(n22379) );
  IV U41042 ( .A(n22394), .Z(n39406) );
  XOR U41043 ( .A(n39414), .B(n39415), .Z(n22394) );
  XNOR U41044 ( .A(n22411), .B(n22392), .Z(n39415) );
  XNOR U41045 ( .A(q[1]), .B(DB[2326]), .Z(n22392) );
  XOR U41046 ( .A(n39416), .B(n22400), .Z(n22411) );
  XNOR U41047 ( .A(q[8]), .B(DB[2333]), .Z(n22400) );
  IV U41048 ( .A(n22399), .Z(n39416) );
  XNOR U41049 ( .A(n22397), .B(n39417), .Z(n22399) );
  XNOR U41050 ( .A(q[7]), .B(DB[2332]), .Z(n39417) );
  XNOR U41051 ( .A(q[6]), .B(DB[2331]), .Z(n22397) );
  IV U41052 ( .A(n22410), .Z(n39414) );
  XOR U41053 ( .A(n39418), .B(n39419), .Z(n22410) );
  XNOR U41054 ( .A(n22406), .B(n22408), .Z(n39419) );
  XNOR U41055 ( .A(q[2]), .B(DB[2327]), .Z(n22408) );
  XNOR U41056 ( .A(q[5]), .B(DB[2330]), .Z(n22406) );
  IV U41057 ( .A(n22405), .Z(n39418) );
  XNOR U41058 ( .A(n22403), .B(n39420), .Z(n22405) );
  XNOR U41059 ( .A(q[4]), .B(DB[2329]), .Z(n39420) );
  XNOR U41060 ( .A(q[3]), .B(DB[2328]), .Z(n22403) );
  XOR U41061 ( .A(n39421), .B(n22172), .Z(n22023) );
  XOR U41062 ( .A(n39422), .B(n22148), .Z(n22172) );
  XOR U41063 ( .A(n39423), .B(n22140), .Z(n22148) );
  XOR U41064 ( .A(n39424), .B(n22129), .Z(n22140) );
  XNOR U41065 ( .A(q[30]), .B(DB[2386]), .Z(n22129) );
  IV U41066 ( .A(n22128), .Z(n39424) );
  XNOR U41067 ( .A(n22126), .B(n39425), .Z(n22128) );
  XNOR U41068 ( .A(q[29]), .B(DB[2385]), .Z(n39425) );
  XNOR U41069 ( .A(q[28]), .B(DB[2384]), .Z(n22126) );
  IV U41070 ( .A(n22139), .Z(n39423) );
  XOR U41071 ( .A(n39426), .B(n39427), .Z(n22139) );
  XNOR U41072 ( .A(n22135), .B(n22137), .Z(n39427) );
  XNOR U41073 ( .A(q[24]), .B(DB[2380]), .Z(n22137) );
  XNOR U41074 ( .A(q[27]), .B(DB[2383]), .Z(n22135) );
  IV U41075 ( .A(n22134), .Z(n39426) );
  XNOR U41076 ( .A(n22132), .B(n39428), .Z(n22134) );
  XNOR U41077 ( .A(q[26]), .B(DB[2382]), .Z(n39428) );
  XNOR U41078 ( .A(q[25]), .B(DB[2381]), .Z(n22132) );
  IV U41079 ( .A(n22147), .Z(n39422) );
  XOR U41080 ( .A(n39429), .B(n39430), .Z(n22147) );
  XNOR U41081 ( .A(n22164), .B(n22145), .Z(n39430) );
  XNOR U41082 ( .A(q[16]), .B(DB[2372]), .Z(n22145) );
  XOR U41083 ( .A(n39431), .B(n22153), .Z(n22164) );
  XNOR U41084 ( .A(q[23]), .B(DB[2379]), .Z(n22153) );
  IV U41085 ( .A(n22152), .Z(n39431) );
  XNOR U41086 ( .A(n22150), .B(n39432), .Z(n22152) );
  XNOR U41087 ( .A(q[22]), .B(DB[2378]), .Z(n39432) );
  XNOR U41088 ( .A(q[21]), .B(DB[2377]), .Z(n22150) );
  IV U41089 ( .A(n22163), .Z(n39429) );
  XOR U41090 ( .A(n39433), .B(n39434), .Z(n22163) );
  XNOR U41091 ( .A(n22159), .B(n22161), .Z(n39434) );
  XNOR U41092 ( .A(q[17]), .B(DB[2373]), .Z(n22161) );
  XNOR U41093 ( .A(q[20]), .B(DB[2376]), .Z(n22159) );
  IV U41094 ( .A(n22158), .Z(n39433) );
  XNOR U41095 ( .A(n22156), .B(n39435), .Z(n22158) );
  XNOR U41096 ( .A(q[19]), .B(DB[2375]), .Z(n39435) );
  XNOR U41097 ( .A(q[18]), .B(DB[2374]), .Z(n22156) );
  IV U41098 ( .A(n22171), .Z(n39421) );
  XOR U41099 ( .A(n39436), .B(n39437), .Z(n22171) );
  XNOR U41100 ( .A(n22198), .B(n22169), .Z(n39437) );
  XNOR U41101 ( .A(q[0]), .B(DB[2356]), .Z(n22169) );
  XOR U41102 ( .A(n39438), .B(n22190), .Z(n22198) );
  XOR U41103 ( .A(n39439), .B(n22178), .Z(n22190) );
  XNOR U41104 ( .A(q[15]), .B(DB[2371]), .Z(n22178) );
  IV U41105 ( .A(n22177), .Z(n39439) );
  XNOR U41106 ( .A(n22175), .B(n39440), .Z(n22177) );
  XNOR U41107 ( .A(q[14]), .B(DB[2370]), .Z(n39440) );
  XNOR U41108 ( .A(q[13]), .B(DB[2369]), .Z(n22175) );
  IV U41109 ( .A(n22189), .Z(n39438) );
  XOR U41110 ( .A(n39441), .B(n39442), .Z(n22189) );
  XNOR U41111 ( .A(n22185), .B(n22187), .Z(n39442) );
  XNOR U41112 ( .A(q[9]), .B(DB[2365]), .Z(n22187) );
  XNOR U41113 ( .A(q[12]), .B(DB[2368]), .Z(n22185) );
  IV U41114 ( .A(n22184), .Z(n39441) );
  XNOR U41115 ( .A(n22182), .B(n39443), .Z(n22184) );
  XNOR U41116 ( .A(q[11]), .B(DB[2367]), .Z(n39443) );
  XNOR U41117 ( .A(q[10]), .B(DB[2366]), .Z(n22182) );
  IV U41118 ( .A(n22197), .Z(n39436) );
  XOR U41119 ( .A(n39444), .B(n39445), .Z(n22197) );
  XNOR U41120 ( .A(n22214), .B(n22195), .Z(n39445) );
  XNOR U41121 ( .A(q[1]), .B(DB[2357]), .Z(n22195) );
  XOR U41122 ( .A(n39446), .B(n22203), .Z(n22214) );
  XNOR U41123 ( .A(q[8]), .B(DB[2364]), .Z(n22203) );
  IV U41124 ( .A(n22202), .Z(n39446) );
  XNOR U41125 ( .A(n22200), .B(n39447), .Z(n22202) );
  XNOR U41126 ( .A(q[7]), .B(DB[2363]), .Z(n39447) );
  XNOR U41127 ( .A(q[6]), .B(DB[2362]), .Z(n22200) );
  IV U41128 ( .A(n22213), .Z(n39444) );
  XOR U41129 ( .A(n39448), .B(n39449), .Z(n22213) );
  XNOR U41130 ( .A(n22209), .B(n22211), .Z(n39449) );
  XNOR U41131 ( .A(q[2]), .B(DB[2358]), .Z(n22211) );
  XNOR U41132 ( .A(q[5]), .B(DB[2361]), .Z(n22209) );
  IV U41133 ( .A(n22208), .Z(n39448) );
  XNOR U41134 ( .A(n22206), .B(n39450), .Z(n22208) );
  XNOR U41135 ( .A(q[4]), .B(DB[2360]), .Z(n39450) );
  XNOR U41136 ( .A(q[3]), .B(DB[2359]), .Z(n22206) );
  XOR U41137 ( .A(n39451), .B(n21975), .Z(n21826) );
  XOR U41138 ( .A(n39452), .B(n21951), .Z(n21975) );
  XOR U41139 ( .A(n39453), .B(n21943), .Z(n21951) );
  XOR U41140 ( .A(n39454), .B(n21932), .Z(n21943) );
  XNOR U41141 ( .A(q[30]), .B(DB[2417]), .Z(n21932) );
  IV U41142 ( .A(n21931), .Z(n39454) );
  XNOR U41143 ( .A(n21929), .B(n39455), .Z(n21931) );
  XNOR U41144 ( .A(q[29]), .B(DB[2416]), .Z(n39455) );
  XNOR U41145 ( .A(q[28]), .B(DB[2415]), .Z(n21929) );
  IV U41146 ( .A(n21942), .Z(n39453) );
  XOR U41147 ( .A(n39456), .B(n39457), .Z(n21942) );
  XNOR U41148 ( .A(n21938), .B(n21940), .Z(n39457) );
  XNOR U41149 ( .A(q[24]), .B(DB[2411]), .Z(n21940) );
  XNOR U41150 ( .A(q[27]), .B(DB[2414]), .Z(n21938) );
  IV U41151 ( .A(n21937), .Z(n39456) );
  XNOR U41152 ( .A(n21935), .B(n39458), .Z(n21937) );
  XNOR U41153 ( .A(q[26]), .B(DB[2413]), .Z(n39458) );
  XNOR U41154 ( .A(q[25]), .B(DB[2412]), .Z(n21935) );
  IV U41155 ( .A(n21950), .Z(n39452) );
  XOR U41156 ( .A(n39459), .B(n39460), .Z(n21950) );
  XNOR U41157 ( .A(n21967), .B(n21948), .Z(n39460) );
  XNOR U41158 ( .A(q[16]), .B(DB[2403]), .Z(n21948) );
  XOR U41159 ( .A(n39461), .B(n21956), .Z(n21967) );
  XNOR U41160 ( .A(q[23]), .B(DB[2410]), .Z(n21956) );
  IV U41161 ( .A(n21955), .Z(n39461) );
  XNOR U41162 ( .A(n21953), .B(n39462), .Z(n21955) );
  XNOR U41163 ( .A(q[22]), .B(DB[2409]), .Z(n39462) );
  XNOR U41164 ( .A(q[21]), .B(DB[2408]), .Z(n21953) );
  IV U41165 ( .A(n21966), .Z(n39459) );
  XOR U41166 ( .A(n39463), .B(n39464), .Z(n21966) );
  XNOR U41167 ( .A(n21962), .B(n21964), .Z(n39464) );
  XNOR U41168 ( .A(q[17]), .B(DB[2404]), .Z(n21964) );
  XNOR U41169 ( .A(q[20]), .B(DB[2407]), .Z(n21962) );
  IV U41170 ( .A(n21961), .Z(n39463) );
  XNOR U41171 ( .A(n21959), .B(n39465), .Z(n21961) );
  XNOR U41172 ( .A(q[19]), .B(DB[2406]), .Z(n39465) );
  XNOR U41173 ( .A(q[18]), .B(DB[2405]), .Z(n21959) );
  IV U41174 ( .A(n21974), .Z(n39451) );
  XOR U41175 ( .A(n39466), .B(n39467), .Z(n21974) );
  XNOR U41176 ( .A(n22001), .B(n21972), .Z(n39467) );
  XNOR U41177 ( .A(q[0]), .B(DB[2387]), .Z(n21972) );
  XOR U41178 ( .A(n39468), .B(n21993), .Z(n22001) );
  XOR U41179 ( .A(n39469), .B(n21981), .Z(n21993) );
  XNOR U41180 ( .A(q[15]), .B(DB[2402]), .Z(n21981) );
  IV U41181 ( .A(n21980), .Z(n39469) );
  XNOR U41182 ( .A(n21978), .B(n39470), .Z(n21980) );
  XNOR U41183 ( .A(q[14]), .B(DB[2401]), .Z(n39470) );
  XNOR U41184 ( .A(q[13]), .B(DB[2400]), .Z(n21978) );
  IV U41185 ( .A(n21992), .Z(n39468) );
  XOR U41186 ( .A(n39471), .B(n39472), .Z(n21992) );
  XNOR U41187 ( .A(n21988), .B(n21990), .Z(n39472) );
  XNOR U41188 ( .A(q[9]), .B(DB[2396]), .Z(n21990) );
  XNOR U41189 ( .A(q[12]), .B(DB[2399]), .Z(n21988) );
  IV U41190 ( .A(n21987), .Z(n39471) );
  XNOR U41191 ( .A(n21985), .B(n39473), .Z(n21987) );
  XNOR U41192 ( .A(q[11]), .B(DB[2398]), .Z(n39473) );
  XNOR U41193 ( .A(q[10]), .B(DB[2397]), .Z(n21985) );
  IV U41194 ( .A(n22000), .Z(n39466) );
  XOR U41195 ( .A(n39474), .B(n39475), .Z(n22000) );
  XNOR U41196 ( .A(n22017), .B(n21998), .Z(n39475) );
  XNOR U41197 ( .A(q[1]), .B(DB[2388]), .Z(n21998) );
  XOR U41198 ( .A(n39476), .B(n22006), .Z(n22017) );
  XNOR U41199 ( .A(q[8]), .B(DB[2395]), .Z(n22006) );
  IV U41200 ( .A(n22005), .Z(n39476) );
  XNOR U41201 ( .A(n22003), .B(n39477), .Z(n22005) );
  XNOR U41202 ( .A(q[7]), .B(DB[2394]), .Z(n39477) );
  XNOR U41203 ( .A(q[6]), .B(DB[2393]), .Z(n22003) );
  IV U41204 ( .A(n22016), .Z(n39474) );
  XOR U41205 ( .A(n39478), .B(n39479), .Z(n22016) );
  XNOR U41206 ( .A(n22012), .B(n22014), .Z(n39479) );
  XNOR U41207 ( .A(q[2]), .B(DB[2389]), .Z(n22014) );
  XNOR U41208 ( .A(q[5]), .B(DB[2392]), .Z(n22012) );
  IV U41209 ( .A(n22011), .Z(n39478) );
  XNOR U41210 ( .A(n22009), .B(n39480), .Z(n22011) );
  XNOR U41211 ( .A(q[4]), .B(DB[2391]), .Z(n39480) );
  XNOR U41212 ( .A(q[3]), .B(DB[2390]), .Z(n22009) );
  XOR U41213 ( .A(n39481), .B(n21778), .Z(n21629) );
  XOR U41214 ( .A(n39482), .B(n21754), .Z(n21778) );
  XOR U41215 ( .A(n39483), .B(n21746), .Z(n21754) );
  XOR U41216 ( .A(n39484), .B(n21735), .Z(n21746) );
  XNOR U41217 ( .A(q[30]), .B(DB[2448]), .Z(n21735) );
  IV U41218 ( .A(n21734), .Z(n39484) );
  XNOR U41219 ( .A(n21732), .B(n39485), .Z(n21734) );
  XNOR U41220 ( .A(q[29]), .B(DB[2447]), .Z(n39485) );
  XNOR U41221 ( .A(q[28]), .B(DB[2446]), .Z(n21732) );
  IV U41222 ( .A(n21745), .Z(n39483) );
  XOR U41223 ( .A(n39486), .B(n39487), .Z(n21745) );
  XNOR U41224 ( .A(n21741), .B(n21743), .Z(n39487) );
  XNOR U41225 ( .A(q[24]), .B(DB[2442]), .Z(n21743) );
  XNOR U41226 ( .A(q[27]), .B(DB[2445]), .Z(n21741) );
  IV U41227 ( .A(n21740), .Z(n39486) );
  XNOR U41228 ( .A(n21738), .B(n39488), .Z(n21740) );
  XNOR U41229 ( .A(q[26]), .B(DB[2444]), .Z(n39488) );
  XNOR U41230 ( .A(q[25]), .B(DB[2443]), .Z(n21738) );
  IV U41231 ( .A(n21753), .Z(n39482) );
  XOR U41232 ( .A(n39489), .B(n39490), .Z(n21753) );
  XNOR U41233 ( .A(n21770), .B(n21751), .Z(n39490) );
  XNOR U41234 ( .A(q[16]), .B(DB[2434]), .Z(n21751) );
  XOR U41235 ( .A(n39491), .B(n21759), .Z(n21770) );
  XNOR U41236 ( .A(q[23]), .B(DB[2441]), .Z(n21759) );
  IV U41237 ( .A(n21758), .Z(n39491) );
  XNOR U41238 ( .A(n21756), .B(n39492), .Z(n21758) );
  XNOR U41239 ( .A(q[22]), .B(DB[2440]), .Z(n39492) );
  XNOR U41240 ( .A(q[21]), .B(DB[2439]), .Z(n21756) );
  IV U41241 ( .A(n21769), .Z(n39489) );
  XOR U41242 ( .A(n39493), .B(n39494), .Z(n21769) );
  XNOR U41243 ( .A(n21765), .B(n21767), .Z(n39494) );
  XNOR U41244 ( .A(q[17]), .B(DB[2435]), .Z(n21767) );
  XNOR U41245 ( .A(q[20]), .B(DB[2438]), .Z(n21765) );
  IV U41246 ( .A(n21764), .Z(n39493) );
  XNOR U41247 ( .A(n21762), .B(n39495), .Z(n21764) );
  XNOR U41248 ( .A(q[19]), .B(DB[2437]), .Z(n39495) );
  XNOR U41249 ( .A(q[18]), .B(DB[2436]), .Z(n21762) );
  IV U41250 ( .A(n21777), .Z(n39481) );
  XOR U41251 ( .A(n39496), .B(n39497), .Z(n21777) );
  XNOR U41252 ( .A(n21804), .B(n21775), .Z(n39497) );
  XNOR U41253 ( .A(q[0]), .B(DB[2418]), .Z(n21775) );
  XOR U41254 ( .A(n39498), .B(n21796), .Z(n21804) );
  XOR U41255 ( .A(n39499), .B(n21784), .Z(n21796) );
  XNOR U41256 ( .A(q[15]), .B(DB[2433]), .Z(n21784) );
  IV U41257 ( .A(n21783), .Z(n39499) );
  XNOR U41258 ( .A(n21781), .B(n39500), .Z(n21783) );
  XNOR U41259 ( .A(q[14]), .B(DB[2432]), .Z(n39500) );
  XNOR U41260 ( .A(q[13]), .B(DB[2431]), .Z(n21781) );
  IV U41261 ( .A(n21795), .Z(n39498) );
  XOR U41262 ( .A(n39501), .B(n39502), .Z(n21795) );
  XNOR U41263 ( .A(n21791), .B(n21793), .Z(n39502) );
  XNOR U41264 ( .A(q[9]), .B(DB[2427]), .Z(n21793) );
  XNOR U41265 ( .A(q[12]), .B(DB[2430]), .Z(n21791) );
  IV U41266 ( .A(n21790), .Z(n39501) );
  XNOR U41267 ( .A(n21788), .B(n39503), .Z(n21790) );
  XNOR U41268 ( .A(q[11]), .B(DB[2429]), .Z(n39503) );
  XNOR U41269 ( .A(q[10]), .B(DB[2428]), .Z(n21788) );
  IV U41270 ( .A(n21803), .Z(n39496) );
  XOR U41271 ( .A(n39504), .B(n39505), .Z(n21803) );
  XNOR U41272 ( .A(n21820), .B(n21801), .Z(n39505) );
  XNOR U41273 ( .A(q[1]), .B(DB[2419]), .Z(n21801) );
  XOR U41274 ( .A(n39506), .B(n21809), .Z(n21820) );
  XNOR U41275 ( .A(q[8]), .B(DB[2426]), .Z(n21809) );
  IV U41276 ( .A(n21808), .Z(n39506) );
  XNOR U41277 ( .A(n21806), .B(n39507), .Z(n21808) );
  XNOR U41278 ( .A(q[7]), .B(DB[2425]), .Z(n39507) );
  XNOR U41279 ( .A(q[6]), .B(DB[2424]), .Z(n21806) );
  IV U41280 ( .A(n21819), .Z(n39504) );
  XOR U41281 ( .A(n39508), .B(n39509), .Z(n21819) );
  XNOR U41282 ( .A(n21815), .B(n21817), .Z(n39509) );
  XNOR U41283 ( .A(q[2]), .B(DB[2420]), .Z(n21817) );
  XNOR U41284 ( .A(q[5]), .B(DB[2423]), .Z(n21815) );
  IV U41285 ( .A(n21814), .Z(n39508) );
  XNOR U41286 ( .A(n21812), .B(n39510), .Z(n21814) );
  XNOR U41287 ( .A(q[4]), .B(DB[2422]), .Z(n39510) );
  XNOR U41288 ( .A(q[3]), .B(DB[2421]), .Z(n21812) );
  XOR U41289 ( .A(n39511), .B(n21581), .Z(n21432) );
  XOR U41290 ( .A(n39512), .B(n21557), .Z(n21581) );
  XOR U41291 ( .A(n39513), .B(n21549), .Z(n21557) );
  XOR U41292 ( .A(n39514), .B(n21538), .Z(n21549) );
  XNOR U41293 ( .A(q[30]), .B(DB[2479]), .Z(n21538) );
  IV U41294 ( .A(n21537), .Z(n39514) );
  XNOR U41295 ( .A(n21535), .B(n39515), .Z(n21537) );
  XNOR U41296 ( .A(q[29]), .B(DB[2478]), .Z(n39515) );
  XNOR U41297 ( .A(q[28]), .B(DB[2477]), .Z(n21535) );
  IV U41298 ( .A(n21548), .Z(n39513) );
  XOR U41299 ( .A(n39516), .B(n39517), .Z(n21548) );
  XNOR U41300 ( .A(n21544), .B(n21546), .Z(n39517) );
  XNOR U41301 ( .A(q[24]), .B(DB[2473]), .Z(n21546) );
  XNOR U41302 ( .A(q[27]), .B(DB[2476]), .Z(n21544) );
  IV U41303 ( .A(n21543), .Z(n39516) );
  XNOR U41304 ( .A(n21541), .B(n39518), .Z(n21543) );
  XNOR U41305 ( .A(q[26]), .B(DB[2475]), .Z(n39518) );
  XNOR U41306 ( .A(q[25]), .B(DB[2474]), .Z(n21541) );
  IV U41307 ( .A(n21556), .Z(n39512) );
  XOR U41308 ( .A(n39519), .B(n39520), .Z(n21556) );
  XNOR U41309 ( .A(n21573), .B(n21554), .Z(n39520) );
  XNOR U41310 ( .A(q[16]), .B(DB[2465]), .Z(n21554) );
  XOR U41311 ( .A(n39521), .B(n21562), .Z(n21573) );
  XNOR U41312 ( .A(q[23]), .B(DB[2472]), .Z(n21562) );
  IV U41313 ( .A(n21561), .Z(n39521) );
  XNOR U41314 ( .A(n21559), .B(n39522), .Z(n21561) );
  XNOR U41315 ( .A(q[22]), .B(DB[2471]), .Z(n39522) );
  XNOR U41316 ( .A(q[21]), .B(DB[2470]), .Z(n21559) );
  IV U41317 ( .A(n21572), .Z(n39519) );
  XOR U41318 ( .A(n39523), .B(n39524), .Z(n21572) );
  XNOR U41319 ( .A(n21568), .B(n21570), .Z(n39524) );
  XNOR U41320 ( .A(q[17]), .B(DB[2466]), .Z(n21570) );
  XNOR U41321 ( .A(q[20]), .B(DB[2469]), .Z(n21568) );
  IV U41322 ( .A(n21567), .Z(n39523) );
  XNOR U41323 ( .A(n21565), .B(n39525), .Z(n21567) );
  XNOR U41324 ( .A(q[19]), .B(DB[2468]), .Z(n39525) );
  XNOR U41325 ( .A(q[18]), .B(DB[2467]), .Z(n21565) );
  IV U41326 ( .A(n21580), .Z(n39511) );
  XOR U41327 ( .A(n39526), .B(n39527), .Z(n21580) );
  XNOR U41328 ( .A(n21607), .B(n21578), .Z(n39527) );
  XNOR U41329 ( .A(q[0]), .B(DB[2449]), .Z(n21578) );
  XOR U41330 ( .A(n39528), .B(n21599), .Z(n21607) );
  XOR U41331 ( .A(n39529), .B(n21587), .Z(n21599) );
  XNOR U41332 ( .A(q[15]), .B(DB[2464]), .Z(n21587) );
  IV U41333 ( .A(n21586), .Z(n39529) );
  XNOR U41334 ( .A(n21584), .B(n39530), .Z(n21586) );
  XNOR U41335 ( .A(q[14]), .B(DB[2463]), .Z(n39530) );
  XNOR U41336 ( .A(q[13]), .B(DB[2462]), .Z(n21584) );
  IV U41337 ( .A(n21598), .Z(n39528) );
  XOR U41338 ( .A(n39531), .B(n39532), .Z(n21598) );
  XNOR U41339 ( .A(n21594), .B(n21596), .Z(n39532) );
  XNOR U41340 ( .A(q[9]), .B(DB[2458]), .Z(n21596) );
  XNOR U41341 ( .A(q[12]), .B(DB[2461]), .Z(n21594) );
  IV U41342 ( .A(n21593), .Z(n39531) );
  XNOR U41343 ( .A(n21591), .B(n39533), .Z(n21593) );
  XNOR U41344 ( .A(q[11]), .B(DB[2460]), .Z(n39533) );
  XNOR U41345 ( .A(q[10]), .B(DB[2459]), .Z(n21591) );
  IV U41346 ( .A(n21606), .Z(n39526) );
  XOR U41347 ( .A(n39534), .B(n39535), .Z(n21606) );
  XNOR U41348 ( .A(n21623), .B(n21604), .Z(n39535) );
  XNOR U41349 ( .A(q[1]), .B(DB[2450]), .Z(n21604) );
  XOR U41350 ( .A(n39536), .B(n21612), .Z(n21623) );
  XNOR U41351 ( .A(q[8]), .B(DB[2457]), .Z(n21612) );
  IV U41352 ( .A(n21611), .Z(n39536) );
  XNOR U41353 ( .A(n21609), .B(n39537), .Z(n21611) );
  XNOR U41354 ( .A(q[7]), .B(DB[2456]), .Z(n39537) );
  XNOR U41355 ( .A(q[6]), .B(DB[2455]), .Z(n21609) );
  IV U41356 ( .A(n21622), .Z(n39534) );
  XOR U41357 ( .A(n39538), .B(n39539), .Z(n21622) );
  XNOR U41358 ( .A(n21618), .B(n21620), .Z(n39539) );
  XNOR U41359 ( .A(q[2]), .B(DB[2451]), .Z(n21620) );
  XNOR U41360 ( .A(q[5]), .B(DB[2454]), .Z(n21618) );
  IV U41361 ( .A(n21617), .Z(n39538) );
  XNOR U41362 ( .A(n21615), .B(n39540), .Z(n21617) );
  XNOR U41363 ( .A(q[4]), .B(DB[2453]), .Z(n39540) );
  XNOR U41364 ( .A(q[3]), .B(DB[2452]), .Z(n21615) );
  XOR U41365 ( .A(n39541), .B(n21384), .Z(n21235) );
  XOR U41366 ( .A(n39542), .B(n21360), .Z(n21384) );
  XOR U41367 ( .A(n39543), .B(n21352), .Z(n21360) );
  XOR U41368 ( .A(n39544), .B(n21341), .Z(n21352) );
  XNOR U41369 ( .A(q[30]), .B(DB[2510]), .Z(n21341) );
  IV U41370 ( .A(n21340), .Z(n39544) );
  XNOR U41371 ( .A(n21338), .B(n39545), .Z(n21340) );
  XNOR U41372 ( .A(q[29]), .B(DB[2509]), .Z(n39545) );
  XNOR U41373 ( .A(q[28]), .B(DB[2508]), .Z(n21338) );
  IV U41374 ( .A(n21351), .Z(n39543) );
  XOR U41375 ( .A(n39546), .B(n39547), .Z(n21351) );
  XNOR U41376 ( .A(n21347), .B(n21349), .Z(n39547) );
  XNOR U41377 ( .A(q[24]), .B(DB[2504]), .Z(n21349) );
  XNOR U41378 ( .A(q[27]), .B(DB[2507]), .Z(n21347) );
  IV U41379 ( .A(n21346), .Z(n39546) );
  XNOR U41380 ( .A(n21344), .B(n39548), .Z(n21346) );
  XNOR U41381 ( .A(q[26]), .B(DB[2506]), .Z(n39548) );
  XNOR U41382 ( .A(q[25]), .B(DB[2505]), .Z(n21344) );
  IV U41383 ( .A(n21359), .Z(n39542) );
  XOR U41384 ( .A(n39549), .B(n39550), .Z(n21359) );
  XNOR U41385 ( .A(n21376), .B(n21357), .Z(n39550) );
  XNOR U41386 ( .A(q[16]), .B(DB[2496]), .Z(n21357) );
  XOR U41387 ( .A(n39551), .B(n21365), .Z(n21376) );
  XNOR U41388 ( .A(q[23]), .B(DB[2503]), .Z(n21365) );
  IV U41389 ( .A(n21364), .Z(n39551) );
  XNOR U41390 ( .A(n21362), .B(n39552), .Z(n21364) );
  XNOR U41391 ( .A(q[22]), .B(DB[2502]), .Z(n39552) );
  XNOR U41392 ( .A(q[21]), .B(DB[2501]), .Z(n21362) );
  IV U41393 ( .A(n21375), .Z(n39549) );
  XOR U41394 ( .A(n39553), .B(n39554), .Z(n21375) );
  XNOR U41395 ( .A(n21371), .B(n21373), .Z(n39554) );
  XNOR U41396 ( .A(q[17]), .B(DB[2497]), .Z(n21373) );
  XNOR U41397 ( .A(q[20]), .B(DB[2500]), .Z(n21371) );
  IV U41398 ( .A(n21370), .Z(n39553) );
  XNOR U41399 ( .A(n21368), .B(n39555), .Z(n21370) );
  XNOR U41400 ( .A(q[19]), .B(DB[2499]), .Z(n39555) );
  XNOR U41401 ( .A(q[18]), .B(DB[2498]), .Z(n21368) );
  IV U41402 ( .A(n21383), .Z(n39541) );
  XOR U41403 ( .A(n39556), .B(n39557), .Z(n21383) );
  XNOR U41404 ( .A(n21410), .B(n21381), .Z(n39557) );
  XNOR U41405 ( .A(q[0]), .B(DB[2480]), .Z(n21381) );
  XOR U41406 ( .A(n39558), .B(n21402), .Z(n21410) );
  XOR U41407 ( .A(n39559), .B(n21390), .Z(n21402) );
  XNOR U41408 ( .A(q[15]), .B(DB[2495]), .Z(n21390) );
  IV U41409 ( .A(n21389), .Z(n39559) );
  XNOR U41410 ( .A(n21387), .B(n39560), .Z(n21389) );
  XNOR U41411 ( .A(q[14]), .B(DB[2494]), .Z(n39560) );
  XNOR U41412 ( .A(q[13]), .B(DB[2493]), .Z(n21387) );
  IV U41413 ( .A(n21401), .Z(n39558) );
  XOR U41414 ( .A(n39561), .B(n39562), .Z(n21401) );
  XNOR U41415 ( .A(n21397), .B(n21399), .Z(n39562) );
  XNOR U41416 ( .A(q[9]), .B(DB[2489]), .Z(n21399) );
  XNOR U41417 ( .A(q[12]), .B(DB[2492]), .Z(n21397) );
  IV U41418 ( .A(n21396), .Z(n39561) );
  XNOR U41419 ( .A(n21394), .B(n39563), .Z(n21396) );
  XNOR U41420 ( .A(q[11]), .B(DB[2491]), .Z(n39563) );
  XNOR U41421 ( .A(q[10]), .B(DB[2490]), .Z(n21394) );
  IV U41422 ( .A(n21409), .Z(n39556) );
  XOR U41423 ( .A(n39564), .B(n39565), .Z(n21409) );
  XNOR U41424 ( .A(n21426), .B(n21407), .Z(n39565) );
  XNOR U41425 ( .A(q[1]), .B(DB[2481]), .Z(n21407) );
  XOR U41426 ( .A(n39566), .B(n21415), .Z(n21426) );
  XNOR U41427 ( .A(q[8]), .B(DB[2488]), .Z(n21415) );
  IV U41428 ( .A(n21414), .Z(n39566) );
  XNOR U41429 ( .A(n21412), .B(n39567), .Z(n21414) );
  XNOR U41430 ( .A(q[7]), .B(DB[2487]), .Z(n39567) );
  XNOR U41431 ( .A(q[6]), .B(DB[2486]), .Z(n21412) );
  IV U41432 ( .A(n21425), .Z(n39564) );
  XOR U41433 ( .A(n39568), .B(n39569), .Z(n21425) );
  XNOR U41434 ( .A(n21421), .B(n21423), .Z(n39569) );
  XNOR U41435 ( .A(q[2]), .B(DB[2482]), .Z(n21423) );
  XNOR U41436 ( .A(q[5]), .B(DB[2485]), .Z(n21421) );
  IV U41437 ( .A(n21420), .Z(n39568) );
  XNOR U41438 ( .A(n21418), .B(n39570), .Z(n21420) );
  XNOR U41439 ( .A(q[4]), .B(DB[2484]), .Z(n39570) );
  XNOR U41440 ( .A(q[3]), .B(DB[2483]), .Z(n21418) );
  XOR U41441 ( .A(n39571), .B(n21187), .Z(n21038) );
  XOR U41442 ( .A(n39572), .B(n21163), .Z(n21187) );
  XOR U41443 ( .A(n39573), .B(n21155), .Z(n21163) );
  XOR U41444 ( .A(n39574), .B(n21144), .Z(n21155) );
  XNOR U41445 ( .A(q[30]), .B(DB[2541]), .Z(n21144) );
  IV U41446 ( .A(n21143), .Z(n39574) );
  XNOR U41447 ( .A(n21141), .B(n39575), .Z(n21143) );
  XNOR U41448 ( .A(q[29]), .B(DB[2540]), .Z(n39575) );
  XNOR U41449 ( .A(q[28]), .B(DB[2539]), .Z(n21141) );
  IV U41450 ( .A(n21154), .Z(n39573) );
  XOR U41451 ( .A(n39576), .B(n39577), .Z(n21154) );
  XNOR U41452 ( .A(n21150), .B(n21152), .Z(n39577) );
  XNOR U41453 ( .A(q[24]), .B(DB[2535]), .Z(n21152) );
  XNOR U41454 ( .A(q[27]), .B(DB[2538]), .Z(n21150) );
  IV U41455 ( .A(n21149), .Z(n39576) );
  XNOR U41456 ( .A(n21147), .B(n39578), .Z(n21149) );
  XNOR U41457 ( .A(q[26]), .B(DB[2537]), .Z(n39578) );
  XNOR U41458 ( .A(q[25]), .B(DB[2536]), .Z(n21147) );
  IV U41459 ( .A(n21162), .Z(n39572) );
  XOR U41460 ( .A(n39579), .B(n39580), .Z(n21162) );
  XNOR U41461 ( .A(n21179), .B(n21160), .Z(n39580) );
  XNOR U41462 ( .A(q[16]), .B(DB[2527]), .Z(n21160) );
  XOR U41463 ( .A(n39581), .B(n21168), .Z(n21179) );
  XNOR U41464 ( .A(q[23]), .B(DB[2534]), .Z(n21168) );
  IV U41465 ( .A(n21167), .Z(n39581) );
  XNOR U41466 ( .A(n21165), .B(n39582), .Z(n21167) );
  XNOR U41467 ( .A(q[22]), .B(DB[2533]), .Z(n39582) );
  XNOR U41468 ( .A(q[21]), .B(DB[2532]), .Z(n21165) );
  IV U41469 ( .A(n21178), .Z(n39579) );
  XOR U41470 ( .A(n39583), .B(n39584), .Z(n21178) );
  XNOR U41471 ( .A(n21174), .B(n21176), .Z(n39584) );
  XNOR U41472 ( .A(q[17]), .B(DB[2528]), .Z(n21176) );
  XNOR U41473 ( .A(q[20]), .B(DB[2531]), .Z(n21174) );
  IV U41474 ( .A(n21173), .Z(n39583) );
  XNOR U41475 ( .A(n21171), .B(n39585), .Z(n21173) );
  XNOR U41476 ( .A(q[19]), .B(DB[2530]), .Z(n39585) );
  XNOR U41477 ( .A(q[18]), .B(DB[2529]), .Z(n21171) );
  IV U41478 ( .A(n21186), .Z(n39571) );
  XOR U41479 ( .A(n39586), .B(n39587), .Z(n21186) );
  XNOR U41480 ( .A(n21213), .B(n21184), .Z(n39587) );
  XNOR U41481 ( .A(q[0]), .B(DB[2511]), .Z(n21184) );
  XOR U41482 ( .A(n39588), .B(n21205), .Z(n21213) );
  XOR U41483 ( .A(n39589), .B(n21193), .Z(n21205) );
  XNOR U41484 ( .A(q[15]), .B(DB[2526]), .Z(n21193) );
  IV U41485 ( .A(n21192), .Z(n39589) );
  XNOR U41486 ( .A(n21190), .B(n39590), .Z(n21192) );
  XNOR U41487 ( .A(q[14]), .B(DB[2525]), .Z(n39590) );
  XNOR U41488 ( .A(q[13]), .B(DB[2524]), .Z(n21190) );
  IV U41489 ( .A(n21204), .Z(n39588) );
  XOR U41490 ( .A(n39591), .B(n39592), .Z(n21204) );
  XNOR U41491 ( .A(n21200), .B(n21202), .Z(n39592) );
  XNOR U41492 ( .A(q[9]), .B(DB[2520]), .Z(n21202) );
  XNOR U41493 ( .A(q[12]), .B(DB[2523]), .Z(n21200) );
  IV U41494 ( .A(n21199), .Z(n39591) );
  XNOR U41495 ( .A(n21197), .B(n39593), .Z(n21199) );
  XNOR U41496 ( .A(q[11]), .B(DB[2522]), .Z(n39593) );
  XNOR U41497 ( .A(q[10]), .B(DB[2521]), .Z(n21197) );
  IV U41498 ( .A(n21212), .Z(n39586) );
  XOR U41499 ( .A(n39594), .B(n39595), .Z(n21212) );
  XNOR U41500 ( .A(n21229), .B(n21210), .Z(n39595) );
  XNOR U41501 ( .A(q[1]), .B(DB[2512]), .Z(n21210) );
  XOR U41502 ( .A(n39596), .B(n21218), .Z(n21229) );
  XNOR U41503 ( .A(q[8]), .B(DB[2519]), .Z(n21218) );
  IV U41504 ( .A(n21217), .Z(n39596) );
  XNOR U41505 ( .A(n21215), .B(n39597), .Z(n21217) );
  XNOR U41506 ( .A(q[7]), .B(DB[2518]), .Z(n39597) );
  XNOR U41507 ( .A(q[6]), .B(DB[2517]), .Z(n21215) );
  IV U41508 ( .A(n21228), .Z(n39594) );
  XOR U41509 ( .A(n39598), .B(n39599), .Z(n21228) );
  XNOR U41510 ( .A(n21224), .B(n21226), .Z(n39599) );
  XNOR U41511 ( .A(q[2]), .B(DB[2513]), .Z(n21226) );
  XNOR U41512 ( .A(q[5]), .B(DB[2516]), .Z(n21224) );
  IV U41513 ( .A(n21223), .Z(n39598) );
  XNOR U41514 ( .A(n21221), .B(n39600), .Z(n21223) );
  XNOR U41515 ( .A(q[4]), .B(DB[2515]), .Z(n39600) );
  XNOR U41516 ( .A(q[3]), .B(DB[2514]), .Z(n21221) );
  XOR U41517 ( .A(n39601), .B(n20990), .Z(n20841) );
  XOR U41518 ( .A(n39602), .B(n20966), .Z(n20990) );
  XOR U41519 ( .A(n39603), .B(n20958), .Z(n20966) );
  XOR U41520 ( .A(n39604), .B(n20947), .Z(n20958) );
  XNOR U41521 ( .A(q[30]), .B(DB[2572]), .Z(n20947) );
  IV U41522 ( .A(n20946), .Z(n39604) );
  XNOR U41523 ( .A(n20944), .B(n39605), .Z(n20946) );
  XNOR U41524 ( .A(q[29]), .B(DB[2571]), .Z(n39605) );
  XNOR U41525 ( .A(q[28]), .B(DB[2570]), .Z(n20944) );
  IV U41526 ( .A(n20957), .Z(n39603) );
  XOR U41527 ( .A(n39606), .B(n39607), .Z(n20957) );
  XNOR U41528 ( .A(n20953), .B(n20955), .Z(n39607) );
  XNOR U41529 ( .A(q[24]), .B(DB[2566]), .Z(n20955) );
  XNOR U41530 ( .A(q[27]), .B(DB[2569]), .Z(n20953) );
  IV U41531 ( .A(n20952), .Z(n39606) );
  XNOR U41532 ( .A(n20950), .B(n39608), .Z(n20952) );
  XNOR U41533 ( .A(q[26]), .B(DB[2568]), .Z(n39608) );
  XNOR U41534 ( .A(q[25]), .B(DB[2567]), .Z(n20950) );
  IV U41535 ( .A(n20965), .Z(n39602) );
  XOR U41536 ( .A(n39609), .B(n39610), .Z(n20965) );
  XNOR U41537 ( .A(n20982), .B(n20963), .Z(n39610) );
  XNOR U41538 ( .A(q[16]), .B(DB[2558]), .Z(n20963) );
  XOR U41539 ( .A(n39611), .B(n20971), .Z(n20982) );
  XNOR U41540 ( .A(q[23]), .B(DB[2565]), .Z(n20971) );
  IV U41541 ( .A(n20970), .Z(n39611) );
  XNOR U41542 ( .A(n20968), .B(n39612), .Z(n20970) );
  XNOR U41543 ( .A(q[22]), .B(DB[2564]), .Z(n39612) );
  XNOR U41544 ( .A(q[21]), .B(DB[2563]), .Z(n20968) );
  IV U41545 ( .A(n20981), .Z(n39609) );
  XOR U41546 ( .A(n39613), .B(n39614), .Z(n20981) );
  XNOR U41547 ( .A(n20977), .B(n20979), .Z(n39614) );
  XNOR U41548 ( .A(q[17]), .B(DB[2559]), .Z(n20979) );
  XNOR U41549 ( .A(q[20]), .B(DB[2562]), .Z(n20977) );
  IV U41550 ( .A(n20976), .Z(n39613) );
  XNOR U41551 ( .A(n20974), .B(n39615), .Z(n20976) );
  XNOR U41552 ( .A(q[19]), .B(DB[2561]), .Z(n39615) );
  XNOR U41553 ( .A(q[18]), .B(DB[2560]), .Z(n20974) );
  IV U41554 ( .A(n20989), .Z(n39601) );
  XOR U41555 ( .A(n39616), .B(n39617), .Z(n20989) );
  XNOR U41556 ( .A(n21016), .B(n20987), .Z(n39617) );
  XNOR U41557 ( .A(q[0]), .B(DB[2542]), .Z(n20987) );
  XOR U41558 ( .A(n39618), .B(n21008), .Z(n21016) );
  XOR U41559 ( .A(n39619), .B(n20996), .Z(n21008) );
  XNOR U41560 ( .A(q[15]), .B(DB[2557]), .Z(n20996) );
  IV U41561 ( .A(n20995), .Z(n39619) );
  XNOR U41562 ( .A(n20993), .B(n39620), .Z(n20995) );
  XNOR U41563 ( .A(q[14]), .B(DB[2556]), .Z(n39620) );
  XNOR U41564 ( .A(q[13]), .B(DB[2555]), .Z(n20993) );
  IV U41565 ( .A(n21007), .Z(n39618) );
  XOR U41566 ( .A(n39621), .B(n39622), .Z(n21007) );
  XNOR U41567 ( .A(n21003), .B(n21005), .Z(n39622) );
  XNOR U41568 ( .A(q[9]), .B(DB[2551]), .Z(n21005) );
  XNOR U41569 ( .A(q[12]), .B(DB[2554]), .Z(n21003) );
  IV U41570 ( .A(n21002), .Z(n39621) );
  XNOR U41571 ( .A(n21000), .B(n39623), .Z(n21002) );
  XNOR U41572 ( .A(q[11]), .B(DB[2553]), .Z(n39623) );
  XNOR U41573 ( .A(q[10]), .B(DB[2552]), .Z(n21000) );
  IV U41574 ( .A(n21015), .Z(n39616) );
  XOR U41575 ( .A(n39624), .B(n39625), .Z(n21015) );
  XNOR U41576 ( .A(n21032), .B(n21013), .Z(n39625) );
  XNOR U41577 ( .A(q[1]), .B(DB[2543]), .Z(n21013) );
  XOR U41578 ( .A(n39626), .B(n21021), .Z(n21032) );
  XNOR U41579 ( .A(q[8]), .B(DB[2550]), .Z(n21021) );
  IV U41580 ( .A(n21020), .Z(n39626) );
  XNOR U41581 ( .A(n21018), .B(n39627), .Z(n21020) );
  XNOR U41582 ( .A(q[7]), .B(DB[2549]), .Z(n39627) );
  XNOR U41583 ( .A(q[6]), .B(DB[2548]), .Z(n21018) );
  IV U41584 ( .A(n21031), .Z(n39624) );
  XOR U41585 ( .A(n39628), .B(n39629), .Z(n21031) );
  XNOR U41586 ( .A(n21027), .B(n21029), .Z(n39629) );
  XNOR U41587 ( .A(q[2]), .B(DB[2544]), .Z(n21029) );
  XNOR U41588 ( .A(q[5]), .B(DB[2547]), .Z(n21027) );
  IV U41589 ( .A(n21026), .Z(n39628) );
  XNOR U41590 ( .A(n21024), .B(n39630), .Z(n21026) );
  XNOR U41591 ( .A(q[4]), .B(DB[2546]), .Z(n39630) );
  XNOR U41592 ( .A(q[3]), .B(DB[2545]), .Z(n21024) );
  XOR U41593 ( .A(n39631), .B(n20793), .Z(n20644) );
  XOR U41594 ( .A(n39632), .B(n20769), .Z(n20793) );
  XOR U41595 ( .A(n39633), .B(n20761), .Z(n20769) );
  XOR U41596 ( .A(n39634), .B(n20750), .Z(n20761) );
  XNOR U41597 ( .A(q[30]), .B(DB[2603]), .Z(n20750) );
  IV U41598 ( .A(n20749), .Z(n39634) );
  XNOR U41599 ( .A(n20747), .B(n39635), .Z(n20749) );
  XNOR U41600 ( .A(q[29]), .B(DB[2602]), .Z(n39635) );
  XNOR U41601 ( .A(q[28]), .B(DB[2601]), .Z(n20747) );
  IV U41602 ( .A(n20760), .Z(n39633) );
  XOR U41603 ( .A(n39636), .B(n39637), .Z(n20760) );
  XNOR U41604 ( .A(n20756), .B(n20758), .Z(n39637) );
  XNOR U41605 ( .A(q[24]), .B(DB[2597]), .Z(n20758) );
  XNOR U41606 ( .A(q[27]), .B(DB[2600]), .Z(n20756) );
  IV U41607 ( .A(n20755), .Z(n39636) );
  XNOR U41608 ( .A(n20753), .B(n39638), .Z(n20755) );
  XNOR U41609 ( .A(q[26]), .B(DB[2599]), .Z(n39638) );
  XNOR U41610 ( .A(q[25]), .B(DB[2598]), .Z(n20753) );
  IV U41611 ( .A(n20768), .Z(n39632) );
  XOR U41612 ( .A(n39639), .B(n39640), .Z(n20768) );
  XNOR U41613 ( .A(n20785), .B(n20766), .Z(n39640) );
  XNOR U41614 ( .A(q[16]), .B(DB[2589]), .Z(n20766) );
  XOR U41615 ( .A(n39641), .B(n20774), .Z(n20785) );
  XNOR U41616 ( .A(q[23]), .B(DB[2596]), .Z(n20774) );
  IV U41617 ( .A(n20773), .Z(n39641) );
  XNOR U41618 ( .A(n20771), .B(n39642), .Z(n20773) );
  XNOR U41619 ( .A(q[22]), .B(DB[2595]), .Z(n39642) );
  XNOR U41620 ( .A(q[21]), .B(DB[2594]), .Z(n20771) );
  IV U41621 ( .A(n20784), .Z(n39639) );
  XOR U41622 ( .A(n39643), .B(n39644), .Z(n20784) );
  XNOR U41623 ( .A(n20780), .B(n20782), .Z(n39644) );
  XNOR U41624 ( .A(q[17]), .B(DB[2590]), .Z(n20782) );
  XNOR U41625 ( .A(q[20]), .B(DB[2593]), .Z(n20780) );
  IV U41626 ( .A(n20779), .Z(n39643) );
  XNOR U41627 ( .A(n20777), .B(n39645), .Z(n20779) );
  XNOR U41628 ( .A(q[19]), .B(DB[2592]), .Z(n39645) );
  XNOR U41629 ( .A(q[18]), .B(DB[2591]), .Z(n20777) );
  IV U41630 ( .A(n20792), .Z(n39631) );
  XOR U41631 ( .A(n39646), .B(n39647), .Z(n20792) );
  XNOR U41632 ( .A(n20819), .B(n20790), .Z(n39647) );
  XNOR U41633 ( .A(q[0]), .B(DB[2573]), .Z(n20790) );
  XOR U41634 ( .A(n39648), .B(n20811), .Z(n20819) );
  XOR U41635 ( .A(n39649), .B(n20799), .Z(n20811) );
  XNOR U41636 ( .A(q[15]), .B(DB[2588]), .Z(n20799) );
  IV U41637 ( .A(n20798), .Z(n39649) );
  XNOR U41638 ( .A(n20796), .B(n39650), .Z(n20798) );
  XNOR U41639 ( .A(q[14]), .B(DB[2587]), .Z(n39650) );
  XNOR U41640 ( .A(q[13]), .B(DB[2586]), .Z(n20796) );
  IV U41641 ( .A(n20810), .Z(n39648) );
  XOR U41642 ( .A(n39651), .B(n39652), .Z(n20810) );
  XNOR U41643 ( .A(n20806), .B(n20808), .Z(n39652) );
  XNOR U41644 ( .A(q[9]), .B(DB[2582]), .Z(n20808) );
  XNOR U41645 ( .A(q[12]), .B(DB[2585]), .Z(n20806) );
  IV U41646 ( .A(n20805), .Z(n39651) );
  XNOR U41647 ( .A(n20803), .B(n39653), .Z(n20805) );
  XNOR U41648 ( .A(q[11]), .B(DB[2584]), .Z(n39653) );
  XNOR U41649 ( .A(q[10]), .B(DB[2583]), .Z(n20803) );
  IV U41650 ( .A(n20818), .Z(n39646) );
  XOR U41651 ( .A(n39654), .B(n39655), .Z(n20818) );
  XNOR U41652 ( .A(n20835), .B(n20816), .Z(n39655) );
  XNOR U41653 ( .A(q[1]), .B(DB[2574]), .Z(n20816) );
  XOR U41654 ( .A(n39656), .B(n20824), .Z(n20835) );
  XNOR U41655 ( .A(q[8]), .B(DB[2581]), .Z(n20824) );
  IV U41656 ( .A(n20823), .Z(n39656) );
  XNOR U41657 ( .A(n20821), .B(n39657), .Z(n20823) );
  XNOR U41658 ( .A(q[7]), .B(DB[2580]), .Z(n39657) );
  XNOR U41659 ( .A(q[6]), .B(DB[2579]), .Z(n20821) );
  IV U41660 ( .A(n20834), .Z(n39654) );
  XOR U41661 ( .A(n39658), .B(n39659), .Z(n20834) );
  XNOR U41662 ( .A(n20830), .B(n20832), .Z(n39659) );
  XNOR U41663 ( .A(q[2]), .B(DB[2575]), .Z(n20832) );
  XNOR U41664 ( .A(q[5]), .B(DB[2578]), .Z(n20830) );
  IV U41665 ( .A(n20829), .Z(n39658) );
  XNOR U41666 ( .A(n20827), .B(n39660), .Z(n20829) );
  XNOR U41667 ( .A(q[4]), .B(DB[2577]), .Z(n39660) );
  XNOR U41668 ( .A(q[3]), .B(DB[2576]), .Z(n20827) );
  XOR U41669 ( .A(n39661), .B(n20596), .Z(n20447) );
  XOR U41670 ( .A(n39662), .B(n20572), .Z(n20596) );
  XOR U41671 ( .A(n39663), .B(n20564), .Z(n20572) );
  XOR U41672 ( .A(n39664), .B(n20553), .Z(n20564) );
  XNOR U41673 ( .A(q[30]), .B(DB[2634]), .Z(n20553) );
  IV U41674 ( .A(n20552), .Z(n39664) );
  XNOR U41675 ( .A(n20550), .B(n39665), .Z(n20552) );
  XNOR U41676 ( .A(q[29]), .B(DB[2633]), .Z(n39665) );
  XNOR U41677 ( .A(q[28]), .B(DB[2632]), .Z(n20550) );
  IV U41678 ( .A(n20563), .Z(n39663) );
  XOR U41679 ( .A(n39666), .B(n39667), .Z(n20563) );
  XNOR U41680 ( .A(n20559), .B(n20561), .Z(n39667) );
  XNOR U41681 ( .A(q[24]), .B(DB[2628]), .Z(n20561) );
  XNOR U41682 ( .A(q[27]), .B(DB[2631]), .Z(n20559) );
  IV U41683 ( .A(n20558), .Z(n39666) );
  XNOR U41684 ( .A(n20556), .B(n39668), .Z(n20558) );
  XNOR U41685 ( .A(q[26]), .B(DB[2630]), .Z(n39668) );
  XNOR U41686 ( .A(q[25]), .B(DB[2629]), .Z(n20556) );
  IV U41687 ( .A(n20571), .Z(n39662) );
  XOR U41688 ( .A(n39669), .B(n39670), .Z(n20571) );
  XNOR U41689 ( .A(n20588), .B(n20569), .Z(n39670) );
  XNOR U41690 ( .A(q[16]), .B(DB[2620]), .Z(n20569) );
  XOR U41691 ( .A(n39671), .B(n20577), .Z(n20588) );
  XNOR U41692 ( .A(q[23]), .B(DB[2627]), .Z(n20577) );
  IV U41693 ( .A(n20576), .Z(n39671) );
  XNOR U41694 ( .A(n20574), .B(n39672), .Z(n20576) );
  XNOR U41695 ( .A(q[22]), .B(DB[2626]), .Z(n39672) );
  XNOR U41696 ( .A(q[21]), .B(DB[2625]), .Z(n20574) );
  IV U41697 ( .A(n20587), .Z(n39669) );
  XOR U41698 ( .A(n39673), .B(n39674), .Z(n20587) );
  XNOR U41699 ( .A(n20583), .B(n20585), .Z(n39674) );
  XNOR U41700 ( .A(q[17]), .B(DB[2621]), .Z(n20585) );
  XNOR U41701 ( .A(q[20]), .B(DB[2624]), .Z(n20583) );
  IV U41702 ( .A(n20582), .Z(n39673) );
  XNOR U41703 ( .A(n20580), .B(n39675), .Z(n20582) );
  XNOR U41704 ( .A(q[19]), .B(DB[2623]), .Z(n39675) );
  XNOR U41705 ( .A(q[18]), .B(DB[2622]), .Z(n20580) );
  IV U41706 ( .A(n20595), .Z(n39661) );
  XOR U41707 ( .A(n39676), .B(n39677), .Z(n20595) );
  XNOR U41708 ( .A(n20622), .B(n20593), .Z(n39677) );
  XNOR U41709 ( .A(q[0]), .B(DB[2604]), .Z(n20593) );
  XOR U41710 ( .A(n39678), .B(n20614), .Z(n20622) );
  XOR U41711 ( .A(n39679), .B(n20602), .Z(n20614) );
  XNOR U41712 ( .A(q[15]), .B(DB[2619]), .Z(n20602) );
  IV U41713 ( .A(n20601), .Z(n39679) );
  XNOR U41714 ( .A(n20599), .B(n39680), .Z(n20601) );
  XNOR U41715 ( .A(q[14]), .B(DB[2618]), .Z(n39680) );
  XNOR U41716 ( .A(q[13]), .B(DB[2617]), .Z(n20599) );
  IV U41717 ( .A(n20613), .Z(n39678) );
  XOR U41718 ( .A(n39681), .B(n39682), .Z(n20613) );
  XNOR U41719 ( .A(n20609), .B(n20611), .Z(n39682) );
  XNOR U41720 ( .A(q[9]), .B(DB[2613]), .Z(n20611) );
  XNOR U41721 ( .A(q[12]), .B(DB[2616]), .Z(n20609) );
  IV U41722 ( .A(n20608), .Z(n39681) );
  XNOR U41723 ( .A(n20606), .B(n39683), .Z(n20608) );
  XNOR U41724 ( .A(q[11]), .B(DB[2615]), .Z(n39683) );
  XNOR U41725 ( .A(q[10]), .B(DB[2614]), .Z(n20606) );
  IV U41726 ( .A(n20621), .Z(n39676) );
  XOR U41727 ( .A(n39684), .B(n39685), .Z(n20621) );
  XNOR U41728 ( .A(n20638), .B(n20619), .Z(n39685) );
  XNOR U41729 ( .A(q[1]), .B(DB[2605]), .Z(n20619) );
  XOR U41730 ( .A(n39686), .B(n20627), .Z(n20638) );
  XNOR U41731 ( .A(q[8]), .B(DB[2612]), .Z(n20627) );
  IV U41732 ( .A(n20626), .Z(n39686) );
  XNOR U41733 ( .A(n20624), .B(n39687), .Z(n20626) );
  XNOR U41734 ( .A(q[7]), .B(DB[2611]), .Z(n39687) );
  XNOR U41735 ( .A(q[6]), .B(DB[2610]), .Z(n20624) );
  IV U41736 ( .A(n20637), .Z(n39684) );
  XOR U41737 ( .A(n39688), .B(n39689), .Z(n20637) );
  XNOR U41738 ( .A(n20633), .B(n20635), .Z(n39689) );
  XNOR U41739 ( .A(q[2]), .B(DB[2606]), .Z(n20635) );
  XNOR U41740 ( .A(q[5]), .B(DB[2609]), .Z(n20633) );
  IV U41741 ( .A(n20632), .Z(n39688) );
  XNOR U41742 ( .A(n20630), .B(n39690), .Z(n20632) );
  XNOR U41743 ( .A(q[4]), .B(DB[2608]), .Z(n39690) );
  XNOR U41744 ( .A(q[3]), .B(DB[2607]), .Z(n20630) );
  XOR U41745 ( .A(n39691), .B(n20399), .Z(n20250) );
  XOR U41746 ( .A(n39692), .B(n20375), .Z(n20399) );
  XOR U41747 ( .A(n39693), .B(n20367), .Z(n20375) );
  XOR U41748 ( .A(n39694), .B(n20356), .Z(n20367) );
  XNOR U41749 ( .A(q[30]), .B(DB[2665]), .Z(n20356) );
  IV U41750 ( .A(n20355), .Z(n39694) );
  XNOR U41751 ( .A(n20353), .B(n39695), .Z(n20355) );
  XNOR U41752 ( .A(q[29]), .B(DB[2664]), .Z(n39695) );
  XNOR U41753 ( .A(q[28]), .B(DB[2663]), .Z(n20353) );
  IV U41754 ( .A(n20366), .Z(n39693) );
  XOR U41755 ( .A(n39696), .B(n39697), .Z(n20366) );
  XNOR U41756 ( .A(n20362), .B(n20364), .Z(n39697) );
  XNOR U41757 ( .A(q[24]), .B(DB[2659]), .Z(n20364) );
  XNOR U41758 ( .A(q[27]), .B(DB[2662]), .Z(n20362) );
  IV U41759 ( .A(n20361), .Z(n39696) );
  XNOR U41760 ( .A(n20359), .B(n39698), .Z(n20361) );
  XNOR U41761 ( .A(q[26]), .B(DB[2661]), .Z(n39698) );
  XNOR U41762 ( .A(q[25]), .B(DB[2660]), .Z(n20359) );
  IV U41763 ( .A(n20374), .Z(n39692) );
  XOR U41764 ( .A(n39699), .B(n39700), .Z(n20374) );
  XNOR U41765 ( .A(n20391), .B(n20372), .Z(n39700) );
  XNOR U41766 ( .A(q[16]), .B(DB[2651]), .Z(n20372) );
  XOR U41767 ( .A(n39701), .B(n20380), .Z(n20391) );
  XNOR U41768 ( .A(q[23]), .B(DB[2658]), .Z(n20380) );
  IV U41769 ( .A(n20379), .Z(n39701) );
  XNOR U41770 ( .A(n20377), .B(n39702), .Z(n20379) );
  XNOR U41771 ( .A(q[22]), .B(DB[2657]), .Z(n39702) );
  XNOR U41772 ( .A(q[21]), .B(DB[2656]), .Z(n20377) );
  IV U41773 ( .A(n20390), .Z(n39699) );
  XOR U41774 ( .A(n39703), .B(n39704), .Z(n20390) );
  XNOR U41775 ( .A(n20386), .B(n20388), .Z(n39704) );
  XNOR U41776 ( .A(q[17]), .B(DB[2652]), .Z(n20388) );
  XNOR U41777 ( .A(q[20]), .B(DB[2655]), .Z(n20386) );
  IV U41778 ( .A(n20385), .Z(n39703) );
  XNOR U41779 ( .A(n20383), .B(n39705), .Z(n20385) );
  XNOR U41780 ( .A(q[19]), .B(DB[2654]), .Z(n39705) );
  XNOR U41781 ( .A(q[18]), .B(DB[2653]), .Z(n20383) );
  IV U41782 ( .A(n20398), .Z(n39691) );
  XOR U41783 ( .A(n39706), .B(n39707), .Z(n20398) );
  XNOR U41784 ( .A(n20425), .B(n20396), .Z(n39707) );
  XNOR U41785 ( .A(q[0]), .B(DB[2635]), .Z(n20396) );
  XOR U41786 ( .A(n39708), .B(n20417), .Z(n20425) );
  XOR U41787 ( .A(n39709), .B(n20405), .Z(n20417) );
  XNOR U41788 ( .A(q[15]), .B(DB[2650]), .Z(n20405) );
  IV U41789 ( .A(n20404), .Z(n39709) );
  XNOR U41790 ( .A(n20402), .B(n39710), .Z(n20404) );
  XNOR U41791 ( .A(q[14]), .B(DB[2649]), .Z(n39710) );
  XNOR U41792 ( .A(q[13]), .B(DB[2648]), .Z(n20402) );
  IV U41793 ( .A(n20416), .Z(n39708) );
  XOR U41794 ( .A(n39711), .B(n39712), .Z(n20416) );
  XNOR U41795 ( .A(n20412), .B(n20414), .Z(n39712) );
  XNOR U41796 ( .A(q[9]), .B(DB[2644]), .Z(n20414) );
  XNOR U41797 ( .A(q[12]), .B(DB[2647]), .Z(n20412) );
  IV U41798 ( .A(n20411), .Z(n39711) );
  XNOR U41799 ( .A(n20409), .B(n39713), .Z(n20411) );
  XNOR U41800 ( .A(q[11]), .B(DB[2646]), .Z(n39713) );
  XNOR U41801 ( .A(q[10]), .B(DB[2645]), .Z(n20409) );
  IV U41802 ( .A(n20424), .Z(n39706) );
  XOR U41803 ( .A(n39714), .B(n39715), .Z(n20424) );
  XNOR U41804 ( .A(n20441), .B(n20422), .Z(n39715) );
  XNOR U41805 ( .A(q[1]), .B(DB[2636]), .Z(n20422) );
  XOR U41806 ( .A(n39716), .B(n20430), .Z(n20441) );
  XNOR U41807 ( .A(q[8]), .B(DB[2643]), .Z(n20430) );
  IV U41808 ( .A(n20429), .Z(n39716) );
  XNOR U41809 ( .A(n20427), .B(n39717), .Z(n20429) );
  XNOR U41810 ( .A(q[7]), .B(DB[2642]), .Z(n39717) );
  XNOR U41811 ( .A(q[6]), .B(DB[2641]), .Z(n20427) );
  IV U41812 ( .A(n20440), .Z(n39714) );
  XOR U41813 ( .A(n39718), .B(n39719), .Z(n20440) );
  XNOR U41814 ( .A(n20436), .B(n20438), .Z(n39719) );
  XNOR U41815 ( .A(q[2]), .B(DB[2637]), .Z(n20438) );
  XNOR U41816 ( .A(q[5]), .B(DB[2640]), .Z(n20436) );
  IV U41817 ( .A(n20435), .Z(n39718) );
  XNOR U41818 ( .A(n20433), .B(n39720), .Z(n20435) );
  XNOR U41819 ( .A(q[4]), .B(DB[2639]), .Z(n39720) );
  XNOR U41820 ( .A(q[3]), .B(DB[2638]), .Z(n20433) );
  XOR U41821 ( .A(n39721), .B(n20202), .Z(n20053) );
  XOR U41822 ( .A(n39722), .B(n20178), .Z(n20202) );
  XOR U41823 ( .A(n39723), .B(n20170), .Z(n20178) );
  XOR U41824 ( .A(n39724), .B(n20159), .Z(n20170) );
  XNOR U41825 ( .A(q[30]), .B(DB[2696]), .Z(n20159) );
  IV U41826 ( .A(n20158), .Z(n39724) );
  XNOR U41827 ( .A(n20156), .B(n39725), .Z(n20158) );
  XNOR U41828 ( .A(q[29]), .B(DB[2695]), .Z(n39725) );
  XNOR U41829 ( .A(q[28]), .B(DB[2694]), .Z(n20156) );
  IV U41830 ( .A(n20169), .Z(n39723) );
  XOR U41831 ( .A(n39726), .B(n39727), .Z(n20169) );
  XNOR U41832 ( .A(n20165), .B(n20167), .Z(n39727) );
  XNOR U41833 ( .A(q[24]), .B(DB[2690]), .Z(n20167) );
  XNOR U41834 ( .A(q[27]), .B(DB[2693]), .Z(n20165) );
  IV U41835 ( .A(n20164), .Z(n39726) );
  XNOR U41836 ( .A(n20162), .B(n39728), .Z(n20164) );
  XNOR U41837 ( .A(q[26]), .B(DB[2692]), .Z(n39728) );
  XNOR U41838 ( .A(q[25]), .B(DB[2691]), .Z(n20162) );
  IV U41839 ( .A(n20177), .Z(n39722) );
  XOR U41840 ( .A(n39729), .B(n39730), .Z(n20177) );
  XNOR U41841 ( .A(n20194), .B(n20175), .Z(n39730) );
  XNOR U41842 ( .A(q[16]), .B(DB[2682]), .Z(n20175) );
  XOR U41843 ( .A(n39731), .B(n20183), .Z(n20194) );
  XNOR U41844 ( .A(q[23]), .B(DB[2689]), .Z(n20183) );
  IV U41845 ( .A(n20182), .Z(n39731) );
  XNOR U41846 ( .A(n20180), .B(n39732), .Z(n20182) );
  XNOR U41847 ( .A(q[22]), .B(DB[2688]), .Z(n39732) );
  XNOR U41848 ( .A(q[21]), .B(DB[2687]), .Z(n20180) );
  IV U41849 ( .A(n20193), .Z(n39729) );
  XOR U41850 ( .A(n39733), .B(n39734), .Z(n20193) );
  XNOR U41851 ( .A(n20189), .B(n20191), .Z(n39734) );
  XNOR U41852 ( .A(q[17]), .B(DB[2683]), .Z(n20191) );
  XNOR U41853 ( .A(q[20]), .B(DB[2686]), .Z(n20189) );
  IV U41854 ( .A(n20188), .Z(n39733) );
  XNOR U41855 ( .A(n20186), .B(n39735), .Z(n20188) );
  XNOR U41856 ( .A(q[19]), .B(DB[2685]), .Z(n39735) );
  XNOR U41857 ( .A(q[18]), .B(DB[2684]), .Z(n20186) );
  IV U41858 ( .A(n20201), .Z(n39721) );
  XOR U41859 ( .A(n39736), .B(n39737), .Z(n20201) );
  XNOR U41860 ( .A(n20228), .B(n20199), .Z(n39737) );
  XNOR U41861 ( .A(q[0]), .B(DB[2666]), .Z(n20199) );
  XOR U41862 ( .A(n39738), .B(n20220), .Z(n20228) );
  XOR U41863 ( .A(n39739), .B(n20208), .Z(n20220) );
  XNOR U41864 ( .A(q[15]), .B(DB[2681]), .Z(n20208) );
  IV U41865 ( .A(n20207), .Z(n39739) );
  XNOR U41866 ( .A(n20205), .B(n39740), .Z(n20207) );
  XNOR U41867 ( .A(q[14]), .B(DB[2680]), .Z(n39740) );
  XNOR U41868 ( .A(q[13]), .B(DB[2679]), .Z(n20205) );
  IV U41869 ( .A(n20219), .Z(n39738) );
  XOR U41870 ( .A(n39741), .B(n39742), .Z(n20219) );
  XNOR U41871 ( .A(n20215), .B(n20217), .Z(n39742) );
  XNOR U41872 ( .A(q[9]), .B(DB[2675]), .Z(n20217) );
  XNOR U41873 ( .A(q[12]), .B(DB[2678]), .Z(n20215) );
  IV U41874 ( .A(n20214), .Z(n39741) );
  XNOR U41875 ( .A(n20212), .B(n39743), .Z(n20214) );
  XNOR U41876 ( .A(q[11]), .B(DB[2677]), .Z(n39743) );
  XNOR U41877 ( .A(q[10]), .B(DB[2676]), .Z(n20212) );
  IV U41878 ( .A(n20227), .Z(n39736) );
  XOR U41879 ( .A(n39744), .B(n39745), .Z(n20227) );
  XNOR U41880 ( .A(n20244), .B(n20225), .Z(n39745) );
  XNOR U41881 ( .A(q[1]), .B(DB[2667]), .Z(n20225) );
  XOR U41882 ( .A(n39746), .B(n20233), .Z(n20244) );
  XNOR U41883 ( .A(q[8]), .B(DB[2674]), .Z(n20233) );
  IV U41884 ( .A(n20232), .Z(n39746) );
  XNOR U41885 ( .A(n20230), .B(n39747), .Z(n20232) );
  XNOR U41886 ( .A(q[7]), .B(DB[2673]), .Z(n39747) );
  XNOR U41887 ( .A(q[6]), .B(DB[2672]), .Z(n20230) );
  IV U41888 ( .A(n20243), .Z(n39744) );
  XOR U41889 ( .A(n39748), .B(n39749), .Z(n20243) );
  XNOR U41890 ( .A(n20239), .B(n20241), .Z(n39749) );
  XNOR U41891 ( .A(q[2]), .B(DB[2668]), .Z(n20241) );
  XNOR U41892 ( .A(q[5]), .B(DB[2671]), .Z(n20239) );
  IV U41893 ( .A(n20238), .Z(n39748) );
  XNOR U41894 ( .A(n20236), .B(n39750), .Z(n20238) );
  XNOR U41895 ( .A(q[4]), .B(DB[2670]), .Z(n39750) );
  XNOR U41896 ( .A(q[3]), .B(DB[2669]), .Z(n20236) );
  XOR U41897 ( .A(n39751), .B(n20005), .Z(n19856) );
  XOR U41898 ( .A(n39752), .B(n19981), .Z(n20005) );
  XOR U41899 ( .A(n39753), .B(n19973), .Z(n19981) );
  XOR U41900 ( .A(n39754), .B(n19962), .Z(n19973) );
  XNOR U41901 ( .A(q[30]), .B(DB[2727]), .Z(n19962) );
  IV U41902 ( .A(n19961), .Z(n39754) );
  XNOR U41903 ( .A(n19959), .B(n39755), .Z(n19961) );
  XNOR U41904 ( .A(q[29]), .B(DB[2726]), .Z(n39755) );
  XNOR U41905 ( .A(q[28]), .B(DB[2725]), .Z(n19959) );
  IV U41906 ( .A(n19972), .Z(n39753) );
  XOR U41907 ( .A(n39756), .B(n39757), .Z(n19972) );
  XNOR U41908 ( .A(n19968), .B(n19970), .Z(n39757) );
  XNOR U41909 ( .A(q[24]), .B(DB[2721]), .Z(n19970) );
  XNOR U41910 ( .A(q[27]), .B(DB[2724]), .Z(n19968) );
  IV U41911 ( .A(n19967), .Z(n39756) );
  XNOR U41912 ( .A(n19965), .B(n39758), .Z(n19967) );
  XNOR U41913 ( .A(q[26]), .B(DB[2723]), .Z(n39758) );
  XNOR U41914 ( .A(q[25]), .B(DB[2722]), .Z(n19965) );
  IV U41915 ( .A(n19980), .Z(n39752) );
  XOR U41916 ( .A(n39759), .B(n39760), .Z(n19980) );
  XNOR U41917 ( .A(n19997), .B(n19978), .Z(n39760) );
  XNOR U41918 ( .A(q[16]), .B(DB[2713]), .Z(n19978) );
  XOR U41919 ( .A(n39761), .B(n19986), .Z(n19997) );
  XNOR U41920 ( .A(q[23]), .B(DB[2720]), .Z(n19986) );
  IV U41921 ( .A(n19985), .Z(n39761) );
  XNOR U41922 ( .A(n19983), .B(n39762), .Z(n19985) );
  XNOR U41923 ( .A(q[22]), .B(DB[2719]), .Z(n39762) );
  XNOR U41924 ( .A(q[21]), .B(DB[2718]), .Z(n19983) );
  IV U41925 ( .A(n19996), .Z(n39759) );
  XOR U41926 ( .A(n39763), .B(n39764), .Z(n19996) );
  XNOR U41927 ( .A(n19992), .B(n19994), .Z(n39764) );
  XNOR U41928 ( .A(q[17]), .B(DB[2714]), .Z(n19994) );
  XNOR U41929 ( .A(q[20]), .B(DB[2717]), .Z(n19992) );
  IV U41930 ( .A(n19991), .Z(n39763) );
  XNOR U41931 ( .A(n19989), .B(n39765), .Z(n19991) );
  XNOR U41932 ( .A(q[19]), .B(DB[2716]), .Z(n39765) );
  XNOR U41933 ( .A(q[18]), .B(DB[2715]), .Z(n19989) );
  IV U41934 ( .A(n20004), .Z(n39751) );
  XOR U41935 ( .A(n39766), .B(n39767), .Z(n20004) );
  XNOR U41936 ( .A(n20031), .B(n20002), .Z(n39767) );
  XNOR U41937 ( .A(q[0]), .B(DB[2697]), .Z(n20002) );
  XOR U41938 ( .A(n39768), .B(n20023), .Z(n20031) );
  XOR U41939 ( .A(n39769), .B(n20011), .Z(n20023) );
  XNOR U41940 ( .A(q[15]), .B(DB[2712]), .Z(n20011) );
  IV U41941 ( .A(n20010), .Z(n39769) );
  XNOR U41942 ( .A(n20008), .B(n39770), .Z(n20010) );
  XNOR U41943 ( .A(q[14]), .B(DB[2711]), .Z(n39770) );
  XNOR U41944 ( .A(q[13]), .B(DB[2710]), .Z(n20008) );
  IV U41945 ( .A(n20022), .Z(n39768) );
  XOR U41946 ( .A(n39771), .B(n39772), .Z(n20022) );
  XNOR U41947 ( .A(n20018), .B(n20020), .Z(n39772) );
  XNOR U41948 ( .A(q[9]), .B(DB[2706]), .Z(n20020) );
  XNOR U41949 ( .A(q[12]), .B(DB[2709]), .Z(n20018) );
  IV U41950 ( .A(n20017), .Z(n39771) );
  XNOR U41951 ( .A(n20015), .B(n39773), .Z(n20017) );
  XNOR U41952 ( .A(q[11]), .B(DB[2708]), .Z(n39773) );
  XNOR U41953 ( .A(q[10]), .B(DB[2707]), .Z(n20015) );
  IV U41954 ( .A(n20030), .Z(n39766) );
  XOR U41955 ( .A(n39774), .B(n39775), .Z(n20030) );
  XNOR U41956 ( .A(n20047), .B(n20028), .Z(n39775) );
  XNOR U41957 ( .A(q[1]), .B(DB[2698]), .Z(n20028) );
  XOR U41958 ( .A(n39776), .B(n20036), .Z(n20047) );
  XNOR U41959 ( .A(q[8]), .B(DB[2705]), .Z(n20036) );
  IV U41960 ( .A(n20035), .Z(n39776) );
  XNOR U41961 ( .A(n20033), .B(n39777), .Z(n20035) );
  XNOR U41962 ( .A(q[7]), .B(DB[2704]), .Z(n39777) );
  XNOR U41963 ( .A(q[6]), .B(DB[2703]), .Z(n20033) );
  IV U41964 ( .A(n20046), .Z(n39774) );
  XOR U41965 ( .A(n39778), .B(n39779), .Z(n20046) );
  XNOR U41966 ( .A(n20042), .B(n20044), .Z(n39779) );
  XNOR U41967 ( .A(q[2]), .B(DB[2699]), .Z(n20044) );
  XNOR U41968 ( .A(q[5]), .B(DB[2702]), .Z(n20042) );
  IV U41969 ( .A(n20041), .Z(n39778) );
  XNOR U41970 ( .A(n20039), .B(n39780), .Z(n20041) );
  XNOR U41971 ( .A(q[4]), .B(DB[2701]), .Z(n39780) );
  XNOR U41972 ( .A(q[3]), .B(DB[2700]), .Z(n20039) );
  XOR U41973 ( .A(n39781), .B(n19808), .Z(n19659) );
  XOR U41974 ( .A(n39782), .B(n19784), .Z(n19808) );
  XOR U41975 ( .A(n39783), .B(n19776), .Z(n19784) );
  XOR U41976 ( .A(n39784), .B(n19765), .Z(n19776) );
  XNOR U41977 ( .A(q[30]), .B(DB[2758]), .Z(n19765) );
  IV U41978 ( .A(n19764), .Z(n39784) );
  XNOR U41979 ( .A(n19762), .B(n39785), .Z(n19764) );
  XNOR U41980 ( .A(q[29]), .B(DB[2757]), .Z(n39785) );
  XNOR U41981 ( .A(q[28]), .B(DB[2756]), .Z(n19762) );
  IV U41982 ( .A(n19775), .Z(n39783) );
  XOR U41983 ( .A(n39786), .B(n39787), .Z(n19775) );
  XNOR U41984 ( .A(n19771), .B(n19773), .Z(n39787) );
  XNOR U41985 ( .A(q[24]), .B(DB[2752]), .Z(n19773) );
  XNOR U41986 ( .A(q[27]), .B(DB[2755]), .Z(n19771) );
  IV U41987 ( .A(n19770), .Z(n39786) );
  XNOR U41988 ( .A(n19768), .B(n39788), .Z(n19770) );
  XNOR U41989 ( .A(q[26]), .B(DB[2754]), .Z(n39788) );
  XNOR U41990 ( .A(q[25]), .B(DB[2753]), .Z(n19768) );
  IV U41991 ( .A(n19783), .Z(n39782) );
  XOR U41992 ( .A(n39789), .B(n39790), .Z(n19783) );
  XNOR U41993 ( .A(n19800), .B(n19781), .Z(n39790) );
  XNOR U41994 ( .A(q[16]), .B(DB[2744]), .Z(n19781) );
  XOR U41995 ( .A(n39791), .B(n19789), .Z(n19800) );
  XNOR U41996 ( .A(q[23]), .B(DB[2751]), .Z(n19789) );
  IV U41997 ( .A(n19788), .Z(n39791) );
  XNOR U41998 ( .A(n19786), .B(n39792), .Z(n19788) );
  XNOR U41999 ( .A(q[22]), .B(DB[2750]), .Z(n39792) );
  XNOR U42000 ( .A(q[21]), .B(DB[2749]), .Z(n19786) );
  IV U42001 ( .A(n19799), .Z(n39789) );
  XOR U42002 ( .A(n39793), .B(n39794), .Z(n19799) );
  XNOR U42003 ( .A(n19795), .B(n19797), .Z(n39794) );
  XNOR U42004 ( .A(q[17]), .B(DB[2745]), .Z(n19797) );
  XNOR U42005 ( .A(q[20]), .B(DB[2748]), .Z(n19795) );
  IV U42006 ( .A(n19794), .Z(n39793) );
  XNOR U42007 ( .A(n19792), .B(n39795), .Z(n19794) );
  XNOR U42008 ( .A(q[19]), .B(DB[2747]), .Z(n39795) );
  XNOR U42009 ( .A(q[18]), .B(DB[2746]), .Z(n19792) );
  IV U42010 ( .A(n19807), .Z(n39781) );
  XOR U42011 ( .A(n39796), .B(n39797), .Z(n19807) );
  XNOR U42012 ( .A(n19834), .B(n19805), .Z(n39797) );
  XNOR U42013 ( .A(q[0]), .B(DB[2728]), .Z(n19805) );
  XOR U42014 ( .A(n39798), .B(n19826), .Z(n19834) );
  XOR U42015 ( .A(n39799), .B(n19814), .Z(n19826) );
  XNOR U42016 ( .A(q[15]), .B(DB[2743]), .Z(n19814) );
  IV U42017 ( .A(n19813), .Z(n39799) );
  XNOR U42018 ( .A(n19811), .B(n39800), .Z(n19813) );
  XNOR U42019 ( .A(q[14]), .B(DB[2742]), .Z(n39800) );
  XNOR U42020 ( .A(q[13]), .B(DB[2741]), .Z(n19811) );
  IV U42021 ( .A(n19825), .Z(n39798) );
  XOR U42022 ( .A(n39801), .B(n39802), .Z(n19825) );
  XNOR U42023 ( .A(n19821), .B(n19823), .Z(n39802) );
  XNOR U42024 ( .A(q[9]), .B(DB[2737]), .Z(n19823) );
  XNOR U42025 ( .A(q[12]), .B(DB[2740]), .Z(n19821) );
  IV U42026 ( .A(n19820), .Z(n39801) );
  XNOR U42027 ( .A(n19818), .B(n39803), .Z(n19820) );
  XNOR U42028 ( .A(q[11]), .B(DB[2739]), .Z(n39803) );
  XNOR U42029 ( .A(q[10]), .B(DB[2738]), .Z(n19818) );
  IV U42030 ( .A(n19833), .Z(n39796) );
  XOR U42031 ( .A(n39804), .B(n39805), .Z(n19833) );
  XNOR U42032 ( .A(n19850), .B(n19831), .Z(n39805) );
  XNOR U42033 ( .A(q[1]), .B(DB[2729]), .Z(n19831) );
  XOR U42034 ( .A(n39806), .B(n19839), .Z(n19850) );
  XNOR U42035 ( .A(q[8]), .B(DB[2736]), .Z(n19839) );
  IV U42036 ( .A(n19838), .Z(n39806) );
  XNOR U42037 ( .A(n19836), .B(n39807), .Z(n19838) );
  XNOR U42038 ( .A(q[7]), .B(DB[2735]), .Z(n39807) );
  XNOR U42039 ( .A(q[6]), .B(DB[2734]), .Z(n19836) );
  IV U42040 ( .A(n19849), .Z(n39804) );
  XOR U42041 ( .A(n39808), .B(n39809), .Z(n19849) );
  XNOR U42042 ( .A(n19845), .B(n19847), .Z(n39809) );
  XNOR U42043 ( .A(q[2]), .B(DB[2730]), .Z(n19847) );
  XNOR U42044 ( .A(q[5]), .B(DB[2733]), .Z(n19845) );
  IV U42045 ( .A(n19844), .Z(n39808) );
  XNOR U42046 ( .A(n19842), .B(n39810), .Z(n19844) );
  XNOR U42047 ( .A(q[4]), .B(DB[2732]), .Z(n39810) );
  XNOR U42048 ( .A(q[3]), .B(DB[2731]), .Z(n19842) );
  XOR U42049 ( .A(n39811), .B(n19611), .Z(n19462) );
  XOR U42050 ( .A(n39812), .B(n19587), .Z(n19611) );
  XOR U42051 ( .A(n39813), .B(n19579), .Z(n19587) );
  XOR U42052 ( .A(n39814), .B(n19568), .Z(n19579) );
  XNOR U42053 ( .A(q[30]), .B(DB[2789]), .Z(n19568) );
  IV U42054 ( .A(n19567), .Z(n39814) );
  XNOR U42055 ( .A(n19565), .B(n39815), .Z(n19567) );
  XNOR U42056 ( .A(q[29]), .B(DB[2788]), .Z(n39815) );
  XNOR U42057 ( .A(q[28]), .B(DB[2787]), .Z(n19565) );
  IV U42058 ( .A(n19578), .Z(n39813) );
  XOR U42059 ( .A(n39816), .B(n39817), .Z(n19578) );
  XNOR U42060 ( .A(n19574), .B(n19576), .Z(n39817) );
  XNOR U42061 ( .A(q[24]), .B(DB[2783]), .Z(n19576) );
  XNOR U42062 ( .A(q[27]), .B(DB[2786]), .Z(n19574) );
  IV U42063 ( .A(n19573), .Z(n39816) );
  XNOR U42064 ( .A(n19571), .B(n39818), .Z(n19573) );
  XNOR U42065 ( .A(q[26]), .B(DB[2785]), .Z(n39818) );
  XNOR U42066 ( .A(q[25]), .B(DB[2784]), .Z(n19571) );
  IV U42067 ( .A(n19586), .Z(n39812) );
  XOR U42068 ( .A(n39819), .B(n39820), .Z(n19586) );
  XNOR U42069 ( .A(n19603), .B(n19584), .Z(n39820) );
  XNOR U42070 ( .A(q[16]), .B(DB[2775]), .Z(n19584) );
  XOR U42071 ( .A(n39821), .B(n19592), .Z(n19603) );
  XNOR U42072 ( .A(q[23]), .B(DB[2782]), .Z(n19592) );
  IV U42073 ( .A(n19591), .Z(n39821) );
  XNOR U42074 ( .A(n19589), .B(n39822), .Z(n19591) );
  XNOR U42075 ( .A(q[22]), .B(DB[2781]), .Z(n39822) );
  XNOR U42076 ( .A(q[21]), .B(DB[2780]), .Z(n19589) );
  IV U42077 ( .A(n19602), .Z(n39819) );
  XOR U42078 ( .A(n39823), .B(n39824), .Z(n19602) );
  XNOR U42079 ( .A(n19598), .B(n19600), .Z(n39824) );
  XNOR U42080 ( .A(q[17]), .B(DB[2776]), .Z(n19600) );
  XNOR U42081 ( .A(q[20]), .B(DB[2779]), .Z(n19598) );
  IV U42082 ( .A(n19597), .Z(n39823) );
  XNOR U42083 ( .A(n19595), .B(n39825), .Z(n19597) );
  XNOR U42084 ( .A(q[19]), .B(DB[2778]), .Z(n39825) );
  XNOR U42085 ( .A(q[18]), .B(DB[2777]), .Z(n19595) );
  IV U42086 ( .A(n19610), .Z(n39811) );
  XOR U42087 ( .A(n39826), .B(n39827), .Z(n19610) );
  XNOR U42088 ( .A(n19637), .B(n19608), .Z(n39827) );
  XNOR U42089 ( .A(q[0]), .B(DB[2759]), .Z(n19608) );
  XOR U42090 ( .A(n39828), .B(n19629), .Z(n19637) );
  XOR U42091 ( .A(n39829), .B(n19617), .Z(n19629) );
  XNOR U42092 ( .A(q[15]), .B(DB[2774]), .Z(n19617) );
  IV U42093 ( .A(n19616), .Z(n39829) );
  XNOR U42094 ( .A(n19614), .B(n39830), .Z(n19616) );
  XNOR U42095 ( .A(q[14]), .B(DB[2773]), .Z(n39830) );
  XNOR U42096 ( .A(q[13]), .B(DB[2772]), .Z(n19614) );
  IV U42097 ( .A(n19628), .Z(n39828) );
  XOR U42098 ( .A(n39831), .B(n39832), .Z(n19628) );
  XNOR U42099 ( .A(n19624), .B(n19626), .Z(n39832) );
  XNOR U42100 ( .A(q[9]), .B(DB[2768]), .Z(n19626) );
  XNOR U42101 ( .A(q[12]), .B(DB[2771]), .Z(n19624) );
  IV U42102 ( .A(n19623), .Z(n39831) );
  XNOR U42103 ( .A(n19621), .B(n39833), .Z(n19623) );
  XNOR U42104 ( .A(q[11]), .B(DB[2770]), .Z(n39833) );
  XNOR U42105 ( .A(q[10]), .B(DB[2769]), .Z(n19621) );
  IV U42106 ( .A(n19636), .Z(n39826) );
  XOR U42107 ( .A(n39834), .B(n39835), .Z(n19636) );
  XNOR U42108 ( .A(n19653), .B(n19634), .Z(n39835) );
  XNOR U42109 ( .A(q[1]), .B(DB[2760]), .Z(n19634) );
  XOR U42110 ( .A(n39836), .B(n19642), .Z(n19653) );
  XNOR U42111 ( .A(q[8]), .B(DB[2767]), .Z(n19642) );
  IV U42112 ( .A(n19641), .Z(n39836) );
  XNOR U42113 ( .A(n19639), .B(n39837), .Z(n19641) );
  XNOR U42114 ( .A(q[7]), .B(DB[2766]), .Z(n39837) );
  XNOR U42115 ( .A(q[6]), .B(DB[2765]), .Z(n19639) );
  IV U42116 ( .A(n19652), .Z(n39834) );
  XOR U42117 ( .A(n39838), .B(n39839), .Z(n19652) );
  XNOR U42118 ( .A(n19648), .B(n19650), .Z(n39839) );
  XNOR U42119 ( .A(q[2]), .B(DB[2761]), .Z(n19650) );
  XNOR U42120 ( .A(q[5]), .B(DB[2764]), .Z(n19648) );
  IV U42121 ( .A(n19647), .Z(n39838) );
  XNOR U42122 ( .A(n19645), .B(n39840), .Z(n19647) );
  XNOR U42123 ( .A(q[4]), .B(DB[2763]), .Z(n39840) );
  XNOR U42124 ( .A(q[3]), .B(DB[2762]), .Z(n19645) );
  XOR U42125 ( .A(n39841), .B(n19414), .Z(n19265) );
  XOR U42126 ( .A(n39842), .B(n19390), .Z(n19414) );
  XOR U42127 ( .A(n39843), .B(n19382), .Z(n19390) );
  XOR U42128 ( .A(n39844), .B(n19371), .Z(n19382) );
  XNOR U42129 ( .A(q[30]), .B(DB[2820]), .Z(n19371) );
  IV U42130 ( .A(n19370), .Z(n39844) );
  XNOR U42131 ( .A(n19368), .B(n39845), .Z(n19370) );
  XNOR U42132 ( .A(q[29]), .B(DB[2819]), .Z(n39845) );
  XNOR U42133 ( .A(q[28]), .B(DB[2818]), .Z(n19368) );
  IV U42134 ( .A(n19381), .Z(n39843) );
  XOR U42135 ( .A(n39846), .B(n39847), .Z(n19381) );
  XNOR U42136 ( .A(n19377), .B(n19379), .Z(n39847) );
  XNOR U42137 ( .A(q[24]), .B(DB[2814]), .Z(n19379) );
  XNOR U42138 ( .A(q[27]), .B(DB[2817]), .Z(n19377) );
  IV U42139 ( .A(n19376), .Z(n39846) );
  XNOR U42140 ( .A(n19374), .B(n39848), .Z(n19376) );
  XNOR U42141 ( .A(q[26]), .B(DB[2816]), .Z(n39848) );
  XNOR U42142 ( .A(q[25]), .B(DB[2815]), .Z(n19374) );
  IV U42143 ( .A(n19389), .Z(n39842) );
  XOR U42144 ( .A(n39849), .B(n39850), .Z(n19389) );
  XNOR U42145 ( .A(n19406), .B(n19387), .Z(n39850) );
  XNOR U42146 ( .A(q[16]), .B(DB[2806]), .Z(n19387) );
  XOR U42147 ( .A(n39851), .B(n19395), .Z(n19406) );
  XNOR U42148 ( .A(q[23]), .B(DB[2813]), .Z(n19395) );
  IV U42149 ( .A(n19394), .Z(n39851) );
  XNOR U42150 ( .A(n19392), .B(n39852), .Z(n19394) );
  XNOR U42151 ( .A(q[22]), .B(DB[2812]), .Z(n39852) );
  XNOR U42152 ( .A(q[21]), .B(DB[2811]), .Z(n19392) );
  IV U42153 ( .A(n19405), .Z(n39849) );
  XOR U42154 ( .A(n39853), .B(n39854), .Z(n19405) );
  XNOR U42155 ( .A(n19401), .B(n19403), .Z(n39854) );
  XNOR U42156 ( .A(q[17]), .B(DB[2807]), .Z(n19403) );
  XNOR U42157 ( .A(q[20]), .B(DB[2810]), .Z(n19401) );
  IV U42158 ( .A(n19400), .Z(n39853) );
  XNOR U42159 ( .A(n19398), .B(n39855), .Z(n19400) );
  XNOR U42160 ( .A(q[19]), .B(DB[2809]), .Z(n39855) );
  XNOR U42161 ( .A(q[18]), .B(DB[2808]), .Z(n19398) );
  IV U42162 ( .A(n19413), .Z(n39841) );
  XOR U42163 ( .A(n39856), .B(n39857), .Z(n19413) );
  XNOR U42164 ( .A(n19440), .B(n19411), .Z(n39857) );
  XNOR U42165 ( .A(q[0]), .B(DB[2790]), .Z(n19411) );
  XOR U42166 ( .A(n39858), .B(n19432), .Z(n19440) );
  XOR U42167 ( .A(n39859), .B(n19420), .Z(n19432) );
  XNOR U42168 ( .A(q[15]), .B(DB[2805]), .Z(n19420) );
  IV U42169 ( .A(n19419), .Z(n39859) );
  XNOR U42170 ( .A(n19417), .B(n39860), .Z(n19419) );
  XNOR U42171 ( .A(q[14]), .B(DB[2804]), .Z(n39860) );
  XNOR U42172 ( .A(q[13]), .B(DB[2803]), .Z(n19417) );
  IV U42173 ( .A(n19431), .Z(n39858) );
  XOR U42174 ( .A(n39861), .B(n39862), .Z(n19431) );
  XNOR U42175 ( .A(n19427), .B(n19429), .Z(n39862) );
  XNOR U42176 ( .A(q[9]), .B(DB[2799]), .Z(n19429) );
  XNOR U42177 ( .A(q[12]), .B(DB[2802]), .Z(n19427) );
  IV U42178 ( .A(n19426), .Z(n39861) );
  XNOR U42179 ( .A(n19424), .B(n39863), .Z(n19426) );
  XNOR U42180 ( .A(q[11]), .B(DB[2801]), .Z(n39863) );
  XNOR U42181 ( .A(q[10]), .B(DB[2800]), .Z(n19424) );
  IV U42182 ( .A(n19439), .Z(n39856) );
  XOR U42183 ( .A(n39864), .B(n39865), .Z(n19439) );
  XNOR U42184 ( .A(n19456), .B(n19437), .Z(n39865) );
  XNOR U42185 ( .A(q[1]), .B(DB[2791]), .Z(n19437) );
  XOR U42186 ( .A(n39866), .B(n19445), .Z(n19456) );
  XNOR U42187 ( .A(q[8]), .B(DB[2798]), .Z(n19445) );
  IV U42188 ( .A(n19444), .Z(n39866) );
  XNOR U42189 ( .A(n19442), .B(n39867), .Z(n19444) );
  XNOR U42190 ( .A(q[7]), .B(DB[2797]), .Z(n39867) );
  XNOR U42191 ( .A(q[6]), .B(DB[2796]), .Z(n19442) );
  IV U42192 ( .A(n19455), .Z(n39864) );
  XOR U42193 ( .A(n39868), .B(n39869), .Z(n19455) );
  XNOR U42194 ( .A(n19451), .B(n19453), .Z(n39869) );
  XNOR U42195 ( .A(q[2]), .B(DB[2792]), .Z(n19453) );
  XNOR U42196 ( .A(q[5]), .B(DB[2795]), .Z(n19451) );
  IV U42197 ( .A(n19450), .Z(n39868) );
  XNOR U42198 ( .A(n19448), .B(n39870), .Z(n19450) );
  XNOR U42199 ( .A(q[4]), .B(DB[2794]), .Z(n39870) );
  XNOR U42200 ( .A(q[3]), .B(DB[2793]), .Z(n19448) );
  XOR U42201 ( .A(n39871), .B(n19217), .Z(n19068) );
  XOR U42202 ( .A(n39872), .B(n19193), .Z(n19217) );
  XOR U42203 ( .A(n39873), .B(n19185), .Z(n19193) );
  XOR U42204 ( .A(n39874), .B(n19174), .Z(n19185) );
  XNOR U42205 ( .A(q[30]), .B(DB[2851]), .Z(n19174) );
  IV U42206 ( .A(n19173), .Z(n39874) );
  XNOR U42207 ( .A(n19171), .B(n39875), .Z(n19173) );
  XNOR U42208 ( .A(q[29]), .B(DB[2850]), .Z(n39875) );
  XNOR U42209 ( .A(q[28]), .B(DB[2849]), .Z(n19171) );
  IV U42210 ( .A(n19184), .Z(n39873) );
  XOR U42211 ( .A(n39876), .B(n39877), .Z(n19184) );
  XNOR U42212 ( .A(n19180), .B(n19182), .Z(n39877) );
  XNOR U42213 ( .A(q[24]), .B(DB[2845]), .Z(n19182) );
  XNOR U42214 ( .A(q[27]), .B(DB[2848]), .Z(n19180) );
  IV U42215 ( .A(n19179), .Z(n39876) );
  XNOR U42216 ( .A(n19177), .B(n39878), .Z(n19179) );
  XNOR U42217 ( .A(q[26]), .B(DB[2847]), .Z(n39878) );
  XNOR U42218 ( .A(q[25]), .B(DB[2846]), .Z(n19177) );
  IV U42219 ( .A(n19192), .Z(n39872) );
  XOR U42220 ( .A(n39879), .B(n39880), .Z(n19192) );
  XNOR U42221 ( .A(n19209), .B(n19190), .Z(n39880) );
  XNOR U42222 ( .A(q[16]), .B(DB[2837]), .Z(n19190) );
  XOR U42223 ( .A(n39881), .B(n19198), .Z(n19209) );
  XNOR U42224 ( .A(q[23]), .B(DB[2844]), .Z(n19198) );
  IV U42225 ( .A(n19197), .Z(n39881) );
  XNOR U42226 ( .A(n19195), .B(n39882), .Z(n19197) );
  XNOR U42227 ( .A(q[22]), .B(DB[2843]), .Z(n39882) );
  XNOR U42228 ( .A(q[21]), .B(DB[2842]), .Z(n19195) );
  IV U42229 ( .A(n19208), .Z(n39879) );
  XOR U42230 ( .A(n39883), .B(n39884), .Z(n19208) );
  XNOR U42231 ( .A(n19204), .B(n19206), .Z(n39884) );
  XNOR U42232 ( .A(q[17]), .B(DB[2838]), .Z(n19206) );
  XNOR U42233 ( .A(q[20]), .B(DB[2841]), .Z(n19204) );
  IV U42234 ( .A(n19203), .Z(n39883) );
  XNOR U42235 ( .A(n19201), .B(n39885), .Z(n19203) );
  XNOR U42236 ( .A(q[19]), .B(DB[2840]), .Z(n39885) );
  XNOR U42237 ( .A(q[18]), .B(DB[2839]), .Z(n19201) );
  IV U42238 ( .A(n19216), .Z(n39871) );
  XOR U42239 ( .A(n39886), .B(n39887), .Z(n19216) );
  XNOR U42240 ( .A(n19243), .B(n19214), .Z(n39887) );
  XNOR U42241 ( .A(q[0]), .B(DB[2821]), .Z(n19214) );
  XOR U42242 ( .A(n39888), .B(n19235), .Z(n19243) );
  XOR U42243 ( .A(n39889), .B(n19223), .Z(n19235) );
  XNOR U42244 ( .A(q[15]), .B(DB[2836]), .Z(n19223) );
  IV U42245 ( .A(n19222), .Z(n39889) );
  XNOR U42246 ( .A(n19220), .B(n39890), .Z(n19222) );
  XNOR U42247 ( .A(q[14]), .B(DB[2835]), .Z(n39890) );
  XNOR U42248 ( .A(q[13]), .B(DB[2834]), .Z(n19220) );
  IV U42249 ( .A(n19234), .Z(n39888) );
  XOR U42250 ( .A(n39891), .B(n39892), .Z(n19234) );
  XNOR U42251 ( .A(n19230), .B(n19232), .Z(n39892) );
  XNOR U42252 ( .A(q[9]), .B(DB[2830]), .Z(n19232) );
  XNOR U42253 ( .A(q[12]), .B(DB[2833]), .Z(n19230) );
  IV U42254 ( .A(n19229), .Z(n39891) );
  XNOR U42255 ( .A(n19227), .B(n39893), .Z(n19229) );
  XNOR U42256 ( .A(q[11]), .B(DB[2832]), .Z(n39893) );
  XNOR U42257 ( .A(q[10]), .B(DB[2831]), .Z(n19227) );
  IV U42258 ( .A(n19242), .Z(n39886) );
  XOR U42259 ( .A(n39894), .B(n39895), .Z(n19242) );
  XNOR U42260 ( .A(n19259), .B(n19240), .Z(n39895) );
  XNOR U42261 ( .A(q[1]), .B(DB[2822]), .Z(n19240) );
  XOR U42262 ( .A(n39896), .B(n19248), .Z(n19259) );
  XNOR U42263 ( .A(q[8]), .B(DB[2829]), .Z(n19248) );
  IV U42264 ( .A(n19247), .Z(n39896) );
  XNOR U42265 ( .A(n19245), .B(n39897), .Z(n19247) );
  XNOR U42266 ( .A(q[7]), .B(DB[2828]), .Z(n39897) );
  XNOR U42267 ( .A(q[6]), .B(DB[2827]), .Z(n19245) );
  IV U42268 ( .A(n19258), .Z(n39894) );
  XOR U42269 ( .A(n39898), .B(n39899), .Z(n19258) );
  XNOR U42270 ( .A(n19254), .B(n19256), .Z(n39899) );
  XNOR U42271 ( .A(q[2]), .B(DB[2823]), .Z(n19256) );
  XNOR U42272 ( .A(q[5]), .B(DB[2826]), .Z(n19254) );
  IV U42273 ( .A(n19253), .Z(n39898) );
  XNOR U42274 ( .A(n19251), .B(n39900), .Z(n19253) );
  XNOR U42275 ( .A(q[4]), .B(DB[2825]), .Z(n39900) );
  XNOR U42276 ( .A(q[3]), .B(DB[2824]), .Z(n19251) );
  XOR U42277 ( .A(n39901), .B(n19020), .Z(n18871) );
  XOR U42278 ( .A(n39902), .B(n18996), .Z(n19020) );
  XOR U42279 ( .A(n39903), .B(n18988), .Z(n18996) );
  XOR U42280 ( .A(n39904), .B(n18977), .Z(n18988) );
  XNOR U42281 ( .A(q[30]), .B(DB[2882]), .Z(n18977) );
  IV U42282 ( .A(n18976), .Z(n39904) );
  XNOR U42283 ( .A(n18974), .B(n39905), .Z(n18976) );
  XNOR U42284 ( .A(q[29]), .B(DB[2881]), .Z(n39905) );
  XNOR U42285 ( .A(q[28]), .B(DB[2880]), .Z(n18974) );
  IV U42286 ( .A(n18987), .Z(n39903) );
  XOR U42287 ( .A(n39906), .B(n39907), .Z(n18987) );
  XNOR U42288 ( .A(n18983), .B(n18985), .Z(n39907) );
  XNOR U42289 ( .A(q[24]), .B(DB[2876]), .Z(n18985) );
  XNOR U42290 ( .A(q[27]), .B(DB[2879]), .Z(n18983) );
  IV U42291 ( .A(n18982), .Z(n39906) );
  XNOR U42292 ( .A(n18980), .B(n39908), .Z(n18982) );
  XNOR U42293 ( .A(q[26]), .B(DB[2878]), .Z(n39908) );
  XNOR U42294 ( .A(q[25]), .B(DB[2877]), .Z(n18980) );
  IV U42295 ( .A(n18995), .Z(n39902) );
  XOR U42296 ( .A(n39909), .B(n39910), .Z(n18995) );
  XNOR U42297 ( .A(n19012), .B(n18993), .Z(n39910) );
  XNOR U42298 ( .A(q[16]), .B(DB[2868]), .Z(n18993) );
  XOR U42299 ( .A(n39911), .B(n19001), .Z(n19012) );
  XNOR U42300 ( .A(q[23]), .B(DB[2875]), .Z(n19001) );
  IV U42301 ( .A(n19000), .Z(n39911) );
  XNOR U42302 ( .A(n18998), .B(n39912), .Z(n19000) );
  XNOR U42303 ( .A(q[22]), .B(DB[2874]), .Z(n39912) );
  XNOR U42304 ( .A(q[21]), .B(DB[2873]), .Z(n18998) );
  IV U42305 ( .A(n19011), .Z(n39909) );
  XOR U42306 ( .A(n39913), .B(n39914), .Z(n19011) );
  XNOR U42307 ( .A(n19007), .B(n19009), .Z(n39914) );
  XNOR U42308 ( .A(q[17]), .B(DB[2869]), .Z(n19009) );
  XNOR U42309 ( .A(q[20]), .B(DB[2872]), .Z(n19007) );
  IV U42310 ( .A(n19006), .Z(n39913) );
  XNOR U42311 ( .A(n19004), .B(n39915), .Z(n19006) );
  XNOR U42312 ( .A(q[19]), .B(DB[2871]), .Z(n39915) );
  XNOR U42313 ( .A(q[18]), .B(DB[2870]), .Z(n19004) );
  IV U42314 ( .A(n19019), .Z(n39901) );
  XOR U42315 ( .A(n39916), .B(n39917), .Z(n19019) );
  XNOR U42316 ( .A(n19046), .B(n19017), .Z(n39917) );
  XNOR U42317 ( .A(q[0]), .B(DB[2852]), .Z(n19017) );
  XOR U42318 ( .A(n39918), .B(n19038), .Z(n19046) );
  XOR U42319 ( .A(n39919), .B(n19026), .Z(n19038) );
  XNOR U42320 ( .A(q[15]), .B(DB[2867]), .Z(n19026) );
  IV U42321 ( .A(n19025), .Z(n39919) );
  XNOR U42322 ( .A(n19023), .B(n39920), .Z(n19025) );
  XNOR U42323 ( .A(q[14]), .B(DB[2866]), .Z(n39920) );
  XNOR U42324 ( .A(q[13]), .B(DB[2865]), .Z(n19023) );
  IV U42325 ( .A(n19037), .Z(n39918) );
  XOR U42326 ( .A(n39921), .B(n39922), .Z(n19037) );
  XNOR U42327 ( .A(n19033), .B(n19035), .Z(n39922) );
  XNOR U42328 ( .A(q[9]), .B(DB[2861]), .Z(n19035) );
  XNOR U42329 ( .A(q[12]), .B(DB[2864]), .Z(n19033) );
  IV U42330 ( .A(n19032), .Z(n39921) );
  XNOR U42331 ( .A(n19030), .B(n39923), .Z(n19032) );
  XNOR U42332 ( .A(q[11]), .B(DB[2863]), .Z(n39923) );
  XNOR U42333 ( .A(q[10]), .B(DB[2862]), .Z(n19030) );
  IV U42334 ( .A(n19045), .Z(n39916) );
  XOR U42335 ( .A(n39924), .B(n39925), .Z(n19045) );
  XNOR U42336 ( .A(n19062), .B(n19043), .Z(n39925) );
  XNOR U42337 ( .A(q[1]), .B(DB[2853]), .Z(n19043) );
  XOR U42338 ( .A(n39926), .B(n19051), .Z(n19062) );
  XNOR U42339 ( .A(q[8]), .B(DB[2860]), .Z(n19051) );
  IV U42340 ( .A(n19050), .Z(n39926) );
  XNOR U42341 ( .A(n19048), .B(n39927), .Z(n19050) );
  XNOR U42342 ( .A(q[7]), .B(DB[2859]), .Z(n39927) );
  XNOR U42343 ( .A(q[6]), .B(DB[2858]), .Z(n19048) );
  IV U42344 ( .A(n19061), .Z(n39924) );
  XOR U42345 ( .A(n39928), .B(n39929), .Z(n19061) );
  XNOR U42346 ( .A(n19057), .B(n19059), .Z(n39929) );
  XNOR U42347 ( .A(q[2]), .B(DB[2854]), .Z(n19059) );
  XNOR U42348 ( .A(q[5]), .B(DB[2857]), .Z(n19057) );
  IV U42349 ( .A(n19056), .Z(n39928) );
  XNOR U42350 ( .A(n19054), .B(n39930), .Z(n19056) );
  XNOR U42351 ( .A(q[4]), .B(DB[2856]), .Z(n39930) );
  XNOR U42352 ( .A(q[3]), .B(DB[2855]), .Z(n19054) );
  XOR U42353 ( .A(n39931), .B(n18823), .Z(n18674) );
  XOR U42354 ( .A(n39932), .B(n18799), .Z(n18823) );
  XOR U42355 ( .A(n39933), .B(n18791), .Z(n18799) );
  XOR U42356 ( .A(n39934), .B(n18780), .Z(n18791) );
  XNOR U42357 ( .A(q[30]), .B(DB[2913]), .Z(n18780) );
  IV U42358 ( .A(n18779), .Z(n39934) );
  XNOR U42359 ( .A(n18777), .B(n39935), .Z(n18779) );
  XNOR U42360 ( .A(q[29]), .B(DB[2912]), .Z(n39935) );
  XNOR U42361 ( .A(q[28]), .B(DB[2911]), .Z(n18777) );
  IV U42362 ( .A(n18790), .Z(n39933) );
  XOR U42363 ( .A(n39936), .B(n39937), .Z(n18790) );
  XNOR U42364 ( .A(n18786), .B(n18788), .Z(n39937) );
  XNOR U42365 ( .A(q[24]), .B(DB[2907]), .Z(n18788) );
  XNOR U42366 ( .A(q[27]), .B(DB[2910]), .Z(n18786) );
  IV U42367 ( .A(n18785), .Z(n39936) );
  XNOR U42368 ( .A(n18783), .B(n39938), .Z(n18785) );
  XNOR U42369 ( .A(q[26]), .B(DB[2909]), .Z(n39938) );
  XNOR U42370 ( .A(q[25]), .B(DB[2908]), .Z(n18783) );
  IV U42371 ( .A(n18798), .Z(n39932) );
  XOR U42372 ( .A(n39939), .B(n39940), .Z(n18798) );
  XNOR U42373 ( .A(n18815), .B(n18796), .Z(n39940) );
  XNOR U42374 ( .A(q[16]), .B(DB[2899]), .Z(n18796) );
  XOR U42375 ( .A(n39941), .B(n18804), .Z(n18815) );
  XNOR U42376 ( .A(q[23]), .B(DB[2906]), .Z(n18804) );
  IV U42377 ( .A(n18803), .Z(n39941) );
  XNOR U42378 ( .A(n18801), .B(n39942), .Z(n18803) );
  XNOR U42379 ( .A(q[22]), .B(DB[2905]), .Z(n39942) );
  XNOR U42380 ( .A(q[21]), .B(DB[2904]), .Z(n18801) );
  IV U42381 ( .A(n18814), .Z(n39939) );
  XOR U42382 ( .A(n39943), .B(n39944), .Z(n18814) );
  XNOR U42383 ( .A(n18810), .B(n18812), .Z(n39944) );
  XNOR U42384 ( .A(q[17]), .B(DB[2900]), .Z(n18812) );
  XNOR U42385 ( .A(q[20]), .B(DB[2903]), .Z(n18810) );
  IV U42386 ( .A(n18809), .Z(n39943) );
  XNOR U42387 ( .A(n18807), .B(n39945), .Z(n18809) );
  XNOR U42388 ( .A(q[19]), .B(DB[2902]), .Z(n39945) );
  XNOR U42389 ( .A(q[18]), .B(DB[2901]), .Z(n18807) );
  IV U42390 ( .A(n18822), .Z(n39931) );
  XOR U42391 ( .A(n39946), .B(n39947), .Z(n18822) );
  XNOR U42392 ( .A(n18849), .B(n18820), .Z(n39947) );
  XNOR U42393 ( .A(q[0]), .B(DB[2883]), .Z(n18820) );
  XOR U42394 ( .A(n39948), .B(n18841), .Z(n18849) );
  XOR U42395 ( .A(n39949), .B(n18829), .Z(n18841) );
  XNOR U42396 ( .A(q[15]), .B(DB[2898]), .Z(n18829) );
  IV U42397 ( .A(n18828), .Z(n39949) );
  XNOR U42398 ( .A(n18826), .B(n39950), .Z(n18828) );
  XNOR U42399 ( .A(q[14]), .B(DB[2897]), .Z(n39950) );
  XNOR U42400 ( .A(q[13]), .B(DB[2896]), .Z(n18826) );
  IV U42401 ( .A(n18840), .Z(n39948) );
  XOR U42402 ( .A(n39951), .B(n39952), .Z(n18840) );
  XNOR U42403 ( .A(n18836), .B(n18838), .Z(n39952) );
  XNOR U42404 ( .A(q[9]), .B(DB[2892]), .Z(n18838) );
  XNOR U42405 ( .A(q[12]), .B(DB[2895]), .Z(n18836) );
  IV U42406 ( .A(n18835), .Z(n39951) );
  XNOR U42407 ( .A(n18833), .B(n39953), .Z(n18835) );
  XNOR U42408 ( .A(q[11]), .B(DB[2894]), .Z(n39953) );
  XNOR U42409 ( .A(q[10]), .B(DB[2893]), .Z(n18833) );
  IV U42410 ( .A(n18848), .Z(n39946) );
  XOR U42411 ( .A(n39954), .B(n39955), .Z(n18848) );
  XNOR U42412 ( .A(n18865), .B(n18846), .Z(n39955) );
  XNOR U42413 ( .A(q[1]), .B(DB[2884]), .Z(n18846) );
  XOR U42414 ( .A(n39956), .B(n18854), .Z(n18865) );
  XNOR U42415 ( .A(q[8]), .B(DB[2891]), .Z(n18854) );
  IV U42416 ( .A(n18853), .Z(n39956) );
  XNOR U42417 ( .A(n18851), .B(n39957), .Z(n18853) );
  XNOR U42418 ( .A(q[7]), .B(DB[2890]), .Z(n39957) );
  XNOR U42419 ( .A(q[6]), .B(DB[2889]), .Z(n18851) );
  IV U42420 ( .A(n18864), .Z(n39954) );
  XOR U42421 ( .A(n39958), .B(n39959), .Z(n18864) );
  XNOR U42422 ( .A(n18860), .B(n18862), .Z(n39959) );
  XNOR U42423 ( .A(q[2]), .B(DB[2885]), .Z(n18862) );
  XNOR U42424 ( .A(q[5]), .B(DB[2888]), .Z(n18860) );
  IV U42425 ( .A(n18859), .Z(n39958) );
  XNOR U42426 ( .A(n18857), .B(n39960), .Z(n18859) );
  XNOR U42427 ( .A(q[4]), .B(DB[2887]), .Z(n39960) );
  XNOR U42428 ( .A(q[3]), .B(DB[2886]), .Z(n18857) );
  XOR U42429 ( .A(n39961), .B(n18626), .Z(n18477) );
  XOR U42430 ( .A(n39962), .B(n18602), .Z(n18626) );
  XOR U42431 ( .A(n39963), .B(n18594), .Z(n18602) );
  XOR U42432 ( .A(n39964), .B(n18583), .Z(n18594) );
  XNOR U42433 ( .A(q[30]), .B(DB[2944]), .Z(n18583) );
  IV U42434 ( .A(n18582), .Z(n39964) );
  XNOR U42435 ( .A(n18580), .B(n39965), .Z(n18582) );
  XNOR U42436 ( .A(q[29]), .B(DB[2943]), .Z(n39965) );
  XNOR U42437 ( .A(q[28]), .B(DB[2942]), .Z(n18580) );
  IV U42438 ( .A(n18593), .Z(n39963) );
  XOR U42439 ( .A(n39966), .B(n39967), .Z(n18593) );
  XNOR U42440 ( .A(n18589), .B(n18591), .Z(n39967) );
  XNOR U42441 ( .A(q[24]), .B(DB[2938]), .Z(n18591) );
  XNOR U42442 ( .A(q[27]), .B(DB[2941]), .Z(n18589) );
  IV U42443 ( .A(n18588), .Z(n39966) );
  XNOR U42444 ( .A(n18586), .B(n39968), .Z(n18588) );
  XNOR U42445 ( .A(q[26]), .B(DB[2940]), .Z(n39968) );
  XNOR U42446 ( .A(q[25]), .B(DB[2939]), .Z(n18586) );
  IV U42447 ( .A(n18601), .Z(n39962) );
  XOR U42448 ( .A(n39969), .B(n39970), .Z(n18601) );
  XNOR U42449 ( .A(n18618), .B(n18599), .Z(n39970) );
  XNOR U42450 ( .A(q[16]), .B(DB[2930]), .Z(n18599) );
  XOR U42451 ( .A(n39971), .B(n18607), .Z(n18618) );
  XNOR U42452 ( .A(q[23]), .B(DB[2937]), .Z(n18607) );
  IV U42453 ( .A(n18606), .Z(n39971) );
  XNOR U42454 ( .A(n18604), .B(n39972), .Z(n18606) );
  XNOR U42455 ( .A(q[22]), .B(DB[2936]), .Z(n39972) );
  XNOR U42456 ( .A(q[21]), .B(DB[2935]), .Z(n18604) );
  IV U42457 ( .A(n18617), .Z(n39969) );
  XOR U42458 ( .A(n39973), .B(n39974), .Z(n18617) );
  XNOR U42459 ( .A(n18613), .B(n18615), .Z(n39974) );
  XNOR U42460 ( .A(q[17]), .B(DB[2931]), .Z(n18615) );
  XNOR U42461 ( .A(q[20]), .B(DB[2934]), .Z(n18613) );
  IV U42462 ( .A(n18612), .Z(n39973) );
  XNOR U42463 ( .A(n18610), .B(n39975), .Z(n18612) );
  XNOR U42464 ( .A(q[19]), .B(DB[2933]), .Z(n39975) );
  XNOR U42465 ( .A(q[18]), .B(DB[2932]), .Z(n18610) );
  IV U42466 ( .A(n18625), .Z(n39961) );
  XOR U42467 ( .A(n39976), .B(n39977), .Z(n18625) );
  XNOR U42468 ( .A(n18652), .B(n18623), .Z(n39977) );
  XNOR U42469 ( .A(q[0]), .B(DB[2914]), .Z(n18623) );
  XOR U42470 ( .A(n39978), .B(n18644), .Z(n18652) );
  XOR U42471 ( .A(n39979), .B(n18632), .Z(n18644) );
  XNOR U42472 ( .A(q[15]), .B(DB[2929]), .Z(n18632) );
  IV U42473 ( .A(n18631), .Z(n39979) );
  XNOR U42474 ( .A(n18629), .B(n39980), .Z(n18631) );
  XNOR U42475 ( .A(q[14]), .B(DB[2928]), .Z(n39980) );
  XNOR U42476 ( .A(q[13]), .B(DB[2927]), .Z(n18629) );
  IV U42477 ( .A(n18643), .Z(n39978) );
  XOR U42478 ( .A(n39981), .B(n39982), .Z(n18643) );
  XNOR U42479 ( .A(n18639), .B(n18641), .Z(n39982) );
  XNOR U42480 ( .A(q[9]), .B(DB[2923]), .Z(n18641) );
  XNOR U42481 ( .A(q[12]), .B(DB[2926]), .Z(n18639) );
  IV U42482 ( .A(n18638), .Z(n39981) );
  XNOR U42483 ( .A(n18636), .B(n39983), .Z(n18638) );
  XNOR U42484 ( .A(q[11]), .B(DB[2925]), .Z(n39983) );
  XNOR U42485 ( .A(q[10]), .B(DB[2924]), .Z(n18636) );
  IV U42486 ( .A(n18651), .Z(n39976) );
  XOR U42487 ( .A(n39984), .B(n39985), .Z(n18651) );
  XNOR U42488 ( .A(n18668), .B(n18649), .Z(n39985) );
  XNOR U42489 ( .A(q[1]), .B(DB[2915]), .Z(n18649) );
  XOR U42490 ( .A(n39986), .B(n18657), .Z(n18668) );
  XNOR U42491 ( .A(q[8]), .B(DB[2922]), .Z(n18657) );
  IV U42492 ( .A(n18656), .Z(n39986) );
  XNOR U42493 ( .A(n18654), .B(n39987), .Z(n18656) );
  XNOR U42494 ( .A(q[7]), .B(DB[2921]), .Z(n39987) );
  XNOR U42495 ( .A(q[6]), .B(DB[2920]), .Z(n18654) );
  IV U42496 ( .A(n18667), .Z(n39984) );
  XOR U42497 ( .A(n39988), .B(n39989), .Z(n18667) );
  XNOR U42498 ( .A(n18663), .B(n18665), .Z(n39989) );
  XNOR U42499 ( .A(q[2]), .B(DB[2916]), .Z(n18665) );
  XNOR U42500 ( .A(q[5]), .B(DB[2919]), .Z(n18663) );
  IV U42501 ( .A(n18662), .Z(n39988) );
  XNOR U42502 ( .A(n18660), .B(n39990), .Z(n18662) );
  XNOR U42503 ( .A(q[4]), .B(DB[2918]), .Z(n39990) );
  XNOR U42504 ( .A(q[3]), .B(DB[2917]), .Z(n18660) );
  XOR U42505 ( .A(n39991), .B(n18429), .Z(n18280) );
  XOR U42506 ( .A(n39992), .B(n18405), .Z(n18429) );
  XOR U42507 ( .A(n39993), .B(n18397), .Z(n18405) );
  XOR U42508 ( .A(n39994), .B(n18386), .Z(n18397) );
  XNOR U42509 ( .A(q[30]), .B(DB[2975]), .Z(n18386) );
  IV U42510 ( .A(n18385), .Z(n39994) );
  XNOR U42511 ( .A(n18383), .B(n39995), .Z(n18385) );
  XNOR U42512 ( .A(q[29]), .B(DB[2974]), .Z(n39995) );
  XNOR U42513 ( .A(q[28]), .B(DB[2973]), .Z(n18383) );
  IV U42514 ( .A(n18396), .Z(n39993) );
  XOR U42515 ( .A(n39996), .B(n39997), .Z(n18396) );
  XNOR U42516 ( .A(n18392), .B(n18394), .Z(n39997) );
  XNOR U42517 ( .A(q[24]), .B(DB[2969]), .Z(n18394) );
  XNOR U42518 ( .A(q[27]), .B(DB[2972]), .Z(n18392) );
  IV U42519 ( .A(n18391), .Z(n39996) );
  XNOR U42520 ( .A(n18389), .B(n39998), .Z(n18391) );
  XNOR U42521 ( .A(q[26]), .B(DB[2971]), .Z(n39998) );
  XNOR U42522 ( .A(q[25]), .B(DB[2970]), .Z(n18389) );
  IV U42523 ( .A(n18404), .Z(n39992) );
  XOR U42524 ( .A(n39999), .B(n40000), .Z(n18404) );
  XNOR U42525 ( .A(n18421), .B(n18402), .Z(n40000) );
  XNOR U42526 ( .A(q[16]), .B(DB[2961]), .Z(n18402) );
  XOR U42527 ( .A(n40001), .B(n18410), .Z(n18421) );
  XNOR U42528 ( .A(q[23]), .B(DB[2968]), .Z(n18410) );
  IV U42529 ( .A(n18409), .Z(n40001) );
  XNOR U42530 ( .A(n18407), .B(n40002), .Z(n18409) );
  XNOR U42531 ( .A(q[22]), .B(DB[2967]), .Z(n40002) );
  XNOR U42532 ( .A(q[21]), .B(DB[2966]), .Z(n18407) );
  IV U42533 ( .A(n18420), .Z(n39999) );
  XOR U42534 ( .A(n40003), .B(n40004), .Z(n18420) );
  XNOR U42535 ( .A(n18416), .B(n18418), .Z(n40004) );
  XNOR U42536 ( .A(q[17]), .B(DB[2962]), .Z(n18418) );
  XNOR U42537 ( .A(q[20]), .B(DB[2965]), .Z(n18416) );
  IV U42538 ( .A(n18415), .Z(n40003) );
  XNOR U42539 ( .A(n18413), .B(n40005), .Z(n18415) );
  XNOR U42540 ( .A(q[19]), .B(DB[2964]), .Z(n40005) );
  XNOR U42541 ( .A(q[18]), .B(DB[2963]), .Z(n18413) );
  IV U42542 ( .A(n18428), .Z(n39991) );
  XOR U42543 ( .A(n40006), .B(n40007), .Z(n18428) );
  XNOR U42544 ( .A(n18455), .B(n18426), .Z(n40007) );
  XNOR U42545 ( .A(q[0]), .B(DB[2945]), .Z(n18426) );
  XOR U42546 ( .A(n40008), .B(n18447), .Z(n18455) );
  XOR U42547 ( .A(n40009), .B(n18435), .Z(n18447) );
  XNOR U42548 ( .A(q[15]), .B(DB[2960]), .Z(n18435) );
  IV U42549 ( .A(n18434), .Z(n40009) );
  XNOR U42550 ( .A(n18432), .B(n40010), .Z(n18434) );
  XNOR U42551 ( .A(q[14]), .B(DB[2959]), .Z(n40010) );
  XNOR U42552 ( .A(q[13]), .B(DB[2958]), .Z(n18432) );
  IV U42553 ( .A(n18446), .Z(n40008) );
  XOR U42554 ( .A(n40011), .B(n40012), .Z(n18446) );
  XNOR U42555 ( .A(n18442), .B(n18444), .Z(n40012) );
  XNOR U42556 ( .A(q[9]), .B(DB[2954]), .Z(n18444) );
  XNOR U42557 ( .A(q[12]), .B(DB[2957]), .Z(n18442) );
  IV U42558 ( .A(n18441), .Z(n40011) );
  XNOR U42559 ( .A(n18439), .B(n40013), .Z(n18441) );
  XNOR U42560 ( .A(q[11]), .B(DB[2956]), .Z(n40013) );
  XNOR U42561 ( .A(q[10]), .B(DB[2955]), .Z(n18439) );
  IV U42562 ( .A(n18454), .Z(n40006) );
  XOR U42563 ( .A(n40014), .B(n40015), .Z(n18454) );
  XNOR U42564 ( .A(n18471), .B(n18452), .Z(n40015) );
  XNOR U42565 ( .A(q[1]), .B(DB[2946]), .Z(n18452) );
  XOR U42566 ( .A(n40016), .B(n18460), .Z(n18471) );
  XNOR U42567 ( .A(q[8]), .B(DB[2953]), .Z(n18460) );
  IV U42568 ( .A(n18459), .Z(n40016) );
  XNOR U42569 ( .A(n18457), .B(n40017), .Z(n18459) );
  XNOR U42570 ( .A(q[7]), .B(DB[2952]), .Z(n40017) );
  XNOR U42571 ( .A(q[6]), .B(DB[2951]), .Z(n18457) );
  IV U42572 ( .A(n18470), .Z(n40014) );
  XOR U42573 ( .A(n40018), .B(n40019), .Z(n18470) );
  XNOR U42574 ( .A(n18466), .B(n18468), .Z(n40019) );
  XNOR U42575 ( .A(q[2]), .B(DB[2947]), .Z(n18468) );
  XNOR U42576 ( .A(q[5]), .B(DB[2950]), .Z(n18466) );
  IV U42577 ( .A(n18465), .Z(n40018) );
  XNOR U42578 ( .A(n18463), .B(n40020), .Z(n18465) );
  XNOR U42579 ( .A(q[4]), .B(DB[2949]), .Z(n40020) );
  XNOR U42580 ( .A(q[3]), .B(DB[2948]), .Z(n18463) );
  XOR U42581 ( .A(n40021), .B(n18232), .Z(n18083) );
  XOR U42582 ( .A(n40022), .B(n18208), .Z(n18232) );
  XOR U42583 ( .A(n40023), .B(n18200), .Z(n18208) );
  XOR U42584 ( .A(n40024), .B(n18189), .Z(n18200) );
  XNOR U42585 ( .A(q[30]), .B(DB[3006]), .Z(n18189) );
  IV U42586 ( .A(n18188), .Z(n40024) );
  XNOR U42587 ( .A(n18186), .B(n40025), .Z(n18188) );
  XNOR U42588 ( .A(q[29]), .B(DB[3005]), .Z(n40025) );
  XNOR U42589 ( .A(q[28]), .B(DB[3004]), .Z(n18186) );
  IV U42590 ( .A(n18199), .Z(n40023) );
  XOR U42591 ( .A(n40026), .B(n40027), .Z(n18199) );
  XNOR U42592 ( .A(n18195), .B(n18197), .Z(n40027) );
  XNOR U42593 ( .A(q[24]), .B(DB[3000]), .Z(n18197) );
  XNOR U42594 ( .A(q[27]), .B(DB[3003]), .Z(n18195) );
  IV U42595 ( .A(n18194), .Z(n40026) );
  XNOR U42596 ( .A(n18192), .B(n40028), .Z(n18194) );
  XNOR U42597 ( .A(q[26]), .B(DB[3002]), .Z(n40028) );
  XNOR U42598 ( .A(q[25]), .B(DB[3001]), .Z(n18192) );
  IV U42599 ( .A(n18207), .Z(n40022) );
  XOR U42600 ( .A(n40029), .B(n40030), .Z(n18207) );
  XNOR U42601 ( .A(n18224), .B(n18205), .Z(n40030) );
  XNOR U42602 ( .A(q[16]), .B(DB[2992]), .Z(n18205) );
  XOR U42603 ( .A(n40031), .B(n18213), .Z(n18224) );
  XNOR U42604 ( .A(q[23]), .B(DB[2999]), .Z(n18213) );
  IV U42605 ( .A(n18212), .Z(n40031) );
  XNOR U42606 ( .A(n18210), .B(n40032), .Z(n18212) );
  XNOR U42607 ( .A(q[22]), .B(DB[2998]), .Z(n40032) );
  XNOR U42608 ( .A(q[21]), .B(DB[2997]), .Z(n18210) );
  IV U42609 ( .A(n18223), .Z(n40029) );
  XOR U42610 ( .A(n40033), .B(n40034), .Z(n18223) );
  XNOR U42611 ( .A(n18219), .B(n18221), .Z(n40034) );
  XNOR U42612 ( .A(q[17]), .B(DB[2993]), .Z(n18221) );
  XNOR U42613 ( .A(q[20]), .B(DB[2996]), .Z(n18219) );
  IV U42614 ( .A(n18218), .Z(n40033) );
  XNOR U42615 ( .A(n18216), .B(n40035), .Z(n18218) );
  XNOR U42616 ( .A(q[19]), .B(DB[2995]), .Z(n40035) );
  XNOR U42617 ( .A(q[18]), .B(DB[2994]), .Z(n18216) );
  IV U42618 ( .A(n18231), .Z(n40021) );
  XOR U42619 ( .A(n40036), .B(n40037), .Z(n18231) );
  XNOR U42620 ( .A(n18258), .B(n18229), .Z(n40037) );
  XNOR U42621 ( .A(q[0]), .B(DB[2976]), .Z(n18229) );
  XOR U42622 ( .A(n40038), .B(n18250), .Z(n18258) );
  XOR U42623 ( .A(n40039), .B(n18238), .Z(n18250) );
  XNOR U42624 ( .A(q[15]), .B(DB[2991]), .Z(n18238) );
  IV U42625 ( .A(n18237), .Z(n40039) );
  XNOR U42626 ( .A(n18235), .B(n40040), .Z(n18237) );
  XNOR U42627 ( .A(q[14]), .B(DB[2990]), .Z(n40040) );
  XNOR U42628 ( .A(q[13]), .B(DB[2989]), .Z(n18235) );
  IV U42629 ( .A(n18249), .Z(n40038) );
  XOR U42630 ( .A(n40041), .B(n40042), .Z(n18249) );
  XNOR U42631 ( .A(n18245), .B(n18247), .Z(n40042) );
  XNOR U42632 ( .A(q[9]), .B(DB[2985]), .Z(n18247) );
  XNOR U42633 ( .A(q[12]), .B(DB[2988]), .Z(n18245) );
  IV U42634 ( .A(n18244), .Z(n40041) );
  XNOR U42635 ( .A(n18242), .B(n40043), .Z(n18244) );
  XNOR U42636 ( .A(q[11]), .B(DB[2987]), .Z(n40043) );
  XNOR U42637 ( .A(q[10]), .B(DB[2986]), .Z(n18242) );
  IV U42638 ( .A(n18257), .Z(n40036) );
  XOR U42639 ( .A(n40044), .B(n40045), .Z(n18257) );
  XNOR U42640 ( .A(n18274), .B(n18255), .Z(n40045) );
  XNOR U42641 ( .A(q[1]), .B(DB[2977]), .Z(n18255) );
  XOR U42642 ( .A(n40046), .B(n18263), .Z(n18274) );
  XNOR U42643 ( .A(q[8]), .B(DB[2984]), .Z(n18263) );
  IV U42644 ( .A(n18262), .Z(n40046) );
  XNOR U42645 ( .A(n18260), .B(n40047), .Z(n18262) );
  XNOR U42646 ( .A(q[7]), .B(DB[2983]), .Z(n40047) );
  XNOR U42647 ( .A(q[6]), .B(DB[2982]), .Z(n18260) );
  IV U42648 ( .A(n18273), .Z(n40044) );
  XOR U42649 ( .A(n40048), .B(n40049), .Z(n18273) );
  XNOR U42650 ( .A(n18269), .B(n18271), .Z(n40049) );
  XNOR U42651 ( .A(q[2]), .B(DB[2978]), .Z(n18271) );
  XNOR U42652 ( .A(q[5]), .B(DB[2981]), .Z(n18269) );
  IV U42653 ( .A(n18268), .Z(n40048) );
  XNOR U42654 ( .A(n18266), .B(n40050), .Z(n18268) );
  XNOR U42655 ( .A(q[4]), .B(DB[2980]), .Z(n40050) );
  XNOR U42656 ( .A(q[3]), .B(DB[2979]), .Z(n18266) );
  XOR U42657 ( .A(n40051), .B(n18035), .Z(n17886) );
  XOR U42658 ( .A(n40052), .B(n18011), .Z(n18035) );
  XOR U42659 ( .A(n40053), .B(n18003), .Z(n18011) );
  XOR U42660 ( .A(n40054), .B(n17992), .Z(n18003) );
  XNOR U42661 ( .A(q[30]), .B(DB[3037]), .Z(n17992) );
  IV U42662 ( .A(n17991), .Z(n40054) );
  XNOR U42663 ( .A(n17989), .B(n40055), .Z(n17991) );
  XNOR U42664 ( .A(q[29]), .B(DB[3036]), .Z(n40055) );
  XNOR U42665 ( .A(q[28]), .B(DB[3035]), .Z(n17989) );
  IV U42666 ( .A(n18002), .Z(n40053) );
  XOR U42667 ( .A(n40056), .B(n40057), .Z(n18002) );
  XNOR U42668 ( .A(n17998), .B(n18000), .Z(n40057) );
  XNOR U42669 ( .A(q[24]), .B(DB[3031]), .Z(n18000) );
  XNOR U42670 ( .A(q[27]), .B(DB[3034]), .Z(n17998) );
  IV U42671 ( .A(n17997), .Z(n40056) );
  XNOR U42672 ( .A(n17995), .B(n40058), .Z(n17997) );
  XNOR U42673 ( .A(q[26]), .B(DB[3033]), .Z(n40058) );
  XNOR U42674 ( .A(q[25]), .B(DB[3032]), .Z(n17995) );
  IV U42675 ( .A(n18010), .Z(n40052) );
  XOR U42676 ( .A(n40059), .B(n40060), .Z(n18010) );
  XNOR U42677 ( .A(n18027), .B(n18008), .Z(n40060) );
  XNOR U42678 ( .A(q[16]), .B(DB[3023]), .Z(n18008) );
  XOR U42679 ( .A(n40061), .B(n18016), .Z(n18027) );
  XNOR U42680 ( .A(q[23]), .B(DB[3030]), .Z(n18016) );
  IV U42681 ( .A(n18015), .Z(n40061) );
  XNOR U42682 ( .A(n18013), .B(n40062), .Z(n18015) );
  XNOR U42683 ( .A(q[22]), .B(DB[3029]), .Z(n40062) );
  XNOR U42684 ( .A(q[21]), .B(DB[3028]), .Z(n18013) );
  IV U42685 ( .A(n18026), .Z(n40059) );
  XOR U42686 ( .A(n40063), .B(n40064), .Z(n18026) );
  XNOR U42687 ( .A(n18022), .B(n18024), .Z(n40064) );
  XNOR U42688 ( .A(q[17]), .B(DB[3024]), .Z(n18024) );
  XNOR U42689 ( .A(q[20]), .B(DB[3027]), .Z(n18022) );
  IV U42690 ( .A(n18021), .Z(n40063) );
  XNOR U42691 ( .A(n18019), .B(n40065), .Z(n18021) );
  XNOR U42692 ( .A(q[19]), .B(DB[3026]), .Z(n40065) );
  XNOR U42693 ( .A(q[18]), .B(DB[3025]), .Z(n18019) );
  IV U42694 ( .A(n18034), .Z(n40051) );
  XOR U42695 ( .A(n40066), .B(n40067), .Z(n18034) );
  XNOR U42696 ( .A(n18061), .B(n18032), .Z(n40067) );
  XNOR U42697 ( .A(q[0]), .B(DB[3007]), .Z(n18032) );
  XOR U42698 ( .A(n40068), .B(n18053), .Z(n18061) );
  XOR U42699 ( .A(n40069), .B(n18041), .Z(n18053) );
  XNOR U42700 ( .A(q[15]), .B(DB[3022]), .Z(n18041) );
  IV U42701 ( .A(n18040), .Z(n40069) );
  XNOR U42702 ( .A(n18038), .B(n40070), .Z(n18040) );
  XNOR U42703 ( .A(q[14]), .B(DB[3021]), .Z(n40070) );
  XNOR U42704 ( .A(q[13]), .B(DB[3020]), .Z(n18038) );
  IV U42705 ( .A(n18052), .Z(n40068) );
  XOR U42706 ( .A(n40071), .B(n40072), .Z(n18052) );
  XNOR U42707 ( .A(n18048), .B(n18050), .Z(n40072) );
  XNOR U42708 ( .A(q[9]), .B(DB[3016]), .Z(n18050) );
  XNOR U42709 ( .A(q[12]), .B(DB[3019]), .Z(n18048) );
  IV U42710 ( .A(n18047), .Z(n40071) );
  XNOR U42711 ( .A(n18045), .B(n40073), .Z(n18047) );
  XNOR U42712 ( .A(q[11]), .B(DB[3018]), .Z(n40073) );
  XNOR U42713 ( .A(q[10]), .B(DB[3017]), .Z(n18045) );
  IV U42714 ( .A(n18060), .Z(n40066) );
  XOR U42715 ( .A(n40074), .B(n40075), .Z(n18060) );
  XNOR U42716 ( .A(n18077), .B(n18058), .Z(n40075) );
  XNOR U42717 ( .A(q[1]), .B(DB[3008]), .Z(n18058) );
  XOR U42718 ( .A(n40076), .B(n18066), .Z(n18077) );
  XNOR U42719 ( .A(q[8]), .B(DB[3015]), .Z(n18066) );
  IV U42720 ( .A(n18065), .Z(n40076) );
  XNOR U42721 ( .A(n18063), .B(n40077), .Z(n18065) );
  XNOR U42722 ( .A(q[7]), .B(DB[3014]), .Z(n40077) );
  XNOR U42723 ( .A(q[6]), .B(DB[3013]), .Z(n18063) );
  IV U42724 ( .A(n18076), .Z(n40074) );
  XOR U42725 ( .A(n40078), .B(n40079), .Z(n18076) );
  XNOR U42726 ( .A(n18072), .B(n18074), .Z(n40079) );
  XNOR U42727 ( .A(q[2]), .B(DB[3009]), .Z(n18074) );
  XNOR U42728 ( .A(q[5]), .B(DB[3012]), .Z(n18072) );
  IV U42729 ( .A(n18071), .Z(n40078) );
  XNOR U42730 ( .A(n18069), .B(n40080), .Z(n18071) );
  XNOR U42731 ( .A(q[4]), .B(DB[3011]), .Z(n40080) );
  XNOR U42732 ( .A(q[3]), .B(DB[3010]), .Z(n18069) );
  XOR U42733 ( .A(n40081), .B(n17838), .Z(n17689) );
  XOR U42734 ( .A(n40082), .B(n17814), .Z(n17838) );
  XOR U42735 ( .A(n40083), .B(n17806), .Z(n17814) );
  XOR U42736 ( .A(n40084), .B(n17795), .Z(n17806) );
  XNOR U42737 ( .A(q[30]), .B(DB[3068]), .Z(n17795) );
  IV U42738 ( .A(n17794), .Z(n40084) );
  XNOR U42739 ( .A(n17792), .B(n40085), .Z(n17794) );
  XNOR U42740 ( .A(q[29]), .B(DB[3067]), .Z(n40085) );
  XNOR U42741 ( .A(q[28]), .B(DB[3066]), .Z(n17792) );
  IV U42742 ( .A(n17805), .Z(n40083) );
  XOR U42743 ( .A(n40086), .B(n40087), .Z(n17805) );
  XNOR U42744 ( .A(n17801), .B(n17803), .Z(n40087) );
  XNOR U42745 ( .A(q[24]), .B(DB[3062]), .Z(n17803) );
  XNOR U42746 ( .A(q[27]), .B(DB[3065]), .Z(n17801) );
  IV U42747 ( .A(n17800), .Z(n40086) );
  XNOR U42748 ( .A(n17798), .B(n40088), .Z(n17800) );
  XNOR U42749 ( .A(q[26]), .B(DB[3064]), .Z(n40088) );
  XNOR U42750 ( .A(q[25]), .B(DB[3063]), .Z(n17798) );
  IV U42751 ( .A(n17813), .Z(n40082) );
  XOR U42752 ( .A(n40089), .B(n40090), .Z(n17813) );
  XNOR U42753 ( .A(n17830), .B(n17811), .Z(n40090) );
  XNOR U42754 ( .A(q[16]), .B(DB[3054]), .Z(n17811) );
  XOR U42755 ( .A(n40091), .B(n17819), .Z(n17830) );
  XNOR U42756 ( .A(q[23]), .B(DB[3061]), .Z(n17819) );
  IV U42757 ( .A(n17818), .Z(n40091) );
  XNOR U42758 ( .A(n17816), .B(n40092), .Z(n17818) );
  XNOR U42759 ( .A(q[22]), .B(DB[3060]), .Z(n40092) );
  XNOR U42760 ( .A(q[21]), .B(DB[3059]), .Z(n17816) );
  IV U42761 ( .A(n17829), .Z(n40089) );
  XOR U42762 ( .A(n40093), .B(n40094), .Z(n17829) );
  XNOR U42763 ( .A(n17825), .B(n17827), .Z(n40094) );
  XNOR U42764 ( .A(q[17]), .B(DB[3055]), .Z(n17827) );
  XNOR U42765 ( .A(q[20]), .B(DB[3058]), .Z(n17825) );
  IV U42766 ( .A(n17824), .Z(n40093) );
  XNOR U42767 ( .A(n17822), .B(n40095), .Z(n17824) );
  XNOR U42768 ( .A(q[19]), .B(DB[3057]), .Z(n40095) );
  XNOR U42769 ( .A(q[18]), .B(DB[3056]), .Z(n17822) );
  IV U42770 ( .A(n17837), .Z(n40081) );
  XOR U42771 ( .A(n40096), .B(n40097), .Z(n17837) );
  XNOR U42772 ( .A(n17864), .B(n17835), .Z(n40097) );
  XNOR U42773 ( .A(q[0]), .B(DB[3038]), .Z(n17835) );
  XOR U42774 ( .A(n40098), .B(n17856), .Z(n17864) );
  XOR U42775 ( .A(n40099), .B(n17844), .Z(n17856) );
  XNOR U42776 ( .A(q[15]), .B(DB[3053]), .Z(n17844) );
  IV U42777 ( .A(n17843), .Z(n40099) );
  XNOR U42778 ( .A(n17841), .B(n40100), .Z(n17843) );
  XNOR U42779 ( .A(q[14]), .B(DB[3052]), .Z(n40100) );
  XNOR U42780 ( .A(q[13]), .B(DB[3051]), .Z(n17841) );
  IV U42781 ( .A(n17855), .Z(n40098) );
  XOR U42782 ( .A(n40101), .B(n40102), .Z(n17855) );
  XNOR U42783 ( .A(n17851), .B(n17853), .Z(n40102) );
  XNOR U42784 ( .A(q[9]), .B(DB[3047]), .Z(n17853) );
  XNOR U42785 ( .A(q[12]), .B(DB[3050]), .Z(n17851) );
  IV U42786 ( .A(n17850), .Z(n40101) );
  XNOR U42787 ( .A(n17848), .B(n40103), .Z(n17850) );
  XNOR U42788 ( .A(q[11]), .B(DB[3049]), .Z(n40103) );
  XNOR U42789 ( .A(q[10]), .B(DB[3048]), .Z(n17848) );
  IV U42790 ( .A(n17863), .Z(n40096) );
  XOR U42791 ( .A(n40104), .B(n40105), .Z(n17863) );
  XNOR U42792 ( .A(n17880), .B(n17861), .Z(n40105) );
  XNOR U42793 ( .A(q[1]), .B(DB[3039]), .Z(n17861) );
  XOR U42794 ( .A(n40106), .B(n17869), .Z(n17880) );
  XNOR U42795 ( .A(q[8]), .B(DB[3046]), .Z(n17869) );
  IV U42796 ( .A(n17868), .Z(n40106) );
  XNOR U42797 ( .A(n17866), .B(n40107), .Z(n17868) );
  XNOR U42798 ( .A(q[7]), .B(DB[3045]), .Z(n40107) );
  XNOR U42799 ( .A(q[6]), .B(DB[3044]), .Z(n17866) );
  IV U42800 ( .A(n17879), .Z(n40104) );
  XOR U42801 ( .A(n40108), .B(n40109), .Z(n17879) );
  XNOR U42802 ( .A(n17875), .B(n17877), .Z(n40109) );
  XNOR U42803 ( .A(q[2]), .B(DB[3040]), .Z(n17877) );
  XNOR U42804 ( .A(q[5]), .B(DB[3043]), .Z(n17875) );
  IV U42805 ( .A(n17874), .Z(n40108) );
  XNOR U42806 ( .A(n17872), .B(n40110), .Z(n17874) );
  XNOR U42807 ( .A(q[4]), .B(DB[3042]), .Z(n40110) );
  XNOR U42808 ( .A(q[3]), .B(DB[3041]), .Z(n17872) );
  XOR U42809 ( .A(n40111), .B(n17641), .Z(n17492) );
  XOR U42810 ( .A(n40112), .B(n17617), .Z(n17641) );
  XOR U42811 ( .A(n40113), .B(n17609), .Z(n17617) );
  XOR U42812 ( .A(n40114), .B(n17598), .Z(n17609) );
  XNOR U42813 ( .A(q[30]), .B(DB[3099]), .Z(n17598) );
  IV U42814 ( .A(n17597), .Z(n40114) );
  XNOR U42815 ( .A(n17595), .B(n40115), .Z(n17597) );
  XNOR U42816 ( .A(q[29]), .B(DB[3098]), .Z(n40115) );
  XNOR U42817 ( .A(q[28]), .B(DB[3097]), .Z(n17595) );
  IV U42818 ( .A(n17608), .Z(n40113) );
  XOR U42819 ( .A(n40116), .B(n40117), .Z(n17608) );
  XNOR U42820 ( .A(n17604), .B(n17606), .Z(n40117) );
  XNOR U42821 ( .A(q[24]), .B(DB[3093]), .Z(n17606) );
  XNOR U42822 ( .A(q[27]), .B(DB[3096]), .Z(n17604) );
  IV U42823 ( .A(n17603), .Z(n40116) );
  XNOR U42824 ( .A(n17601), .B(n40118), .Z(n17603) );
  XNOR U42825 ( .A(q[26]), .B(DB[3095]), .Z(n40118) );
  XNOR U42826 ( .A(q[25]), .B(DB[3094]), .Z(n17601) );
  IV U42827 ( .A(n17616), .Z(n40112) );
  XOR U42828 ( .A(n40119), .B(n40120), .Z(n17616) );
  XNOR U42829 ( .A(n17633), .B(n17614), .Z(n40120) );
  XNOR U42830 ( .A(q[16]), .B(DB[3085]), .Z(n17614) );
  XOR U42831 ( .A(n40121), .B(n17622), .Z(n17633) );
  XNOR U42832 ( .A(q[23]), .B(DB[3092]), .Z(n17622) );
  IV U42833 ( .A(n17621), .Z(n40121) );
  XNOR U42834 ( .A(n17619), .B(n40122), .Z(n17621) );
  XNOR U42835 ( .A(q[22]), .B(DB[3091]), .Z(n40122) );
  XNOR U42836 ( .A(q[21]), .B(DB[3090]), .Z(n17619) );
  IV U42837 ( .A(n17632), .Z(n40119) );
  XOR U42838 ( .A(n40123), .B(n40124), .Z(n17632) );
  XNOR U42839 ( .A(n17628), .B(n17630), .Z(n40124) );
  XNOR U42840 ( .A(q[17]), .B(DB[3086]), .Z(n17630) );
  XNOR U42841 ( .A(q[20]), .B(DB[3089]), .Z(n17628) );
  IV U42842 ( .A(n17627), .Z(n40123) );
  XNOR U42843 ( .A(n17625), .B(n40125), .Z(n17627) );
  XNOR U42844 ( .A(q[19]), .B(DB[3088]), .Z(n40125) );
  XNOR U42845 ( .A(q[18]), .B(DB[3087]), .Z(n17625) );
  IV U42846 ( .A(n17640), .Z(n40111) );
  XOR U42847 ( .A(n40126), .B(n40127), .Z(n17640) );
  XNOR U42848 ( .A(n17667), .B(n17638), .Z(n40127) );
  XNOR U42849 ( .A(q[0]), .B(DB[3069]), .Z(n17638) );
  XOR U42850 ( .A(n40128), .B(n17659), .Z(n17667) );
  XOR U42851 ( .A(n40129), .B(n17647), .Z(n17659) );
  XNOR U42852 ( .A(q[15]), .B(DB[3084]), .Z(n17647) );
  IV U42853 ( .A(n17646), .Z(n40129) );
  XNOR U42854 ( .A(n17644), .B(n40130), .Z(n17646) );
  XNOR U42855 ( .A(q[14]), .B(DB[3083]), .Z(n40130) );
  XNOR U42856 ( .A(q[13]), .B(DB[3082]), .Z(n17644) );
  IV U42857 ( .A(n17658), .Z(n40128) );
  XOR U42858 ( .A(n40131), .B(n40132), .Z(n17658) );
  XNOR U42859 ( .A(n17654), .B(n17656), .Z(n40132) );
  XNOR U42860 ( .A(q[9]), .B(DB[3078]), .Z(n17656) );
  XNOR U42861 ( .A(q[12]), .B(DB[3081]), .Z(n17654) );
  IV U42862 ( .A(n17653), .Z(n40131) );
  XNOR U42863 ( .A(n17651), .B(n40133), .Z(n17653) );
  XNOR U42864 ( .A(q[11]), .B(DB[3080]), .Z(n40133) );
  XNOR U42865 ( .A(q[10]), .B(DB[3079]), .Z(n17651) );
  IV U42866 ( .A(n17666), .Z(n40126) );
  XOR U42867 ( .A(n40134), .B(n40135), .Z(n17666) );
  XNOR U42868 ( .A(n17683), .B(n17664), .Z(n40135) );
  XNOR U42869 ( .A(q[1]), .B(DB[3070]), .Z(n17664) );
  XOR U42870 ( .A(n40136), .B(n17672), .Z(n17683) );
  XNOR U42871 ( .A(q[8]), .B(DB[3077]), .Z(n17672) );
  IV U42872 ( .A(n17671), .Z(n40136) );
  XNOR U42873 ( .A(n17669), .B(n40137), .Z(n17671) );
  XNOR U42874 ( .A(q[7]), .B(DB[3076]), .Z(n40137) );
  XNOR U42875 ( .A(q[6]), .B(DB[3075]), .Z(n17669) );
  IV U42876 ( .A(n17682), .Z(n40134) );
  XOR U42877 ( .A(n40138), .B(n40139), .Z(n17682) );
  XNOR U42878 ( .A(n17678), .B(n17680), .Z(n40139) );
  XNOR U42879 ( .A(q[2]), .B(DB[3071]), .Z(n17680) );
  XNOR U42880 ( .A(q[5]), .B(DB[3074]), .Z(n17678) );
  IV U42881 ( .A(n17677), .Z(n40138) );
  XNOR U42882 ( .A(n17675), .B(n40140), .Z(n17677) );
  XNOR U42883 ( .A(q[4]), .B(DB[3073]), .Z(n40140) );
  XNOR U42884 ( .A(q[3]), .B(DB[3072]), .Z(n17675) );
  XOR U42885 ( .A(n40141), .B(n17444), .Z(n17295) );
  XOR U42886 ( .A(n40142), .B(n17420), .Z(n17444) );
  XOR U42887 ( .A(n40143), .B(n17412), .Z(n17420) );
  XOR U42888 ( .A(n40144), .B(n17401), .Z(n17412) );
  XNOR U42889 ( .A(q[30]), .B(DB[3130]), .Z(n17401) );
  IV U42890 ( .A(n17400), .Z(n40144) );
  XNOR U42891 ( .A(n17398), .B(n40145), .Z(n17400) );
  XNOR U42892 ( .A(q[29]), .B(DB[3129]), .Z(n40145) );
  XNOR U42893 ( .A(q[28]), .B(DB[3128]), .Z(n17398) );
  IV U42894 ( .A(n17411), .Z(n40143) );
  XOR U42895 ( .A(n40146), .B(n40147), .Z(n17411) );
  XNOR U42896 ( .A(n17407), .B(n17409), .Z(n40147) );
  XNOR U42897 ( .A(q[24]), .B(DB[3124]), .Z(n17409) );
  XNOR U42898 ( .A(q[27]), .B(DB[3127]), .Z(n17407) );
  IV U42899 ( .A(n17406), .Z(n40146) );
  XNOR U42900 ( .A(n17404), .B(n40148), .Z(n17406) );
  XNOR U42901 ( .A(q[26]), .B(DB[3126]), .Z(n40148) );
  XNOR U42902 ( .A(q[25]), .B(DB[3125]), .Z(n17404) );
  IV U42903 ( .A(n17419), .Z(n40142) );
  XOR U42904 ( .A(n40149), .B(n40150), .Z(n17419) );
  XNOR U42905 ( .A(n17436), .B(n17417), .Z(n40150) );
  XNOR U42906 ( .A(q[16]), .B(DB[3116]), .Z(n17417) );
  XOR U42907 ( .A(n40151), .B(n17425), .Z(n17436) );
  XNOR U42908 ( .A(q[23]), .B(DB[3123]), .Z(n17425) );
  IV U42909 ( .A(n17424), .Z(n40151) );
  XNOR U42910 ( .A(n17422), .B(n40152), .Z(n17424) );
  XNOR U42911 ( .A(q[22]), .B(DB[3122]), .Z(n40152) );
  XNOR U42912 ( .A(q[21]), .B(DB[3121]), .Z(n17422) );
  IV U42913 ( .A(n17435), .Z(n40149) );
  XOR U42914 ( .A(n40153), .B(n40154), .Z(n17435) );
  XNOR U42915 ( .A(n17431), .B(n17433), .Z(n40154) );
  XNOR U42916 ( .A(q[17]), .B(DB[3117]), .Z(n17433) );
  XNOR U42917 ( .A(q[20]), .B(DB[3120]), .Z(n17431) );
  IV U42918 ( .A(n17430), .Z(n40153) );
  XNOR U42919 ( .A(n17428), .B(n40155), .Z(n17430) );
  XNOR U42920 ( .A(q[19]), .B(DB[3119]), .Z(n40155) );
  XNOR U42921 ( .A(q[18]), .B(DB[3118]), .Z(n17428) );
  IV U42922 ( .A(n17443), .Z(n40141) );
  XOR U42923 ( .A(n40156), .B(n40157), .Z(n17443) );
  XNOR U42924 ( .A(n17470), .B(n17441), .Z(n40157) );
  XNOR U42925 ( .A(q[0]), .B(DB[3100]), .Z(n17441) );
  XOR U42926 ( .A(n40158), .B(n17462), .Z(n17470) );
  XOR U42927 ( .A(n40159), .B(n17450), .Z(n17462) );
  XNOR U42928 ( .A(q[15]), .B(DB[3115]), .Z(n17450) );
  IV U42929 ( .A(n17449), .Z(n40159) );
  XNOR U42930 ( .A(n17447), .B(n40160), .Z(n17449) );
  XNOR U42931 ( .A(q[14]), .B(DB[3114]), .Z(n40160) );
  XNOR U42932 ( .A(q[13]), .B(DB[3113]), .Z(n17447) );
  IV U42933 ( .A(n17461), .Z(n40158) );
  XOR U42934 ( .A(n40161), .B(n40162), .Z(n17461) );
  XNOR U42935 ( .A(n17457), .B(n17459), .Z(n40162) );
  XNOR U42936 ( .A(q[9]), .B(DB[3109]), .Z(n17459) );
  XNOR U42937 ( .A(q[12]), .B(DB[3112]), .Z(n17457) );
  IV U42938 ( .A(n17456), .Z(n40161) );
  XNOR U42939 ( .A(n17454), .B(n40163), .Z(n17456) );
  XNOR U42940 ( .A(q[11]), .B(DB[3111]), .Z(n40163) );
  XNOR U42941 ( .A(q[10]), .B(DB[3110]), .Z(n17454) );
  IV U42942 ( .A(n17469), .Z(n40156) );
  XOR U42943 ( .A(n40164), .B(n40165), .Z(n17469) );
  XNOR U42944 ( .A(n17486), .B(n17467), .Z(n40165) );
  XNOR U42945 ( .A(q[1]), .B(DB[3101]), .Z(n17467) );
  XOR U42946 ( .A(n40166), .B(n17475), .Z(n17486) );
  XNOR U42947 ( .A(q[8]), .B(DB[3108]), .Z(n17475) );
  IV U42948 ( .A(n17474), .Z(n40166) );
  XNOR U42949 ( .A(n17472), .B(n40167), .Z(n17474) );
  XNOR U42950 ( .A(q[7]), .B(DB[3107]), .Z(n40167) );
  XNOR U42951 ( .A(q[6]), .B(DB[3106]), .Z(n17472) );
  IV U42952 ( .A(n17485), .Z(n40164) );
  XOR U42953 ( .A(n40168), .B(n40169), .Z(n17485) );
  XNOR U42954 ( .A(n17481), .B(n17483), .Z(n40169) );
  XNOR U42955 ( .A(q[2]), .B(DB[3102]), .Z(n17483) );
  XNOR U42956 ( .A(q[5]), .B(DB[3105]), .Z(n17481) );
  IV U42957 ( .A(n17480), .Z(n40168) );
  XNOR U42958 ( .A(n17478), .B(n40170), .Z(n17480) );
  XNOR U42959 ( .A(q[4]), .B(DB[3104]), .Z(n40170) );
  XNOR U42960 ( .A(q[3]), .B(DB[3103]), .Z(n17478) );
  XOR U42961 ( .A(n40171), .B(n17247), .Z(n17098) );
  XOR U42962 ( .A(n40172), .B(n17223), .Z(n17247) );
  XOR U42963 ( .A(n40173), .B(n17215), .Z(n17223) );
  XOR U42964 ( .A(n40174), .B(n17204), .Z(n17215) );
  XNOR U42965 ( .A(q[30]), .B(DB[3161]), .Z(n17204) );
  IV U42966 ( .A(n17203), .Z(n40174) );
  XNOR U42967 ( .A(n17201), .B(n40175), .Z(n17203) );
  XNOR U42968 ( .A(q[29]), .B(DB[3160]), .Z(n40175) );
  XNOR U42969 ( .A(q[28]), .B(DB[3159]), .Z(n17201) );
  IV U42970 ( .A(n17214), .Z(n40173) );
  XOR U42971 ( .A(n40176), .B(n40177), .Z(n17214) );
  XNOR U42972 ( .A(n17210), .B(n17212), .Z(n40177) );
  XNOR U42973 ( .A(q[24]), .B(DB[3155]), .Z(n17212) );
  XNOR U42974 ( .A(q[27]), .B(DB[3158]), .Z(n17210) );
  IV U42975 ( .A(n17209), .Z(n40176) );
  XNOR U42976 ( .A(n17207), .B(n40178), .Z(n17209) );
  XNOR U42977 ( .A(q[26]), .B(DB[3157]), .Z(n40178) );
  XNOR U42978 ( .A(q[25]), .B(DB[3156]), .Z(n17207) );
  IV U42979 ( .A(n17222), .Z(n40172) );
  XOR U42980 ( .A(n40179), .B(n40180), .Z(n17222) );
  XNOR U42981 ( .A(n17239), .B(n17220), .Z(n40180) );
  XNOR U42982 ( .A(q[16]), .B(DB[3147]), .Z(n17220) );
  XOR U42983 ( .A(n40181), .B(n17228), .Z(n17239) );
  XNOR U42984 ( .A(q[23]), .B(DB[3154]), .Z(n17228) );
  IV U42985 ( .A(n17227), .Z(n40181) );
  XNOR U42986 ( .A(n17225), .B(n40182), .Z(n17227) );
  XNOR U42987 ( .A(q[22]), .B(DB[3153]), .Z(n40182) );
  XNOR U42988 ( .A(q[21]), .B(DB[3152]), .Z(n17225) );
  IV U42989 ( .A(n17238), .Z(n40179) );
  XOR U42990 ( .A(n40183), .B(n40184), .Z(n17238) );
  XNOR U42991 ( .A(n17234), .B(n17236), .Z(n40184) );
  XNOR U42992 ( .A(q[17]), .B(DB[3148]), .Z(n17236) );
  XNOR U42993 ( .A(q[20]), .B(DB[3151]), .Z(n17234) );
  IV U42994 ( .A(n17233), .Z(n40183) );
  XNOR U42995 ( .A(n17231), .B(n40185), .Z(n17233) );
  XNOR U42996 ( .A(q[19]), .B(DB[3150]), .Z(n40185) );
  XNOR U42997 ( .A(q[18]), .B(DB[3149]), .Z(n17231) );
  IV U42998 ( .A(n17246), .Z(n40171) );
  XOR U42999 ( .A(n40186), .B(n40187), .Z(n17246) );
  XNOR U43000 ( .A(n17273), .B(n17244), .Z(n40187) );
  XNOR U43001 ( .A(q[0]), .B(DB[3131]), .Z(n17244) );
  XOR U43002 ( .A(n40188), .B(n17265), .Z(n17273) );
  XOR U43003 ( .A(n40189), .B(n17253), .Z(n17265) );
  XNOR U43004 ( .A(q[15]), .B(DB[3146]), .Z(n17253) );
  IV U43005 ( .A(n17252), .Z(n40189) );
  XNOR U43006 ( .A(n17250), .B(n40190), .Z(n17252) );
  XNOR U43007 ( .A(q[14]), .B(DB[3145]), .Z(n40190) );
  XNOR U43008 ( .A(q[13]), .B(DB[3144]), .Z(n17250) );
  IV U43009 ( .A(n17264), .Z(n40188) );
  XOR U43010 ( .A(n40191), .B(n40192), .Z(n17264) );
  XNOR U43011 ( .A(n17260), .B(n17262), .Z(n40192) );
  XNOR U43012 ( .A(q[9]), .B(DB[3140]), .Z(n17262) );
  XNOR U43013 ( .A(q[12]), .B(DB[3143]), .Z(n17260) );
  IV U43014 ( .A(n17259), .Z(n40191) );
  XNOR U43015 ( .A(n17257), .B(n40193), .Z(n17259) );
  XNOR U43016 ( .A(q[11]), .B(DB[3142]), .Z(n40193) );
  XNOR U43017 ( .A(q[10]), .B(DB[3141]), .Z(n17257) );
  IV U43018 ( .A(n17272), .Z(n40186) );
  XOR U43019 ( .A(n40194), .B(n40195), .Z(n17272) );
  XNOR U43020 ( .A(n17289), .B(n17270), .Z(n40195) );
  XNOR U43021 ( .A(q[1]), .B(DB[3132]), .Z(n17270) );
  XOR U43022 ( .A(n40196), .B(n17278), .Z(n17289) );
  XNOR U43023 ( .A(q[8]), .B(DB[3139]), .Z(n17278) );
  IV U43024 ( .A(n17277), .Z(n40196) );
  XNOR U43025 ( .A(n17275), .B(n40197), .Z(n17277) );
  XNOR U43026 ( .A(q[7]), .B(DB[3138]), .Z(n40197) );
  XNOR U43027 ( .A(q[6]), .B(DB[3137]), .Z(n17275) );
  IV U43028 ( .A(n17288), .Z(n40194) );
  XOR U43029 ( .A(n40198), .B(n40199), .Z(n17288) );
  XNOR U43030 ( .A(n17284), .B(n17286), .Z(n40199) );
  XNOR U43031 ( .A(q[2]), .B(DB[3133]), .Z(n17286) );
  XNOR U43032 ( .A(q[5]), .B(DB[3136]), .Z(n17284) );
  IV U43033 ( .A(n17283), .Z(n40198) );
  XNOR U43034 ( .A(n17281), .B(n40200), .Z(n17283) );
  XNOR U43035 ( .A(q[4]), .B(DB[3135]), .Z(n40200) );
  XNOR U43036 ( .A(q[3]), .B(DB[3134]), .Z(n17281) );
  XOR U43037 ( .A(n40201), .B(n17050), .Z(n16901) );
  XOR U43038 ( .A(n40202), .B(n17026), .Z(n17050) );
  XOR U43039 ( .A(n40203), .B(n17018), .Z(n17026) );
  XOR U43040 ( .A(n40204), .B(n17007), .Z(n17018) );
  XNOR U43041 ( .A(q[30]), .B(DB[3192]), .Z(n17007) );
  IV U43042 ( .A(n17006), .Z(n40204) );
  XNOR U43043 ( .A(n17004), .B(n40205), .Z(n17006) );
  XNOR U43044 ( .A(q[29]), .B(DB[3191]), .Z(n40205) );
  XNOR U43045 ( .A(q[28]), .B(DB[3190]), .Z(n17004) );
  IV U43046 ( .A(n17017), .Z(n40203) );
  XOR U43047 ( .A(n40206), .B(n40207), .Z(n17017) );
  XNOR U43048 ( .A(n17013), .B(n17015), .Z(n40207) );
  XNOR U43049 ( .A(q[24]), .B(DB[3186]), .Z(n17015) );
  XNOR U43050 ( .A(q[27]), .B(DB[3189]), .Z(n17013) );
  IV U43051 ( .A(n17012), .Z(n40206) );
  XNOR U43052 ( .A(n17010), .B(n40208), .Z(n17012) );
  XNOR U43053 ( .A(q[26]), .B(DB[3188]), .Z(n40208) );
  XNOR U43054 ( .A(q[25]), .B(DB[3187]), .Z(n17010) );
  IV U43055 ( .A(n17025), .Z(n40202) );
  XOR U43056 ( .A(n40209), .B(n40210), .Z(n17025) );
  XNOR U43057 ( .A(n17042), .B(n17023), .Z(n40210) );
  XNOR U43058 ( .A(q[16]), .B(DB[3178]), .Z(n17023) );
  XOR U43059 ( .A(n40211), .B(n17031), .Z(n17042) );
  XNOR U43060 ( .A(q[23]), .B(DB[3185]), .Z(n17031) );
  IV U43061 ( .A(n17030), .Z(n40211) );
  XNOR U43062 ( .A(n17028), .B(n40212), .Z(n17030) );
  XNOR U43063 ( .A(q[22]), .B(DB[3184]), .Z(n40212) );
  XNOR U43064 ( .A(q[21]), .B(DB[3183]), .Z(n17028) );
  IV U43065 ( .A(n17041), .Z(n40209) );
  XOR U43066 ( .A(n40213), .B(n40214), .Z(n17041) );
  XNOR U43067 ( .A(n17037), .B(n17039), .Z(n40214) );
  XNOR U43068 ( .A(q[17]), .B(DB[3179]), .Z(n17039) );
  XNOR U43069 ( .A(q[20]), .B(DB[3182]), .Z(n17037) );
  IV U43070 ( .A(n17036), .Z(n40213) );
  XNOR U43071 ( .A(n17034), .B(n40215), .Z(n17036) );
  XNOR U43072 ( .A(q[19]), .B(DB[3181]), .Z(n40215) );
  XNOR U43073 ( .A(q[18]), .B(DB[3180]), .Z(n17034) );
  IV U43074 ( .A(n17049), .Z(n40201) );
  XOR U43075 ( .A(n40216), .B(n40217), .Z(n17049) );
  XNOR U43076 ( .A(n17076), .B(n17047), .Z(n40217) );
  XNOR U43077 ( .A(q[0]), .B(DB[3162]), .Z(n17047) );
  XOR U43078 ( .A(n40218), .B(n17068), .Z(n17076) );
  XOR U43079 ( .A(n40219), .B(n17056), .Z(n17068) );
  XNOR U43080 ( .A(q[15]), .B(DB[3177]), .Z(n17056) );
  IV U43081 ( .A(n17055), .Z(n40219) );
  XNOR U43082 ( .A(n17053), .B(n40220), .Z(n17055) );
  XNOR U43083 ( .A(q[14]), .B(DB[3176]), .Z(n40220) );
  XNOR U43084 ( .A(q[13]), .B(DB[3175]), .Z(n17053) );
  IV U43085 ( .A(n17067), .Z(n40218) );
  XOR U43086 ( .A(n40221), .B(n40222), .Z(n17067) );
  XNOR U43087 ( .A(n17063), .B(n17065), .Z(n40222) );
  XNOR U43088 ( .A(q[9]), .B(DB[3171]), .Z(n17065) );
  XNOR U43089 ( .A(q[12]), .B(DB[3174]), .Z(n17063) );
  IV U43090 ( .A(n17062), .Z(n40221) );
  XNOR U43091 ( .A(n17060), .B(n40223), .Z(n17062) );
  XNOR U43092 ( .A(q[11]), .B(DB[3173]), .Z(n40223) );
  XNOR U43093 ( .A(q[10]), .B(DB[3172]), .Z(n17060) );
  IV U43094 ( .A(n17075), .Z(n40216) );
  XOR U43095 ( .A(n40224), .B(n40225), .Z(n17075) );
  XNOR U43096 ( .A(n17092), .B(n17073), .Z(n40225) );
  XNOR U43097 ( .A(q[1]), .B(DB[3163]), .Z(n17073) );
  XOR U43098 ( .A(n40226), .B(n17081), .Z(n17092) );
  XNOR U43099 ( .A(q[8]), .B(DB[3170]), .Z(n17081) );
  IV U43100 ( .A(n17080), .Z(n40226) );
  XNOR U43101 ( .A(n17078), .B(n40227), .Z(n17080) );
  XNOR U43102 ( .A(q[7]), .B(DB[3169]), .Z(n40227) );
  XNOR U43103 ( .A(q[6]), .B(DB[3168]), .Z(n17078) );
  IV U43104 ( .A(n17091), .Z(n40224) );
  XOR U43105 ( .A(n40228), .B(n40229), .Z(n17091) );
  XNOR U43106 ( .A(n17087), .B(n17089), .Z(n40229) );
  XNOR U43107 ( .A(q[2]), .B(DB[3164]), .Z(n17089) );
  XNOR U43108 ( .A(q[5]), .B(DB[3167]), .Z(n17087) );
  IV U43109 ( .A(n17086), .Z(n40228) );
  XNOR U43110 ( .A(n17084), .B(n40230), .Z(n17086) );
  XNOR U43111 ( .A(q[4]), .B(DB[3166]), .Z(n40230) );
  XNOR U43112 ( .A(q[3]), .B(DB[3165]), .Z(n17084) );
  XOR U43113 ( .A(n40231), .B(n16853), .Z(n16704) );
  XOR U43114 ( .A(n40232), .B(n16829), .Z(n16853) );
  XOR U43115 ( .A(n40233), .B(n16821), .Z(n16829) );
  XOR U43116 ( .A(n40234), .B(n16810), .Z(n16821) );
  XNOR U43117 ( .A(q[30]), .B(DB[3223]), .Z(n16810) );
  IV U43118 ( .A(n16809), .Z(n40234) );
  XNOR U43119 ( .A(n16807), .B(n40235), .Z(n16809) );
  XNOR U43120 ( .A(q[29]), .B(DB[3222]), .Z(n40235) );
  XNOR U43121 ( .A(q[28]), .B(DB[3221]), .Z(n16807) );
  IV U43122 ( .A(n16820), .Z(n40233) );
  XOR U43123 ( .A(n40236), .B(n40237), .Z(n16820) );
  XNOR U43124 ( .A(n16816), .B(n16818), .Z(n40237) );
  XNOR U43125 ( .A(q[24]), .B(DB[3217]), .Z(n16818) );
  XNOR U43126 ( .A(q[27]), .B(DB[3220]), .Z(n16816) );
  IV U43127 ( .A(n16815), .Z(n40236) );
  XNOR U43128 ( .A(n16813), .B(n40238), .Z(n16815) );
  XNOR U43129 ( .A(q[26]), .B(DB[3219]), .Z(n40238) );
  XNOR U43130 ( .A(q[25]), .B(DB[3218]), .Z(n16813) );
  IV U43131 ( .A(n16828), .Z(n40232) );
  XOR U43132 ( .A(n40239), .B(n40240), .Z(n16828) );
  XNOR U43133 ( .A(n16845), .B(n16826), .Z(n40240) );
  XNOR U43134 ( .A(q[16]), .B(DB[3209]), .Z(n16826) );
  XOR U43135 ( .A(n40241), .B(n16834), .Z(n16845) );
  XNOR U43136 ( .A(q[23]), .B(DB[3216]), .Z(n16834) );
  IV U43137 ( .A(n16833), .Z(n40241) );
  XNOR U43138 ( .A(n16831), .B(n40242), .Z(n16833) );
  XNOR U43139 ( .A(q[22]), .B(DB[3215]), .Z(n40242) );
  XNOR U43140 ( .A(q[21]), .B(DB[3214]), .Z(n16831) );
  IV U43141 ( .A(n16844), .Z(n40239) );
  XOR U43142 ( .A(n40243), .B(n40244), .Z(n16844) );
  XNOR U43143 ( .A(n16840), .B(n16842), .Z(n40244) );
  XNOR U43144 ( .A(q[17]), .B(DB[3210]), .Z(n16842) );
  XNOR U43145 ( .A(q[20]), .B(DB[3213]), .Z(n16840) );
  IV U43146 ( .A(n16839), .Z(n40243) );
  XNOR U43147 ( .A(n16837), .B(n40245), .Z(n16839) );
  XNOR U43148 ( .A(q[19]), .B(DB[3212]), .Z(n40245) );
  XNOR U43149 ( .A(q[18]), .B(DB[3211]), .Z(n16837) );
  IV U43150 ( .A(n16852), .Z(n40231) );
  XOR U43151 ( .A(n40246), .B(n40247), .Z(n16852) );
  XNOR U43152 ( .A(n16879), .B(n16850), .Z(n40247) );
  XNOR U43153 ( .A(q[0]), .B(DB[3193]), .Z(n16850) );
  XOR U43154 ( .A(n40248), .B(n16871), .Z(n16879) );
  XOR U43155 ( .A(n40249), .B(n16859), .Z(n16871) );
  XNOR U43156 ( .A(q[15]), .B(DB[3208]), .Z(n16859) );
  IV U43157 ( .A(n16858), .Z(n40249) );
  XNOR U43158 ( .A(n16856), .B(n40250), .Z(n16858) );
  XNOR U43159 ( .A(q[14]), .B(DB[3207]), .Z(n40250) );
  XNOR U43160 ( .A(q[13]), .B(DB[3206]), .Z(n16856) );
  IV U43161 ( .A(n16870), .Z(n40248) );
  XOR U43162 ( .A(n40251), .B(n40252), .Z(n16870) );
  XNOR U43163 ( .A(n16866), .B(n16868), .Z(n40252) );
  XNOR U43164 ( .A(q[9]), .B(DB[3202]), .Z(n16868) );
  XNOR U43165 ( .A(q[12]), .B(DB[3205]), .Z(n16866) );
  IV U43166 ( .A(n16865), .Z(n40251) );
  XNOR U43167 ( .A(n16863), .B(n40253), .Z(n16865) );
  XNOR U43168 ( .A(q[11]), .B(DB[3204]), .Z(n40253) );
  XNOR U43169 ( .A(q[10]), .B(DB[3203]), .Z(n16863) );
  IV U43170 ( .A(n16878), .Z(n40246) );
  XOR U43171 ( .A(n40254), .B(n40255), .Z(n16878) );
  XNOR U43172 ( .A(n16895), .B(n16876), .Z(n40255) );
  XNOR U43173 ( .A(q[1]), .B(DB[3194]), .Z(n16876) );
  XOR U43174 ( .A(n40256), .B(n16884), .Z(n16895) );
  XNOR U43175 ( .A(q[8]), .B(DB[3201]), .Z(n16884) );
  IV U43176 ( .A(n16883), .Z(n40256) );
  XNOR U43177 ( .A(n16881), .B(n40257), .Z(n16883) );
  XNOR U43178 ( .A(q[7]), .B(DB[3200]), .Z(n40257) );
  XNOR U43179 ( .A(q[6]), .B(DB[3199]), .Z(n16881) );
  IV U43180 ( .A(n16894), .Z(n40254) );
  XOR U43181 ( .A(n40258), .B(n40259), .Z(n16894) );
  XNOR U43182 ( .A(n16890), .B(n16892), .Z(n40259) );
  XNOR U43183 ( .A(q[2]), .B(DB[3195]), .Z(n16892) );
  XNOR U43184 ( .A(q[5]), .B(DB[3198]), .Z(n16890) );
  IV U43185 ( .A(n16889), .Z(n40258) );
  XNOR U43186 ( .A(n16887), .B(n40260), .Z(n16889) );
  XNOR U43187 ( .A(q[4]), .B(DB[3197]), .Z(n40260) );
  XNOR U43188 ( .A(q[3]), .B(DB[3196]), .Z(n16887) );
  XOR U43189 ( .A(n40261), .B(n16656), .Z(n16507) );
  XOR U43190 ( .A(n40262), .B(n16632), .Z(n16656) );
  XOR U43191 ( .A(n40263), .B(n16624), .Z(n16632) );
  XOR U43192 ( .A(n40264), .B(n16613), .Z(n16624) );
  XNOR U43193 ( .A(q[30]), .B(DB[3254]), .Z(n16613) );
  IV U43194 ( .A(n16612), .Z(n40264) );
  XNOR U43195 ( .A(n16610), .B(n40265), .Z(n16612) );
  XNOR U43196 ( .A(q[29]), .B(DB[3253]), .Z(n40265) );
  XNOR U43197 ( .A(q[28]), .B(DB[3252]), .Z(n16610) );
  IV U43198 ( .A(n16623), .Z(n40263) );
  XOR U43199 ( .A(n40266), .B(n40267), .Z(n16623) );
  XNOR U43200 ( .A(n16619), .B(n16621), .Z(n40267) );
  XNOR U43201 ( .A(q[24]), .B(DB[3248]), .Z(n16621) );
  XNOR U43202 ( .A(q[27]), .B(DB[3251]), .Z(n16619) );
  IV U43203 ( .A(n16618), .Z(n40266) );
  XNOR U43204 ( .A(n16616), .B(n40268), .Z(n16618) );
  XNOR U43205 ( .A(q[26]), .B(DB[3250]), .Z(n40268) );
  XNOR U43206 ( .A(q[25]), .B(DB[3249]), .Z(n16616) );
  IV U43207 ( .A(n16631), .Z(n40262) );
  XOR U43208 ( .A(n40269), .B(n40270), .Z(n16631) );
  XNOR U43209 ( .A(n16648), .B(n16629), .Z(n40270) );
  XNOR U43210 ( .A(q[16]), .B(DB[3240]), .Z(n16629) );
  XOR U43211 ( .A(n40271), .B(n16637), .Z(n16648) );
  XNOR U43212 ( .A(q[23]), .B(DB[3247]), .Z(n16637) );
  IV U43213 ( .A(n16636), .Z(n40271) );
  XNOR U43214 ( .A(n16634), .B(n40272), .Z(n16636) );
  XNOR U43215 ( .A(q[22]), .B(DB[3246]), .Z(n40272) );
  XNOR U43216 ( .A(q[21]), .B(DB[3245]), .Z(n16634) );
  IV U43217 ( .A(n16647), .Z(n40269) );
  XOR U43218 ( .A(n40273), .B(n40274), .Z(n16647) );
  XNOR U43219 ( .A(n16643), .B(n16645), .Z(n40274) );
  XNOR U43220 ( .A(q[17]), .B(DB[3241]), .Z(n16645) );
  XNOR U43221 ( .A(q[20]), .B(DB[3244]), .Z(n16643) );
  IV U43222 ( .A(n16642), .Z(n40273) );
  XNOR U43223 ( .A(n16640), .B(n40275), .Z(n16642) );
  XNOR U43224 ( .A(q[19]), .B(DB[3243]), .Z(n40275) );
  XNOR U43225 ( .A(q[18]), .B(DB[3242]), .Z(n16640) );
  IV U43226 ( .A(n16655), .Z(n40261) );
  XOR U43227 ( .A(n40276), .B(n40277), .Z(n16655) );
  XNOR U43228 ( .A(n16682), .B(n16653), .Z(n40277) );
  XNOR U43229 ( .A(q[0]), .B(DB[3224]), .Z(n16653) );
  XOR U43230 ( .A(n40278), .B(n16674), .Z(n16682) );
  XOR U43231 ( .A(n40279), .B(n16662), .Z(n16674) );
  XNOR U43232 ( .A(q[15]), .B(DB[3239]), .Z(n16662) );
  IV U43233 ( .A(n16661), .Z(n40279) );
  XNOR U43234 ( .A(n16659), .B(n40280), .Z(n16661) );
  XNOR U43235 ( .A(q[14]), .B(DB[3238]), .Z(n40280) );
  XNOR U43236 ( .A(q[13]), .B(DB[3237]), .Z(n16659) );
  IV U43237 ( .A(n16673), .Z(n40278) );
  XOR U43238 ( .A(n40281), .B(n40282), .Z(n16673) );
  XNOR U43239 ( .A(n16669), .B(n16671), .Z(n40282) );
  XNOR U43240 ( .A(q[9]), .B(DB[3233]), .Z(n16671) );
  XNOR U43241 ( .A(q[12]), .B(DB[3236]), .Z(n16669) );
  IV U43242 ( .A(n16668), .Z(n40281) );
  XNOR U43243 ( .A(n16666), .B(n40283), .Z(n16668) );
  XNOR U43244 ( .A(q[11]), .B(DB[3235]), .Z(n40283) );
  XNOR U43245 ( .A(q[10]), .B(DB[3234]), .Z(n16666) );
  IV U43246 ( .A(n16681), .Z(n40276) );
  XOR U43247 ( .A(n40284), .B(n40285), .Z(n16681) );
  XNOR U43248 ( .A(n16698), .B(n16679), .Z(n40285) );
  XNOR U43249 ( .A(q[1]), .B(DB[3225]), .Z(n16679) );
  XOR U43250 ( .A(n40286), .B(n16687), .Z(n16698) );
  XNOR U43251 ( .A(q[8]), .B(DB[3232]), .Z(n16687) );
  IV U43252 ( .A(n16686), .Z(n40286) );
  XNOR U43253 ( .A(n16684), .B(n40287), .Z(n16686) );
  XNOR U43254 ( .A(q[7]), .B(DB[3231]), .Z(n40287) );
  XNOR U43255 ( .A(q[6]), .B(DB[3230]), .Z(n16684) );
  IV U43256 ( .A(n16697), .Z(n40284) );
  XOR U43257 ( .A(n40288), .B(n40289), .Z(n16697) );
  XNOR U43258 ( .A(n16693), .B(n16695), .Z(n40289) );
  XNOR U43259 ( .A(q[2]), .B(DB[3226]), .Z(n16695) );
  XNOR U43260 ( .A(q[5]), .B(DB[3229]), .Z(n16693) );
  IV U43261 ( .A(n16692), .Z(n40288) );
  XNOR U43262 ( .A(n16690), .B(n40290), .Z(n16692) );
  XNOR U43263 ( .A(q[4]), .B(DB[3228]), .Z(n40290) );
  XNOR U43264 ( .A(q[3]), .B(DB[3227]), .Z(n16690) );
  XOR U43265 ( .A(n40291), .B(n16459), .Z(n16310) );
  XOR U43266 ( .A(n40292), .B(n16435), .Z(n16459) );
  XOR U43267 ( .A(n40293), .B(n16427), .Z(n16435) );
  XOR U43268 ( .A(n40294), .B(n16416), .Z(n16427) );
  XNOR U43269 ( .A(q[30]), .B(DB[3285]), .Z(n16416) );
  IV U43270 ( .A(n16415), .Z(n40294) );
  XNOR U43271 ( .A(n16413), .B(n40295), .Z(n16415) );
  XNOR U43272 ( .A(q[29]), .B(DB[3284]), .Z(n40295) );
  XNOR U43273 ( .A(q[28]), .B(DB[3283]), .Z(n16413) );
  IV U43274 ( .A(n16426), .Z(n40293) );
  XOR U43275 ( .A(n40296), .B(n40297), .Z(n16426) );
  XNOR U43276 ( .A(n16422), .B(n16424), .Z(n40297) );
  XNOR U43277 ( .A(q[24]), .B(DB[3279]), .Z(n16424) );
  XNOR U43278 ( .A(q[27]), .B(DB[3282]), .Z(n16422) );
  IV U43279 ( .A(n16421), .Z(n40296) );
  XNOR U43280 ( .A(n16419), .B(n40298), .Z(n16421) );
  XNOR U43281 ( .A(q[26]), .B(DB[3281]), .Z(n40298) );
  XNOR U43282 ( .A(q[25]), .B(DB[3280]), .Z(n16419) );
  IV U43283 ( .A(n16434), .Z(n40292) );
  XOR U43284 ( .A(n40299), .B(n40300), .Z(n16434) );
  XNOR U43285 ( .A(n16451), .B(n16432), .Z(n40300) );
  XNOR U43286 ( .A(q[16]), .B(DB[3271]), .Z(n16432) );
  XOR U43287 ( .A(n40301), .B(n16440), .Z(n16451) );
  XNOR U43288 ( .A(q[23]), .B(DB[3278]), .Z(n16440) );
  IV U43289 ( .A(n16439), .Z(n40301) );
  XNOR U43290 ( .A(n16437), .B(n40302), .Z(n16439) );
  XNOR U43291 ( .A(q[22]), .B(DB[3277]), .Z(n40302) );
  XNOR U43292 ( .A(q[21]), .B(DB[3276]), .Z(n16437) );
  IV U43293 ( .A(n16450), .Z(n40299) );
  XOR U43294 ( .A(n40303), .B(n40304), .Z(n16450) );
  XNOR U43295 ( .A(n16446), .B(n16448), .Z(n40304) );
  XNOR U43296 ( .A(q[17]), .B(DB[3272]), .Z(n16448) );
  XNOR U43297 ( .A(q[20]), .B(DB[3275]), .Z(n16446) );
  IV U43298 ( .A(n16445), .Z(n40303) );
  XNOR U43299 ( .A(n16443), .B(n40305), .Z(n16445) );
  XNOR U43300 ( .A(q[19]), .B(DB[3274]), .Z(n40305) );
  XNOR U43301 ( .A(q[18]), .B(DB[3273]), .Z(n16443) );
  IV U43302 ( .A(n16458), .Z(n40291) );
  XOR U43303 ( .A(n40306), .B(n40307), .Z(n16458) );
  XNOR U43304 ( .A(n16485), .B(n16456), .Z(n40307) );
  XNOR U43305 ( .A(q[0]), .B(DB[3255]), .Z(n16456) );
  XOR U43306 ( .A(n40308), .B(n16477), .Z(n16485) );
  XOR U43307 ( .A(n40309), .B(n16465), .Z(n16477) );
  XNOR U43308 ( .A(q[15]), .B(DB[3270]), .Z(n16465) );
  IV U43309 ( .A(n16464), .Z(n40309) );
  XNOR U43310 ( .A(n16462), .B(n40310), .Z(n16464) );
  XNOR U43311 ( .A(q[14]), .B(DB[3269]), .Z(n40310) );
  XNOR U43312 ( .A(q[13]), .B(DB[3268]), .Z(n16462) );
  IV U43313 ( .A(n16476), .Z(n40308) );
  XOR U43314 ( .A(n40311), .B(n40312), .Z(n16476) );
  XNOR U43315 ( .A(n16472), .B(n16474), .Z(n40312) );
  XNOR U43316 ( .A(q[9]), .B(DB[3264]), .Z(n16474) );
  XNOR U43317 ( .A(q[12]), .B(DB[3267]), .Z(n16472) );
  IV U43318 ( .A(n16471), .Z(n40311) );
  XNOR U43319 ( .A(n16469), .B(n40313), .Z(n16471) );
  XNOR U43320 ( .A(q[11]), .B(DB[3266]), .Z(n40313) );
  XNOR U43321 ( .A(q[10]), .B(DB[3265]), .Z(n16469) );
  IV U43322 ( .A(n16484), .Z(n40306) );
  XOR U43323 ( .A(n40314), .B(n40315), .Z(n16484) );
  XNOR U43324 ( .A(n16501), .B(n16482), .Z(n40315) );
  XNOR U43325 ( .A(q[1]), .B(DB[3256]), .Z(n16482) );
  XOR U43326 ( .A(n40316), .B(n16490), .Z(n16501) );
  XNOR U43327 ( .A(q[8]), .B(DB[3263]), .Z(n16490) );
  IV U43328 ( .A(n16489), .Z(n40316) );
  XNOR U43329 ( .A(n16487), .B(n40317), .Z(n16489) );
  XNOR U43330 ( .A(q[7]), .B(DB[3262]), .Z(n40317) );
  XNOR U43331 ( .A(q[6]), .B(DB[3261]), .Z(n16487) );
  IV U43332 ( .A(n16500), .Z(n40314) );
  XOR U43333 ( .A(n40318), .B(n40319), .Z(n16500) );
  XNOR U43334 ( .A(n16496), .B(n16498), .Z(n40319) );
  XNOR U43335 ( .A(q[2]), .B(DB[3257]), .Z(n16498) );
  XNOR U43336 ( .A(q[5]), .B(DB[3260]), .Z(n16496) );
  IV U43337 ( .A(n16495), .Z(n40318) );
  XNOR U43338 ( .A(n16493), .B(n40320), .Z(n16495) );
  XNOR U43339 ( .A(q[4]), .B(DB[3259]), .Z(n40320) );
  XNOR U43340 ( .A(q[3]), .B(DB[3258]), .Z(n16493) );
  XOR U43341 ( .A(n40321), .B(n16262), .Z(n16113) );
  XOR U43342 ( .A(n40322), .B(n16238), .Z(n16262) );
  XOR U43343 ( .A(n40323), .B(n16230), .Z(n16238) );
  XOR U43344 ( .A(n40324), .B(n16219), .Z(n16230) );
  XNOR U43345 ( .A(q[30]), .B(DB[3316]), .Z(n16219) );
  IV U43346 ( .A(n16218), .Z(n40324) );
  XNOR U43347 ( .A(n16216), .B(n40325), .Z(n16218) );
  XNOR U43348 ( .A(q[29]), .B(DB[3315]), .Z(n40325) );
  XNOR U43349 ( .A(q[28]), .B(DB[3314]), .Z(n16216) );
  IV U43350 ( .A(n16229), .Z(n40323) );
  XOR U43351 ( .A(n40326), .B(n40327), .Z(n16229) );
  XNOR U43352 ( .A(n16225), .B(n16227), .Z(n40327) );
  XNOR U43353 ( .A(q[24]), .B(DB[3310]), .Z(n16227) );
  XNOR U43354 ( .A(q[27]), .B(DB[3313]), .Z(n16225) );
  IV U43355 ( .A(n16224), .Z(n40326) );
  XNOR U43356 ( .A(n16222), .B(n40328), .Z(n16224) );
  XNOR U43357 ( .A(q[26]), .B(DB[3312]), .Z(n40328) );
  XNOR U43358 ( .A(q[25]), .B(DB[3311]), .Z(n16222) );
  IV U43359 ( .A(n16237), .Z(n40322) );
  XOR U43360 ( .A(n40329), .B(n40330), .Z(n16237) );
  XNOR U43361 ( .A(n16254), .B(n16235), .Z(n40330) );
  XNOR U43362 ( .A(q[16]), .B(DB[3302]), .Z(n16235) );
  XOR U43363 ( .A(n40331), .B(n16243), .Z(n16254) );
  XNOR U43364 ( .A(q[23]), .B(DB[3309]), .Z(n16243) );
  IV U43365 ( .A(n16242), .Z(n40331) );
  XNOR U43366 ( .A(n16240), .B(n40332), .Z(n16242) );
  XNOR U43367 ( .A(q[22]), .B(DB[3308]), .Z(n40332) );
  XNOR U43368 ( .A(q[21]), .B(DB[3307]), .Z(n16240) );
  IV U43369 ( .A(n16253), .Z(n40329) );
  XOR U43370 ( .A(n40333), .B(n40334), .Z(n16253) );
  XNOR U43371 ( .A(n16249), .B(n16251), .Z(n40334) );
  XNOR U43372 ( .A(q[17]), .B(DB[3303]), .Z(n16251) );
  XNOR U43373 ( .A(q[20]), .B(DB[3306]), .Z(n16249) );
  IV U43374 ( .A(n16248), .Z(n40333) );
  XNOR U43375 ( .A(n16246), .B(n40335), .Z(n16248) );
  XNOR U43376 ( .A(q[19]), .B(DB[3305]), .Z(n40335) );
  XNOR U43377 ( .A(q[18]), .B(DB[3304]), .Z(n16246) );
  IV U43378 ( .A(n16261), .Z(n40321) );
  XOR U43379 ( .A(n40336), .B(n40337), .Z(n16261) );
  XNOR U43380 ( .A(n16288), .B(n16259), .Z(n40337) );
  XNOR U43381 ( .A(q[0]), .B(DB[3286]), .Z(n16259) );
  XOR U43382 ( .A(n40338), .B(n16280), .Z(n16288) );
  XOR U43383 ( .A(n40339), .B(n16268), .Z(n16280) );
  XNOR U43384 ( .A(q[15]), .B(DB[3301]), .Z(n16268) );
  IV U43385 ( .A(n16267), .Z(n40339) );
  XNOR U43386 ( .A(n16265), .B(n40340), .Z(n16267) );
  XNOR U43387 ( .A(q[14]), .B(DB[3300]), .Z(n40340) );
  XNOR U43388 ( .A(q[13]), .B(DB[3299]), .Z(n16265) );
  IV U43389 ( .A(n16279), .Z(n40338) );
  XOR U43390 ( .A(n40341), .B(n40342), .Z(n16279) );
  XNOR U43391 ( .A(n16275), .B(n16277), .Z(n40342) );
  XNOR U43392 ( .A(q[9]), .B(DB[3295]), .Z(n16277) );
  XNOR U43393 ( .A(q[12]), .B(DB[3298]), .Z(n16275) );
  IV U43394 ( .A(n16274), .Z(n40341) );
  XNOR U43395 ( .A(n16272), .B(n40343), .Z(n16274) );
  XNOR U43396 ( .A(q[11]), .B(DB[3297]), .Z(n40343) );
  XNOR U43397 ( .A(q[10]), .B(DB[3296]), .Z(n16272) );
  IV U43398 ( .A(n16287), .Z(n40336) );
  XOR U43399 ( .A(n40344), .B(n40345), .Z(n16287) );
  XNOR U43400 ( .A(n16304), .B(n16285), .Z(n40345) );
  XNOR U43401 ( .A(q[1]), .B(DB[3287]), .Z(n16285) );
  XOR U43402 ( .A(n40346), .B(n16293), .Z(n16304) );
  XNOR U43403 ( .A(q[8]), .B(DB[3294]), .Z(n16293) );
  IV U43404 ( .A(n16292), .Z(n40346) );
  XNOR U43405 ( .A(n16290), .B(n40347), .Z(n16292) );
  XNOR U43406 ( .A(q[7]), .B(DB[3293]), .Z(n40347) );
  XNOR U43407 ( .A(q[6]), .B(DB[3292]), .Z(n16290) );
  IV U43408 ( .A(n16303), .Z(n40344) );
  XOR U43409 ( .A(n40348), .B(n40349), .Z(n16303) );
  XNOR U43410 ( .A(n16299), .B(n16301), .Z(n40349) );
  XNOR U43411 ( .A(q[2]), .B(DB[3288]), .Z(n16301) );
  XNOR U43412 ( .A(q[5]), .B(DB[3291]), .Z(n16299) );
  IV U43413 ( .A(n16298), .Z(n40348) );
  XNOR U43414 ( .A(n16296), .B(n40350), .Z(n16298) );
  XNOR U43415 ( .A(q[4]), .B(DB[3290]), .Z(n40350) );
  XNOR U43416 ( .A(q[3]), .B(DB[3289]), .Z(n16296) );
  XOR U43417 ( .A(n40351), .B(n16065), .Z(n15916) );
  XOR U43418 ( .A(n40352), .B(n16041), .Z(n16065) );
  XOR U43419 ( .A(n40353), .B(n16033), .Z(n16041) );
  XOR U43420 ( .A(n40354), .B(n16022), .Z(n16033) );
  XNOR U43421 ( .A(q[30]), .B(DB[3347]), .Z(n16022) );
  IV U43422 ( .A(n16021), .Z(n40354) );
  XNOR U43423 ( .A(n16019), .B(n40355), .Z(n16021) );
  XNOR U43424 ( .A(q[29]), .B(DB[3346]), .Z(n40355) );
  XNOR U43425 ( .A(q[28]), .B(DB[3345]), .Z(n16019) );
  IV U43426 ( .A(n16032), .Z(n40353) );
  XOR U43427 ( .A(n40356), .B(n40357), .Z(n16032) );
  XNOR U43428 ( .A(n16028), .B(n16030), .Z(n40357) );
  XNOR U43429 ( .A(q[24]), .B(DB[3341]), .Z(n16030) );
  XNOR U43430 ( .A(q[27]), .B(DB[3344]), .Z(n16028) );
  IV U43431 ( .A(n16027), .Z(n40356) );
  XNOR U43432 ( .A(n16025), .B(n40358), .Z(n16027) );
  XNOR U43433 ( .A(q[26]), .B(DB[3343]), .Z(n40358) );
  XNOR U43434 ( .A(q[25]), .B(DB[3342]), .Z(n16025) );
  IV U43435 ( .A(n16040), .Z(n40352) );
  XOR U43436 ( .A(n40359), .B(n40360), .Z(n16040) );
  XNOR U43437 ( .A(n16057), .B(n16038), .Z(n40360) );
  XNOR U43438 ( .A(q[16]), .B(DB[3333]), .Z(n16038) );
  XOR U43439 ( .A(n40361), .B(n16046), .Z(n16057) );
  XNOR U43440 ( .A(q[23]), .B(DB[3340]), .Z(n16046) );
  IV U43441 ( .A(n16045), .Z(n40361) );
  XNOR U43442 ( .A(n16043), .B(n40362), .Z(n16045) );
  XNOR U43443 ( .A(q[22]), .B(DB[3339]), .Z(n40362) );
  XNOR U43444 ( .A(q[21]), .B(DB[3338]), .Z(n16043) );
  IV U43445 ( .A(n16056), .Z(n40359) );
  XOR U43446 ( .A(n40363), .B(n40364), .Z(n16056) );
  XNOR U43447 ( .A(n16052), .B(n16054), .Z(n40364) );
  XNOR U43448 ( .A(q[17]), .B(DB[3334]), .Z(n16054) );
  XNOR U43449 ( .A(q[20]), .B(DB[3337]), .Z(n16052) );
  IV U43450 ( .A(n16051), .Z(n40363) );
  XNOR U43451 ( .A(n16049), .B(n40365), .Z(n16051) );
  XNOR U43452 ( .A(q[19]), .B(DB[3336]), .Z(n40365) );
  XNOR U43453 ( .A(q[18]), .B(DB[3335]), .Z(n16049) );
  IV U43454 ( .A(n16064), .Z(n40351) );
  XOR U43455 ( .A(n40366), .B(n40367), .Z(n16064) );
  XNOR U43456 ( .A(n16091), .B(n16062), .Z(n40367) );
  XNOR U43457 ( .A(q[0]), .B(DB[3317]), .Z(n16062) );
  XOR U43458 ( .A(n40368), .B(n16083), .Z(n16091) );
  XOR U43459 ( .A(n40369), .B(n16071), .Z(n16083) );
  XNOR U43460 ( .A(q[15]), .B(DB[3332]), .Z(n16071) );
  IV U43461 ( .A(n16070), .Z(n40369) );
  XNOR U43462 ( .A(n16068), .B(n40370), .Z(n16070) );
  XNOR U43463 ( .A(q[14]), .B(DB[3331]), .Z(n40370) );
  XNOR U43464 ( .A(q[13]), .B(DB[3330]), .Z(n16068) );
  IV U43465 ( .A(n16082), .Z(n40368) );
  XOR U43466 ( .A(n40371), .B(n40372), .Z(n16082) );
  XNOR U43467 ( .A(n16078), .B(n16080), .Z(n40372) );
  XNOR U43468 ( .A(q[9]), .B(DB[3326]), .Z(n16080) );
  XNOR U43469 ( .A(q[12]), .B(DB[3329]), .Z(n16078) );
  IV U43470 ( .A(n16077), .Z(n40371) );
  XNOR U43471 ( .A(n16075), .B(n40373), .Z(n16077) );
  XNOR U43472 ( .A(q[11]), .B(DB[3328]), .Z(n40373) );
  XNOR U43473 ( .A(q[10]), .B(DB[3327]), .Z(n16075) );
  IV U43474 ( .A(n16090), .Z(n40366) );
  XOR U43475 ( .A(n40374), .B(n40375), .Z(n16090) );
  XNOR U43476 ( .A(n16107), .B(n16088), .Z(n40375) );
  XNOR U43477 ( .A(q[1]), .B(DB[3318]), .Z(n16088) );
  XOR U43478 ( .A(n40376), .B(n16096), .Z(n16107) );
  XNOR U43479 ( .A(q[8]), .B(DB[3325]), .Z(n16096) );
  IV U43480 ( .A(n16095), .Z(n40376) );
  XNOR U43481 ( .A(n16093), .B(n40377), .Z(n16095) );
  XNOR U43482 ( .A(q[7]), .B(DB[3324]), .Z(n40377) );
  XNOR U43483 ( .A(q[6]), .B(DB[3323]), .Z(n16093) );
  IV U43484 ( .A(n16106), .Z(n40374) );
  XOR U43485 ( .A(n40378), .B(n40379), .Z(n16106) );
  XNOR U43486 ( .A(n16102), .B(n16104), .Z(n40379) );
  XNOR U43487 ( .A(q[2]), .B(DB[3319]), .Z(n16104) );
  XNOR U43488 ( .A(q[5]), .B(DB[3322]), .Z(n16102) );
  IV U43489 ( .A(n16101), .Z(n40378) );
  XNOR U43490 ( .A(n16099), .B(n40380), .Z(n16101) );
  XNOR U43491 ( .A(q[4]), .B(DB[3321]), .Z(n40380) );
  XNOR U43492 ( .A(q[3]), .B(DB[3320]), .Z(n16099) );
  XOR U43493 ( .A(n40381), .B(n15868), .Z(n15719) );
  XOR U43494 ( .A(n40382), .B(n15844), .Z(n15868) );
  XOR U43495 ( .A(n40383), .B(n15836), .Z(n15844) );
  XOR U43496 ( .A(n40384), .B(n15825), .Z(n15836) );
  XNOR U43497 ( .A(q[30]), .B(DB[3378]), .Z(n15825) );
  IV U43498 ( .A(n15824), .Z(n40384) );
  XNOR U43499 ( .A(n15822), .B(n40385), .Z(n15824) );
  XNOR U43500 ( .A(q[29]), .B(DB[3377]), .Z(n40385) );
  XNOR U43501 ( .A(q[28]), .B(DB[3376]), .Z(n15822) );
  IV U43502 ( .A(n15835), .Z(n40383) );
  XOR U43503 ( .A(n40386), .B(n40387), .Z(n15835) );
  XNOR U43504 ( .A(n15831), .B(n15833), .Z(n40387) );
  XNOR U43505 ( .A(q[24]), .B(DB[3372]), .Z(n15833) );
  XNOR U43506 ( .A(q[27]), .B(DB[3375]), .Z(n15831) );
  IV U43507 ( .A(n15830), .Z(n40386) );
  XNOR U43508 ( .A(n15828), .B(n40388), .Z(n15830) );
  XNOR U43509 ( .A(q[26]), .B(DB[3374]), .Z(n40388) );
  XNOR U43510 ( .A(q[25]), .B(DB[3373]), .Z(n15828) );
  IV U43511 ( .A(n15843), .Z(n40382) );
  XOR U43512 ( .A(n40389), .B(n40390), .Z(n15843) );
  XNOR U43513 ( .A(n15860), .B(n15841), .Z(n40390) );
  XNOR U43514 ( .A(q[16]), .B(DB[3364]), .Z(n15841) );
  XOR U43515 ( .A(n40391), .B(n15849), .Z(n15860) );
  XNOR U43516 ( .A(q[23]), .B(DB[3371]), .Z(n15849) );
  IV U43517 ( .A(n15848), .Z(n40391) );
  XNOR U43518 ( .A(n15846), .B(n40392), .Z(n15848) );
  XNOR U43519 ( .A(q[22]), .B(DB[3370]), .Z(n40392) );
  XNOR U43520 ( .A(q[21]), .B(DB[3369]), .Z(n15846) );
  IV U43521 ( .A(n15859), .Z(n40389) );
  XOR U43522 ( .A(n40393), .B(n40394), .Z(n15859) );
  XNOR U43523 ( .A(n15855), .B(n15857), .Z(n40394) );
  XNOR U43524 ( .A(q[17]), .B(DB[3365]), .Z(n15857) );
  XNOR U43525 ( .A(q[20]), .B(DB[3368]), .Z(n15855) );
  IV U43526 ( .A(n15854), .Z(n40393) );
  XNOR U43527 ( .A(n15852), .B(n40395), .Z(n15854) );
  XNOR U43528 ( .A(q[19]), .B(DB[3367]), .Z(n40395) );
  XNOR U43529 ( .A(q[18]), .B(DB[3366]), .Z(n15852) );
  IV U43530 ( .A(n15867), .Z(n40381) );
  XOR U43531 ( .A(n40396), .B(n40397), .Z(n15867) );
  XNOR U43532 ( .A(n15894), .B(n15865), .Z(n40397) );
  XNOR U43533 ( .A(q[0]), .B(DB[3348]), .Z(n15865) );
  XOR U43534 ( .A(n40398), .B(n15886), .Z(n15894) );
  XOR U43535 ( .A(n40399), .B(n15874), .Z(n15886) );
  XNOR U43536 ( .A(q[15]), .B(DB[3363]), .Z(n15874) );
  IV U43537 ( .A(n15873), .Z(n40399) );
  XNOR U43538 ( .A(n15871), .B(n40400), .Z(n15873) );
  XNOR U43539 ( .A(q[14]), .B(DB[3362]), .Z(n40400) );
  XNOR U43540 ( .A(q[13]), .B(DB[3361]), .Z(n15871) );
  IV U43541 ( .A(n15885), .Z(n40398) );
  XOR U43542 ( .A(n40401), .B(n40402), .Z(n15885) );
  XNOR U43543 ( .A(n15881), .B(n15883), .Z(n40402) );
  XNOR U43544 ( .A(q[9]), .B(DB[3357]), .Z(n15883) );
  XNOR U43545 ( .A(q[12]), .B(DB[3360]), .Z(n15881) );
  IV U43546 ( .A(n15880), .Z(n40401) );
  XNOR U43547 ( .A(n15878), .B(n40403), .Z(n15880) );
  XNOR U43548 ( .A(q[11]), .B(DB[3359]), .Z(n40403) );
  XNOR U43549 ( .A(q[10]), .B(DB[3358]), .Z(n15878) );
  IV U43550 ( .A(n15893), .Z(n40396) );
  XOR U43551 ( .A(n40404), .B(n40405), .Z(n15893) );
  XNOR U43552 ( .A(n15910), .B(n15891), .Z(n40405) );
  XNOR U43553 ( .A(q[1]), .B(DB[3349]), .Z(n15891) );
  XOR U43554 ( .A(n40406), .B(n15899), .Z(n15910) );
  XNOR U43555 ( .A(q[8]), .B(DB[3356]), .Z(n15899) );
  IV U43556 ( .A(n15898), .Z(n40406) );
  XNOR U43557 ( .A(n15896), .B(n40407), .Z(n15898) );
  XNOR U43558 ( .A(q[7]), .B(DB[3355]), .Z(n40407) );
  XNOR U43559 ( .A(q[6]), .B(DB[3354]), .Z(n15896) );
  IV U43560 ( .A(n15909), .Z(n40404) );
  XOR U43561 ( .A(n40408), .B(n40409), .Z(n15909) );
  XNOR U43562 ( .A(n15905), .B(n15907), .Z(n40409) );
  XNOR U43563 ( .A(q[2]), .B(DB[3350]), .Z(n15907) );
  XNOR U43564 ( .A(q[5]), .B(DB[3353]), .Z(n15905) );
  IV U43565 ( .A(n15904), .Z(n40408) );
  XNOR U43566 ( .A(n15902), .B(n40410), .Z(n15904) );
  XNOR U43567 ( .A(q[4]), .B(DB[3352]), .Z(n40410) );
  XNOR U43568 ( .A(q[3]), .B(DB[3351]), .Z(n15902) );
  XOR U43569 ( .A(n40411), .B(n15671), .Z(n15522) );
  XOR U43570 ( .A(n40412), .B(n15647), .Z(n15671) );
  XOR U43571 ( .A(n40413), .B(n15639), .Z(n15647) );
  XOR U43572 ( .A(n40414), .B(n15628), .Z(n15639) );
  XNOR U43573 ( .A(q[30]), .B(DB[3409]), .Z(n15628) );
  IV U43574 ( .A(n15627), .Z(n40414) );
  XNOR U43575 ( .A(n15625), .B(n40415), .Z(n15627) );
  XNOR U43576 ( .A(q[29]), .B(DB[3408]), .Z(n40415) );
  XNOR U43577 ( .A(q[28]), .B(DB[3407]), .Z(n15625) );
  IV U43578 ( .A(n15638), .Z(n40413) );
  XOR U43579 ( .A(n40416), .B(n40417), .Z(n15638) );
  XNOR U43580 ( .A(n15634), .B(n15636), .Z(n40417) );
  XNOR U43581 ( .A(q[24]), .B(DB[3403]), .Z(n15636) );
  XNOR U43582 ( .A(q[27]), .B(DB[3406]), .Z(n15634) );
  IV U43583 ( .A(n15633), .Z(n40416) );
  XNOR U43584 ( .A(n15631), .B(n40418), .Z(n15633) );
  XNOR U43585 ( .A(q[26]), .B(DB[3405]), .Z(n40418) );
  XNOR U43586 ( .A(q[25]), .B(DB[3404]), .Z(n15631) );
  IV U43587 ( .A(n15646), .Z(n40412) );
  XOR U43588 ( .A(n40419), .B(n40420), .Z(n15646) );
  XNOR U43589 ( .A(n15663), .B(n15644), .Z(n40420) );
  XNOR U43590 ( .A(q[16]), .B(DB[3395]), .Z(n15644) );
  XOR U43591 ( .A(n40421), .B(n15652), .Z(n15663) );
  XNOR U43592 ( .A(q[23]), .B(DB[3402]), .Z(n15652) );
  IV U43593 ( .A(n15651), .Z(n40421) );
  XNOR U43594 ( .A(n15649), .B(n40422), .Z(n15651) );
  XNOR U43595 ( .A(q[22]), .B(DB[3401]), .Z(n40422) );
  XNOR U43596 ( .A(q[21]), .B(DB[3400]), .Z(n15649) );
  IV U43597 ( .A(n15662), .Z(n40419) );
  XOR U43598 ( .A(n40423), .B(n40424), .Z(n15662) );
  XNOR U43599 ( .A(n15658), .B(n15660), .Z(n40424) );
  XNOR U43600 ( .A(q[17]), .B(DB[3396]), .Z(n15660) );
  XNOR U43601 ( .A(q[20]), .B(DB[3399]), .Z(n15658) );
  IV U43602 ( .A(n15657), .Z(n40423) );
  XNOR U43603 ( .A(n15655), .B(n40425), .Z(n15657) );
  XNOR U43604 ( .A(q[19]), .B(DB[3398]), .Z(n40425) );
  XNOR U43605 ( .A(q[18]), .B(DB[3397]), .Z(n15655) );
  IV U43606 ( .A(n15670), .Z(n40411) );
  XOR U43607 ( .A(n40426), .B(n40427), .Z(n15670) );
  XNOR U43608 ( .A(n15697), .B(n15668), .Z(n40427) );
  XNOR U43609 ( .A(q[0]), .B(DB[3379]), .Z(n15668) );
  XOR U43610 ( .A(n40428), .B(n15689), .Z(n15697) );
  XOR U43611 ( .A(n40429), .B(n15677), .Z(n15689) );
  XNOR U43612 ( .A(q[15]), .B(DB[3394]), .Z(n15677) );
  IV U43613 ( .A(n15676), .Z(n40429) );
  XNOR U43614 ( .A(n15674), .B(n40430), .Z(n15676) );
  XNOR U43615 ( .A(q[14]), .B(DB[3393]), .Z(n40430) );
  XNOR U43616 ( .A(q[13]), .B(DB[3392]), .Z(n15674) );
  IV U43617 ( .A(n15688), .Z(n40428) );
  XOR U43618 ( .A(n40431), .B(n40432), .Z(n15688) );
  XNOR U43619 ( .A(n15684), .B(n15686), .Z(n40432) );
  XNOR U43620 ( .A(q[9]), .B(DB[3388]), .Z(n15686) );
  XNOR U43621 ( .A(q[12]), .B(DB[3391]), .Z(n15684) );
  IV U43622 ( .A(n15683), .Z(n40431) );
  XNOR U43623 ( .A(n15681), .B(n40433), .Z(n15683) );
  XNOR U43624 ( .A(q[11]), .B(DB[3390]), .Z(n40433) );
  XNOR U43625 ( .A(q[10]), .B(DB[3389]), .Z(n15681) );
  IV U43626 ( .A(n15696), .Z(n40426) );
  XOR U43627 ( .A(n40434), .B(n40435), .Z(n15696) );
  XNOR U43628 ( .A(n15713), .B(n15694), .Z(n40435) );
  XNOR U43629 ( .A(q[1]), .B(DB[3380]), .Z(n15694) );
  XOR U43630 ( .A(n40436), .B(n15702), .Z(n15713) );
  XNOR U43631 ( .A(q[8]), .B(DB[3387]), .Z(n15702) );
  IV U43632 ( .A(n15701), .Z(n40436) );
  XNOR U43633 ( .A(n15699), .B(n40437), .Z(n15701) );
  XNOR U43634 ( .A(q[7]), .B(DB[3386]), .Z(n40437) );
  XNOR U43635 ( .A(q[6]), .B(DB[3385]), .Z(n15699) );
  IV U43636 ( .A(n15712), .Z(n40434) );
  XOR U43637 ( .A(n40438), .B(n40439), .Z(n15712) );
  XNOR U43638 ( .A(n15708), .B(n15710), .Z(n40439) );
  XNOR U43639 ( .A(q[2]), .B(DB[3381]), .Z(n15710) );
  XNOR U43640 ( .A(q[5]), .B(DB[3384]), .Z(n15708) );
  IV U43641 ( .A(n15707), .Z(n40438) );
  XNOR U43642 ( .A(n15705), .B(n40440), .Z(n15707) );
  XNOR U43643 ( .A(q[4]), .B(DB[3383]), .Z(n40440) );
  XNOR U43644 ( .A(q[3]), .B(DB[3382]), .Z(n15705) );
  XOR U43645 ( .A(n40441), .B(n15474), .Z(n15325) );
  XOR U43646 ( .A(n40442), .B(n15450), .Z(n15474) );
  XOR U43647 ( .A(n40443), .B(n15442), .Z(n15450) );
  XOR U43648 ( .A(n40444), .B(n15431), .Z(n15442) );
  XNOR U43649 ( .A(q[30]), .B(DB[3440]), .Z(n15431) );
  IV U43650 ( .A(n15430), .Z(n40444) );
  XNOR U43651 ( .A(n15428), .B(n40445), .Z(n15430) );
  XNOR U43652 ( .A(q[29]), .B(DB[3439]), .Z(n40445) );
  XNOR U43653 ( .A(q[28]), .B(DB[3438]), .Z(n15428) );
  IV U43654 ( .A(n15441), .Z(n40443) );
  XOR U43655 ( .A(n40446), .B(n40447), .Z(n15441) );
  XNOR U43656 ( .A(n15437), .B(n15439), .Z(n40447) );
  XNOR U43657 ( .A(q[24]), .B(DB[3434]), .Z(n15439) );
  XNOR U43658 ( .A(q[27]), .B(DB[3437]), .Z(n15437) );
  IV U43659 ( .A(n15436), .Z(n40446) );
  XNOR U43660 ( .A(n15434), .B(n40448), .Z(n15436) );
  XNOR U43661 ( .A(q[26]), .B(DB[3436]), .Z(n40448) );
  XNOR U43662 ( .A(q[25]), .B(DB[3435]), .Z(n15434) );
  IV U43663 ( .A(n15449), .Z(n40442) );
  XOR U43664 ( .A(n40449), .B(n40450), .Z(n15449) );
  XNOR U43665 ( .A(n15466), .B(n15447), .Z(n40450) );
  XNOR U43666 ( .A(q[16]), .B(DB[3426]), .Z(n15447) );
  XOR U43667 ( .A(n40451), .B(n15455), .Z(n15466) );
  XNOR U43668 ( .A(q[23]), .B(DB[3433]), .Z(n15455) );
  IV U43669 ( .A(n15454), .Z(n40451) );
  XNOR U43670 ( .A(n15452), .B(n40452), .Z(n15454) );
  XNOR U43671 ( .A(q[22]), .B(DB[3432]), .Z(n40452) );
  XNOR U43672 ( .A(q[21]), .B(DB[3431]), .Z(n15452) );
  IV U43673 ( .A(n15465), .Z(n40449) );
  XOR U43674 ( .A(n40453), .B(n40454), .Z(n15465) );
  XNOR U43675 ( .A(n15461), .B(n15463), .Z(n40454) );
  XNOR U43676 ( .A(q[17]), .B(DB[3427]), .Z(n15463) );
  XNOR U43677 ( .A(q[20]), .B(DB[3430]), .Z(n15461) );
  IV U43678 ( .A(n15460), .Z(n40453) );
  XNOR U43679 ( .A(n15458), .B(n40455), .Z(n15460) );
  XNOR U43680 ( .A(q[19]), .B(DB[3429]), .Z(n40455) );
  XNOR U43681 ( .A(q[18]), .B(DB[3428]), .Z(n15458) );
  IV U43682 ( .A(n15473), .Z(n40441) );
  XOR U43683 ( .A(n40456), .B(n40457), .Z(n15473) );
  XNOR U43684 ( .A(n15500), .B(n15471), .Z(n40457) );
  XNOR U43685 ( .A(q[0]), .B(DB[3410]), .Z(n15471) );
  XOR U43686 ( .A(n40458), .B(n15492), .Z(n15500) );
  XOR U43687 ( .A(n40459), .B(n15480), .Z(n15492) );
  XNOR U43688 ( .A(q[15]), .B(DB[3425]), .Z(n15480) );
  IV U43689 ( .A(n15479), .Z(n40459) );
  XNOR U43690 ( .A(n15477), .B(n40460), .Z(n15479) );
  XNOR U43691 ( .A(q[14]), .B(DB[3424]), .Z(n40460) );
  XNOR U43692 ( .A(q[13]), .B(DB[3423]), .Z(n15477) );
  IV U43693 ( .A(n15491), .Z(n40458) );
  XOR U43694 ( .A(n40461), .B(n40462), .Z(n15491) );
  XNOR U43695 ( .A(n15487), .B(n15489), .Z(n40462) );
  XNOR U43696 ( .A(q[9]), .B(DB[3419]), .Z(n15489) );
  XNOR U43697 ( .A(q[12]), .B(DB[3422]), .Z(n15487) );
  IV U43698 ( .A(n15486), .Z(n40461) );
  XNOR U43699 ( .A(n15484), .B(n40463), .Z(n15486) );
  XNOR U43700 ( .A(q[11]), .B(DB[3421]), .Z(n40463) );
  XNOR U43701 ( .A(q[10]), .B(DB[3420]), .Z(n15484) );
  IV U43702 ( .A(n15499), .Z(n40456) );
  XOR U43703 ( .A(n40464), .B(n40465), .Z(n15499) );
  XNOR U43704 ( .A(n15516), .B(n15497), .Z(n40465) );
  XNOR U43705 ( .A(q[1]), .B(DB[3411]), .Z(n15497) );
  XOR U43706 ( .A(n40466), .B(n15505), .Z(n15516) );
  XNOR U43707 ( .A(q[8]), .B(DB[3418]), .Z(n15505) );
  IV U43708 ( .A(n15504), .Z(n40466) );
  XNOR U43709 ( .A(n15502), .B(n40467), .Z(n15504) );
  XNOR U43710 ( .A(q[7]), .B(DB[3417]), .Z(n40467) );
  XNOR U43711 ( .A(q[6]), .B(DB[3416]), .Z(n15502) );
  IV U43712 ( .A(n15515), .Z(n40464) );
  XOR U43713 ( .A(n40468), .B(n40469), .Z(n15515) );
  XNOR U43714 ( .A(n15511), .B(n15513), .Z(n40469) );
  XNOR U43715 ( .A(q[2]), .B(DB[3412]), .Z(n15513) );
  XNOR U43716 ( .A(q[5]), .B(DB[3415]), .Z(n15511) );
  IV U43717 ( .A(n15510), .Z(n40468) );
  XNOR U43718 ( .A(n15508), .B(n40470), .Z(n15510) );
  XNOR U43719 ( .A(q[4]), .B(DB[3414]), .Z(n40470) );
  XNOR U43720 ( .A(q[3]), .B(DB[3413]), .Z(n15508) );
  XOR U43721 ( .A(n40471), .B(n15277), .Z(n15128) );
  XOR U43722 ( .A(n40472), .B(n15253), .Z(n15277) );
  XOR U43723 ( .A(n40473), .B(n15245), .Z(n15253) );
  XOR U43724 ( .A(n40474), .B(n15234), .Z(n15245) );
  XNOR U43725 ( .A(q[30]), .B(DB[3471]), .Z(n15234) );
  IV U43726 ( .A(n15233), .Z(n40474) );
  XNOR U43727 ( .A(n15231), .B(n40475), .Z(n15233) );
  XNOR U43728 ( .A(q[29]), .B(DB[3470]), .Z(n40475) );
  XNOR U43729 ( .A(q[28]), .B(DB[3469]), .Z(n15231) );
  IV U43730 ( .A(n15244), .Z(n40473) );
  XOR U43731 ( .A(n40476), .B(n40477), .Z(n15244) );
  XNOR U43732 ( .A(n15240), .B(n15242), .Z(n40477) );
  XNOR U43733 ( .A(q[24]), .B(DB[3465]), .Z(n15242) );
  XNOR U43734 ( .A(q[27]), .B(DB[3468]), .Z(n15240) );
  IV U43735 ( .A(n15239), .Z(n40476) );
  XNOR U43736 ( .A(n15237), .B(n40478), .Z(n15239) );
  XNOR U43737 ( .A(q[26]), .B(DB[3467]), .Z(n40478) );
  XNOR U43738 ( .A(q[25]), .B(DB[3466]), .Z(n15237) );
  IV U43739 ( .A(n15252), .Z(n40472) );
  XOR U43740 ( .A(n40479), .B(n40480), .Z(n15252) );
  XNOR U43741 ( .A(n15269), .B(n15250), .Z(n40480) );
  XNOR U43742 ( .A(q[16]), .B(DB[3457]), .Z(n15250) );
  XOR U43743 ( .A(n40481), .B(n15258), .Z(n15269) );
  XNOR U43744 ( .A(q[23]), .B(DB[3464]), .Z(n15258) );
  IV U43745 ( .A(n15257), .Z(n40481) );
  XNOR U43746 ( .A(n15255), .B(n40482), .Z(n15257) );
  XNOR U43747 ( .A(q[22]), .B(DB[3463]), .Z(n40482) );
  XNOR U43748 ( .A(q[21]), .B(DB[3462]), .Z(n15255) );
  IV U43749 ( .A(n15268), .Z(n40479) );
  XOR U43750 ( .A(n40483), .B(n40484), .Z(n15268) );
  XNOR U43751 ( .A(n15264), .B(n15266), .Z(n40484) );
  XNOR U43752 ( .A(q[17]), .B(DB[3458]), .Z(n15266) );
  XNOR U43753 ( .A(q[20]), .B(DB[3461]), .Z(n15264) );
  IV U43754 ( .A(n15263), .Z(n40483) );
  XNOR U43755 ( .A(n15261), .B(n40485), .Z(n15263) );
  XNOR U43756 ( .A(q[19]), .B(DB[3460]), .Z(n40485) );
  XNOR U43757 ( .A(q[18]), .B(DB[3459]), .Z(n15261) );
  IV U43758 ( .A(n15276), .Z(n40471) );
  XOR U43759 ( .A(n40486), .B(n40487), .Z(n15276) );
  XNOR U43760 ( .A(n15303), .B(n15274), .Z(n40487) );
  XNOR U43761 ( .A(q[0]), .B(DB[3441]), .Z(n15274) );
  XOR U43762 ( .A(n40488), .B(n15295), .Z(n15303) );
  XOR U43763 ( .A(n40489), .B(n15283), .Z(n15295) );
  XNOR U43764 ( .A(q[15]), .B(DB[3456]), .Z(n15283) );
  IV U43765 ( .A(n15282), .Z(n40489) );
  XNOR U43766 ( .A(n15280), .B(n40490), .Z(n15282) );
  XNOR U43767 ( .A(q[14]), .B(DB[3455]), .Z(n40490) );
  XNOR U43768 ( .A(q[13]), .B(DB[3454]), .Z(n15280) );
  IV U43769 ( .A(n15294), .Z(n40488) );
  XOR U43770 ( .A(n40491), .B(n40492), .Z(n15294) );
  XNOR U43771 ( .A(n15290), .B(n15292), .Z(n40492) );
  XNOR U43772 ( .A(q[9]), .B(DB[3450]), .Z(n15292) );
  XNOR U43773 ( .A(q[12]), .B(DB[3453]), .Z(n15290) );
  IV U43774 ( .A(n15289), .Z(n40491) );
  XNOR U43775 ( .A(n15287), .B(n40493), .Z(n15289) );
  XNOR U43776 ( .A(q[11]), .B(DB[3452]), .Z(n40493) );
  XNOR U43777 ( .A(q[10]), .B(DB[3451]), .Z(n15287) );
  IV U43778 ( .A(n15302), .Z(n40486) );
  XOR U43779 ( .A(n40494), .B(n40495), .Z(n15302) );
  XNOR U43780 ( .A(n15319), .B(n15300), .Z(n40495) );
  XNOR U43781 ( .A(q[1]), .B(DB[3442]), .Z(n15300) );
  XOR U43782 ( .A(n40496), .B(n15308), .Z(n15319) );
  XNOR U43783 ( .A(q[8]), .B(DB[3449]), .Z(n15308) );
  IV U43784 ( .A(n15307), .Z(n40496) );
  XNOR U43785 ( .A(n15305), .B(n40497), .Z(n15307) );
  XNOR U43786 ( .A(q[7]), .B(DB[3448]), .Z(n40497) );
  XNOR U43787 ( .A(q[6]), .B(DB[3447]), .Z(n15305) );
  IV U43788 ( .A(n15318), .Z(n40494) );
  XOR U43789 ( .A(n40498), .B(n40499), .Z(n15318) );
  XNOR U43790 ( .A(n15314), .B(n15316), .Z(n40499) );
  XNOR U43791 ( .A(q[2]), .B(DB[3443]), .Z(n15316) );
  XNOR U43792 ( .A(q[5]), .B(DB[3446]), .Z(n15314) );
  IV U43793 ( .A(n15313), .Z(n40498) );
  XNOR U43794 ( .A(n15311), .B(n40500), .Z(n15313) );
  XNOR U43795 ( .A(q[4]), .B(DB[3445]), .Z(n40500) );
  XNOR U43796 ( .A(q[3]), .B(DB[3444]), .Z(n15311) );
  XOR U43797 ( .A(n40501), .B(n15080), .Z(n14931) );
  XOR U43798 ( .A(n40502), .B(n15056), .Z(n15080) );
  XOR U43799 ( .A(n40503), .B(n15048), .Z(n15056) );
  XOR U43800 ( .A(n40504), .B(n15037), .Z(n15048) );
  XNOR U43801 ( .A(q[30]), .B(DB[3502]), .Z(n15037) );
  IV U43802 ( .A(n15036), .Z(n40504) );
  XNOR U43803 ( .A(n15034), .B(n40505), .Z(n15036) );
  XNOR U43804 ( .A(q[29]), .B(DB[3501]), .Z(n40505) );
  XNOR U43805 ( .A(q[28]), .B(DB[3500]), .Z(n15034) );
  IV U43806 ( .A(n15047), .Z(n40503) );
  XOR U43807 ( .A(n40506), .B(n40507), .Z(n15047) );
  XNOR U43808 ( .A(n15043), .B(n15045), .Z(n40507) );
  XNOR U43809 ( .A(q[24]), .B(DB[3496]), .Z(n15045) );
  XNOR U43810 ( .A(q[27]), .B(DB[3499]), .Z(n15043) );
  IV U43811 ( .A(n15042), .Z(n40506) );
  XNOR U43812 ( .A(n15040), .B(n40508), .Z(n15042) );
  XNOR U43813 ( .A(q[26]), .B(DB[3498]), .Z(n40508) );
  XNOR U43814 ( .A(q[25]), .B(DB[3497]), .Z(n15040) );
  IV U43815 ( .A(n15055), .Z(n40502) );
  XOR U43816 ( .A(n40509), .B(n40510), .Z(n15055) );
  XNOR U43817 ( .A(n15072), .B(n15053), .Z(n40510) );
  XNOR U43818 ( .A(q[16]), .B(DB[3488]), .Z(n15053) );
  XOR U43819 ( .A(n40511), .B(n15061), .Z(n15072) );
  XNOR U43820 ( .A(q[23]), .B(DB[3495]), .Z(n15061) );
  IV U43821 ( .A(n15060), .Z(n40511) );
  XNOR U43822 ( .A(n15058), .B(n40512), .Z(n15060) );
  XNOR U43823 ( .A(q[22]), .B(DB[3494]), .Z(n40512) );
  XNOR U43824 ( .A(q[21]), .B(DB[3493]), .Z(n15058) );
  IV U43825 ( .A(n15071), .Z(n40509) );
  XOR U43826 ( .A(n40513), .B(n40514), .Z(n15071) );
  XNOR U43827 ( .A(n15067), .B(n15069), .Z(n40514) );
  XNOR U43828 ( .A(q[17]), .B(DB[3489]), .Z(n15069) );
  XNOR U43829 ( .A(q[20]), .B(DB[3492]), .Z(n15067) );
  IV U43830 ( .A(n15066), .Z(n40513) );
  XNOR U43831 ( .A(n15064), .B(n40515), .Z(n15066) );
  XNOR U43832 ( .A(q[19]), .B(DB[3491]), .Z(n40515) );
  XNOR U43833 ( .A(q[18]), .B(DB[3490]), .Z(n15064) );
  IV U43834 ( .A(n15079), .Z(n40501) );
  XOR U43835 ( .A(n40516), .B(n40517), .Z(n15079) );
  XNOR U43836 ( .A(n15106), .B(n15077), .Z(n40517) );
  XNOR U43837 ( .A(q[0]), .B(DB[3472]), .Z(n15077) );
  XOR U43838 ( .A(n40518), .B(n15098), .Z(n15106) );
  XOR U43839 ( .A(n40519), .B(n15086), .Z(n15098) );
  XNOR U43840 ( .A(q[15]), .B(DB[3487]), .Z(n15086) );
  IV U43841 ( .A(n15085), .Z(n40519) );
  XNOR U43842 ( .A(n15083), .B(n40520), .Z(n15085) );
  XNOR U43843 ( .A(q[14]), .B(DB[3486]), .Z(n40520) );
  XNOR U43844 ( .A(q[13]), .B(DB[3485]), .Z(n15083) );
  IV U43845 ( .A(n15097), .Z(n40518) );
  XOR U43846 ( .A(n40521), .B(n40522), .Z(n15097) );
  XNOR U43847 ( .A(n15093), .B(n15095), .Z(n40522) );
  XNOR U43848 ( .A(q[9]), .B(DB[3481]), .Z(n15095) );
  XNOR U43849 ( .A(q[12]), .B(DB[3484]), .Z(n15093) );
  IV U43850 ( .A(n15092), .Z(n40521) );
  XNOR U43851 ( .A(n15090), .B(n40523), .Z(n15092) );
  XNOR U43852 ( .A(q[11]), .B(DB[3483]), .Z(n40523) );
  XNOR U43853 ( .A(q[10]), .B(DB[3482]), .Z(n15090) );
  IV U43854 ( .A(n15105), .Z(n40516) );
  XOR U43855 ( .A(n40524), .B(n40525), .Z(n15105) );
  XNOR U43856 ( .A(n15122), .B(n15103), .Z(n40525) );
  XNOR U43857 ( .A(q[1]), .B(DB[3473]), .Z(n15103) );
  XOR U43858 ( .A(n40526), .B(n15111), .Z(n15122) );
  XNOR U43859 ( .A(q[8]), .B(DB[3480]), .Z(n15111) );
  IV U43860 ( .A(n15110), .Z(n40526) );
  XNOR U43861 ( .A(n15108), .B(n40527), .Z(n15110) );
  XNOR U43862 ( .A(q[7]), .B(DB[3479]), .Z(n40527) );
  XNOR U43863 ( .A(q[6]), .B(DB[3478]), .Z(n15108) );
  IV U43864 ( .A(n15121), .Z(n40524) );
  XOR U43865 ( .A(n40528), .B(n40529), .Z(n15121) );
  XNOR U43866 ( .A(n15117), .B(n15119), .Z(n40529) );
  XNOR U43867 ( .A(q[2]), .B(DB[3474]), .Z(n15119) );
  XNOR U43868 ( .A(q[5]), .B(DB[3477]), .Z(n15117) );
  IV U43869 ( .A(n15116), .Z(n40528) );
  XNOR U43870 ( .A(n15114), .B(n40530), .Z(n15116) );
  XNOR U43871 ( .A(q[4]), .B(DB[3476]), .Z(n40530) );
  XNOR U43872 ( .A(q[3]), .B(DB[3475]), .Z(n15114) );
  XOR U43873 ( .A(n40531), .B(n14883), .Z(n14734) );
  XOR U43874 ( .A(n40532), .B(n14859), .Z(n14883) );
  XOR U43875 ( .A(n40533), .B(n14851), .Z(n14859) );
  XOR U43876 ( .A(n40534), .B(n14840), .Z(n14851) );
  XNOR U43877 ( .A(q[30]), .B(DB[3533]), .Z(n14840) );
  IV U43878 ( .A(n14839), .Z(n40534) );
  XNOR U43879 ( .A(n14837), .B(n40535), .Z(n14839) );
  XNOR U43880 ( .A(q[29]), .B(DB[3532]), .Z(n40535) );
  XNOR U43881 ( .A(q[28]), .B(DB[3531]), .Z(n14837) );
  IV U43882 ( .A(n14850), .Z(n40533) );
  XOR U43883 ( .A(n40536), .B(n40537), .Z(n14850) );
  XNOR U43884 ( .A(n14846), .B(n14848), .Z(n40537) );
  XNOR U43885 ( .A(q[24]), .B(DB[3527]), .Z(n14848) );
  XNOR U43886 ( .A(q[27]), .B(DB[3530]), .Z(n14846) );
  IV U43887 ( .A(n14845), .Z(n40536) );
  XNOR U43888 ( .A(n14843), .B(n40538), .Z(n14845) );
  XNOR U43889 ( .A(q[26]), .B(DB[3529]), .Z(n40538) );
  XNOR U43890 ( .A(q[25]), .B(DB[3528]), .Z(n14843) );
  IV U43891 ( .A(n14858), .Z(n40532) );
  XOR U43892 ( .A(n40539), .B(n40540), .Z(n14858) );
  XNOR U43893 ( .A(n14875), .B(n14856), .Z(n40540) );
  XNOR U43894 ( .A(q[16]), .B(DB[3519]), .Z(n14856) );
  XOR U43895 ( .A(n40541), .B(n14864), .Z(n14875) );
  XNOR U43896 ( .A(q[23]), .B(DB[3526]), .Z(n14864) );
  IV U43897 ( .A(n14863), .Z(n40541) );
  XNOR U43898 ( .A(n14861), .B(n40542), .Z(n14863) );
  XNOR U43899 ( .A(q[22]), .B(DB[3525]), .Z(n40542) );
  XNOR U43900 ( .A(q[21]), .B(DB[3524]), .Z(n14861) );
  IV U43901 ( .A(n14874), .Z(n40539) );
  XOR U43902 ( .A(n40543), .B(n40544), .Z(n14874) );
  XNOR U43903 ( .A(n14870), .B(n14872), .Z(n40544) );
  XNOR U43904 ( .A(q[17]), .B(DB[3520]), .Z(n14872) );
  XNOR U43905 ( .A(q[20]), .B(DB[3523]), .Z(n14870) );
  IV U43906 ( .A(n14869), .Z(n40543) );
  XNOR U43907 ( .A(n14867), .B(n40545), .Z(n14869) );
  XNOR U43908 ( .A(q[19]), .B(DB[3522]), .Z(n40545) );
  XNOR U43909 ( .A(q[18]), .B(DB[3521]), .Z(n14867) );
  IV U43910 ( .A(n14882), .Z(n40531) );
  XOR U43911 ( .A(n40546), .B(n40547), .Z(n14882) );
  XNOR U43912 ( .A(n14909), .B(n14880), .Z(n40547) );
  XNOR U43913 ( .A(q[0]), .B(DB[3503]), .Z(n14880) );
  XOR U43914 ( .A(n40548), .B(n14901), .Z(n14909) );
  XOR U43915 ( .A(n40549), .B(n14889), .Z(n14901) );
  XNOR U43916 ( .A(q[15]), .B(DB[3518]), .Z(n14889) );
  IV U43917 ( .A(n14888), .Z(n40549) );
  XNOR U43918 ( .A(n14886), .B(n40550), .Z(n14888) );
  XNOR U43919 ( .A(q[14]), .B(DB[3517]), .Z(n40550) );
  XNOR U43920 ( .A(q[13]), .B(DB[3516]), .Z(n14886) );
  IV U43921 ( .A(n14900), .Z(n40548) );
  XOR U43922 ( .A(n40551), .B(n40552), .Z(n14900) );
  XNOR U43923 ( .A(n14896), .B(n14898), .Z(n40552) );
  XNOR U43924 ( .A(q[9]), .B(DB[3512]), .Z(n14898) );
  XNOR U43925 ( .A(q[12]), .B(DB[3515]), .Z(n14896) );
  IV U43926 ( .A(n14895), .Z(n40551) );
  XNOR U43927 ( .A(n14893), .B(n40553), .Z(n14895) );
  XNOR U43928 ( .A(q[11]), .B(DB[3514]), .Z(n40553) );
  XNOR U43929 ( .A(q[10]), .B(DB[3513]), .Z(n14893) );
  IV U43930 ( .A(n14908), .Z(n40546) );
  XOR U43931 ( .A(n40554), .B(n40555), .Z(n14908) );
  XNOR U43932 ( .A(n14925), .B(n14906), .Z(n40555) );
  XNOR U43933 ( .A(q[1]), .B(DB[3504]), .Z(n14906) );
  XOR U43934 ( .A(n40556), .B(n14914), .Z(n14925) );
  XNOR U43935 ( .A(q[8]), .B(DB[3511]), .Z(n14914) );
  IV U43936 ( .A(n14913), .Z(n40556) );
  XNOR U43937 ( .A(n14911), .B(n40557), .Z(n14913) );
  XNOR U43938 ( .A(q[7]), .B(DB[3510]), .Z(n40557) );
  XNOR U43939 ( .A(q[6]), .B(DB[3509]), .Z(n14911) );
  IV U43940 ( .A(n14924), .Z(n40554) );
  XOR U43941 ( .A(n40558), .B(n40559), .Z(n14924) );
  XNOR U43942 ( .A(n14920), .B(n14922), .Z(n40559) );
  XNOR U43943 ( .A(q[2]), .B(DB[3505]), .Z(n14922) );
  XNOR U43944 ( .A(q[5]), .B(DB[3508]), .Z(n14920) );
  IV U43945 ( .A(n14919), .Z(n40558) );
  XNOR U43946 ( .A(n14917), .B(n40560), .Z(n14919) );
  XNOR U43947 ( .A(q[4]), .B(DB[3507]), .Z(n40560) );
  XNOR U43948 ( .A(q[3]), .B(DB[3506]), .Z(n14917) );
  XOR U43949 ( .A(n40561), .B(n14686), .Z(n14537) );
  XOR U43950 ( .A(n40562), .B(n14662), .Z(n14686) );
  XOR U43951 ( .A(n40563), .B(n14654), .Z(n14662) );
  XOR U43952 ( .A(n40564), .B(n14643), .Z(n14654) );
  XNOR U43953 ( .A(q[30]), .B(DB[3564]), .Z(n14643) );
  IV U43954 ( .A(n14642), .Z(n40564) );
  XNOR U43955 ( .A(n14640), .B(n40565), .Z(n14642) );
  XNOR U43956 ( .A(q[29]), .B(DB[3563]), .Z(n40565) );
  XNOR U43957 ( .A(q[28]), .B(DB[3562]), .Z(n14640) );
  IV U43958 ( .A(n14653), .Z(n40563) );
  XOR U43959 ( .A(n40566), .B(n40567), .Z(n14653) );
  XNOR U43960 ( .A(n14649), .B(n14651), .Z(n40567) );
  XNOR U43961 ( .A(q[24]), .B(DB[3558]), .Z(n14651) );
  XNOR U43962 ( .A(q[27]), .B(DB[3561]), .Z(n14649) );
  IV U43963 ( .A(n14648), .Z(n40566) );
  XNOR U43964 ( .A(n14646), .B(n40568), .Z(n14648) );
  XNOR U43965 ( .A(q[26]), .B(DB[3560]), .Z(n40568) );
  XNOR U43966 ( .A(q[25]), .B(DB[3559]), .Z(n14646) );
  IV U43967 ( .A(n14661), .Z(n40562) );
  XOR U43968 ( .A(n40569), .B(n40570), .Z(n14661) );
  XNOR U43969 ( .A(n14678), .B(n14659), .Z(n40570) );
  XNOR U43970 ( .A(q[16]), .B(DB[3550]), .Z(n14659) );
  XOR U43971 ( .A(n40571), .B(n14667), .Z(n14678) );
  XNOR U43972 ( .A(q[23]), .B(DB[3557]), .Z(n14667) );
  IV U43973 ( .A(n14666), .Z(n40571) );
  XNOR U43974 ( .A(n14664), .B(n40572), .Z(n14666) );
  XNOR U43975 ( .A(q[22]), .B(DB[3556]), .Z(n40572) );
  XNOR U43976 ( .A(q[21]), .B(DB[3555]), .Z(n14664) );
  IV U43977 ( .A(n14677), .Z(n40569) );
  XOR U43978 ( .A(n40573), .B(n40574), .Z(n14677) );
  XNOR U43979 ( .A(n14673), .B(n14675), .Z(n40574) );
  XNOR U43980 ( .A(q[17]), .B(DB[3551]), .Z(n14675) );
  XNOR U43981 ( .A(q[20]), .B(DB[3554]), .Z(n14673) );
  IV U43982 ( .A(n14672), .Z(n40573) );
  XNOR U43983 ( .A(n14670), .B(n40575), .Z(n14672) );
  XNOR U43984 ( .A(q[19]), .B(DB[3553]), .Z(n40575) );
  XNOR U43985 ( .A(q[18]), .B(DB[3552]), .Z(n14670) );
  IV U43986 ( .A(n14685), .Z(n40561) );
  XOR U43987 ( .A(n40576), .B(n40577), .Z(n14685) );
  XNOR U43988 ( .A(n14712), .B(n14683), .Z(n40577) );
  XNOR U43989 ( .A(q[0]), .B(DB[3534]), .Z(n14683) );
  XOR U43990 ( .A(n40578), .B(n14704), .Z(n14712) );
  XOR U43991 ( .A(n40579), .B(n14692), .Z(n14704) );
  XNOR U43992 ( .A(q[15]), .B(DB[3549]), .Z(n14692) );
  IV U43993 ( .A(n14691), .Z(n40579) );
  XNOR U43994 ( .A(n14689), .B(n40580), .Z(n14691) );
  XNOR U43995 ( .A(q[14]), .B(DB[3548]), .Z(n40580) );
  XNOR U43996 ( .A(q[13]), .B(DB[3547]), .Z(n14689) );
  IV U43997 ( .A(n14703), .Z(n40578) );
  XOR U43998 ( .A(n40581), .B(n40582), .Z(n14703) );
  XNOR U43999 ( .A(n14699), .B(n14701), .Z(n40582) );
  XNOR U44000 ( .A(q[9]), .B(DB[3543]), .Z(n14701) );
  XNOR U44001 ( .A(q[12]), .B(DB[3546]), .Z(n14699) );
  IV U44002 ( .A(n14698), .Z(n40581) );
  XNOR U44003 ( .A(n14696), .B(n40583), .Z(n14698) );
  XNOR U44004 ( .A(q[11]), .B(DB[3545]), .Z(n40583) );
  XNOR U44005 ( .A(q[10]), .B(DB[3544]), .Z(n14696) );
  IV U44006 ( .A(n14711), .Z(n40576) );
  XOR U44007 ( .A(n40584), .B(n40585), .Z(n14711) );
  XNOR U44008 ( .A(n14728), .B(n14709), .Z(n40585) );
  XNOR U44009 ( .A(q[1]), .B(DB[3535]), .Z(n14709) );
  XOR U44010 ( .A(n40586), .B(n14717), .Z(n14728) );
  XNOR U44011 ( .A(q[8]), .B(DB[3542]), .Z(n14717) );
  IV U44012 ( .A(n14716), .Z(n40586) );
  XNOR U44013 ( .A(n14714), .B(n40587), .Z(n14716) );
  XNOR U44014 ( .A(q[7]), .B(DB[3541]), .Z(n40587) );
  XNOR U44015 ( .A(q[6]), .B(DB[3540]), .Z(n14714) );
  IV U44016 ( .A(n14727), .Z(n40584) );
  XOR U44017 ( .A(n40588), .B(n40589), .Z(n14727) );
  XNOR U44018 ( .A(n14723), .B(n14725), .Z(n40589) );
  XNOR U44019 ( .A(q[2]), .B(DB[3536]), .Z(n14725) );
  XNOR U44020 ( .A(q[5]), .B(DB[3539]), .Z(n14723) );
  IV U44021 ( .A(n14722), .Z(n40588) );
  XNOR U44022 ( .A(n14720), .B(n40590), .Z(n14722) );
  XNOR U44023 ( .A(q[4]), .B(DB[3538]), .Z(n40590) );
  XNOR U44024 ( .A(q[3]), .B(DB[3537]), .Z(n14720) );
  XOR U44025 ( .A(n40591), .B(n14489), .Z(n14340) );
  XOR U44026 ( .A(n40592), .B(n14465), .Z(n14489) );
  XOR U44027 ( .A(n40593), .B(n14457), .Z(n14465) );
  XOR U44028 ( .A(n40594), .B(n14446), .Z(n14457) );
  XNOR U44029 ( .A(q[30]), .B(DB[3595]), .Z(n14446) );
  IV U44030 ( .A(n14445), .Z(n40594) );
  XNOR U44031 ( .A(n14443), .B(n40595), .Z(n14445) );
  XNOR U44032 ( .A(q[29]), .B(DB[3594]), .Z(n40595) );
  XNOR U44033 ( .A(q[28]), .B(DB[3593]), .Z(n14443) );
  IV U44034 ( .A(n14456), .Z(n40593) );
  XOR U44035 ( .A(n40596), .B(n40597), .Z(n14456) );
  XNOR U44036 ( .A(n14452), .B(n14454), .Z(n40597) );
  XNOR U44037 ( .A(q[24]), .B(DB[3589]), .Z(n14454) );
  XNOR U44038 ( .A(q[27]), .B(DB[3592]), .Z(n14452) );
  IV U44039 ( .A(n14451), .Z(n40596) );
  XNOR U44040 ( .A(n14449), .B(n40598), .Z(n14451) );
  XNOR U44041 ( .A(q[26]), .B(DB[3591]), .Z(n40598) );
  XNOR U44042 ( .A(q[25]), .B(DB[3590]), .Z(n14449) );
  IV U44043 ( .A(n14464), .Z(n40592) );
  XOR U44044 ( .A(n40599), .B(n40600), .Z(n14464) );
  XNOR U44045 ( .A(n14481), .B(n14462), .Z(n40600) );
  XNOR U44046 ( .A(q[16]), .B(DB[3581]), .Z(n14462) );
  XOR U44047 ( .A(n40601), .B(n14470), .Z(n14481) );
  XNOR U44048 ( .A(q[23]), .B(DB[3588]), .Z(n14470) );
  IV U44049 ( .A(n14469), .Z(n40601) );
  XNOR U44050 ( .A(n14467), .B(n40602), .Z(n14469) );
  XNOR U44051 ( .A(q[22]), .B(DB[3587]), .Z(n40602) );
  XNOR U44052 ( .A(q[21]), .B(DB[3586]), .Z(n14467) );
  IV U44053 ( .A(n14480), .Z(n40599) );
  XOR U44054 ( .A(n40603), .B(n40604), .Z(n14480) );
  XNOR U44055 ( .A(n14476), .B(n14478), .Z(n40604) );
  XNOR U44056 ( .A(q[17]), .B(DB[3582]), .Z(n14478) );
  XNOR U44057 ( .A(q[20]), .B(DB[3585]), .Z(n14476) );
  IV U44058 ( .A(n14475), .Z(n40603) );
  XNOR U44059 ( .A(n14473), .B(n40605), .Z(n14475) );
  XNOR U44060 ( .A(q[19]), .B(DB[3584]), .Z(n40605) );
  XNOR U44061 ( .A(q[18]), .B(DB[3583]), .Z(n14473) );
  IV U44062 ( .A(n14488), .Z(n40591) );
  XOR U44063 ( .A(n40606), .B(n40607), .Z(n14488) );
  XNOR U44064 ( .A(n14515), .B(n14486), .Z(n40607) );
  XNOR U44065 ( .A(q[0]), .B(DB[3565]), .Z(n14486) );
  XOR U44066 ( .A(n40608), .B(n14507), .Z(n14515) );
  XOR U44067 ( .A(n40609), .B(n14495), .Z(n14507) );
  XNOR U44068 ( .A(q[15]), .B(DB[3580]), .Z(n14495) );
  IV U44069 ( .A(n14494), .Z(n40609) );
  XNOR U44070 ( .A(n14492), .B(n40610), .Z(n14494) );
  XNOR U44071 ( .A(q[14]), .B(DB[3579]), .Z(n40610) );
  XNOR U44072 ( .A(q[13]), .B(DB[3578]), .Z(n14492) );
  IV U44073 ( .A(n14506), .Z(n40608) );
  XOR U44074 ( .A(n40611), .B(n40612), .Z(n14506) );
  XNOR U44075 ( .A(n14502), .B(n14504), .Z(n40612) );
  XNOR U44076 ( .A(q[9]), .B(DB[3574]), .Z(n14504) );
  XNOR U44077 ( .A(q[12]), .B(DB[3577]), .Z(n14502) );
  IV U44078 ( .A(n14501), .Z(n40611) );
  XNOR U44079 ( .A(n14499), .B(n40613), .Z(n14501) );
  XNOR U44080 ( .A(q[11]), .B(DB[3576]), .Z(n40613) );
  XNOR U44081 ( .A(q[10]), .B(DB[3575]), .Z(n14499) );
  IV U44082 ( .A(n14514), .Z(n40606) );
  XOR U44083 ( .A(n40614), .B(n40615), .Z(n14514) );
  XNOR U44084 ( .A(n14531), .B(n14512), .Z(n40615) );
  XNOR U44085 ( .A(q[1]), .B(DB[3566]), .Z(n14512) );
  XOR U44086 ( .A(n40616), .B(n14520), .Z(n14531) );
  XNOR U44087 ( .A(q[8]), .B(DB[3573]), .Z(n14520) );
  IV U44088 ( .A(n14519), .Z(n40616) );
  XNOR U44089 ( .A(n14517), .B(n40617), .Z(n14519) );
  XNOR U44090 ( .A(q[7]), .B(DB[3572]), .Z(n40617) );
  XNOR U44091 ( .A(q[6]), .B(DB[3571]), .Z(n14517) );
  IV U44092 ( .A(n14530), .Z(n40614) );
  XOR U44093 ( .A(n40618), .B(n40619), .Z(n14530) );
  XNOR U44094 ( .A(n14526), .B(n14528), .Z(n40619) );
  XNOR U44095 ( .A(q[2]), .B(DB[3567]), .Z(n14528) );
  XNOR U44096 ( .A(q[5]), .B(DB[3570]), .Z(n14526) );
  IV U44097 ( .A(n14525), .Z(n40618) );
  XNOR U44098 ( .A(n14523), .B(n40620), .Z(n14525) );
  XNOR U44099 ( .A(q[4]), .B(DB[3569]), .Z(n40620) );
  XNOR U44100 ( .A(q[3]), .B(DB[3568]), .Z(n14523) );
  XOR U44101 ( .A(n40621), .B(n14292), .Z(n14143) );
  XOR U44102 ( .A(n40622), .B(n14268), .Z(n14292) );
  XOR U44103 ( .A(n40623), .B(n14260), .Z(n14268) );
  XOR U44104 ( .A(n40624), .B(n14249), .Z(n14260) );
  XNOR U44105 ( .A(q[30]), .B(DB[3626]), .Z(n14249) );
  IV U44106 ( .A(n14248), .Z(n40624) );
  XNOR U44107 ( .A(n14246), .B(n40625), .Z(n14248) );
  XNOR U44108 ( .A(q[29]), .B(DB[3625]), .Z(n40625) );
  XNOR U44109 ( .A(q[28]), .B(DB[3624]), .Z(n14246) );
  IV U44110 ( .A(n14259), .Z(n40623) );
  XOR U44111 ( .A(n40626), .B(n40627), .Z(n14259) );
  XNOR U44112 ( .A(n14255), .B(n14257), .Z(n40627) );
  XNOR U44113 ( .A(q[24]), .B(DB[3620]), .Z(n14257) );
  XNOR U44114 ( .A(q[27]), .B(DB[3623]), .Z(n14255) );
  IV U44115 ( .A(n14254), .Z(n40626) );
  XNOR U44116 ( .A(n14252), .B(n40628), .Z(n14254) );
  XNOR U44117 ( .A(q[26]), .B(DB[3622]), .Z(n40628) );
  XNOR U44118 ( .A(q[25]), .B(DB[3621]), .Z(n14252) );
  IV U44119 ( .A(n14267), .Z(n40622) );
  XOR U44120 ( .A(n40629), .B(n40630), .Z(n14267) );
  XNOR U44121 ( .A(n14284), .B(n14265), .Z(n40630) );
  XNOR U44122 ( .A(q[16]), .B(DB[3612]), .Z(n14265) );
  XOR U44123 ( .A(n40631), .B(n14273), .Z(n14284) );
  XNOR U44124 ( .A(q[23]), .B(DB[3619]), .Z(n14273) );
  IV U44125 ( .A(n14272), .Z(n40631) );
  XNOR U44126 ( .A(n14270), .B(n40632), .Z(n14272) );
  XNOR U44127 ( .A(q[22]), .B(DB[3618]), .Z(n40632) );
  XNOR U44128 ( .A(q[21]), .B(DB[3617]), .Z(n14270) );
  IV U44129 ( .A(n14283), .Z(n40629) );
  XOR U44130 ( .A(n40633), .B(n40634), .Z(n14283) );
  XNOR U44131 ( .A(n14279), .B(n14281), .Z(n40634) );
  XNOR U44132 ( .A(q[17]), .B(DB[3613]), .Z(n14281) );
  XNOR U44133 ( .A(q[20]), .B(DB[3616]), .Z(n14279) );
  IV U44134 ( .A(n14278), .Z(n40633) );
  XNOR U44135 ( .A(n14276), .B(n40635), .Z(n14278) );
  XNOR U44136 ( .A(q[19]), .B(DB[3615]), .Z(n40635) );
  XNOR U44137 ( .A(q[18]), .B(DB[3614]), .Z(n14276) );
  IV U44138 ( .A(n14291), .Z(n40621) );
  XOR U44139 ( .A(n40636), .B(n40637), .Z(n14291) );
  XNOR U44140 ( .A(n14318), .B(n14289), .Z(n40637) );
  XNOR U44141 ( .A(q[0]), .B(DB[3596]), .Z(n14289) );
  XOR U44142 ( .A(n40638), .B(n14310), .Z(n14318) );
  XOR U44143 ( .A(n40639), .B(n14298), .Z(n14310) );
  XNOR U44144 ( .A(q[15]), .B(DB[3611]), .Z(n14298) );
  IV U44145 ( .A(n14297), .Z(n40639) );
  XNOR U44146 ( .A(n14295), .B(n40640), .Z(n14297) );
  XNOR U44147 ( .A(q[14]), .B(DB[3610]), .Z(n40640) );
  XNOR U44148 ( .A(q[13]), .B(DB[3609]), .Z(n14295) );
  IV U44149 ( .A(n14309), .Z(n40638) );
  XOR U44150 ( .A(n40641), .B(n40642), .Z(n14309) );
  XNOR U44151 ( .A(n14305), .B(n14307), .Z(n40642) );
  XNOR U44152 ( .A(q[9]), .B(DB[3605]), .Z(n14307) );
  XNOR U44153 ( .A(q[12]), .B(DB[3608]), .Z(n14305) );
  IV U44154 ( .A(n14304), .Z(n40641) );
  XNOR U44155 ( .A(n14302), .B(n40643), .Z(n14304) );
  XNOR U44156 ( .A(q[11]), .B(DB[3607]), .Z(n40643) );
  XNOR U44157 ( .A(q[10]), .B(DB[3606]), .Z(n14302) );
  IV U44158 ( .A(n14317), .Z(n40636) );
  XOR U44159 ( .A(n40644), .B(n40645), .Z(n14317) );
  XNOR U44160 ( .A(n14334), .B(n14315), .Z(n40645) );
  XNOR U44161 ( .A(q[1]), .B(DB[3597]), .Z(n14315) );
  XOR U44162 ( .A(n40646), .B(n14323), .Z(n14334) );
  XNOR U44163 ( .A(q[8]), .B(DB[3604]), .Z(n14323) );
  IV U44164 ( .A(n14322), .Z(n40646) );
  XNOR U44165 ( .A(n14320), .B(n40647), .Z(n14322) );
  XNOR U44166 ( .A(q[7]), .B(DB[3603]), .Z(n40647) );
  XNOR U44167 ( .A(q[6]), .B(DB[3602]), .Z(n14320) );
  IV U44168 ( .A(n14333), .Z(n40644) );
  XOR U44169 ( .A(n40648), .B(n40649), .Z(n14333) );
  XNOR U44170 ( .A(n14329), .B(n14331), .Z(n40649) );
  XNOR U44171 ( .A(q[2]), .B(DB[3598]), .Z(n14331) );
  XNOR U44172 ( .A(q[5]), .B(DB[3601]), .Z(n14329) );
  IV U44173 ( .A(n14328), .Z(n40648) );
  XNOR U44174 ( .A(n14326), .B(n40650), .Z(n14328) );
  XNOR U44175 ( .A(q[4]), .B(DB[3600]), .Z(n40650) );
  XNOR U44176 ( .A(q[3]), .B(DB[3599]), .Z(n14326) );
  XOR U44177 ( .A(n40651), .B(n14095), .Z(n13946) );
  XOR U44178 ( .A(n40652), .B(n14071), .Z(n14095) );
  XOR U44179 ( .A(n40653), .B(n14063), .Z(n14071) );
  XOR U44180 ( .A(n40654), .B(n14052), .Z(n14063) );
  XNOR U44181 ( .A(q[30]), .B(DB[3657]), .Z(n14052) );
  IV U44182 ( .A(n14051), .Z(n40654) );
  XNOR U44183 ( .A(n14049), .B(n40655), .Z(n14051) );
  XNOR U44184 ( .A(q[29]), .B(DB[3656]), .Z(n40655) );
  XNOR U44185 ( .A(q[28]), .B(DB[3655]), .Z(n14049) );
  IV U44186 ( .A(n14062), .Z(n40653) );
  XOR U44187 ( .A(n40656), .B(n40657), .Z(n14062) );
  XNOR U44188 ( .A(n14058), .B(n14060), .Z(n40657) );
  XNOR U44189 ( .A(q[24]), .B(DB[3651]), .Z(n14060) );
  XNOR U44190 ( .A(q[27]), .B(DB[3654]), .Z(n14058) );
  IV U44191 ( .A(n14057), .Z(n40656) );
  XNOR U44192 ( .A(n14055), .B(n40658), .Z(n14057) );
  XNOR U44193 ( .A(q[26]), .B(DB[3653]), .Z(n40658) );
  XNOR U44194 ( .A(q[25]), .B(DB[3652]), .Z(n14055) );
  IV U44195 ( .A(n14070), .Z(n40652) );
  XOR U44196 ( .A(n40659), .B(n40660), .Z(n14070) );
  XNOR U44197 ( .A(n14087), .B(n14068), .Z(n40660) );
  XNOR U44198 ( .A(q[16]), .B(DB[3643]), .Z(n14068) );
  XOR U44199 ( .A(n40661), .B(n14076), .Z(n14087) );
  XNOR U44200 ( .A(q[23]), .B(DB[3650]), .Z(n14076) );
  IV U44201 ( .A(n14075), .Z(n40661) );
  XNOR U44202 ( .A(n14073), .B(n40662), .Z(n14075) );
  XNOR U44203 ( .A(q[22]), .B(DB[3649]), .Z(n40662) );
  XNOR U44204 ( .A(q[21]), .B(DB[3648]), .Z(n14073) );
  IV U44205 ( .A(n14086), .Z(n40659) );
  XOR U44206 ( .A(n40663), .B(n40664), .Z(n14086) );
  XNOR U44207 ( .A(n14082), .B(n14084), .Z(n40664) );
  XNOR U44208 ( .A(q[17]), .B(DB[3644]), .Z(n14084) );
  XNOR U44209 ( .A(q[20]), .B(DB[3647]), .Z(n14082) );
  IV U44210 ( .A(n14081), .Z(n40663) );
  XNOR U44211 ( .A(n14079), .B(n40665), .Z(n14081) );
  XNOR U44212 ( .A(q[19]), .B(DB[3646]), .Z(n40665) );
  XNOR U44213 ( .A(q[18]), .B(DB[3645]), .Z(n14079) );
  IV U44214 ( .A(n14094), .Z(n40651) );
  XOR U44215 ( .A(n40666), .B(n40667), .Z(n14094) );
  XNOR U44216 ( .A(n14121), .B(n14092), .Z(n40667) );
  XNOR U44217 ( .A(q[0]), .B(DB[3627]), .Z(n14092) );
  XOR U44218 ( .A(n40668), .B(n14113), .Z(n14121) );
  XOR U44219 ( .A(n40669), .B(n14101), .Z(n14113) );
  XNOR U44220 ( .A(q[15]), .B(DB[3642]), .Z(n14101) );
  IV U44221 ( .A(n14100), .Z(n40669) );
  XNOR U44222 ( .A(n14098), .B(n40670), .Z(n14100) );
  XNOR U44223 ( .A(q[14]), .B(DB[3641]), .Z(n40670) );
  XNOR U44224 ( .A(q[13]), .B(DB[3640]), .Z(n14098) );
  IV U44225 ( .A(n14112), .Z(n40668) );
  XOR U44226 ( .A(n40671), .B(n40672), .Z(n14112) );
  XNOR U44227 ( .A(n14108), .B(n14110), .Z(n40672) );
  XNOR U44228 ( .A(q[9]), .B(DB[3636]), .Z(n14110) );
  XNOR U44229 ( .A(q[12]), .B(DB[3639]), .Z(n14108) );
  IV U44230 ( .A(n14107), .Z(n40671) );
  XNOR U44231 ( .A(n14105), .B(n40673), .Z(n14107) );
  XNOR U44232 ( .A(q[11]), .B(DB[3638]), .Z(n40673) );
  XNOR U44233 ( .A(q[10]), .B(DB[3637]), .Z(n14105) );
  IV U44234 ( .A(n14120), .Z(n40666) );
  XOR U44235 ( .A(n40674), .B(n40675), .Z(n14120) );
  XNOR U44236 ( .A(n14137), .B(n14118), .Z(n40675) );
  XNOR U44237 ( .A(q[1]), .B(DB[3628]), .Z(n14118) );
  XOR U44238 ( .A(n40676), .B(n14126), .Z(n14137) );
  XNOR U44239 ( .A(q[8]), .B(DB[3635]), .Z(n14126) );
  IV U44240 ( .A(n14125), .Z(n40676) );
  XNOR U44241 ( .A(n14123), .B(n40677), .Z(n14125) );
  XNOR U44242 ( .A(q[7]), .B(DB[3634]), .Z(n40677) );
  XNOR U44243 ( .A(q[6]), .B(DB[3633]), .Z(n14123) );
  IV U44244 ( .A(n14136), .Z(n40674) );
  XOR U44245 ( .A(n40678), .B(n40679), .Z(n14136) );
  XNOR U44246 ( .A(n14132), .B(n14134), .Z(n40679) );
  XNOR U44247 ( .A(q[2]), .B(DB[3629]), .Z(n14134) );
  XNOR U44248 ( .A(q[5]), .B(DB[3632]), .Z(n14132) );
  IV U44249 ( .A(n14131), .Z(n40678) );
  XNOR U44250 ( .A(n14129), .B(n40680), .Z(n14131) );
  XNOR U44251 ( .A(q[4]), .B(DB[3631]), .Z(n40680) );
  XNOR U44252 ( .A(q[3]), .B(DB[3630]), .Z(n14129) );
  XOR U44253 ( .A(n40681), .B(n13898), .Z(n13749) );
  XOR U44254 ( .A(n40682), .B(n13874), .Z(n13898) );
  XOR U44255 ( .A(n40683), .B(n13866), .Z(n13874) );
  XOR U44256 ( .A(n40684), .B(n13855), .Z(n13866) );
  XNOR U44257 ( .A(q[30]), .B(DB[3688]), .Z(n13855) );
  IV U44258 ( .A(n13854), .Z(n40684) );
  XNOR U44259 ( .A(n13852), .B(n40685), .Z(n13854) );
  XNOR U44260 ( .A(q[29]), .B(DB[3687]), .Z(n40685) );
  XNOR U44261 ( .A(q[28]), .B(DB[3686]), .Z(n13852) );
  IV U44262 ( .A(n13865), .Z(n40683) );
  XOR U44263 ( .A(n40686), .B(n40687), .Z(n13865) );
  XNOR U44264 ( .A(n13861), .B(n13863), .Z(n40687) );
  XNOR U44265 ( .A(q[24]), .B(DB[3682]), .Z(n13863) );
  XNOR U44266 ( .A(q[27]), .B(DB[3685]), .Z(n13861) );
  IV U44267 ( .A(n13860), .Z(n40686) );
  XNOR U44268 ( .A(n13858), .B(n40688), .Z(n13860) );
  XNOR U44269 ( .A(q[26]), .B(DB[3684]), .Z(n40688) );
  XNOR U44270 ( .A(q[25]), .B(DB[3683]), .Z(n13858) );
  IV U44271 ( .A(n13873), .Z(n40682) );
  XOR U44272 ( .A(n40689), .B(n40690), .Z(n13873) );
  XNOR U44273 ( .A(n13890), .B(n13871), .Z(n40690) );
  XNOR U44274 ( .A(q[16]), .B(DB[3674]), .Z(n13871) );
  XOR U44275 ( .A(n40691), .B(n13879), .Z(n13890) );
  XNOR U44276 ( .A(q[23]), .B(DB[3681]), .Z(n13879) );
  IV U44277 ( .A(n13878), .Z(n40691) );
  XNOR U44278 ( .A(n13876), .B(n40692), .Z(n13878) );
  XNOR U44279 ( .A(q[22]), .B(DB[3680]), .Z(n40692) );
  XNOR U44280 ( .A(q[21]), .B(DB[3679]), .Z(n13876) );
  IV U44281 ( .A(n13889), .Z(n40689) );
  XOR U44282 ( .A(n40693), .B(n40694), .Z(n13889) );
  XNOR U44283 ( .A(n13885), .B(n13887), .Z(n40694) );
  XNOR U44284 ( .A(q[17]), .B(DB[3675]), .Z(n13887) );
  XNOR U44285 ( .A(q[20]), .B(DB[3678]), .Z(n13885) );
  IV U44286 ( .A(n13884), .Z(n40693) );
  XNOR U44287 ( .A(n13882), .B(n40695), .Z(n13884) );
  XNOR U44288 ( .A(q[19]), .B(DB[3677]), .Z(n40695) );
  XNOR U44289 ( .A(q[18]), .B(DB[3676]), .Z(n13882) );
  IV U44290 ( .A(n13897), .Z(n40681) );
  XOR U44291 ( .A(n40696), .B(n40697), .Z(n13897) );
  XNOR U44292 ( .A(n13924), .B(n13895), .Z(n40697) );
  XNOR U44293 ( .A(q[0]), .B(DB[3658]), .Z(n13895) );
  XOR U44294 ( .A(n40698), .B(n13916), .Z(n13924) );
  XOR U44295 ( .A(n40699), .B(n13904), .Z(n13916) );
  XNOR U44296 ( .A(q[15]), .B(DB[3673]), .Z(n13904) );
  IV U44297 ( .A(n13903), .Z(n40699) );
  XNOR U44298 ( .A(n13901), .B(n40700), .Z(n13903) );
  XNOR U44299 ( .A(q[14]), .B(DB[3672]), .Z(n40700) );
  XNOR U44300 ( .A(q[13]), .B(DB[3671]), .Z(n13901) );
  IV U44301 ( .A(n13915), .Z(n40698) );
  XOR U44302 ( .A(n40701), .B(n40702), .Z(n13915) );
  XNOR U44303 ( .A(n13911), .B(n13913), .Z(n40702) );
  XNOR U44304 ( .A(q[9]), .B(DB[3667]), .Z(n13913) );
  XNOR U44305 ( .A(q[12]), .B(DB[3670]), .Z(n13911) );
  IV U44306 ( .A(n13910), .Z(n40701) );
  XNOR U44307 ( .A(n13908), .B(n40703), .Z(n13910) );
  XNOR U44308 ( .A(q[11]), .B(DB[3669]), .Z(n40703) );
  XNOR U44309 ( .A(q[10]), .B(DB[3668]), .Z(n13908) );
  IV U44310 ( .A(n13923), .Z(n40696) );
  XOR U44311 ( .A(n40704), .B(n40705), .Z(n13923) );
  XNOR U44312 ( .A(n13940), .B(n13921), .Z(n40705) );
  XNOR U44313 ( .A(q[1]), .B(DB[3659]), .Z(n13921) );
  XOR U44314 ( .A(n40706), .B(n13929), .Z(n13940) );
  XNOR U44315 ( .A(q[8]), .B(DB[3666]), .Z(n13929) );
  IV U44316 ( .A(n13928), .Z(n40706) );
  XNOR U44317 ( .A(n13926), .B(n40707), .Z(n13928) );
  XNOR U44318 ( .A(q[7]), .B(DB[3665]), .Z(n40707) );
  XNOR U44319 ( .A(q[6]), .B(DB[3664]), .Z(n13926) );
  IV U44320 ( .A(n13939), .Z(n40704) );
  XOR U44321 ( .A(n40708), .B(n40709), .Z(n13939) );
  XNOR U44322 ( .A(n13935), .B(n13937), .Z(n40709) );
  XNOR U44323 ( .A(q[2]), .B(DB[3660]), .Z(n13937) );
  XNOR U44324 ( .A(q[5]), .B(DB[3663]), .Z(n13935) );
  IV U44325 ( .A(n13934), .Z(n40708) );
  XNOR U44326 ( .A(n13932), .B(n40710), .Z(n13934) );
  XNOR U44327 ( .A(q[4]), .B(DB[3662]), .Z(n40710) );
  XNOR U44328 ( .A(q[3]), .B(DB[3661]), .Z(n13932) );
  XOR U44329 ( .A(n40711), .B(n13701), .Z(n13552) );
  XOR U44330 ( .A(n40712), .B(n13677), .Z(n13701) );
  XOR U44331 ( .A(n40713), .B(n13669), .Z(n13677) );
  XOR U44332 ( .A(n40714), .B(n13658), .Z(n13669) );
  XNOR U44333 ( .A(q[30]), .B(DB[3719]), .Z(n13658) );
  IV U44334 ( .A(n13657), .Z(n40714) );
  XNOR U44335 ( .A(n13655), .B(n40715), .Z(n13657) );
  XNOR U44336 ( .A(q[29]), .B(DB[3718]), .Z(n40715) );
  XNOR U44337 ( .A(q[28]), .B(DB[3717]), .Z(n13655) );
  IV U44338 ( .A(n13668), .Z(n40713) );
  XOR U44339 ( .A(n40716), .B(n40717), .Z(n13668) );
  XNOR U44340 ( .A(n13664), .B(n13666), .Z(n40717) );
  XNOR U44341 ( .A(q[24]), .B(DB[3713]), .Z(n13666) );
  XNOR U44342 ( .A(q[27]), .B(DB[3716]), .Z(n13664) );
  IV U44343 ( .A(n13663), .Z(n40716) );
  XNOR U44344 ( .A(n13661), .B(n40718), .Z(n13663) );
  XNOR U44345 ( .A(q[26]), .B(DB[3715]), .Z(n40718) );
  XNOR U44346 ( .A(q[25]), .B(DB[3714]), .Z(n13661) );
  IV U44347 ( .A(n13676), .Z(n40712) );
  XOR U44348 ( .A(n40719), .B(n40720), .Z(n13676) );
  XNOR U44349 ( .A(n13693), .B(n13674), .Z(n40720) );
  XNOR U44350 ( .A(q[16]), .B(DB[3705]), .Z(n13674) );
  XOR U44351 ( .A(n40721), .B(n13682), .Z(n13693) );
  XNOR U44352 ( .A(q[23]), .B(DB[3712]), .Z(n13682) );
  IV U44353 ( .A(n13681), .Z(n40721) );
  XNOR U44354 ( .A(n13679), .B(n40722), .Z(n13681) );
  XNOR U44355 ( .A(q[22]), .B(DB[3711]), .Z(n40722) );
  XNOR U44356 ( .A(q[21]), .B(DB[3710]), .Z(n13679) );
  IV U44357 ( .A(n13692), .Z(n40719) );
  XOR U44358 ( .A(n40723), .B(n40724), .Z(n13692) );
  XNOR U44359 ( .A(n13688), .B(n13690), .Z(n40724) );
  XNOR U44360 ( .A(q[17]), .B(DB[3706]), .Z(n13690) );
  XNOR U44361 ( .A(q[20]), .B(DB[3709]), .Z(n13688) );
  IV U44362 ( .A(n13687), .Z(n40723) );
  XNOR U44363 ( .A(n13685), .B(n40725), .Z(n13687) );
  XNOR U44364 ( .A(q[19]), .B(DB[3708]), .Z(n40725) );
  XNOR U44365 ( .A(q[18]), .B(DB[3707]), .Z(n13685) );
  IV U44366 ( .A(n13700), .Z(n40711) );
  XOR U44367 ( .A(n40726), .B(n40727), .Z(n13700) );
  XNOR U44368 ( .A(n13727), .B(n13698), .Z(n40727) );
  XNOR U44369 ( .A(q[0]), .B(DB[3689]), .Z(n13698) );
  XOR U44370 ( .A(n40728), .B(n13719), .Z(n13727) );
  XOR U44371 ( .A(n40729), .B(n13707), .Z(n13719) );
  XNOR U44372 ( .A(q[15]), .B(DB[3704]), .Z(n13707) );
  IV U44373 ( .A(n13706), .Z(n40729) );
  XNOR U44374 ( .A(n13704), .B(n40730), .Z(n13706) );
  XNOR U44375 ( .A(q[14]), .B(DB[3703]), .Z(n40730) );
  XNOR U44376 ( .A(q[13]), .B(DB[3702]), .Z(n13704) );
  IV U44377 ( .A(n13718), .Z(n40728) );
  XOR U44378 ( .A(n40731), .B(n40732), .Z(n13718) );
  XNOR U44379 ( .A(n13714), .B(n13716), .Z(n40732) );
  XNOR U44380 ( .A(q[9]), .B(DB[3698]), .Z(n13716) );
  XNOR U44381 ( .A(q[12]), .B(DB[3701]), .Z(n13714) );
  IV U44382 ( .A(n13713), .Z(n40731) );
  XNOR U44383 ( .A(n13711), .B(n40733), .Z(n13713) );
  XNOR U44384 ( .A(q[11]), .B(DB[3700]), .Z(n40733) );
  XNOR U44385 ( .A(q[10]), .B(DB[3699]), .Z(n13711) );
  IV U44386 ( .A(n13726), .Z(n40726) );
  XOR U44387 ( .A(n40734), .B(n40735), .Z(n13726) );
  XNOR U44388 ( .A(n13743), .B(n13724), .Z(n40735) );
  XNOR U44389 ( .A(q[1]), .B(DB[3690]), .Z(n13724) );
  XOR U44390 ( .A(n40736), .B(n13732), .Z(n13743) );
  XNOR U44391 ( .A(q[8]), .B(DB[3697]), .Z(n13732) );
  IV U44392 ( .A(n13731), .Z(n40736) );
  XNOR U44393 ( .A(n13729), .B(n40737), .Z(n13731) );
  XNOR U44394 ( .A(q[7]), .B(DB[3696]), .Z(n40737) );
  XNOR U44395 ( .A(q[6]), .B(DB[3695]), .Z(n13729) );
  IV U44396 ( .A(n13742), .Z(n40734) );
  XOR U44397 ( .A(n40738), .B(n40739), .Z(n13742) );
  XNOR U44398 ( .A(n13738), .B(n13740), .Z(n40739) );
  XNOR U44399 ( .A(q[2]), .B(DB[3691]), .Z(n13740) );
  XNOR U44400 ( .A(q[5]), .B(DB[3694]), .Z(n13738) );
  IV U44401 ( .A(n13737), .Z(n40738) );
  XNOR U44402 ( .A(n13735), .B(n40740), .Z(n13737) );
  XNOR U44403 ( .A(q[4]), .B(DB[3693]), .Z(n40740) );
  XNOR U44404 ( .A(q[3]), .B(DB[3692]), .Z(n13735) );
  XOR U44405 ( .A(n40741), .B(n13504), .Z(n13355) );
  XOR U44406 ( .A(n40742), .B(n13480), .Z(n13504) );
  XOR U44407 ( .A(n40743), .B(n13472), .Z(n13480) );
  XOR U44408 ( .A(n40744), .B(n13461), .Z(n13472) );
  XNOR U44409 ( .A(q[30]), .B(DB[3750]), .Z(n13461) );
  IV U44410 ( .A(n13460), .Z(n40744) );
  XNOR U44411 ( .A(n13458), .B(n40745), .Z(n13460) );
  XNOR U44412 ( .A(q[29]), .B(DB[3749]), .Z(n40745) );
  XNOR U44413 ( .A(q[28]), .B(DB[3748]), .Z(n13458) );
  IV U44414 ( .A(n13471), .Z(n40743) );
  XOR U44415 ( .A(n40746), .B(n40747), .Z(n13471) );
  XNOR U44416 ( .A(n13467), .B(n13469), .Z(n40747) );
  XNOR U44417 ( .A(q[24]), .B(DB[3744]), .Z(n13469) );
  XNOR U44418 ( .A(q[27]), .B(DB[3747]), .Z(n13467) );
  IV U44419 ( .A(n13466), .Z(n40746) );
  XNOR U44420 ( .A(n13464), .B(n40748), .Z(n13466) );
  XNOR U44421 ( .A(q[26]), .B(DB[3746]), .Z(n40748) );
  XNOR U44422 ( .A(q[25]), .B(DB[3745]), .Z(n13464) );
  IV U44423 ( .A(n13479), .Z(n40742) );
  XOR U44424 ( .A(n40749), .B(n40750), .Z(n13479) );
  XNOR U44425 ( .A(n13496), .B(n13477), .Z(n40750) );
  XNOR U44426 ( .A(q[16]), .B(DB[3736]), .Z(n13477) );
  XOR U44427 ( .A(n40751), .B(n13485), .Z(n13496) );
  XNOR U44428 ( .A(q[23]), .B(DB[3743]), .Z(n13485) );
  IV U44429 ( .A(n13484), .Z(n40751) );
  XNOR U44430 ( .A(n13482), .B(n40752), .Z(n13484) );
  XNOR U44431 ( .A(q[22]), .B(DB[3742]), .Z(n40752) );
  XNOR U44432 ( .A(q[21]), .B(DB[3741]), .Z(n13482) );
  IV U44433 ( .A(n13495), .Z(n40749) );
  XOR U44434 ( .A(n40753), .B(n40754), .Z(n13495) );
  XNOR U44435 ( .A(n13491), .B(n13493), .Z(n40754) );
  XNOR U44436 ( .A(q[17]), .B(DB[3737]), .Z(n13493) );
  XNOR U44437 ( .A(q[20]), .B(DB[3740]), .Z(n13491) );
  IV U44438 ( .A(n13490), .Z(n40753) );
  XNOR U44439 ( .A(n13488), .B(n40755), .Z(n13490) );
  XNOR U44440 ( .A(q[19]), .B(DB[3739]), .Z(n40755) );
  XNOR U44441 ( .A(q[18]), .B(DB[3738]), .Z(n13488) );
  IV U44442 ( .A(n13503), .Z(n40741) );
  XOR U44443 ( .A(n40756), .B(n40757), .Z(n13503) );
  XNOR U44444 ( .A(n13530), .B(n13501), .Z(n40757) );
  XNOR U44445 ( .A(q[0]), .B(DB[3720]), .Z(n13501) );
  XOR U44446 ( .A(n40758), .B(n13522), .Z(n13530) );
  XOR U44447 ( .A(n40759), .B(n13510), .Z(n13522) );
  XNOR U44448 ( .A(q[15]), .B(DB[3735]), .Z(n13510) );
  IV U44449 ( .A(n13509), .Z(n40759) );
  XNOR U44450 ( .A(n13507), .B(n40760), .Z(n13509) );
  XNOR U44451 ( .A(q[14]), .B(DB[3734]), .Z(n40760) );
  XNOR U44452 ( .A(q[13]), .B(DB[3733]), .Z(n13507) );
  IV U44453 ( .A(n13521), .Z(n40758) );
  XOR U44454 ( .A(n40761), .B(n40762), .Z(n13521) );
  XNOR U44455 ( .A(n13517), .B(n13519), .Z(n40762) );
  XNOR U44456 ( .A(q[9]), .B(DB[3729]), .Z(n13519) );
  XNOR U44457 ( .A(q[12]), .B(DB[3732]), .Z(n13517) );
  IV U44458 ( .A(n13516), .Z(n40761) );
  XNOR U44459 ( .A(n13514), .B(n40763), .Z(n13516) );
  XNOR U44460 ( .A(q[11]), .B(DB[3731]), .Z(n40763) );
  XNOR U44461 ( .A(q[10]), .B(DB[3730]), .Z(n13514) );
  IV U44462 ( .A(n13529), .Z(n40756) );
  XOR U44463 ( .A(n40764), .B(n40765), .Z(n13529) );
  XNOR U44464 ( .A(n13546), .B(n13527), .Z(n40765) );
  XNOR U44465 ( .A(q[1]), .B(DB[3721]), .Z(n13527) );
  XOR U44466 ( .A(n40766), .B(n13535), .Z(n13546) );
  XNOR U44467 ( .A(q[8]), .B(DB[3728]), .Z(n13535) );
  IV U44468 ( .A(n13534), .Z(n40766) );
  XNOR U44469 ( .A(n13532), .B(n40767), .Z(n13534) );
  XNOR U44470 ( .A(q[7]), .B(DB[3727]), .Z(n40767) );
  XNOR U44471 ( .A(q[6]), .B(DB[3726]), .Z(n13532) );
  IV U44472 ( .A(n13545), .Z(n40764) );
  XOR U44473 ( .A(n40768), .B(n40769), .Z(n13545) );
  XNOR U44474 ( .A(n13541), .B(n13543), .Z(n40769) );
  XNOR U44475 ( .A(q[2]), .B(DB[3722]), .Z(n13543) );
  XNOR U44476 ( .A(q[5]), .B(DB[3725]), .Z(n13541) );
  IV U44477 ( .A(n13540), .Z(n40768) );
  XNOR U44478 ( .A(n13538), .B(n40770), .Z(n13540) );
  XNOR U44479 ( .A(q[4]), .B(DB[3724]), .Z(n40770) );
  XNOR U44480 ( .A(q[3]), .B(DB[3723]), .Z(n13538) );
  XOR U44481 ( .A(n40771), .B(n13307), .Z(n13158) );
  XOR U44482 ( .A(n40772), .B(n13283), .Z(n13307) );
  XOR U44483 ( .A(n40773), .B(n13275), .Z(n13283) );
  XOR U44484 ( .A(n40774), .B(n13264), .Z(n13275) );
  XNOR U44485 ( .A(q[30]), .B(DB[3781]), .Z(n13264) );
  IV U44486 ( .A(n13263), .Z(n40774) );
  XNOR U44487 ( .A(n13261), .B(n40775), .Z(n13263) );
  XNOR U44488 ( .A(q[29]), .B(DB[3780]), .Z(n40775) );
  XNOR U44489 ( .A(q[28]), .B(DB[3779]), .Z(n13261) );
  IV U44490 ( .A(n13274), .Z(n40773) );
  XOR U44491 ( .A(n40776), .B(n40777), .Z(n13274) );
  XNOR U44492 ( .A(n13270), .B(n13272), .Z(n40777) );
  XNOR U44493 ( .A(q[24]), .B(DB[3775]), .Z(n13272) );
  XNOR U44494 ( .A(q[27]), .B(DB[3778]), .Z(n13270) );
  IV U44495 ( .A(n13269), .Z(n40776) );
  XNOR U44496 ( .A(n13267), .B(n40778), .Z(n13269) );
  XNOR U44497 ( .A(q[26]), .B(DB[3777]), .Z(n40778) );
  XNOR U44498 ( .A(q[25]), .B(DB[3776]), .Z(n13267) );
  IV U44499 ( .A(n13282), .Z(n40772) );
  XOR U44500 ( .A(n40779), .B(n40780), .Z(n13282) );
  XNOR U44501 ( .A(n13299), .B(n13280), .Z(n40780) );
  XNOR U44502 ( .A(q[16]), .B(DB[3767]), .Z(n13280) );
  XOR U44503 ( .A(n40781), .B(n13288), .Z(n13299) );
  XNOR U44504 ( .A(q[23]), .B(DB[3774]), .Z(n13288) );
  IV U44505 ( .A(n13287), .Z(n40781) );
  XNOR U44506 ( .A(n13285), .B(n40782), .Z(n13287) );
  XNOR U44507 ( .A(q[22]), .B(DB[3773]), .Z(n40782) );
  XNOR U44508 ( .A(q[21]), .B(DB[3772]), .Z(n13285) );
  IV U44509 ( .A(n13298), .Z(n40779) );
  XOR U44510 ( .A(n40783), .B(n40784), .Z(n13298) );
  XNOR U44511 ( .A(n13294), .B(n13296), .Z(n40784) );
  XNOR U44512 ( .A(q[17]), .B(DB[3768]), .Z(n13296) );
  XNOR U44513 ( .A(q[20]), .B(DB[3771]), .Z(n13294) );
  IV U44514 ( .A(n13293), .Z(n40783) );
  XNOR U44515 ( .A(n13291), .B(n40785), .Z(n13293) );
  XNOR U44516 ( .A(q[19]), .B(DB[3770]), .Z(n40785) );
  XNOR U44517 ( .A(q[18]), .B(DB[3769]), .Z(n13291) );
  IV U44518 ( .A(n13306), .Z(n40771) );
  XOR U44519 ( .A(n40786), .B(n40787), .Z(n13306) );
  XNOR U44520 ( .A(n13333), .B(n13304), .Z(n40787) );
  XNOR U44521 ( .A(q[0]), .B(DB[3751]), .Z(n13304) );
  XOR U44522 ( .A(n40788), .B(n13325), .Z(n13333) );
  XOR U44523 ( .A(n40789), .B(n13313), .Z(n13325) );
  XNOR U44524 ( .A(q[15]), .B(DB[3766]), .Z(n13313) );
  IV U44525 ( .A(n13312), .Z(n40789) );
  XNOR U44526 ( .A(n13310), .B(n40790), .Z(n13312) );
  XNOR U44527 ( .A(q[14]), .B(DB[3765]), .Z(n40790) );
  XNOR U44528 ( .A(q[13]), .B(DB[3764]), .Z(n13310) );
  IV U44529 ( .A(n13324), .Z(n40788) );
  XOR U44530 ( .A(n40791), .B(n40792), .Z(n13324) );
  XNOR U44531 ( .A(n13320), .B(n13322), .Z(n40792) );
  XNOR U44532 ( .A(q[9]), .B(DB[3760]), .Z(n13322) );
  XNOR U44533 ( .A(q[12]), .B(DB[3763]), .Z(n13320) );
  IV U44534 ( .A(n13319), .Z(n40791) );
  XNOR U44535 ( .A(n13317), .B(n40793), .Z(n13319) );
  XNOR U44536 ( .A(q[11]), .B(DB[3762]), .Z(n40793) );
  XNOR U44537 ( .A(q[10]), .B(DB[3761]), .Z(n13317) );
  IV U44538 ( .A(n13332), .Z(n40786) );
  XOR U44539 ( .A(n40794), .B(n40795), .Z(n13332) );
  XNOR U44540 ( .A(n13349), .B(n13330), .Z(n40795) );
  XNOR U44541 ( .A(q[1]), .B(DB[3752]), .Z(n13330) );
  XOR U44542 ( .A(n40796), .B(n13338), .Z(n13349) );
  XNOR U44543 ( .A(q[8]), .B(DB[3759]), .Z(n13338) );
  IV U44544 ( .A(n13337), .Z(n40796) );
  XNOR U44545 ( .A(n13335), .B(n40797), .Z(n13337) );
  XNOR U44546 ( .A(q[7]), .B(DB[3758]), .Z(n40797) );
  XNOR U44547 ( .A(q[6]), .B(DB[3757]), .Z(n13335) );
  IV U44548 ( .A(n13348), .Z(n40794) );
  XOR U44549 ( .A(n40798), .B(n40799), .Z(n13348) );
  XNOR U44550 ( .A(n13344), .B(n13346), .Z(n40799) );
  XNOR U44551 ( .A(q[2]), .B(DB[3753]), .Z(n13346) );
  XNOR U44552 ( .A(q[5]), .B(DB[3756]), .Z(n13344) );
  IV U44553 ( .A(n13343), .Z(n40798) );
  XNOR U44554 ( .A(n13341), .B(n40800), .Z(n13343) );
  XNOR U44555 ( .A(q[4]), .B(DB[3755]), .Z(n40800) );
  XNOR U44556 ( .A(q[3]), .B(DB[3754]), .Z(n13341) );
  XOR U44557 ( .A(n40801), .B(n13110), .Z(n12961) );
  XOR U44558 ( .A(n40802), .B(n13086), .Z(n13110) );
  XOR U44559 ( .A(n40803), .B(n13078), .Z(n13086) );
  XOR U44560 ( .A(n40804), .B(n13067), .Z(n13078) );
  XNOR U44561 ( .A(q[30]), .B(DB[3812]), .Z(n13067) );
  IV U44562 ( .A(n13066), .Z(n40804) );
  XNOR U44563 ( .A(n13064), .B(n40805), .Z(n13066) );
  XNOR U44564 ( .A(q[29]), .B(DB[3811]), .Z(n40805) );
  XNOR U44565 ( .A(q[28]), .B(DB[3810]), .Z(n13064) );
  IV U44566 ( .A(n13077), .Z(n40803) );
  XOR U44567 ( .A(n40806), .B(n40807), .Z(n13077) );
  XNOR U44568 ( .A(n13073), .B(n13075), .Z(n40807) );
  XNOR U44569 ( .A(q[24]), .B(DB[3806]), .Z(n13075) );
  XNOR U44570 ( .A(q[27]), .B(DB[3809]), .Z(n13073) );
  IV U44571 ( .A(n13072), .Z(n40806) );
  XNOR U44572 ( .A(n13070), .B(n40808), .Z(n13072) );
  XNOR U44573 ( .A(q[26]), .B(DB[3808]), .Z(n40808) );
  XNOR U44574 ( .A(q[25]), .B(DB[3807]), .Z(n13070) );
  IV U44575 ( .A(n13085), .Z(n40802) );
  XOR U44576 ( .A(n40809), .B(n40810), .Z(n13085) );
  XNOR U44577 ( .A(n13102), .B(n13083), .Z(n40810) );
  XNOR U44578 ( .A(q[16]), .B(DB[3798]), .Z(n13083) );
  XOR U44579 ( .A(n40811), .B(n13091), .Z(n13102) );
  XNOR U44580 ( .A(q[23]), .B(DB[3805]), .Z(n13091) );
  IV U44581 ( .A(n13090), .Z(n40811) );
  XNOR U44582 ( .A(n13088), .B(n40812), .Z(n13090) );
  XNOR U44583 ( .A(q[22]), .B(DB[3804]), .Z(n40812) );
  XNOR U44584 ( .A(q[21]), .B(DB[3803]), .Z(n13088) );
  IV U44585 ( .A(n13101), .Z(n40809) );
  XOR U44586 ( .A(n40813), .B(n40814), .Z(n13101) );
  XNOR U44587 ( .A(n13097), .B(n13099), .Z(n40814) );
  XNOR U44588 ( .A(q[17]), .B(DB[3799]), .Z(n13099) );
  XNOR U44589 ( .A(q[20]), .B(DB[3802]), .Z(n13097) );
  IV U44590 ( .A(n13096), .Z(n40813) );
  XNOR U44591 ( .A(n13094), .B(n40815), .Z(n13096) );
  XNOR U44592 ( .A(q[19]), .B(DB[3801]), .Z(n40815) );
  XNOR U44593 ( .A(q[18]), .B(DB[3800]), .Z(n13094) );
  IV U44594 ( .A(n13109), .Z(n40801) );
  XOR U44595 ( .A(n40816), .B(n40817), .Z(n13109) );
  XNOR U44596 ( .A(n13136), .B(n13107), .Z(n40817) );
  XNOR U44597 ( .A(q[0]), .B(DB[3782]), .Z(n13107) );
  XOR U44598 ( .A(n40818), .B(n13128), .Z(n13136) );
  XOR U44599 ( .A(n40819), .B(n13116), .Z(n13128) );
  XNOR U44600 ( .A(q[15]), .B(DB[3797]), .Z(n13116) );
  IV U44601 ( .A(n13115), .Z(n40819) );
  XNOR U44602 ( .A(n13113), .B(n40820), .Z(n13115) );
  XNOR U44603 ( .A(q[14]), .B(DB[3796]), .Z(n40820) );
  XNOR U44604 ( .A(q[13]), .B(DB[3795]), .Z(n13113) );
  IV U44605 ( .A(n13127), .Z(n40818) );
  XOR U44606 ( .A(n40821), .B(n40822), .Z(n13127) );
  XNOR U44607 ( .A(n13123), .B(n13125), .Z(n40822) );
  XNOR U44608 ( .A(q[9]), .B(DB[3791]), .Z(n13125) );
  XNOR U44609 ( .A(q[12]), .B(DB[3794]), .Z(n13123) );
  IV U44610 ( .A(n13122), .Z(n40821) );
  XNOR U44611 ( .A(n13120), .B(n40823), .Z(n13122) );
  XNOR U44612 ( .A(q[11]), .B(DB[3793]), .Z(n40823) );
  XNOR U44613 ( .A(q[10]), .B(DB[3792]), .Z(n13120) );
  IV U44614 ( .A(n13135), .Z(n40816) );
  XOR U44615 ( .A(n40824), .B(n40825), .Z(n13135) );
  XNOR U44616 ( .A(n13152), .B(n13133), .Z(n40825) );
  XNOR U44617 ( .A(q[1]), .B(DB[3783]), .Z(n13133) );
  XOR U44618 ( .A(n40826), .B(n13141), .Z(n13152) );
  XNOR U44619 ( .A(q[8]), .B(DB[3790]), .Z(n13141) );
  IV U44620 ( .A(n13140), .Z(n40826) );
  XNOR U44621 ( .A(n13138), .B(n40827), .Z(n13140) );
  XNOR U44622 ( .A(q[7]), .B(DB[3789]), .Z(n40827) );
  XNOR U44623 ( .A(q[6]), .B(DB[3788]), .Z(n13138) );
  IV U44624 ( .A(n13151), .Z(n40824) );
  XOR U44625 ( .A(n40828), .B(n40829), .Z(n13151) );
  XNOR U44626 ( .A(n13147), .B(n13149), .Z(n40829) );
  XNOR U44627 ( .A(q[2]), .B(DB[3784]), .Z(n13149) );
  XNOR U44628 ( .A(q[5]), .B(DB[3787]), .Z(n13147) );
  IV U44629 ( .A(n13146), .Z(n40828) );
  XNOR U44630 ( .A(n13144), .B(n40830), .Z(n13146) );
  XNOR U44631 ( .A(q[4]), .B(DB[3786]), .Z(n40830) );
  XNOR U44632 ( .A(q[3]), .B(DB[3785]), .Z(n13144) );
  XOR U44633 ( .A(n40831), .B(n12913), .Z(n12764) );
  XOR U44634 ( .A(n40832), .B(n12889), .Z(n12913) );
  XOR U44635 ( .A(n40833), .B(n12881), .Z(n12889) );
  XOR U44636 ( .A(n40834), .B(n12870), .Z(n12881) );
  XNOR U44637 ( .A(q[30]), .B(DB[3843]), .Z(n12870) );
  IV U44638 ( .A(n12869), .Z(n40834) );
  XNOR U44639 ( .A(n12867), .B(n40835), .Z(n12869) );
  XNOR U44640 ( .A(q[29]), .B(DB[3842]), .Z(n40835) );
  XNOR U44641 ( .A(q[28]), .B(DB[3841]), .Z(n12867) );
  IV U44642 ( .A(n12880), .Z(n40833) );
  XOR U44643 ( .A(n40836), .B(n40837), .Z(n12880) );
  XNOR U44644 ( .A(n12876), .B(n12878), .Z(n40837) );
  XNOR U44645 ( .A(q[24]), .B(DB[3837]), .Z(n12878) );
  XNOR U44646 ( .A(q[27]), .B(DB[3840]), .Z(n12876) );
  IV U44647 ( .A(n12875), .Z(n40836) );
  XNOR U44648 ( .A(n12873), .B(n40838), .Z(n12875) );
  XNOR U44649 ( .A(q[26]), .B(DB[3839]), .Z(n40838) );
  XNOR U44650 ( .A(q[25]), .B(DB[3838]), .Z(n12873) );
  IV U44651 ( .A(n12888), .Z(n40832) );
  XOR U44652 ( .A(n40839), .B(n40840), .Z(n12888) );
  XNOR U44653 ( .A(n12905), .B(n12886), .Z(n40840) );
  XNOR U44654 ( .A(q[16]), .B(DB[3829]), .Z(n12886) );
  XOR U44655 ( .A(n40841), .B(n12894), .Z(n12905) );
  XNOR U44656 ( .A(q[23]), .B(DB[3836]), .Z(n12894) );
  IV U44657 ( .A(n12893), .Z(n40841) );
  XNOR U44658 ( .A(n12891), .B(n40842), .Z(n12893) );
  XNOR U44659 ( .A(q[22]), .B(DB[3835]), .Z(n40842) );
  XNOR U44660 ( .A(q[21]), .B(DB[3834]), .Z(n12891) );
  IV U44661 ( .A(n12904), .Z(n40839) );
  XOR U44662 ( .A(n40843), .B(n40844), .Z(n12904) );
  XNOR U44663 ( .A(n12900), .B(n12902), .Z(n40844) );
  XNOR U44664 ( .A(q[17]), .B(DB[3830]), .Z(n12902) );
  XNOR U44665 ( .A(q[20]), .B(DB[3833]), .Z(n12900) );
  IV U44666 ( .A(n12899), .Z(n40843) );
  XNOR U44667 ( .A(n12897), .B(n40845), .Z(n12899) );
  XNOR U44668 ( .A(q[19]), .B(DB[3832]), .Z(n40845) );
  XNOR U44669 ( .A(q[18]), .B(DB[3831]), .Z(n12897) );
  IV U44670 ( .A(n12912), .Z(n40831) );
  XOR U44671 ( .A(n40846), .B(n40847), .Z(n12912) );
  XNOR U44672 ( .A(n12939), .B(n12910), .Z(n40847) );
  XNOR U44673 ( .A(q[0]), .B(DB[3813]), .Z(n12910) );
  XOR U44674 ( .A(n40848), .B(n12931), .Z(n12939) );
  XOR U44675 ( .A(n40849), .B(n12919), .Z(n12931) );
  XNOR U44676 ( .A(q[15]), .B(DB[3828]), .Z(n12919) );
  IV U44677 ( .A(n12918), .Z(n40849) );
  XNOR U44678 ( .A(n12916), .B(n40850), .Z(n12918) );
  XNOR U44679 ( .A(q[14]), .B(DB[3827]), .Z(n40850) );
  XNOR U44680 ( .A(q[13]), .B(DB[3826]), .Z(n12916) );
  IV U44681 ( .A(n12930), .Z(n40848) );
  XOR U44682 ( .A(n40851), .B(n40852), .Z(n12930) );
  XNOR U44683 ( .A(n12926), .B(n12928), .Z(n40852) );
  XNOR U44684 ( .A(q[9]), .B(DB[3822]), .Z(n12928) );
  XNOR U44685 ( .A(q[12]), .B(DB[3825]), .Z(n12926) );
  IV U44686 ( .A(n12925), .Z(n40851) );
  XNOR U44687 ( .A(n12923), .B(n40853), .Z(n12925) );
  XNOR U44688 ( .A(q[11]), .B(DB[3824]), .Z(n40853) );
  XNOR U44689 ( .A(q[10]), .B(DB[3823]), .Z(n12923) );
  IV U44690 ( .A(n12938), .Z(n40846) );
  XOR U44691 ( .A(n40854), .B(n40855), .Z(n12938) );
  XNOR U44692 ( .A(n12955), .B(n12936), .Z(n40855) );
  XNOR U44693 ( .A(q[1]), .B(DB[3814]), .Z(n12936) );
  XOR U44694 ( .A(n40856), .B(n12944), .Z(n12955) );
  XNOR U44695 ( .A(q[8]), .B(DB[3821]), .Z(n12944) );
  IV U44696 ( .A(n12943), .Z(n40856) );
  XNOR U44697 ( .A(n12941), .B(n40857), .Z(n12943) );
  XNOR U44698 ( .A(q[7]), .B(DB[3820]), .Z(n40857) );
  XNOR U44699 ( .A(q[6]), .B(DB[3819]), .Z(n12941) );
  IV U44700 ( .A(n12954), .Z(n40854) );
  XOR U44701 ( .A(n40858), .B(n40859), .Z(n12954) );
  XNOR U44702 ( .A(n12950), .B(n12952), .Z(n40859) );
  XNOR U44703 ( .A(q[2]), .B(DB[3815]), .Z(n12952) );
  XNOR U44704 ( .A(q[5]), .B(DB[3818]), .Z(n12950) );
  IV U44705 ( .A(n12949), .Z(n40858) );
  XNOR U44706 ( .A(n12947), .B(n40860), .Z(n12949) );
  XNOR U44707 ( .A(q[4]), .B(DB[3817]), .Z(n40860) );
  XNOR U44708 ( .A(q[3]), .B(DB[3816]), .Z(n12947) );
  XOR U44709 ( .A(n40861), .B(n12716), .Z(n12567) );
  XOR U44710 ( .A(n40862), .B(n12692), .Z(n12716) );
  XOR U44711 ( .A(n40863), .B(n12684), .Z(n12692) );
  XOR U44712 ( .A(n40864), .B(n12673), .Z(n12684) );
  XNOR U44713 ( .A(q[30]), .B(DB[3874]), .Z(n12673) );
  IV U44714 ( .A(n12672), .Z(n40864) );
  XNOR U44715 ( .A(n12670), .B(n40865), .Z(n12672) );
  XNOR U44716 ( .A(q[29]), .B(DB[3873]), .Z(n40865) );
  XNOR U44717 ( .A(q[28]), .B(DB[3872]), .Z(n12670) );
  IV U44718 ( .A(n12683), .Z(n40863) );
  XOR U44719 ( .A(n40866), .B(n40867), .Z(n12683) );
  XNOR U44720 ( .A(n12679), .B(n12681), .Z(n40867) );
  XNOR U44721 ( .A(q[24]), .B(DB[3868]), .Z(n12681) );
  XNOR U44722 ( .A(q[27]), .B(DB[3871]), .Z(n12679) );
  IV U44723 ( .A(n12678), .Z(n40866) );
  XNOR U44724 ( .A(n12676), .B(n40868), .Z(n12678) );
  XNOR U44725 ( .A(q[26]), .B(DB[3870]), .Z(n40868) );
  XNOR U44726 ( .A(q[25]), .B(DB[3869]), .Z(n12676) );
  IV U44727 ( .A(n12691), .Z(n40862) );
  XOR U44728 ( .A(n40869), .B(n40870), .Z(n12691) );
  XNOR U44729 ( .A(n12708), .B(n12689), .Z(n40870) );
  XNOR U44730 ( .A(q[16]), .B(DB[3860]), .Z(n12689) );
  XOR U44731 ( .A(n40871), .B(n12697), .Z(n12708) );
  XNOR U44732 ( .A(q[23]), .B(DB[3867]), .Z(n12697) );
  IV U44733 ( .A(n12696), .Z(n40871) );
  XNOR U44734 ( .A(n12694), .B(n40872), .Z(n12696) );
  XNOR U44735 ( .A(q[22]), .B(DB[3866]), .Z(n40872) );
  XNOR U44736 ( .A(q[21]), .B(DB[3865]), .Z(n12694) );
  IV U44737 ( .A(n12707), .Z(n40869) );
  XOR U44738 ( .A(n40873), .B(n40874), .Z(n12707) );
  XNOR U44739 ( .A(n12703), .B(n12705), .Z(n40874) );
  XNOR U44740 ( .A(q[17]), .B(DB[3861]), .Z(n12705) );
  XNOR U44741 ( .A(q[20]), .B(DB[3864]), .Z(n12703) );
  IV U44742 ( .A(n12702), .Z(n40873) );
  XNOR U44743 ( .A(n12700), .B(n40875), .Z(n12702) );
  XNOR U44744 ( .A(q[19]), .B(DB[3863]), .Z(n40875) );
  XNOR U44745 ( .A(q[18]), .B(DB[3862]), .Z(n12700) );
  IV U44746 ( .A(n12715), .Z(n40861) );
  XOR U44747 ( .A(n40876), .B(n40877), .Z(n12715) );
  XNOR U44748 ( .A(n12742), .B(n12713), .Z(n40877) );
  XNOR U44749 ( .A(q[0]), .B(DB[3844]), .Z(n12713) );
  XOR U44750 ( .A(n40878), .B(n12734), .Z(n12742) );
  XOR U44751 ( .A(n40879), .B(n12722), .Z(n12734) );
  XNOR U44752 ( .A(q[15]), .B(DB[3859]), .Z(n12722) );
  IV U44753 ( .A(n12721), .Z(n40879) );
  XNOR U44754 ( .A(n12719), .B(n40880), .Z(n12721) );
  XNOR U44755 ( .A(q[14]), .B(DB[3858]), .Z(n40880) );
  XNOR U44756 ( .A(q[13]), .B(DB[3857]), .Z(n12719) );
  IV U44757 ( .A(n12733), .Z(n40878) );
  XOR U44758 ( .A(n40881), .B(n40882), .Z(n12733) );
  XNOR U44759 ( .A(n12729), .B(n12731), .Z(n40882) );
  XNOR U44760 ( .A(q[9]), .B(DB[3853]), .Z(n12731) );
  XNOR U44761 ( .A(q[12]), .B(DB[3856]), .Z(n12729) );
  IV U44762 ( .A(n12728), .Z(n40881) );
  XNOR U44763 ( .A(n12726), .B(n40883), .Z(n12728) );
  XNOR U44764 ( .A(q[11]), .B(DB[3855]), .Z(n40883) );
  XNOR U44765 ( .A(q[10]), .B(DB[3854]), .Z(n12726) );
  IV U44766 ( .A(n12741), .Z(n40876) );
  XOR U44767 ( .A(n40884), .B(n40885), .Z(n12741) );
  XNOR U44768 ( .A(n12758), .B(n12739), .Z(n40885) );
  XNOR U44769 ( .A(q[1]), .B(DB[3845]), .Z(n12739) );
  XOR U44770 ( .A(n40886), .B(n12747), .Z(n12758) );
  XNOR U44771 ( .A(q[8]), .B(DB[3852]), .Z(n12747) );
  IV U44772 ( .A(n12746), .Z(n40886) );
  XNOR U44773 ( .A(n12744), .B(n40887), .Z(n12746) );
  XNOR U44774 ( .A(q[7]), .B(DB[3851]), .Z(n40887) );
  XNOR U44775 ( .A(q[6]), .B(DB[3850]), .Z(n12744) );
  IV U44776 ( .A(n12757), .Z(n40884) );
  XOR U44777 ( .A(n40888), .B(n40889), .Z(n12757) );
  XNOR U44778 ( .A(n12753), .B(n12755), .Z(n40889) );
  XNOR U44779 ( .A(q[2]), .B(DB[3846]), .Z(n12755) );
  XNOR U44780 ( .A(q[5]), .B(DB[3849]), .Z(n12753) );
  IV U44781 ( .A(n12752), .Z(n40888) );
  XNOR U44782 ( .A(n12750), .B(n40890), .Z(n12752) );
  XNOR U44783 ( .A(q[4]), .B(DB[3848]), .Z(n40890) );
  XNOR U44784 ( .A(q[3]), .B(DB[3847]), .Z(n12750) );
  XOR U44785 ( .A(n40891), .B(n12519), .Z(n12370) );
  XOR U44786 ( .A(n40892), .B(n12495), .Z(n12519) );
  XOR U44787 ( .A(n40893), .B(n12487), .Z(n12495) );
  XOR U44788 ( .A(n40894), .B(n12476), .Z(n12487) );
  XNOR U44789 ( .A(q[30]), .B(DB[3905]), .Z(n12476) );
  IV U44790 ( .A(n12475), .Z(n40894) );
  XNOR U44791 ( .A(n12473), .B(n40895), .Z(n12475) );
  XNOR U44792 ( .A(q[29]), .B(DB[3904]), .Z(n40895) );
  XNOR U44793 ( .A(q[28]), .B(DB[3903]), .Z(n12473) );
  IV U44794 ( .A(n12486), .Z(n40893) );
  XOR U44795 ( .A(n40896), .B(n40897), .Z(n12486) );
  XNOR U44796 ( .A(n12482), .B(n12484), .Z(n40897) );
  XNOR U44797 ( .A(q[24]), .B(DB[3899]), .Z(n12484) );
  XNOR U44798 ( .A(q[27]), .B(DB[3902]), .Z(n12482) );
  IV U44799 ( .A(n12481), .Z(n40896) );
  XNOR U44800 ( .A(n12479), .B(n40898), .Z(n12481) );
  XNOR U44801 ( .A(q[26]), .B(DB[3901]), .Z(n40898) );
  XNOR U44802 ( .A(q[25]), .B(DB[3900]), .Z(n12479) );
  IV U44803 ( .A(n12494), .Z(n40892) );
  XOR U44804 ( .A(n40899), .B(n40900), .Z(n12494) );
  XNOR U44805 ( .A(n12511), .B(n12492), .Z(n40900) );
  XNOR U44806 ( .A(q[16]), .B(DB[3891]), .Z(n12492) );
  XOR U44807 ( .A(n40901), .B(n12500), .Z(n12511) );
  XNOR U44808 ( .A(q[23]), .B(DB[3898]), .Z(n12500) );
  IV U44809 ( .A(n12499), .Z(n40901) );
  XNOR U44810 ( .A(n12497), .B(n40902), .Z(n12499) );
  XNOR U44811 ( .A(q[22]), .B(DB[3897]), .Z(n40902) );
  XNOR U44812 ( .A(q[21]), .B(DB[3896]), .Z(n12497) );
  IV U44813 ( .A(n12510), .Z(n40899) );
  XOR U44814 ( .A(n40903), .B(n40904), .Z(n12510) );
  XNOR U44815 ( .A(n12506), .B(n12508), .Z(n40904) );
  XNOR U44816 ( .A(q[17]), .B(DB[3892]), .Z(n12508) );
  XNOR U44817 ( .A(q[20]), .B(DB[3895]), .Z(n12506) );
  IV U44818 ( .A(n12505), .Z(n40903) );
  XNOR U44819 ( .A(n12503), .B(n40905), .Z(n12505) );
  XNOR U44820 ( .A(q[19]), .B(DB[3894]), .Z(n40905) );
  XNOR U44821 ( .A(q[18]), .B(DB[3893]), .Z(n12503) );
  IV U44822 ( .A(n12518), .Z(n40891) );
  XOR U44823 ( .A(n40906), .B(n40907), .Z(n12518) );
  XNOR U44824 ( .A(n12545), .B(n12516), .Z(n40907) );
  XNOR U44825 ( .A(q[0]), .B(DB[3875]), .Z(n12516) );
  XOR U44826 ( .A(n40908), .B(n12537), .Z(n12545) );
  XOR U44827 ( .A(n40909), .B(n12525), .Z(n12537) );
  XNOR U44828 ( .A(q[15]), .B(DB[3890]), .Z(n12525) );
  IV U44829 ( .A(n12524), .Z(n40909) );
  XNOR U44830 ( .A(n12522), .B(n40910), .Z(n12524) );
  XNOR U44831 ( .A(q[14]), .B(DB[3889]), .Z(n40910) );
  XNOR U44832 ( .A(q[13]), .B(DB[3888]), .Z(n12522) );
  IV U44833 ( .A(n12536), .Z(n40908) );
  XOR U44834 ( .A(n40911), .B(n40912), .Z(n12536) );
  XNOR U44835 ( .A(n12532), .B(n12534), .Z(n40912) );
  XNOR U44836 ( .A(q[9]), .B(DB[3884]), .Z(n12534) );
  XNOR U44837 ( .A(q[12]), .B(DB[3887]), .Z(n12532) );
  IV U44838 ( .A(n12531), .Z(n40911) );
  XNOR U44839 ( .A(n12529), .B(n40913), .Z(n12531) );
  XNOR U44840 ( .A(q[11]), .B(DB[3886]), .Z(n40913) );
  XNOR U44841 ( .A(q[10]), .B(DB[3885]), .Z(n12529) );
  IV U44842 ( .A(n12544), .Z(n40906) );
  XOR U44843 ( .A(n40914), .B(n40915), .Z(n12544) );
  XNOR U44844 ( .A(n12561), .B(n12542), .Z(n40915) );
  XNOR U44845 ( .A(q[1]), .B(DB[3876]), .Z(n12542) );
  XOR U44846 ( .A(n40916), .B(n12550), .Z(n12561) );
  XNOR U44847 ( .A(q[8]), .B(DB[3883]), .Z(n12550) );
  IV U44848 ( .A(n12549), .Z(n40916) );
  XNOR U44849 ( .A(n12547), .B(n40917), .Z(n12549) );
  XNOR U44850 ( .A(q[7]), .B(DB[3882]), .Z(n40917) );
  XNOR U44851 ( .A(q[6]), .B(DB[3881]), .Z(n12547) );
  IV U44852 ( .A(n12560), .Z(n40914) );
  XOR U44853 ( .A(n40918), .B(n40919), .Z(n12560) );
  XNOR U44854 ( .A(n12556), .B(n12558), .Z(n40919) );
  XNOR U44855 ( .A(q[2]), .B(DB[3877]), .Z(n12558) );
  XNOR U44856 ( .A(q[5]), .B(DB[3880]), .Z(n12556) );
  IV U44857 ( .A(n12555), .Z(n40918) );
  XNOR U44858 ( .A(n12553), .B(n40920), .Z(n12555) );
  XNOR U44859 ( .A(q[4]), .B(DB[3879]), .Z(n40920) );
  XNOR U44860 ( .A(q[3]), .B(DB[3878]), .Z(n12553) );
  XOR U44861 ( .A(n40921), .B(n12322), .Z(n12170) );
  XOR U44862 ( .A(n40922), .B(n12298), .Z(n12322) );
  XOR U44863 ( .A(n40923), .B(n12290), .Z(n12298) );
  XOR U44864 ( .A(n40924), .B(n12279), .Z(n12290) );
  XNOR U44865 ( .A(q[30]), .B(DB[3936]), .Z(n12279) );
  IV U44866 ( .A(n12278), .Z(n40924) );
  XNOR U44867 ( .A(n12276), .B(n40925), .Z(n12278) );
  XNOR U44868 ( .A(q[29]), .B(DB[3935]), .Z(n40925) );
  XOR U44869 ( .A(q[28]), .B(n3935), .Z(n12276) );
  IV U44870 ( .A(DB[3934]), .Z(n3935) );
  IV U44871 ( .A(n12289), .Z(n40923) );
  XOR U44872 ( .A(n40926), .B(n40927), .Z(n12289) );
  XNOR U44873 ( .A(n12285), .B(n12287), .Z(n40927) );
  XOR U44874 ( .A(q[24]), .B(n5461), .Z(n12287) );
  IV U44875 ( .A(DB[3930]), .Z(n5461) );
  XOR U44876 ( .A(q[27]), .B(n4317), .Z(n12285) );
  IV U44877 ( .A(DB[3933]), .Z(n4317) );
  IV U44878 ( .A(n12284), .Z(n40926) );
  XNOR U44879 ( .A(n12282), .B(n40928), .Z(n12284) );
  XNOR U44880 ( .A(q[26]), .B(DB[3932]), .Z(n40928) );
  XOR U44881 ( .A(q[25]), .B(n5079), .Z(n12282) );
  IV U44882 ( .A(DB[3931]), .Z(n5079) );
  IV U44883 ( .A(n12297), .Z(n40922) );
  XOR U44884 ( .A(n40929), .B(n40930), .Z(n12297) );
  XNOR U44885 ( .A(n12314), .B(n12295), .Z(n40930) );
  XOR U44886 ( .A(q[16]), .B(n8891), .Z(n12295) );
  IV U44887 ( .A(DB[3922]), .Z(n8891) );
  XOR U44888 ( .A(n40931), .B(n12303), .Z(n12314) );
  XNOR U44889 ( .A(q[23]), .B(DB[3929]), .Z(n12303) );
  IV U44890 ( .A(n12302), .Z(n40931) );
  XNOR U44891 ( .A(n12300), .B(n40932), .Z(n12302) );
  XNOR U44892 ( .A(q[22]), .B(DB[3928]), .Z(n40932) );
  XOR U44893 ( .A(q[21]), .B(n6603), .Z(n12300) );
  IV U44894 ( .A(DB[3927]), .Z(n6603) );
  IV U44895 ( .A(n12313), .Z(n40929) );
  XOR U44896 ( .A(n40933), .B(n40934), .Z(n12313) );
  XNOR U44897 ( .A(n12309), .B(n12311), .Z(n40934) );
  XOR U44898 ( .A(q[17]), .B(n8509), .Z(n12311) );
  IV U44899 ( .A(DB[3923]), .Z(n8509) );
  XOR U44900 ( .A(q[20]), .B(n6985), .Z(n12309) );
  IV U44901 ( .A(DB[3926]), .Z(n6985) );
  IV U44902 ( .A(n12308), .Z(n40933) );
  XNOR U44903 ( .A(n12306), .B(n40935), .Z(n12308) );
  XNOR U44904 ( .A(q[19]), .B(DB[3925]), .Z(n40935) );
  XOR U44905 ( .A(q[18]), .B(n8127), .Z(n12306) );
  IV U44906 ( .A(DB[3924]), .Z(n8127) );
  IV U44907 ( .A(n12321), .Z(n40921) );
  XOR U44908 ( .A(n40936), .B(n40937), .Z(n12321) );
  XNOR U44909 ( .A(n12348), .B(n12319), .Z(n40937) );
  XNOR U44910 ( .A(q[0]), .B(DB[3906]), .Z(n12319) );
  XOR U44911 ( .A(n40938), .B(n12340), .Z(n12348) );
  XOR U44912 ( .A(n40939), .B(n12328), .Z(n12340) );
  XNOR U44913 ( .A(q[15]), .B(DB[3921]), .Z(n12328) );
  IV U44914 ( .A(n12327), .Z(n40939) );
  XNOR U44915 ( .A(n12325), .B(n40940), .Z(n12327) );
  XNOR U44916 ( .A(q[14]), .B(DB[3920]), .Z(n40940) );
  XOR U44917 ( .A(q[13]), .B(n10033), .Z(n12325) );
  IV U44918 ( .A(DB[3919]), .Z(n10033) );
  IV U44919 ( .A(n12339), .Z(n40938) );
  XOR U44920 ( .A(n40941), .B(n40942), .Z(n12339) );
  XNOR U44921 ( .A(n12335), .B(n12337), .Z(n40942) );
  XOR U44922 ( .A(q[9]), .B(n7), .Z(n12337) );
  IV U44923 ( .A(DB[3915]), .Z(n7) );
  XOR U44924 ( .A(q[12]), .B(n10415), .Z(n12335) );
  IV U44925 ( .A(DB[3918]), .Z(n10415) );
  IV U44926 ( .A(n12334), .Z(n40941) );
  XNOR U44927 ( .A(n12332), .B(n40943), .Z(n12334) );
  XNOR U44928 ( .A(q[11]), .B(DB[3917]), .Z(n40943) );
  XOR U44929 ( .A(q[10]), .B(n11177), .Z(n12332) );
  IV U44930 ( .A(DB[3916]), .Z(n11177) );
  IV U44931 ( .A(n12347), .Z(n40936) );
  XOR U44932 ( .A(n40944), .B(n40945), .Z(n12347) );
  XNOR U44933 ( .A(n12364), .B(n12345), .Z(n40945) );
  XNOR U44934 ( .A(q[1]), .B(DB[3907]), .Z(n12345) );
  XOR U44935 ( .A(n40946), .B(n12353), .Z(n12364) );
  XNOR U44936 ( .A(q[8]), .B(DB[3914]), .Z(n12353) );
  IV U44937 ( .A(n12352), .Z(n40946) );
  XNOR U44938 ( .A(n12350), .B(n40947), .Z(n12352) );
  XNOR U44939 ( .A(q[7]), .B(DB[3913]), .Z(n40947) );
  XNOR U44940 ( .A(q[6]), .B(DB[3912]), .Z(n12350) );
  IV U44941 ( .A(n12363), .Z(n40944) );
  XOR U44942 ( .A(n40948), .B(n40949), .Z(n12363) );
  XNOR U44943 ( .A(n12359), .B(n12361), .Z(n40949) );
  XNOR U44944 ( .A(q[2]), .B(DB[3908]), .Z(n12361) );
  XNOR U44945 ( .A(q[5]), .B(DB[3911]), .Z(n12359) );
  IV U44946 ( .A(n12358), .Z(n40948) );
  XNOR U44947 ( .A(n12356), .B(n40950), .Z(n12358) );
  XNOR U44948 ( .A(q[4]), .B(DB[3910]), .Z(n40950) );
  XNOR U44949 ( .A(q[3]), .B(DB[3909]), .Z(n12356) );
endmodule

