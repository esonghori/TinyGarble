
module hamming_N160_CC8 ( clk, rst, x, y, o );
  input [19:0] x;
  input [19:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  OR U23 ( .A(n36), .B(n35), .Z(n1) );
  NANDN U24 ( .A(n38), .B(n37), .Z(n2) );
  AND U25 ( .A(n1), .B(n2), .Z(n89) );
  OR U26 ( .A(n61), .B(n60), .Z(n3) );
  NANDN U27 ( .A(n63), .B(n62), .Z(n4) );
  AND U28 ( .A(n3), .B(n4), .Z(n77) );
  OR U29 ( .A(n32), .B(n31), .Z(n5) );
  NANDN U30 ( .A(n34), .B(n33), .Z(n6) );
  NAND U31 ( .A(n5), .B(n6), .Z(n88) );
  OR U32 ( .A(n28), .B(n27), .Z(n7) );
  NANDN U33 ( .A(n30), .B(n29), .Z(n8) );
  NAND U34 ( .A(n7), .B(n8), .Z(n82) );
  OR U35 ( .A(n57), .B(n56), .Z(n9) );
  NANDN U36 ( .A(n59), .B(n58), .Z(n10) );
  NAND U37 ( .A(n9), .B(n10), .Z(n76) );
  NAND U38 ( .A(oglobal[1]), .B(n88), .Z(n11) );
  XOR U39 ( .A(n88), .B(oglobal[1]), .Z(n12) );
  NANDN U40 ( .A(n89), .B(n12), .Z(n13) );
  NAND U41 ( .A(n11), .B(n13), .Z(n90) );
  OR U42 ( .A(n53), .B(n52), .Z(n14) );
  NANDN U43 ( .A(n55), .B(n54), .Z(n15) );
  NAND U44 ( .A(n14), .B(n15), .Z(n79) );
  NANDN U45 ( .A(n21), .B(n20), .Z(n16) );
  NANDN U46 ( .A(n18), .B(n19), .Z(n17) );
  NAND U47 ( .A(n16), .B(n17), .Z(n64) );
  XNOR U48 ( .A(x[14]), .B(y[14]), .Z(n30) );
  XNOR U49 ( .A(x[18]), .B(y[18]), .Z(n28) );
  XNOR U50 ( .A(x[16]), .B(y[16]), .Z(n27) );
  XOR U51 ( .A(n28), .B(n27), .Z(n29) );
  XOR U52 ( .A(n30), .B(n29), .Z(n18) );
  XNOR U53 ( .A(x[10]), .B(y[10]), .Z(n24) );
  XOR U54 ( .A(x[12]), .B(y[12]), .Z(n22) );
  XNOR U55 ( .A(oglobal[0]), .B(n22), .Z(n23) );
  XOR U56 ( .A(n24), .B(n23), .Z(n46) );
  XNOR U57 ( .A(x[4]), .B(y[4]), .Z(n59) );
  XNOR U58 ( .A(x[8]), .B(y[8]), .Z(n57) );
  XNOR U59 ( .A(x[6]), .B(y[6]), .Z(n56) );
  XOR U60 ( .A(n57), .B(n56), .Z(n58) );
  XNOR U61 ( .A(n59), .B(n58), .Z(n47) );
  XNOR U62 ( .A(n46), .B(n47), .Z(n49) );
  XNOR U63 ( .A(x[17]), .B(y[17]), .Z(n63) );
  XNOR U64 ( .A(x[19]), .B(y[19]), .Z(n61) );
  XNOR U65 ( .A(x[15]), .B(y[15]), .Z(n60) );
  XOR U66 ( .A(n61), .B(n60), .Z(n62) );
  XNOR U67 ( .A(n63), .B(n62), .Z(n48) );
  XNOR U68 ( .A(n49), .B(n48), .Z(n19) );
  XNOR U69 ( .A(n18), .B(n19), .Z(n20) );
  XNOR U70 ( .A(x[1]), .B(y[1]), .Z(n55) );
  XNOR U71 ( .A(x[2]), .B(y[2]), .Z(n53) );
  XNOR U72 ( .A(x[0]), .B(y[0]), .Z(n52) );
  XOR U73 ( .A(n53), .B(n52), .Z(n54) );
  XNOR U74 ( .A(n55), .B(n54), .Z(n40) );
  XNOR U75 ( .A(x[13]), .B(y[13]), .Z(n38) );
  XNOR U76 ( .A(x[11]), .B(y[11]), .Z(n36) );
  XNOR U77 ( .A(x[9]), .B(y[9]), .Z(n35) );
  XOR U78 ( .A(n36), .B(n35), .Z(n37) );
  XNOR U79 ( .A(n38), .B(n37), .Z(n41) );
  XNOR U80 ( .A(n40), .B(n41), .Z(n43) );
  XNOR U81 ( .A(x[7]), .B(y[7]), .Z(n34) );
  XNOR U82 ( .A(x[5]), .B(y[5]), .Z(n32) );
  XNOR U83 ( .A(x[3]), .B(y[3]), .Z(n31) );
  XOR U84 ( .A(n32), .B(n31), .Z(n33) );
  XNOR U85 ( .A(n34), .B(n33), .Z(n42) );
  XOR U86 ( .A(n43), .B(n42), .Z(n21) );
  XNOR U87 ( .A(n20), .B(n21), .Z(o[0]) );
  NAND U88 ( .A(n22), .B(oglobal[0]), .Z(n26) );
  OR U89 ( .A(n24), .B(n23), .Z(n25) );
  NAND U90 ( .A(n26), .B(n25), .Z(n85) );
  XOR U91 ( .A(n88), .B(n89), .Z(n39) );
  XOR U92 ( .A(oglobal[1]), .B(n39), .Z(n83) );
  XNOR U93 ( .A(n82), .B(n83), .Z(n84) );
  XNOR U94 ( .A(n85), .B(n84), .Z(n65) );
  XNOR U95 ( .A(n64), .B(n65), .Z(n66) );
  OR U96 ( .A(n41), .B(n40), .Z(n45) );
  OR U97 ( .A(n43), .B(n42), .Z(n44) );
  NAND U98 ( .A(n45), .B(n44), .Z(n71) );
  OR U99 ( .A(n47), .B(n46), .Z(n51) );
  OR U100 ( .A(n49), .B(n48), .Z(n50) );
  NAND U101 ( .A(n51), .B(n50), .Z(n70) );
  XOR U102 ( .A(n71), .B(n70), .Z(n72) );
  XNOR U103 ( .A(n76), .B(n77), .Z(n78) );
  XNOR U104 ( .A(n79), .B(n78), .Z(n73) );
  XOR U105 ( .A(n72), .B(n73), .Z(n67) );
  XNOR U106 ( .A(n66), .B(n67), .Z(o[1]) );
  NANDN U107 ( .A(n65), .B(n64), .Z(n69) );
  NANDN U108 ( .A(n67), .B(n66), .Z(n68) );
  NAND U109 ( .A(n69), .B(n68), .Z(n97) );
  OR U110 ( .A(n71), .B(n70), .Z(n75) );
  NANDN U111 ( .A(n73), .B(n72), .Z(n74) );
  AND U112 ( .A(n75), .B(n74), .Z(n98) );
  XNOR U113 ( .A(n97), .B(n98), .Z(n99) );
  NANDN U114 ( .A(n77), .B(n76), .Z(n81) );
  NAND U115 ( .A(n79), .B(n78), .Z(n80) );
  NAND U116 ( .A(n81), .B(n80), .Z(n94) );
  NANDN U117 ( .A(n83), .B(n82), .Z(n87) );
  NAND U118 ( .A(n85), .B(n84), .Z(n86) );
  NAND U119 ( .A(n87), .B(n86), .Z(n91) );
  XNOR U120 ( .A(n90), .B(oglobal[2]), .Z(n92) );
  XNOR U121 ( .A(n91), .B(n92), .Z(n93) );
  XNOR U122 ( .A(n94), .B(n93), .Z(n100) );
  XNOR U123 ( .A(n99), .B(n100), .Z(o[2]) );
  NAND U124 ( .A(n90), .B(oglobal[2]), .Z(n103) );
  XOR U125 ( .A(oglobal[3]), .B(n103), .Z(n105) );
  NANDN U126 ( .A(n92), .B(n91), .Z(n96) );
  NAND U127 ( .A(n94), .B(n93), .Z(n95) );
  NAND U128 ( .A(n96), .B(n95), .Z(n104) );
  XNOR U129 ( .A(n105), .B(n104), .Z(n106) );
  NANDN U130 ( .A(n98), .B(n97), .Z(n102) );
  NANDN U131 ( .A(n100), .B(n99), .Z(n101) );
  AND U132 ( .A(n102), .B(n101), .Z(n107) );
  XNOR U133 ( .A(n106), .B(n107), .Z(o[3]) );
  NANDN U134 ( .A(n103), .B(oglobal[3]), .Z(n110) );
  XOR U135 ( .A(oglobal[4]), .B(n110), .Z(n112) );
  NANDN U136 ( .A(n105), .B(n104), .Z(n109) );
  NANDN U137 ( .A(n107), .B(n106), .Z(n108) );
  AND U138 ( .A(n109), .B(n108), .Z(n111) );
  XOR U139 ( .A(n112), .B(n111), .Z(o[4]) );
  NANDN U140 ( .A(n110), .B(oglobal[4]), .Z(n114) );
  OR U141 ( .A(n112), .B(n111), .Z(n113) );
  AND U142 ( .A(n114), .B(n113), .Z(n115) );
  XNOR U143 ( .A(oglobal[5]), .B(n115), .Z(o[5]) );
  NANDN U144 ( .A(n115), .B(oglobal[5]), .Z(n116) );
  XNOR U145 ( .A(oglobal[6]), .B(n116), .Z(o[6]) );
  NANDN U146 ( .A(n116), .B(oglobal[6]), .Z(n117) );
  XNOR U147 ( .A(oglobal[7]), .B(n117), .Z(o[7]) );
endmodule

