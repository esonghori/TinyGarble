
module modmult_step_N64_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [65:0] A;
  input [65:0] B;
  output [65:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320;

  IV U1 ( .A(n319), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(DIFF[8]) );
  XOR U6 ( .A(B[8]), .B(A[8]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[7]) );
  XOR U8 ( .A(B[7]), .B(A[7]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[6]) );
  XOR U10 ( .A(B[6]), .B(A[6]), .Z(n10) );
  XOR U11 ( .A(A[65]), .B(n11), .Z(DIFF[65]) );
  ANDN U12 ( .B(n12), .A(A[64]), .Z(n11) );
  XOR U13 ( .A(A[64]), .B(n12), .Z(DIFF[64]) );
  AND U14 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U15 ( .A(B[63]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(A[63]), .B(n16), .Z(n15) );
  NANDN U17 ( .A(n16), .B(A[63]), .Z(n13) );
  XOR U18 ( .A(n16), .B(n17), .Z(DIFF[63]) );
  XOR U19 ( .A(B[63]), .B(A[63]), .Z(n17) );
  AND U20 ( .A(n18), .B(n19), .Z(n16) );
  NANDN U21 ( .A(B[62]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(A[62]), .B(n21), .Z(n20) );
  NANDN U23 ( .A(n21), .B(A[62]), .Z(n18) );
  XOR U24 ( .A(n21), .B(n22), .Z(DIFF[62]) );
  XOR U25 ( .A(B[62]), .B(A[62]), .Z(n22) );
  AND U26 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U27 ( .A(B[61]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(A[61]), .B(n26), .Z(n25) );
  NANDN U29 ( .A(n26), .B(A[61]), .Z(n23) );
  XOR U30 ( .A(n26), .B(n27), .Z(DIFF[61]) );
  XOR U31 ( .A(B[61]), .B(A[61]), .Z(n27) );
  AND U32 ( .A(n28), .B(n29), .Z(n26) );
  NANDN U33 ( .A(B[60]), .B(n30), .Z(n29) );
  NANDN U34 ( .A(A[60]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(n31), .B(A[60]), .Z(n28) );
  XOR U36 ( .A(n31), .B(n32), .Z(DIFF[60]) );
  XOR U37 ( .A(B[60]), .B(A[60]), .Z(n32) );
  AND U38 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U39 ( .A(B[59]), .B(n35), .Z(n34) );
  NANDN U40 ( .A(A[59]), .B(n36), .Z(n35) );
  NANDN U41 ( .A(n36), .B(A[59]), .Z(n33) );
  XOR U42 ( .A(n37), .B(n38), .Z(DIFF[5]) );
  XOR U43 ( .A(B[5]), .B(A[5]), .Z(n38) );
  XOR U44 ( .A(n36), .B(n39), .Z(DIFF[59]) );
  XOR U45 ( .A(B[59]), .B(A[59]), .Z(n39) );
  AND U46 ( .A(n40), .B(n41), .Z(n36) );
  NANDN U47 ( .A(B[58]), .B(n42), .Z(n41) );
  NANDN U48 ( .A(A[58]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(n43), .B(A[58]), .Z(n40) );
  XOR U50 ( .A(n43), .B(n44), .Z(DIFF[58]) );
  XOR U51 ( .A(B[58]), .B(A[58]), .Z(n44) );
  AND U52 ( .A(n45), .B(n46), .Z(n43) );
  NANDN U53 ( .A(B[57]), .B(n47), .Z(n46) );
  NANDN U54 ( .A(A[57]), .B(n48), .Z(n47) );
  NANDN U55 ( .A(n48), .B(A[57]), .Z(n45) );
  XOR U56 ( .A(n48), .B(n49), .Z(DIFF[57]) );
  XOR U57 ( .A(B[57]), .B(A[57]), .Z(n49) );
  AND U58 ( .A(n50), .B(n51), .Z(n48) );
  NANDN U59 ( .A(B[56]), .B(n52), .Z(n51) );
  NANDN U60 ( .A(A[56]), .B(n53), .Z(n52) );
  NANDN U61 ( .A(n53), .B(A[56]), .Z(n50) );
  XOR U62 ( .A(n53), .B(n54), .Z(DIFF[56]) );
  XOR U63 ( .A(B[56]), .B(A[56]), .Z(n54) );
  AND U64 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U65 ( .A(B[55]), .B(n57), .Z(n56) );
  NANDN U66 ( .A(A[55]), .B(n58), .Z(n57) );
  NANDN U67 ( .A(n58), .B(A[55]), .Z(n55) );
  XOR U68 ( .A(n58), .B(n59), .Z(DIFF[55]) );
  XOR U69 ( .A(B[55]), .B(A[55]), .Z(n59) );
  AND U70 ( .A(n60), .B(n61), .Z(n58) );
  NANDN U71 ( .A(B[54]), .B(n62), .Z(n61) );
  NANDN U72 ( .A(A[54]), .B(n63), .Z(n62) );
  NANDN U73 ( .A(n63), .B(A[54]), .Z(n60) );
  XOR U74 ( .A(n63), .B(n64), .Z(DIFF[54]) );
  XOR U75 ( .A(B[54]), .B(A[54]), .Z(n64) );
  AND U76 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U77 ( .A(B[53]), .B(n67), .Z(n66) );
  NANDN U78 ( .A(A[53]), .B(n68), .Z(n67) );
  NANDN U79 ( .A(n68), .B(A[53]), .Z(n65) );
  XOR U80 ( .A(n68), .B(n69), .Z(DIFF[53]) );
  XOR U81 ( .A(B[53]), .B(A[53]), .Z(n69) );
  AND U82 ( .A(n70), .B(n71), .Z(n68) );
  NANDN U83 ( .A(B[52]), .B(n72), .Z(n71) );
  NANDN U84 ( .A(A[52]), .B(n73), .Z(n72) );
  NANDN U85 ( .A(n73), .B(A[52]), .Z(n70) );
  XOR U86 ( .A(n73), .B(n74), .Z(DIFF[52]) );
  XOR U87 ( .A(B[52]), .B(A[52]), .Z(n74) );
  AND U88 ( .A(n75), .B(n76), .Z(n73) );
  NANDN U89 ( .A(B[51]), .B(n77), .Z(n76) );
  NANDN U90 ( .A(A[51]), .B(n78), .Z(n77) );
  NANDN U91 ( .A(n78), .B(A[51]), .Z(n75) );
  XOR U92 ( .A(n78), .B(n79), .Z(DIFF[51]) );
  XOR U93 ( .A(B[51]), .B(A[51]), .Z(n79) );
  AND U94 ( .A(n80), .B(n81), .Z(n78) );
  NANDN U95 ( .A(B[50]), .B(n82), .Z(n81) );
  NANDN U96 ( .A(A[50]), .B(n83), .Z(n82) );
  NANDN U97 ( .A(n83), .B(A[50]), .Z(n80) );
  XOR U98 ( .A(n83), .B(n84), .Z(DIFF[50]) );
  XOR U99 ( .A(B[50]), .B(A[50]), .Z(n84) );
  AND U100 ( .A(n85), .B(n86), .Z(n83) );
  NANDN U101 ( .A(B[49]), .B(n87), .Z(n86) );
  NANDN U102 ( .A(A[49]), .B(n88), .Z(n87) );
  NANDN U103 ( .A(n88), .B(A[49]), .Z(n85) );
  XOR U104 ( .A(n89), .B(n90), .Z(DIFF[4]) );
  XOR U105 ( .A(B[4]), .B(A[4]), .Z(n90) );
  XOR U106 ( .A(n88), .B(n91), .Z(DIFF[49]) );
  XOR U107 ( .A(B[49]), .B(A[49]), .Z(n91) );
  AND U108 ( .A(n92), .B(n93), .Z(n88) );
  NANDN U109 ( .A(B[48]), .B(n94), .Z(n93) );
  NANDN U110 ( .A(A[48]), .B(n95), .Z(n94) );
  NANDN U111 ( .A(n95), .B(A[48]), .Z(n92) );
  XOR U112 ( .A(n95), .B(n96), .Z(DIFF[48]) );
  XOR U113 ( .A(B[48]), .B(A[48]), .Z(n96) );
  AND U114 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U115 ( .A(B[47]), .B(n99), .Z(n98) );
  NANDN U116 ( .A(A[47]), .B(n100), .Z(n99) );
  NANDN U117 ( .A(n100), .B(A[47]), .Z(n97) );
  XOR U118 ( .A(n100), .B(n101), .Z(DIFF[47]) );
  XOR U119 ( .A(B[47]), .B(A[47]), .Z(n101) );
  AND U120 ( .A(n102), .B(n103), .Z(n100) );
  NANDN U121 ( .A(B[46]), .B(n104), .Z(n103) );
  NANDN U122 ( .A(A[46]), .B(n105), .Z(n104) );
  NANDN U123 ( .A(n105), .B(A[46]), .Z(n102) );
  XOR U124 ( .A(n105), .B(n106), .Z(DIFF[46]) );
  XOR U125 ( .A(B[46]), .B(A[46]), .Z(n106) );
  AND U126 ( .A(n107), .B(n108), .Z(n105) );
  NANDN U127 ( .A(B[45]), .B(n109), .Z(n108) );
  NANDN U128 ( .A(A[45]), .B(n110), .Z(n109) );
  NANDN U129 ( .A(n110), .B(A[45]), .Z(n107) );
  XOR U130 ( .A(n110), .B(n111), .Z(DIFF[45]) );
  XOR U131 ( .A(B[45]), .B(A[45]), .Z(n111) );
  AND U132 ( .A(n112), .B(n113), .Z(n110) );
  NANDN U133 ( .A(B[44]), .B(n114), .Z(n113) );
  NANDN U134 ( .A(A[44]), .B(n115), .Z(n114) );
  NANDN U135 ( .A(n115), .B(A[44]), .Z(n112) );
  XOR U136 ( .A(n115), .B(n116), .Z(DIFF[44]) );
  XOR U137 ( .A(B[44]), .B(A[44]), .Z(n116) );
  AND U138 ( .A(n117), .B(n118), .Z(n115) );
  NANDN U139 ( .A(B[43]), .B(n119), .Z(n118) );
  NANDN U140 ( .A(A[43]), .B(n120), .Z(n119) );
  NANDN U141 ( .A(n120), .B(A[43]), .Z(n117) );
  XOR U142 ( .A(n120), .B(n121), .Z(DIFF[43]) );
  XOR U143 ( .A(B[43]), .B(A[43]), .Z(n121) );
  AND U144 ( .A(n122), .B(n123), .Z(n120) );
  NANDN U145 ( .A(B[42]), .B(n124), .Z(n123) );
  NANDN U146 ( .A(A[42]), .B(n125), .Z(n124) );
  NANDN U147 ( .A(n125), .B(A[42]), .Z(n122) );
  XOR U148 ( .A(n125), .B(n126), .Z(DIFF[42]) );
  XOR U149 ( .A(B[42]), .B(A[42]), .Z(n126) );
  AND U150 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U151 ( .A(B[41]), .B(n129), .Z(n128) );
  NANDN U152 ( .A(A[41]), .B(n130), .Z(n129) );
  NANDN U153 ( .A(n130), .B(A[41]), .Z(n127) );
  XOR U154 ( .A(n130), .B(n131), .Z(DIFF[41]) );
  XOR U155 ( .A(B[41]), .B(A[41]), .Z(n131) );
  AND U156 ( .A(n132), .B(n133), .Z(n130) );
  NANDN U157 ( .A(B[40]), .B(n134), .Z(n133) );
  NANDN U158 ( .A(A[40]), .B(n135), .Z(n134) );
  NANDN U159 ( .A(n135), .B(A[40]), .Z(n132) );
  XOR U160 ( .A(n135), .B(n136), .Z(DIFF[40]) );
  XOR U161 ( .A(B[40]), .B(A[40]), .Z(n136) );
  AND U162 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U163 ( .A(B[39]), .B(n139), .Z(n138) );
  NANDN U164 ( .A(A[39]), .B(n140), .Z(n139) );
  NANDN U165 ( .A(n140), .B(A[39]), .Z(n137) );
  XOR U166 ( .A(n141), .B(n142), .Z(DIFF[3]) );
  XOR U167 ( .A(B[3]), .B(A[3]), .Z(n142) );
  XOR U168 ( .A(n140), .B(n143), .Z(DIFF[39]) );
  XOR U169 ( .A(B[39]), .B(A[39]), .Z(n143) );
  AND U170 ( .A(n144), .B(n145), .Z(n140) );
  NANDN U171 ( .A(B[38]), .B(n146), .Z(n145) );
  NANDN U172 ( .A(A[38]), .B(n147), .Z(n146) );
  NANDN U173 ( .A(n147), .B(A[38]), .Z(n144) );
  XOR U174 ( .A(n147), .B(n148), .Z(DIFF[38]) );
  XOR U175 ( .A(B[38]), .B(A[38]), .Z(n148) );
  AND U176 ( .A(n149), .B(n150), .Z(n147) );
  NANDN U177 ( .A(B[37]), .B(n151), .Z(n150) );
  NANDN U178 ( .A(A[37]), .B(n152), .Z(n151) );
  NANDN U179 ( .A(n152), .B(A[37]), .Z(n149) );
  XOR U180 ( .A(n152), .B(n153), .Z(DIFF[37]) );
  XOR U181 ( .A(B[37]), .B(A[37]), .Z(n153) );
  AND U182 ( .A(n154), .B(n155), .Z(n152) );
  NANDN U183 ( .A(B[36]), .B(n156), .Z(n155) );
  NANDN U184 ( .A(A[36]), .B(n157), .Z(n156) );
  NANDN U185 ( .A(n157), .B(A[36]), .Z(n154) );
  XOR U186 ( .A(n157), .B(n158), .Z(DIFF[36]) );
  XOR U187 ( .A(B[36]), .B(A[36]), .Z(n158) );
  AND U188 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U189 ( .A(B[35]), .B(n161), .Z(n160) );
  NANDN U190 ( .A(A[35]), .B(n162), .Z(n161) );
  NANDN U191 ( .A(n162), .B(A[35]), .Z(n159) );
  XOR U192 ( .A(n162), .B(n163), .Z(DIFF[35]) );
  XOR U193 ( .A(B[35]), .B(A[35]), .Z(n163) );
  AND U194 ( .A(n164), .B(n165), .Z(n162) );
  NANDN U195 ( .A(B[34]), .B(n166), .Z(n165) );
  NANDN U196 ( .A(A[34]), .B(n167), .Z(n166) );
  NANDN U197 ( .A(n167), .B(A[34]), .Z(n164) );
  XOR U198 ( .A(n167), .B(n168), .Z(DIFF[34]) );
  XOR U199 ( .A(B[34]), .B(A[34]), .Z(n168) );
  AND U200 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U201 ( .A(B[33]), .B(n171), .Z(n170) );
  NANDN U202 ( .A(A[33]), .B(n172), .Z(n171) );
  NANDN U203 ( .A(n172), .B(A[33]), .Z(n169) );
  XOR U204 ( .A(n172), .B(n173), .Z(DIFF[33]) );
  XOR U205 ( .A(B[33]), .B(A[33]), .Z(n173) );
  AND U206 ( .A(n174), .B(n175), .Z(n172) );
  NANDN U207 ( .A(B[32]), .B(n176), .Z(n175) );
  NANDN U208 ( .A(A[32]), .B(n177), .Z(n176) );
  NANDN U209 ( .A(n177), .B(A[32]), .Z(n174) );
  XOR U210 ( .A(n177), .B(n178), .Z(DIFF[32]) );
  XOR U211 ( .A(B[32]), .B(A[32]), .Z(n178) );
  AND U212 ( .A(n179), .B(n180), .Z(n177) );
  NANDN U213 ( .A(B[31]), .B(n181), .Z(n180) );
  NANDN U214 ( .A(A[31]), .B(n182), .Z(n181) );
  NANDN U215 ( .A(n182), .B(A[31]), .Z(n179) );
  XOR U216 ( .A(n182), .B(n183), .Z(DIFF[31]) );
  XOR U217 ( .A(B[31]), .B(A[31]), .Z(n183) );
  AND U218 ( .A(n184), .B(n185), .Z(n182) );
  NANDN U219 ( .A(B[30]), .B(n186), .Z(n185) );
  NANDN U220 ( .A(A[30]), .B(n187), .Z(n186) );
  NANDN U221 ( .A(n187), .B(A[30]), .Z(n184) );
  XOR U222 ( .A(n187), .B(n188), .Z(DIFF[30]) );
  XOR U223 ( .A(B[30]), .B(A[30]), .Z(n188) );
  AND U224 ( .A(n189), .B(n190), .Z(n187) );
  NANDN U225 ( .A(B[29]), .B(n191), .Z(n190) );
  NANDN U226 ( .A(A[29]), .B(n192), .Z(n191) );
  NANDN U227 ( .A(n192), .B(A[29]), .Z(n189) );
  XOR U228 ( .A(n193), .B(n194), .Z(DIFF[2]) );
  XOR U229 ( .A(B[2]), .B(A[2]), .Z(n194) );
  XOR U230 ( .A(n192), .B(n195), .Z(DIFF[29]) );
  XOR U231 ( .A(B[29]), .B(A[29]), .Z(n195) );
  AND U232 ( .A(n196), .B(n197), .Z(n192) );
  NANDN U233 ( .A(B[28]), .B(n198), .Z(n197) );
  NANDN U234 ( .A(A[28]), .B(n199), .Z(n198) );
  NANDN U235 ( .A(n199), .B(A[28]), .Z(n196) );
  XOR U236 ( .A(n199), .B(n200), .Z(DIFF[28]) );
  XOR U237 ( .A(B[28]), .B(A[28]), .Z(n200) );
  AND U238 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U239 ( .A(B[27]), .B(n203), .Z(n202) );
  NANDN U240 ( .A(A[27]), .B(n204), .Z(n203) );
  NANDN U241 ( .A(n204), .B(A[27]), .Z(n201) );
  XOR U242 ( .A(n204), .B(n205), .Z(DIFF[27]) );
  XOR U243 ( .A(B[27]), .B(A[27]), .Z(n205) );
  AND U244 ( .A(n206), .B(n207), .Z(n204) );
  NANDN U245 ( .A(B[26]), .B(n208), .Z(n207) );
  NANDN U246 ( .A(A[26]), .B(n209), .Z(n208) );
  NANDN U247 ( .A(n209), .B(A[26]), .Z(n206) );
  XOR U248 ( .A(n209), .B(n210), .Z(DIFF[26]) );
  XOR U249 ( .A(B[26]), .B(A[26]), .Z(n210) );
  AND U250 ( .A(n211), .B(n212), .Z(n209) );
  NANDN U251 ( .A(B[25]), .B(n213), .Z(n212) );
  NANDN U252 ( .A(A[25]), .B(n214), .Z(n213) );
  NANDN U253 ( .A(n214), .B(A[25]), .Z(n211) );
  XOR U254 ( .A(n214), .B(n215), .Z(DIFF[25]) );
  XOR U255 ( .A(B[25]), .B(A[25]), .Z(n215) );
  AND U256 ( .A(n216), .B(n217), .Z(n214) );
  NANDN U257 ( .A(B[24]), .B(n218), .Z(n217) );
  NANDN U258 ( .A(A[24]), .B(n219), .Z(n218) );
  NANDN U259 ( .A(n219), .B(A[24]), .Z(n216) );
  XOR U260 ( .A(n219), .B(n220), .Z(DIFF[24]) );
  XOR U261 ( .A(B[24]), .B(A[24]), .Z(n220) );
  AND U262 ( .A(n221), .B(n222), .Z(n219) );
  NANDN U263 ( .A(B[23]), .B(n223), .Z(n222) );
  NANDN U264 ( .A(A[23]), .B(n224), .Z(n223) );
  NANDN U265 ( .A(n224), .B(A[23]), .Z(n221) );
  XOR U266 ( .A(n224), .B(n225), .Z(DIFF[23]) );
  XOR U267 ( .A(B[23]), .B(A[23]), .Z(n225) );
  AND U268 ( .A(n226), .B(n227), .Z(n224) );
  NANDN U269 ( .A(B[22]), .B(n228), .Z(n227) );
  NANDN U270 ( .A(A[22]), .B(n229), .Z(n228) );
  NANDN U271 ( .A(n229), .B(A[22]), .Z(n226) );
  XOR U272 ( .A(n229), .B(n230), .Z(DIFF[22]) );
  XOR U273 ( .A(B[22]), .B(A[22]), .Z(n230) );
  AND U274 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U275 ( .A(B[21]), .B(n233), .Z(n232) );
  NANDN U276 ( .A(A[21]), .B(n234), .Z(n233) );
  NANDN U277 ( .A(n234), .B(A[21]), .Z(n231) );
  XOR U278 ( .A(n234), .B(n235), .Z(DIFF[21]) );
  XOR U279 ( .A(B[21]), .B(A[21]), .Z(n235) );
  AND U280 ( .A(n236), .B(n237), .Z(n234) );
  NANDN U281 ( .A(B[20]), .B(n238), .Z(n237) );
  NANDN U282 ( .A(A[20]), .B(n239), .Z(n238) );
  NANDN U283 ( .A(n239), .B(A[20]), .Z(n236) );
  XOR U284 ( .A(n239), .B(n240), .Z(DIFF[20]) );
  XOR U285 ( .A(B[20]), .B(A[20]), .Z(n240) );
  AND U286 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U287 ( .A(B[19]), .B(n243), .Z(n242) );
  NANDN U288 ( .A(A[19]), .B(n244), .Z(n243) );
  NANDN U289 ( .A(n244), .B(A[19]), .Z(n241) );
  XOR U290 ( .A(n1), .B(n245), .Z(DIFF[1]) );
  XOR U291 ( .A(B[1]), .B(A[1]), .Z(n245) );
  XOR U292 ( .A(n244), .B(n246), .Z(DIFF[19]) );
  XOR U293 ( .A(B[19]), .B(A[19]), .Z(n246) );
  AND U294 ( .A(n247), .B(n248), .Z(n244) );
  NANDN U295 ( .A(B[18]), .B(n249), .Z(n248) );
  NANDN U296 ( .A(A[18]), .B(n250), .Z(n249) );
  NANDN U297 ( .A(n250), .B(A[18]), .Z(n247) );
  XOR U298 ( .A(n250), .B(n251), .Z(DIFF[18]) );
  XOR U299 ( .A(B[18]), .B(A[18]), .Z(n251) );
  AND U300 ( .A(n252), .B(n253), .Z(n250) );
  NANDN U301 ( .A(B[17]), .B(n254), .Z(n253) );
  NANDN U302 ( .A(A[17]), .B(n255), .Z(n254) );
  NANDN U303 ( .A(n255), .B(A[17]), .Z(n252) );
  XOR U304 ( .A(n255), .B(n256), .Z(DIFF[17]) );
  XOR U305 ( .A(B[17]), .B(A[17]), .Z(n256) );
  AND U306 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U307 ( .A(B[16]), .B(n259), .Z(n258) );
  NANDN U308 ( .A(A[16]), .B(n260), .Z(n259) );
  NANDN U309 ( .A(n260), .B(A[16]), .Z(n257) );
  XOR U310 ( .A(n260), .B(n261), .Z(DIFF[16]) );
  XOR U311 ( .A(B[16]), .B(A[16]), .Z(n261) );
  AND U312 ( .A(n262), .B(n263), .Z(n260) );
  NANDN U313 ( .A(B[15]), .B(n264), .Z(n263) );
  NANDN U314 ( .A(A[15]), .B(n265), .Z(n264) );
  NANDN U315 ( .A(n265), .B(A[15]), .Z(n262) );
  XOR U316 ( .A(n265), .B(n266), .Z(DIFF[15]) );
  XOR U317 ( .A(B[15]), .B(A[15]), .Z(n266) );
  AND U318 ( .A(n267), .B(n268), .Z(n265) );
  NANDN U319 ( .A(B[14]), .B(n269), .Z(n268) );
  NANDN U320 ( .A(A[14]), .B(n270), .Z(n269) );
  NANDN U321 ( .A(n270), .B(A[14]), .Z(n267) );
  XOR U322 ( .A(n270), .B(n271), .Z(DIFF[14]) );
  XOR U323 ( .A(B[14]), .B(A[14]), .Z(n271) );
  AND U324 ( .A(n272), .B(n273), .Z(n270) );
  NANDN U325 ( .A(B[13]), .B(n274), .Z(n273) );
  NANDN U326 ( .A(A[13]), .B(n275), .Z(n274) );
  NANDN U327 ( .A(n275), .B(A[13]), .Z(n272) );
  XOR U328 ( .A(n275), .B(n276), .Z(DIFF[13]) );
  XOR U329 ( .A(B[13]), .B(A[13]), .Z(n276) );
  AND U330 ( .A(n277), .B(n278), .Z(n275) );
  NANDN U331 ( .A(B[12]), .B(n279), .Z(n278) );
  NANDN U332 ( .A(A[12]), .B(n280), .Z(n279) );
  NANDN U333 ( .A(n280), .B(A[12]), .Z(n277) );
  XOR U334 ( .A(n280), .B(n281), .Z(DIFF[12]) );
  XOR U335 ( .A(B[12]), .B(A[12]), .Z(n281) );
  AND U336 ( .A(n282), .B(n283), .Z(n280) );
  NANDN U337 ( .A(B[11]), .B(n284), .Z(n283) );
  NANDN U338 ( .A(A[11]), .B(n285), .Z(n284) );
  NANDN U339 ( .A(n285), .B(A[11]), .Z(n282) );
  XOR U340 ( .A(n285), .B(n286), .Z(DIFF[11]) );
  XOR U341 ( .A(B[11]), .B(A[11]), .Z(n286) );
  AND U342 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U343 ( .A(B[10]), .B(n289), .Z(n288) );
  NANDN U344 ( .A(A[10]), .B(n290), .Z(n289) );
  NANDN U345 ( .A(n290), .B(A[10]), .Z(n287) );
  XOR U346 ( .A(n290), .B(n291), .Z(DIFF[10]) );
  XOR U347 ( .A(B[10]), .B(A[10]), .Z(n291) );
  AND U348 ( .A(n292), .B(n293), .Z(n290) );
  NANDN U349 ( .A(B[9]), .B(n294), .Z(n293) );
  OR U350 ( .A(n3), .B(A[9]), .Z(n294) );
  NAND U351 ( .A(A[9]), .B(n3), .Z(n292) );
  NAND U352 ( .A(n295), .B(n296), .Z(n3) );
  NANDN U353 ( .A(B[8]), .B(n297), .Z(n296) );
  NANDN U354 ( .A(A[8]), .B(n5), .Z(n297) );
  NANDN U355 ( .A(n5), .B(A[8]), .Z(n295) );
  AND U356 ( .A(n298), .B(n299), .Z(n5) );
  NANDN U357 ( .A(B[7]), .B(n300), .Z(n299) );
  NANDN U358 ( .A(A[7]), .B(n7), .Z(n300) );
  NANDN U359 ( .A(n7), .B(A[7]), .Z(n298) );
  AND U360 ( .A(n301), .B(n302), .Z(n7) );
  NANDN U361 ( .A(B[6]), .B(n303), .Z(n302) );
  NANDN U362 ( .A(A[6]), .B(n9), .Z(n303) );
  NANDN U363 ( .A(n9), .B(A[6]), .Z(n301) );
  AND U364 ( .A(n304), .B(n305), .Z(n9) );
  NANDN U365 ( .A(B[5]), .B(n306), .Z(n305) );
  NANDN U366 ( .A(A[5]), .B(n37), .Z(n306) );
  NANDN U367 ( .A(n37), .B(A[5]), .Z(n304) );
  AND U368 ( .A(n307), .B(n308), .Z(n37) );
  NANDN U369 ( .A(B[4]), .B(n309), .Z(n308) );
  NANDN U370 ( .A(A[4]), .B(n89), .Z(n309) );
  NANDN U371 ( .A(n89), .B(A[4]), .Z(n307) );
  AND U372 ( .A(n310), .B(n311), .Z(n89) );
  NANDN U373 ( .A(B[3]), .B(n312), .Z(n311) );
  NANDN U374 ( .A(A[3]), .B(n141), .Z(n312) );
  NANDN U375 ( .A(n141), .B(A[3]), .Z(n310) );
  AND U376 ( .A(n313), .B(n314), .Z(n141) );
  NANDN U377 ( .A(B[2]), .B(n315), .Z(n314) );
  NANDN U378 ( .A(A[2]), .B(n193), .Z(n315) );
  NANDN U379 ( .A(n193), .B(A[2]), .Z(n313) );
  AND U380 ( .A(n316), .B(n317), .Z(n193) );
  NANDN U381 ( .A(B[1]), .B(n318), .Z(n317) );
  NAND U382 ( .A(n1), .B(n2), .Z(n318) );
  NAND U383 ( .A(A[1]), .B(n319), .Z(n316) );
  NAND U384 ( .A(n319), .B(n320), .Z(DIFF[0]) );
  NANDN U385 ( .A(B[0]), .B(A[0]), .Z(n320) );
  NANDN U386 ( .A(A[0]), .B(B[0]), .Z(n319) );
endmodule


module modmult_step_N64_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [63:0] A;
  input [0:0] B;
  output [64:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U3 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U4 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U5 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U6 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U7 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U8 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U9 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U10 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U11 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U12 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U13 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U14 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U15 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U16 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U17 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U18 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U19 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U20 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U21 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U22 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U23 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U24 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U25 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U26 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U27 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U28 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U29 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U30 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U31 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U32 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U33 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U34 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U35 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U36 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U37 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U38 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U39 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U40 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U41 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U42 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U43 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U44 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U45 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U46 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U47 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U48 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U49 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U50 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U51 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U52 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U53 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U54 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U55 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U56 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U57 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U58 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U59 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U60 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U61 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U62 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U63 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U64 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U65 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N64_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [65:0] A;
  input [65:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[65]), .B(B[64]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[63]), .B(A[63]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[62]), .B(B[62]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[62]), .B(A[62]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[61]), .B(B[61]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[60]), .B(B[60]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[60]), .B(A[60]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[59]), .B(B[59]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[58]), .B(B[58]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[58]), .B(A[58]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[57]), .B(B[57]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[56]), .B(B[56]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[56]), .B(A[56]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[55]), .B(B[55]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[54]), .B(B[54]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[54]), .B(A[54]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[53]), .B(B[53]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[52]), .B(B[52]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[52]), .B(A[52]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[51]), .B(B[51]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[50]), .B(B[50]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[50]), .B(A[50]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[49]), .B(B[49]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[48]), .B(B[48]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[48]), .B(A[48]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[47]), .B(B[47]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[46]), .B(B[46]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[46]), .B(A[46]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[45]), .B(B[45]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[44]), .B(B[44]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[44]), .B(A[44]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[43]), .B(B[43]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[42]), .B(B[42]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[42]), .B(A[42]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[41]), .B(B[41]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[40]), .B(B[40]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[40]), .B(A[40]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[39]), .B(B[39]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[38]), .B(B[38]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[38]), .B(A[38]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[37]), .B(B[37]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[36]), .B(B[36]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[36]), .B(A[36]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[35]), .B(B[35]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[34]), .B(B[34]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[34]), .B(A[34]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[33]), .B(B[33]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[32]), .B(B[32]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[32]), .B(A[32]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[31]), .B(B[31]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[30]), .B(B[30]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[30]), .B(A[30]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[29]), .B(B[29]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[28]), .B(B[28]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[28]), .B(A[28]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[27]), .B(B[27]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[26]), .B(B[26]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[26]), .B(A[26]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[25]), .B(B[25]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[24]), .B(B[24]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[24]), .B(A[24]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[23]), .B(B[23]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[22]), .B(B[22]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[22]), .B(A[22]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[21]), .B(B[21]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[20]), .B(B[20]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[20]), .B(A[20]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[19]), .B(B[19]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[18]), .B(B[18]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[18]), .B(A[18]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[17]), .B(B[17]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[16]), .B(B[16]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[16]), .B(A[16]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[15]), .B(B[15]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[14]), .B(B[14]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[14]), .B(A[14]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[13]), .B(B[13]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[12]), .B(B[12]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[12]), .B(A[12]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[11]), .B(B[11]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[10]), .B(B[10]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[9]), .B(A[9]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[9]), .B(B[9]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[8]), .B(B[8]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[8]), .B(A[8]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[7]), .B(B[7]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[6]), .B(B[6]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[6]), .B(A[6]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[5]), .B(B[5]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[4]), .B(B[4]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[4]), .B(A[4]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[3]), .B(B[3]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[2]), .B(B[2]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[2]), .B(A[2]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(A[0]), .Z(n252) );
  ANDN U222 ( .B(n254), .A(B[0]), .Z(n253) );
  NANDN U223 ( .A(A[1]), .B(B[1]), .Z(n254) );
  NANDN U224 ( .A(B[1]), .B(A[1]), .Z(n251) );
  NANDN U225 ( .A(B[3]), .B(A[3]), .Z(n243) );
  NANDN U226 ( .A(B[5]), .B(A[5]), .Z(n235) );
  NANDN U227 ( .A(B[7]), .B(A[7]), .Z(n227) );
  NANDN U228 ( .A(B[10]), .B(A[10]), .Z(n219) );
  NANDN U229 ( .A(B[11]), .B(A[11]), .Z(n211) );
  NANDN U230 ( .A(B[13]), .B(A[13]), .Z(n203) );
  NANDN U231 ( .A(B[15]), .B(A[15]), .Z(n195) );
  NANDN U232 ( .A(B[17]), .B(A[17]), .Z(n187) );
  NANDN U233 ( .A(B[19]), .B(A[19]), .Z(n179) );
  NANDN U234 ( .A(B[21]), .B(A[21]), .Z(n171) );
  NANDN U235 ( .A(B[23]), .B(A[23]), .Z(n163) );
  NANDN U236 ( .A(B[25]), .B(A[25]), .Z(n155) );
  NANDN U237 ( .A(B[27]), .B(A[27]), .Z(n147) );
  NANDN U238 ( .A(B[29]), .B(A[29]), .Z(n139) );
  NANDN U239 ( .A(B[31]), .B(A[31]), .Z(n131) );
  NANDN U240 ( .A(B[33]), .B(A[33]), .Z(n123) );
  NANDN U241 ( .A(B[35]), .B(A[35]), .Z(n115) );
  NANDN U242 ( .A(B[37]), .B(A[37]), .Z(n107) );
  NANDN U243 ( .A(B[39]), .B(A[39]), .Z(n99) );
  NANDN U244 ( .A(B[41]), .B(A[41]), .Z(n91) );
  NANDN U245 ( .A(B[43]), .B(A[43]), .Z(n83) );
  NANDN U246 ( .A(B[45]), .B(A[45]), .Z(n75) );
  NANDN U247 ( .A(B[47]), .B(A[47]), .Z(n67) );
  NANDN U248 ( .A(B[49]), .B(A[49]), .Z(n59) );
  NANDN U249 ( .A(B[51]), .B(A[51]), .Z(n51) );
  NANDN U250 ( .A(B[53]), .B(A[53]), .Z(n43) );
  NANDN U251 ( .A(B[55]), .B(A[55]), .Z(n35) );
  NANDN U252 ( .A(B[57]), .B(A[57]), .Z(n27) );
  NANDN U253 ( .A(B[59]), .B(A[59]), .Z(n19) );
  NANDN U254 ( .A(B[61]), .B(A[61]), .Z(n11) );
  NANDN U255 ( .A(A[63]), .B(B[63]), .Z(n3) );
endmodule


module modmult_step_N64_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [65:0] A;
  input [65:0] B;
  output [65:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n319), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(DIFF[8]) );
  XOR U6 ( .A(B[8]), .B(A[8]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[7]) );
  XOR U8 ( .A(B[7]), .B(A[7]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[6]) );
  XOR U10 ( .A(B[6]), .B(A[6]), .Z(n10) );
  XOR U11 ( .A(A[65]), .B(n11), .Z(DIFF[65]) );
  ANDN U12 ( .B(n12), .A(A[64]), .Z(n11) );
  XOR U13 ( .A(A[64]), .B(n12), .Z(DIFF[64]) );
  AND U14 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U15 ( .A(B[63]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(A[63]), .B(n16), .Z(n15) );
  NANDN U17 ( .A(n16), .B(A[63]), .Z(n13) );
  XOR U18 ( .A(n16), .B(n17), .Z(DIFF[63]) );
  XOR U19 ( .A(B[63]), .B(A[63]), .Z(n17) );
  AND U20 ( .A(n18), .B(n19), .Z(n16) );
  NANDN U21 ( .A(B[62]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(A[62]), .B(n21), .Z(n20) );
  NANDN U23 ( .A(n21), .B(A[62]), .Z(n18) );
  XOR U24 ( .A(n21), .B(n22), .Z(DIFF[62]) );
  XOR U25 ( .A(B[62]), .B(A[62]), .Z(n22) );
  AND U26 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U27 ( .A(B[61]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(A[61]), .B(n26), .Z(n25) );
  NANDN U29 ( .A(n26), .B(A[61]), .Z(n23) );
  XOR U30 ( .A(n26), .B(n27), .Z(DIFF[61]) );
  XOR U31 ( .A(B[61]), .B(A[61]), .Z(n27) );
  AND U32 ( .A(n28), .B(n29), .Z(n26) );
  NANDN U33 ( .A(B[60]), .B(n30), .Z(n29) );
  NANDN U34 ( .A(A[60]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(n31), .B(A[60]), .Z(n28) );
  XOR U36 ( .A(n31), .B(n32), .Z(DIFF[60]) );
  XOR U37 ( .A(B[60]), .B(A[60]), .Z(n32) );
  AND U38 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U39 ( .A(B[59]), .B(n35), .Z(n34) );
  NANDN U40 ( .A(A[59]), .B(n36), .Z(n35) );
  NANDN U41 ( .A(n36), .B(A[59]), .Z(n33) );
  XOR U42 ( .A(n37), .B(n38), .Z(DIFF[5]) );
  XOR U43 ( .A(B[5]), .B(A[5]), .Z(n38) );
  XOR U44 ( .A(n36), .B(n39), .Z(DIFF[59]) );
  XOR U45 ( .A(B[59]), .B(A[59]), .Z(n39) );
  AND U46 ( .A(n40), .B(n41), .Z(n36) );
  NANDN U47 ( .A(B[58]), .B(n42), .Z(n41) );
  NANDN U48 ( .A(A[58]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(n43), .B(A[58]), .Z(n40) );
  XOR U50 ( .A(n43), .B(n44), .Z(DIFF[58]) );
  XOR U51 ( .A(B[58]), .B(A[58]), .Z(n44) );
  AND U52 ( .A(n45), .B(n46), .Z(n43) );
  NANDN U53 ( .A(B[57]), .B(n47), .Z(n46) );
  NANDN U54 ( .A(A[57]), .B(n48), .Z(n47) );
  NANDN U55 ( .A(n48), .B(A[57]), .Z(n45) );
  XOR U56 ( .A(n48), .B(n49), .Z(DIFF[57]) );
  XOR U57 ( .A(B[57]), .B(A[57]), .Z(n49) );
  AND U58 ( .A(n50), .B(n51), .Z(n48) );
  NANDN U59 ( .A(B[56]), .B(n52), .Z(n51) );
  NANDN U60 ( .A(A[56]), .B(n53), .Z(n52) );
  NANDN U61 ( .A(n53), .B(A[56]), .Z(n50) );
  XOR U62 ( .A(n53), .B(n54), .Z(DIFF[56]) );
  XOR U63 ( .A(B[56]), .B(A[56]), .Z(n54) );
  AND U64 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U65 ( .A(B[55]), .B(n57), .Z(n56) );
  NANDN U66 ( .A(A[55]), .B(n58), .Z(n57) );
  NANDN U67 ( .A(n58), .B(A[55]), .Z(n55) );
  XOR U68 ( .A(n58), .B(n59), .Z(DIFF[55]) );
  XOR U69 ( .A(B[55]), .B(A[55]), .Z(n59) );
  AND U70 ( .A(n60), .B(n61), .Z(n58) );
  NANDN U71 ( .A(B[54]), .B(n62), .Z(n61) );
  NANDN U72 ( .A(A[54]), .B(n63), .Z(n62) );
  NANDN U73 ( .A(n63), .B(A[54]), .Z(n60) );
  XOR U74 ( .A(n63), .B(n64), .Z(DIFF[54]) );
  XOR U75 ( .A(B[54]), .B(A[54]), .Z(n64) );
  AND U76 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U77 ( .A(B[53]), .B(n67), .Z(n66) );
  NANDN U78 ( .A(A[53]), .B(n68), .Z(n67) );
  NANDN U79 ( .A(n68), .B(A[53]), .Z(n65) );
  XOR U80 ( .A(n68), .B(n69), .Z(DIFF[53]) );
  XOR U81 ( .A(B[53]), .B(A[53]), .Z(n69) );
  AND U82 ( .A(n70), .B(n71), .Z(n68) );
  NANDN U83 ( .A(B[52]), .B(n72), .Z(n71) );
  NANDN U84 ( .A(A[52]), .B(n73), .Z(n72) );
  NANDN U85 ( .A(n73), .B(A[52]), .Z(n70) );
  XOR U86 ( .A(n73), .B(n74), .Z(DIFF[52]) );
  XOR U87 ( .A(B[52]), .B(A[52]), .Z(n74) );
  AND U88 ( .A(n75), .B(n76), .Z(n73) );
  NANDN U89 ( .A(B[51]), .B(n77), .Z(n76) );
  NANDN U90 ( .A(A[51]), .B(n78), .Z(n77) );
  NANDN U91 ( .A(n78), .B(A[51]), .Z(n75) );
  XOR U92 ( .A(n78), .B(n79), .Z(DIFF[51]) );
  XOR U93 ( .A(B[51]), .B(A[51]), .Z(n79) );
  AND U94 ( .A(n80), .B(n81), .Z(n78) );
  NANDN U95 ( .A(B[50]), .B(n82), .Z(n81) );
  NANDN U96 ( .A(A[50]), .B(n83), .Z(n82) );
  NANDN U97 ( .A(n83), .B(A[50]), .Z(n80) );
  XOR U98 ( .A(n83), .B(n84), .Z(DIFF[50]) );
  XOR U99 ( .A(B[50]), .B(A[50]), .Z(n84) );
  AND U100 ( .A(n85), .B(n86), .Z(n83) );
  NANDN U101 ( .A(B[49]), .B(n87), .Z(n86) );
  NANDN U102 ( .A(A[49]), .B(n88), .Z(n87) );
  NANDN U103 ( .A(n88), .B(A[49]), .Z(n85) );
  XOR U104 ( .A(n89), .B(n90), .Z(DIFF[4]) );
  XOR U105 ( .A(B[4]), .B(A[4]), .Z(n90) );
  XOR U106 ( .A(n88), .B(n91), .Z(DIFF[49]) );
  XOR U107 ( .A(B[49]), .B(A[49]), .Z(n91) );
  AND U108 ( .A(n92), .B(n93), .Z(n88) );
  NANDN U109 ( .A(B[48]), .B(n94), .Z(n93) );
  NANDN U110 ( .A(A[48]), .B(n95), .Z(n94) );
  NANDN U111 ( .A(n95), .B(A[48]), .Z(n92) );
  XOR U112 ( .A(n95), .B(n96), .Z(DIFF[48]) );
  XOR U113 ( .A(B[48]), .B(A[48]), .Z(n96) );
  AND U114 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U115 ( .A(B[47]), .B(n99), .Z(n98) );
  NANDN U116 ( .A(A[47]), .B(n100), .Z(n99) );
  NANDN U117 ( .A(n100), .B(A[47]), .Z(n97) );
  XOR U118 ( .A(n100), .B(n101), .Z(DIFF[47]) );
  XOR U119 ( .A(B[47]), .B(A[47]), .Z(n101) );
  AND U120 ( .A(n102), .B(n103), .Z(n100) );
  NANDN U121 ( .A(B[46]), .B(n104), .Z(n103) );
  NANDN U122 ( .A(A[46]), .B(n105), .Z(n104) );
  NANDN U123 ( .A(n105), .B(A[46]), .Z(n102) );
  XOR U124 ( .A(n105), .B(n106), .Z(DIFF[46]) );
  XOR U125 ( .A(B[46]), .B(A[46]), .Z(n106) );
  AND U126 ( .A(n107), .B(n108), .Z(n105) );
  NANDN U127 ( .A(B[45]), .B(n109), .Z(n108) );
  NANDN U128 ( .A(A[45]), .B(n110), .Z(n109) );
  NANDN U129 ( .A(n110), .B(A[45]), .Z(n107) );
  XOR U130 ( .A(n110), .B(n111), .Z(DIFF[45]) );
  XOR U131 ( .A(B[45]), .B(A[45]), .Z(n111) );
  AND U132 ( .A(n112), .B(n113), .Z(n110) );
  NANDN U133 ( .A(B[44]), .B(n114), .Z(n113) );
  NANDN U134 ( .A(A[44]), .B(n115), .Z(n114) );
  NANDN U135 ( .A(n115), .B(A[44]), .Z(n112) );
  XOR U136 ( .A(n115), .B(n116), .Z(DIFF[44]) );
  XOR U137 ( .A(B[44]), .B(A[44]), .Z(n116) );
  AND U138 ( .A(n117), .B(n118), .Z(n115) );
  NANDN U139 ( .A(B[43]), .B(n119), .Z(n118) );
  NANDN U140 ( .A(A[43]), .B(n120), .Z(n119) );
  NANDN U141 ( .A(n120), .B(A[43]), .Z(n117) );
  XOR U142 ( .A(n120), .B(n121), .Z(DIFF[43]) );
  XOR U143 ( .A(B[43]), .B(A[43]), .Z(n121) );
  AND U144 ( .A(n122), .B(n123), .Z(n120) );
  NANDN U145 ( .A(B[42]), .B(n124), .Z(n123) );
  NANDN U146 ( .A(A[42]), .B(n125), .Z(n124) );
  NANDN U147 ( .A(n125), .B(A[42]), .Z(n122) );
  XOR U148 ( .A(n125), .B(n126), .Z(DIFF[42]) );
  XOR U149 ( .A(B[42]), .B(A[42]), .Z(n126) );
  AND U150 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U151 ( .A(B[41]), .B(n129), .Z(n128) );
  NANDN U152 ( .A(A[41]), .B(n130), .Z(n129) );
  NANDN U153 ( .A(n130), .B(A[41]), .Z(n127) );
  XOR U154 ( .A(n130), .B(n131), .Z(DIFF[41]) );
  XOR U155 ( .A(B[41]), .B(A[41]), .Z(n131) );
  AND U156 ( .A(n132), .B(n133), .Z(n130) );
  NANDN U157 ( .A(B[40]), .B(n134), .Z(n133) );
  NANDN U158 ( .A(A[40]), .B(n135), .Z(n134) );
  NANDN U159 ( .A(n135), .B(A[40]), .Z(n132) );
  XOR U160 ( .A(n135), .B(n136), .Z(DIFF[40]) );
  XOR U161 ( .A(B[40]), .B(A[40]), .Z(n136) );
  AND U162 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U163 ( .A(B[39]), .B(n139), .Z(n138) );
  NANDN U164 ( .A(A[39]), .B(n140), .Z(n139) );
  NANDN U165 ( .A(n140), .B(A[39]), .Z(n137) );
  XOR U166 ( .A(n141), .B(n142), .Z(DIFF[3]) );
  XOR U167 ( .A(B[3]), .B(A[3]), .Z(n142) );
  XOR U168 ( .A(n140), .B(n143), .Z(DIFF[39]) );
  XOR U169 ( .A(B[39]), .B(A[39]), .Z(n143) );
  AND U170 ( .A(n144), .B(n145), .Z(n140) );
  NANDN U171 ( .A(B[38]), .B(n146), .Z(n145) );
  NANDN U172 ( .A(A[38]), .B(n147), .Z(n146) );
  NANDN U173 ( .A(n147), .B(A[38]), .Z(n144) );
  XOR U174 ( .A(n147), .B(n148), .Z(DIFF[38]) );
  XOR U175 ( .A(B[38]), .B(A[38]), .Z(n148) );
  AND U176 ( .A(n149), .B(n150), .Z(n147) );
  NANDN U177 ( .A(B[37]), .B(n151), .Z(n150) );
  NANDN U178 ( .A(A[37]), .B(n152), .Z(n151) );
  NANDN U179 ( .A(n152), .B(A[37]), .Z(n149) );
  XOR U180 ( .A(n152), .B(n153), .Z(DIFF[37]) );
  XOR U181 ( .A(B[37]), .B(A[37]), .Z(n153) );
  AND U182 ( .A(n154), .B(n155), .Z(n152) );
  NANDN U183 ( .A(B[36]), .B(n156), .Z(n155) );
  NANDN U184 ( .A(A[36]), .B(n157), .Z(n156) );
  NANDN U185 ( .A(n157), .B(A[36]), .Z(n154) );
  XOR U186 ( .A(n157), .B(n158), .Z(DIFF[36]) );
  XOR U187 ( .A(B[36]), .B(A[36]), .Z(n158) );
  AND U188 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U189 ( .A(B[35]), .B(n161), .Z(n160) );
  NANDN U190 ( .A(A[35]), .B(n162), .Z(n161) );
  NANDN U191 ( .A(n162), .B(A[35]), .Z(n159) );
  XOR U192 ( .A(n162), .B(n163), .Z(DIFF[35]) );
  XOR U193 ( .A(B[35]), .B(A[35]), .Z(n163) );
  AND U194 ( .A(n164), .B(n165), .Z(n162) );
  NANDN U195 ( .A(B[34]), .B(n166), .Z(n165) );
  NANDN U196 ( .A(A[34]), .B(n167), .Z(n166) );
  NANDN U197 ( .A(n167), .B(A[34]), .Z(n164) );
  XOR U198 ( .A(n167), .B(n168), .Z(DIFF[34]) );
  XOR U199 ( .A(B[34]), .B(A[34]), .Z(n168) );
  AND U200 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U201 ( .A(B[33]), .B(n171), .Z(n170) );
  NANDN U202 ( .A(A[33]), .B(n172), .Z(n171) );
  NANDN U203 ( .A(n172), .B(A[33]), .Z(n169) );
  XOR U204 ( .A(n172), .B(n173), .Z(DIFF[33]) );
  XOR U205 ( .A(B[33]), .B(A[33]), .Z(n173) );
  AND U206 ( .A(n174), .B(n175), .Z(n172) );
  NANDN U207 ( .A(B[32]), .B(n176), .Z(n175) );
  NANDN U208 ( .A(A[32]), .B(n177), .Z(n176) );
  NANDN U209 ( .A(n177), .B(A[32]), .Z(n174) );
  XOR U210 ( .A(n177), .B(n178), .Z(DIFF[32]) );
  XOR U211 ( .A(B[32]), .B(A[32]), .Z(n178) );
  AND U212 ( .A(n179), .B(n180), .Z(n177) );
  NANDN U213 ( .A(B[31]), .B(n181), .Z(n180) );
  NANDN U214 ( .A(A[31]), .B(n182), .Z(n181) );
  NANDN U215 ( .A(n182), .B(A[31]), .Z(n179) );
  XOR U216 ( .A(n182), .B(n183), .Z(DIFF[31]) );
  XOR U217 ( .A(B[31]), .B(A[31]), .Z(n183) );
  AND U218 ( .A(n184), .B(n185), .Z(n182) );
  NANDN U219 ( .A(B[30]), .B(n186), .Z(n185) );
  NANDN U220 ( .A(A[30]), .B(n187), .Z(n186) );
  NANDN U221 ( .A(n187), .B(A[30]), .Z(n184) );
  XOR U222 ( .A(n187), .B(n188), .Z(DIFF[30]) );
  XOR U223 ( .A(B[30]), .B(A[30]), .Z(n188) );
  AND U224 ( .A(n189), .B(n190), .Z(n187) );
  NANDN U225 ( .A(B[29]), .B(n191), .Z(n190) );
  NANDN U226 ( .A(A[29]), .B(n192), .Z(n191) );
  NANDN U227 ( .A(n192), .B(A[29]), .Z(n189) );
  XOR U228 ( .A(n193), .B(n194), .Z(DIFF[2]) );
  XOR U229 ( .A(B[2]), .B(A[2]), .Z(n194) );
  XOR U230 ( .A(n192), .B(n195), .Z(DIFF[29]) );
  XOR U231 ( .A(B[29]), .B(A[29]), .Z(n195) );
  AND U232 ( .A(n196), .B(n197), .Z(n192) );
  NANDN U233 ( .A(B[28]), .B(n198), .Z(n197) );
  NANDN U234 ( .A(A[28]), .B(n199), .Z(n198) );
  NANDN U235 ( .A(n199), .B(A[28]), .Z(n196) );
  XOR U236 ( .A(n199), .B(n200), .Z(DIFF[28]) );
  XOR U237 ( .A(B[28]), .B(A[28]), .Z(n200) );
  AND U238 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U239 ( .A(B[27]), .B(n203), .Z(n202) );
  NANDN U240 ( .A(A[27]), .B(n204), .Z(n203) );
  NANDN U241 ( .A(n204), .B(A[27]), .Z(n201) );
  XOR U242 ( .A(n204), .B(n205), .Z(DIFF[27]) );
  XOR U243 ( .A(B[27]), .B(A[27]), .Z(n205) );
  AND U244 ( .A(n206), .B(n207), .Z(n204) );
  NANDN U245 ( .A(B[26]), .B(n208), .Z(n207) );
  NANDN U246 ( .A(A[26]), .B(n209), .Z(n208) );
  NANDN U247 ( .A(n209), .B(A[26]), .Z(n206) );
  XOR U248 ( .A(n209), .B(n210), .Z(DIFF[26]) );
  XOR U249 ( .A(B[26]), .B(A[26]), .Z(n210) );
  AND U250 ( .A(n211), .B(n212), .Z(n209) );
  NANDN U251 ( .A(B[25]), .B(n213), .Z(n212) );
  NANDN U252 ( .A(A[25]), .B(n214), .Z(n213) );
  NANDN U253 ( .A(n214), .B(A[25]), .Z(n211) );
  XOR U254 ( .A(n214), .B(n215), .Z(DIFF[25]) );
  XOR U255 ( .A(B[25]), .B(A[25]), .Z(n215) );
  AND U256 ( .A(n216), .B(n217), .Z(n214) );
  NANDN U257 ( .A(B[24]), .B(n218), .Z(n217) );
  NANDN U258 ( .A(A[24]), .B(n219), .Z(n218) );
  NANDN U259 ( .A(n219), .B(A[24]), .Z(n216) );
  XOR U260 ( .A(n219), .B(n220), .Z(DIFF[24]) );
  XOR U261 ( .A(B[24]), .B(A[24]), .Z(n220) );
  AND U262 ( .A(n221), .B(n222), .Z(n219) );
  NANDN U263 ( .A(B[23]), .B(n223), .Z(n222) );
  NANDN U264 ( .A(A[23]), .B(n224), .Z(n223) );
  NANDN U265 ( .A(n224), .B(A[23]), .Z(n221) );
  XOR U266 ( .A(n224), .B(n225), .Z(DIFF[23]) );
  XOR U267 ( .A(B[23]), .B(A[23]), .Z(n225) );
  AND U268 ( .A(n226), .B(n227), .Z(n224) );
  NANDN U269 ( .A(B[22]), .B(n228), .Z(n227) );
  NANDN U270 ( .A(A[22]), .B(n229), .Z(n228) );
  NANDN U271 ( .A(n229), .B(A[22]), .Z(n226) );
  XOR U272 ( .A(n229), .B(n230), .Z(DIFF[22]) );
  XOR U273 ( .A(B[22]), .B(A[22]), .Z(n230) );
  AND U274 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U275 ( .A(B[21]), .B(n233), .Z(n232) );
  NANDN U276 ( .A(A[21]), .B(n234), .Z(n233) );
  NANDN U277 ( .A(n234), .B(A[21]), .Z(n231) );
  XOR U278 ( .A(n234), .B(n235), .Z(DIFF[21]) );
  XOR U279 ( .A(B[21]), .B(A[21]), .Z(n235) );
  AND U280 ( .A(n236), .B(n237), .Z(n234) );
  NANDN U281 ( .A(B[20]), .B(n238), .Z(n237) );
  NANDN U282 ( .A(A[20]), .B(n239), .Z(n238) );
  NANDN U283 ( .A(n239), .B(A[20]), .Z(n236) );
  XOR U284 ( .A(n239), .B(n240), .Z(DIFF[20]) );
  XOR U285 ( .A(B[20]), .B(A[20]), .Z(n240) );
  AND U286 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U287 ( .A(B[19]), .B(n243), .Z(n242) );
  NANDN U288 ( .A(A[19]), .B(n244), .Z(n243) );
  NANDN U289 ( .A(n244), .B(A[19]), .Z(n241) );
  XOR U290 ( .A(n2), .B(n245), .Z(DIFF[1]) );
  XOR U291 ( .A(B[1]), .B(A[1]), .Z(n245) );
  XOR U292 ( .A(n244), .B(n246), .Z(DIFF[19]) );
  XOR U293 ( .A(B[19]), .B(A[19]), .Z(n246) );
  AND U294 ( .A(n247), .B(n248), .Z(n244) );
  NANDN U295 ( .A(B[18]), .B(n249), .Z(n248) );
  NANDN U296 ( .A(A[18]), .B(n250), .Z(n249) );
  NANDN U297 ( .A(n250), .B(A[18]), .Z(n247) );
  XOR U298 ( .A(n250), .B(n251), .Z(DIFF[18]) );
  XOR U299 ( .A(B[18]), .B(A[18]), .Z(n251) );
  AND U300 ( .A(n252), .B(n253), .Z(n250) );
  NANDN U301 ( .A(B[17]), .B(n254), .Z(n253) );
  NANDN U302 ( .A(A[17]), .B(n255), .Z(n254) );
  NANDN U303 ( .A(n255), .B(A[17]), .Z(n252) );
  XOR U304 ( .A(n255), .B(n256), .Z(DIFF[17]) );
  XOR U305 ( .A(B[17]), .B(A[17]), .Z(n256) );
  AND U306 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U307 ( .A(B[16]), .B(n259), .Z(n258) );
  NANDN U308 ( .A(A[16]), .B(n260), .Z(n259) );
  NANDN U309 ( .A(n260), .B(A[16]), .Z(n257) );
  XOR U310 ( .A(n260), .B(n261), .Z(DIFF[16]) );
  XOR U311 ( .A(B[16]), .B(A[16]), .Z(n261) );
  AND U312 ( .A(n262), .B(n263), .Z(n260) );
  NANDN U313 ( .A(B[15]), .B(n264), .Z(n263) );
  NANDN U314 ( .A(A[15]), .B(n265), .Z(n264) );
  NANDN U315 ( .A(n265), .B(A[15]), .Z(n262) );
  XOR U316 ( .A(n265), .B(n266), .Z(DIFF[15]) );
  XOR U317 ( .A(B[15]), .B(A[15]), .Z(n266) );
  AND U318 ( .A(n267), .B(n268), .Z(n265) );
  NANDN U319 ( .A(B[14]), .B(n269), .Z(n268) );
  NANDN U320 ( .A(A[14]), .B(n270), .Z(n269) );
  NANDN U321 ( .A(n270), .B(A[14]), .Z(n267) );
  XOR U322 ( .A(n270), .B(n271), .Z(DIFF[14]) );
  XOR U323 ( .A(B[14]), .B(A[14]), .Z(n271) );
  AND U324 ( .A(n272), .B(n273), .Z(n270) );
  NANDN U325 ( .A(B[13]), .B(n274), .Z(n273) );
  NANDN U326 ( .A(A[13]), .B(n275), .Z(n274) );
  NANDN U327 ( .A(n275), .B(A[13]), .Z(n272) );
  XOR U328 ( .A(n275), .B(n276), .Z(DIFF[13]) );
  XOR U329 ( .A(B[13]), .B(A[13]), .Z(n276) );
  AND U330 ( .A(n277), .B(n278), .Z(n275) );
  NANDN U331 ( .A(B[12]), .B(n279), .Z(n278) );
  NANDN U332 ( .A(A[12]), .B(n280), .Z(n279) );
  NANDN U333 ( .A(n280), .B(A[12]), .Z(n277) );
  XOR U334 ( .A(n280), .B(n281), .Z(DIFF[12]) );
  XOR U335 ( .A(B[12]), .B(A[12]), .Z(n281) );
  AND U336 ( .A(n282), .B(n283), .Z(n280) );
  NANDN U337 ( .A(B[11]), .B(n284), .Z(n283) );
  NANDN U338 ( .A(A[11]), .B(n285), .Z(n284) );
  NANDN U339 ( .A(n285), .B(A[11]), .Z(n282) );
  XOR U340 ( .A(n285), .B(n286), .Z(DIFF[11]) );
  XOR U341 ( .A(B[11]), .B(A[11]), .Z(n286) );
  AND U342 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U343 ( .A(B[10]), .B(n289), .Z(n288) );
  NANDN U344 ( .A(A[10]), .B(n290), .Z(n289) );
  NANDN U345 ( .A(n290), .B(A[10]), .Z(n287) );
  XOR U346 ( .A(n290), .B(n291), .Z(DIFF[10]) );
  XOR U347 ( .A(B[10]), .B(A[10]), .Z(n291) );
  AND U348 ( .A(n292), .B(n293), .Z(n290) );
  NANDN U349 ( .A(B[9]), .B(n294), .Z(n293) );
  OR U350 ( .A(n3), .B(A[9]), .Z(n294) );
  NAND U351 ( .A(A[9]), .B(n3), .Z(n292) );
  NAND U352 ( .A(n295), .B(n296), .Z(n3) );
  NANDN U353 ( .A(B[8]), .B(n297), .Z(n296) );
  NANDN U354 ( .A(A[8]), .B(n5), .Z(n297) );
  NANDN U355 ( .A(n5), .B(A[8]), .Z(n295) );
  AND U356 ( .A(n298), .B(n299), .Z(n5) );
  NANDN U357 ( .A(B[7]), .B(n300), .Z(n299) );
  NANDN U358 ( .A(A[7]), .B(n7), .Z(n300) );
  NANDN U359 ( .A(n7), .B(A[7]), .Z(n298) );
  AND U360 ( .A(n301), .B(n302), .Z(n7) );
  NANDN U361 ( .A(B[6]), .B(n303), .Z(n302) );
  NANDN U362 ( .A(A[6]), .B(n9), .Z(n303) );
  NANDN U363 ( .A(n9), .B(A[6]), .Z(n301) );
  AND U364 ( .A(n304), .B(n305), .Z(n9) );
  NANDN U365 ( .A(B[5]), .B(n306), .Z(n305) );
  NANDN U366 ( .A(A[5]), .B(n37), .Z(n306) );
  NANDN U367 ( .A(n37), .B(A[5]), .Z(n304) );
  AND U368 ( .A(n307), .B(n308), .Z(n37) );
  NANDN U369 ( .A(B[4]), .B(n309), .Z(n308) );
  NANDN U370 ( .A(A[4]), .B(n89), .Z(n309) );
  NANDN U371 ( .A(n89), .B(A[4]), .Z(n307) );
  AND U372 ( .A(n310), .B(n311), .Z(n89) );
  NANDN U373 ( .A(B[3]), .B(n312), .Z(n311) );
  NANDN U374 ( .A(A[3]), .B(n141), .Z(n312) );
  NANDN U375 ( .A(n141), .B(A[3]), .Z(n310) );
  AND U376 ( .A(n313), .B(n314), .Z(n141) );
  NANDN U377 ( .A(B[2]), .B(n315), .Z(n314) );
  NANDN U378 ( .A(A[2]), .B(n193), .Z(n315) );
  NANDN U379 ( .A(n193), .B(A[2]), .Z(n313) );
  AND U380 ( .A(n316), .B(n317), .Z(n193) );
  NANDN U381 ( .A(B[1]), .B(n318), .Z(n317) );
  NAND U382 ( .A(n2), .B(n1), .Z(n318) );
  NAND U383 ( .A(A[1]), .B(n319), .Z(n316) );
  NAND U384 ( .A(n319), .B(n320), .Z(DIFF[0]) );
  NANDN U385 ( .A(B[0]), .B(A[0]), .Z(n320) );
  NANDN U386 ( .A(A[0]), .B(B[0]), .Z(n319) );
endmodule


module modmult_step_N64_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [65:0] A;
  input [65:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[65]), .B(B[64]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[63]), .B(A[63]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[62]), .B(B[62]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[62]), .B(A[62]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[61]), .B(B[61]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[60]), .B(B[60]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[60]), .B(A[60]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[59]), .B(B[59]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[58]), .B(B[58]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[58]), .B(A[58]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[57]), .B(B[57]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[56]), .B(B[56]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[56]), .B(A[56]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[55]), .B(B[55]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[54]), .B(B[54]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[54]), .B(A[54]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[53]), .B(B[53]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[52]), .B(B[52]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[52]), .B(A[52]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[51]), .B(B[51]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[50]), .B(B[50]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[50]), .B(A[50]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[49]), .B(B[49]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[48]), .B(B[48]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[48]), .B(A[48]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[47]), .B(B[47]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[46]), .B(B[46]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[46]), .B(A[46]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[45]), .B(B[45]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[44]), .B(B[44]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[44]), .B(A[44]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[43]), .B(B[43]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[42]), .B(B[42]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[42]), .B(A[42]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[41]), .B(B[41]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[40]), .B(B[40]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[40]), .B(A[40]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[39]), .B(B[39]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[38]), .B(B[38]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[38]), .B(A[38]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[37]), .B(B[37]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[36]), .B(B[36]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[36]), .B(A[36]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[35]), .B(B[35]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[34]), .B(B[34]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[34]), .B(A[34]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[33]), .B(B[33]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[32]), .B(B[32]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[32]), .B(A[32]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[31]), .B(B[31]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[30]), .B(B[30]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[30]), .B(A[30]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[29]), .B(B[29]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[28]), .B(B[28]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[28]), .B(A[28]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[27]), .B(B[27]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[26]), .B(B[26]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[26]), .B(A[26]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[25]), .B(B[25]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[24]), .B(B[24]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[24]), .B(A[24]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[23]), .B(B[23]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[22]), .B(B[22]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[22]), .B(A[22]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[21]), .B(B[21]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[20]), .B(B[20]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[20]), .B(A[20]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[19]), .B(B[19]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[18]), .B(B[18]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[18]), .B(A[18]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[17]), .B(B[17]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[16]), .B(B[16]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[16]), .B(A[16]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[15]), .B(B[15]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[14]), .B(B[14]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[14]), .B(A[14]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[13]), .B(B[13]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[12]), .B(B[12]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[12]), .B(A[12]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[11]), .B(B[11]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[10]), .B(B[10]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[9]), .B(A[9]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[9]), .B(B[9]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[8]), .B(B[8]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[8]), .B(A[8]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[7]), .B(B[7]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[6]), .B(B[6]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[6]), .B(A[6]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[5]), .B(B[5]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[4]), .B(B[4]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[4]), .B(A[4]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[3]), .B(B[3]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[2]), .B(B[2]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[2]), .B(A[2]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NANDN U221 ( .A(B[1]), .B(n253), .Z(n252) );
  NANDN U222 ( .A(A[1]), .B(n254), .Z(n253) );
  NANDN U223 ( .A(n254), .B(A[1]), .Z(n251) );
  ANDN U224 ( .B(B[0]), .A(A[0]), .Z(n254) );
  NANDN U225 ( .A(B[3]), .B(A[3]), .Z(n243) );
  NANDN U226 ( .A(B[5]), .B(A[5]), .Z(n235) );
  NANDN U227 ( .A(B[7]), .B(A[7]), .Z(n227) );
  NANDN U228 ( .A(B[10]), .B(A[10]), .Z(n219) );
  NANDN U229 ( .A(B[11]), .B(A[11]), .Z(n211) );
  NANDN U230 ( .A(B[13]), .B(A[13]), .Z(n203) );
  NANDN U231 ( .A(B[15]), .B(A[15]), .Z(n195) );
  NANDN U232 ( .A(B[17]), .B(A[17]), .Z(n187) );
  NANDN U233 ( .A(B[19]), .B(A[19]), .Z(n179) );
  NANDN U234 ( .A(B[21]), .B(A[21]), .Z(n171) );
  NANDN U235 ( .A(B[23]), .B(A[23]), .Z(n163) );
  NANDN U236 ( .A(B[25]), .B(A[25]), .Z(n155) );
  NANDN U237 ( .A(B[27]), .B(A[27]), .Z(n147) );
  NANDN U238 ( .A(B[29]), .B(A[29]), .Z(n139) );
  NANDN U239 ( .A(B[31]), .B(A[31]), .Z(n131) );
  NANDN U240 ( .A(B[33]), .B(A[33]), .Z(n123) );
  NANDN U241 ( .A(B[35]), .B(A[35]), .Z(n115) );
  NANDN U242 ( .A(B[37]), .B(A[37]), .Z(n107) );
  NANDN U243 ( .A(B[39]), .B(A[39]), .Z(n99) );
  NANDN U244 ( .A(B[41]), .B(A[41]), .Z(n91) );
  NANDN U245 ( .A(B[43]), .B(A[43]), .Z(n83) );
  NANDN U246 ( .A(B[45]), .B(A[45]), .Z(n75) );
  NANDN U247 ( .A(B[47]), .B(A[47]), .Z(n67) );
  NANDN U248 ( .A(B[49]), .B(A[49]), .Z(n59) );
  NANDN U249 ( .A(B[51]), .B(A[51]), .Z(n51) );
  NANDN U250 ( .A(B[53]), .B(A[53]), .Z(n43) );
  NANDN U251 ( .A(B[55]), .B(A[55]), .Z(n35) );
  NANDN U252 ( .A(B[57]), .B(A[57]), .Z(n27) );
  NANDN U253 ( .A(B[59]), .B(A[59]), .Z(n19) );
  NANDN U254 ( .A(B[61]), .B(A[61]), .Z(n11) );
  NANDN U255 ( .A(A[63]), .B(B[63]), .Z(n3) );
endmodule


module modmult_step_N64_DW01_add_0 ( A, B, CI, SUM, CO );
  input [65:0] A;
  input [65:0] B;
  output [65:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(A[65]), .B(n9), .Z(SUM[65]) );
  AND U10 ( .A(A[64]), .B(n10), .Z(n9) );
  XOR U11 ( .A(A[64]), .B(n10), .Z(SUM[64]) );
  NAND U12 ( .A(n11), .B(n12), .Z(n10) );
  NAND U13 ( .A(B[63]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(A[63]), .B(n14), .Z(n13) );
  NANDN U15 ( .A(n14), .B(A[63]), .Z(n11) );
  XOR U16 ( .A(n14), .B(n15), .Z(SUM[63]) );
  XNOR U17 ( .A(B[63]), .B(A[63]), .Z(n15) );
  AND U18 ( .A(n16), .B(n17), .Z(n14) );
  NAND U19 ( .A(B[62]), .B(n18), .Z(n17) );
  NANDN U20 ( .A(A[62]), .B(n19), .Z(n18) );
  NANDN U21 ( .A(n19), .B(A[62]), .Z(n16) );
  XOR U22 ( .A(n19), .B(n20), .Z(SUM[62]) );
  XNOR U23 ( .A(B[62]), .B(A[62]), .Z(n20) );
  AND U24 ( .A(n21), .B(n22), .Z(n19) );
  NAND U25 ( .A(B[61]), .B(n23), .Z(n22) );
  NANDN U26 ( .A(A[61]), .B(n24), .Z(n23) );
  NANDN U27 ( .A(n24), .B(A[61]), .Z(n21) );
  XOR U28 ( .A(n24), .B(n25), .Z(SUM[61]) );
  XNOR U29 ( .A(B[61]), .B(A[61]), .Z(n25) );
  AND U30 ( .A(n26), .B(n27), .Z(n24) );
  NAND U31 ( .A(B[60]), .B(n28), .Z(n27) );
  NANDN U32 ( .A(A[60]), .B(n29), .Z(n28) );
  NANDN U33 ( .A(n29), .B(A[60]), .Z(n26) );
  XOR U34 ( .A(n29), .B(n30), .Z(SUM[60]) );
  XNOR U35 ( .A(B[60]), .B(A[60]), .Z(n30) );
  AND U36 ( .A(n31), .B(n32), .Z(n29) );
  NAND U37 ( .A(B[59]), .B(n33), .Z(n32) );
  NANDN U38 ( .A(A[59]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(n34), .B(A[59]), .Z(n31) );
  XOR U40 ( .A(n35), .B(n36), .Z(SUM[5]) );
  XNOR U41 ( .A(B[5]), .B(A[5]), .Z(n36) );
  XOR U42 ( .A(n34), .B(n37), .Z(SUM[59]) );
  XNOR U43 ( .A(B[59]), .B(A[59]), .Z(n37) );
  AND U44 ( .A(n38), .B(n39), .Z(n34) );
  NAND U45 ( .A(B[58]), .B(n40), .Z(n39) );
  NANDN U46 ( .A(A[58]), .B(n41), .Z(n40) );
  NANDN U47 ( .A(n41), .B(A[58]), .Z(n38) );
  XOR U48 ( .A(n41), .B(n42), .Z(SUM[58]) );
  XNOR U49 ( .A(B[58]), .B(A[58]), .Z(n42) );
  AND U50 ( .A(n43), .B(n44), .Z(n41) );
  NAND U51 ( .A(B[57]), .B(n45), .Z(n44) );
  NANDN U52 ( .A(A[57]), .B(n46), .Z(n45) );
  NANDN U53 ( .A(n46), .B(A[57]), .Z(n43) );
  XOR U54 ( .A(n46), .B(n47), .Z(SUM[57]) );
  XNOR U55 ( .A(B[57]), .B(A[57]), .Z(n47) );
  AND U56 ( .A(n48), .B(n49), .Z(n46) );
  NAND U57 ( .A(B[56]), .B(n50), .Z(n49) );
  NANDN U58 ( .A(A[56]), .B(n51), .Z(n50) );
  NANDN U59 ( .A(n51), .B(A[56]), .Z(n48) );
  XOR U60 ( .A(n51), .B(n52), .Z(SUM[56]) );
  XNOR U61 ( .A(B[56]), .B(A[56]), .Z(n52) );
  AND U62 ( .A(n53), .B(n54), .Z(n51) );
  NAND U63 ( .A(B[55]), .B(n55), .Z(n54) );
  NANDN U64 ( .A(A[55]), .B(n56), .Z(n55) );
  NANDN U65 ( .A(n56), .B(A[55]), .Z(n53) );
  XOR U66 ( .A(n56), .B(n57), .Z(SUM[55]) );
  XNOR U67 ( .A(B[55]), .B(A[55]), .Z(n57) );
  AND U68 ( .A(n58), .B(n59), .Z(n56) );
  NAND U69 ( .A(B[54]), .B(n60), .Z(n59) );
  NANDN U70 ( .A(A[54]), .B(n61), .Z(n60) );
  NANDN U71 ( .A(n61), .B(A[54]), .Z(n58) );
  XOR U72 ( .A(n61), .B(n62), .Z(SUM[54]) );
  XNOR U73 ( .A(B[54]), .B(A[54]), .Z(n62) );
  AND U74 ( .A(n63), .B(n64), .Z(n61) );
  NAND U75 ( .A(B[53]), .B(n65), .Z(n64) );
  NANDN U76 ( .A(A[53]), .B(n66), .Z(n65) );
  NANDN U77 ( .A(n66), .B(A[53]), .Z(n63) );
  XOR U78 ( .A(n66), .B(n67), .Z(SUM[53]) );
  XNOR U79 ( .A(B[53]), .B(A[53]), .Z(n67) );
  AND U80 ( .A(n68), .B(n69), .Z(n66) );
  NAND U81 ( .A(B[52]), .B(n70), .Z(n69) );
  NANDN U82 ( .A(A[52]), .B(n71), .Z(n70) );
  NANDN U83 ( .A(n71), .B(A[52]), .Z(n68) );
  XOR U84 ( .A(n71), .B(n72), .Z(SUM[52]) );
  XNOR U85 ( .A(B[52]), .B(A[52]), .Z(n72) );
  AND U86 ( .A(n73), .B(n74), .Z(n71) );
  NAND U87 ( .A(B[51]), .B(n75), .Z(n74) );
  NANDN U88 ( .A(A[51]), .B(n76), .Z(n75) );
  NANDN U89 ( .A(n76), .B(A[51]), .Z(n73) );
  XOR U90 ( .A(n76), .B(n77), .Z(SUM[51]) );
  XNOR U91 ( .A(B[51]), .B(A[51]), .Z(n77) );
  AND U92 ( .A(n78), .B(n79), .Z(n76) );
  NAND U93 ( .A(B[50]), .B(n80), .Z(n79) );
  NANDN U94 ( .A(A[50]), .B(n81), .Z(n80) );
  NANDN U95 ( .A(n81), .B(A[50]), .Z(n78) );
  XOR U96 ( .A(n81), .B(n82), .Z(SUM[50]) );
  XNOR U97 ( .A(B[50]), .B(A[50]), .Z(n82) );
  AND U98 ( .A(n83), .B(n84), .Z(n81) );
  NAND U99 ( .A(B[49]), .B(n85), .Z(n84) );
  NANDN U100 ( .A(A[49]), .B(n86), .Z(n85) );
  NANDN U101 ( .A(n86), .B(A[49]), .Z(n83) );
  XOR U102 ( .A(n87), .B(n88), .Z(SUM[4]) );
  XNOR U103 ( .A(B[4]), .B(A[4]), .Z(n88) );
  XOR U104 ( .A(n86), .B(n89), .Z(SUM[49]) );
  XNOR U105 ( .A(B[49]), .B(A[49]), .Z(n89) );
  AND U106 ( .A(n90), .B(n91), .Z(n86) );
  NAND U107 ( .A(B[48]), .B(n92), .Z(n91) );
  NANDN U108 ( .A(A[48]), .B(n93), .Z(n92) );
  NANDN U109 ( .A(n93), .B(A[48]), .Z(n90) );
  XOR U110 ( .A(n93), .B(n94), .Z(SUM[48]) );
  XNOR U111 ( .A(B[48]), .B(A[48]), .Z(n94) );
  AND U112 ( .A(n95), .B(n96), .Z(n93) );
  NAND U113 ( .A(B[47]), .B(n97), .Z(n96) );
  NANDN U114 ( .A(A[47]), .B(n98), .Z(n97) );
  NANDN U115 ( .A(n98), .B(A[47]), .Z(n95) );
  XOR U116 ( .A(n98), .B(n99), .Z(SUM[47]) );
  XNOR U117 ( .A(B[47]), .B(A[47]), .Z(n99) );
  AND U118 ( .A(n100), .B(n101), .Z(n98) );
  NAND U119 ( .A(B[46]), .B(n102), .Z(n101) );
  NANDN U120 ( .A(A[46]), .B(n103), .Z(n102) );
  NANDN U121 ( .A(n103), .B(A[46]), .Z(n100) );
  XOR U122 ( .A(n103), .B(n104), .Z(SUM[46]) );
  XNOR U123 ( .A(B[46]), .B(A[46]), .Z(n104) );
  AND U124 ( .A(n105), .B(n106), .Z(n103) );
  NAND U125 ( .A(B[45]), .B(n107), .Z(n106) );
  NANDN U126 ( .A(A[45]), .B(n108), .Z(n107) );
  NANDN U127 ( .A(n108), .B(A[45]), .Z(n105) );
  XOR U128 ( .A(n108), .B(n109), .Z(SUM[45]) );
  XNOR U129 ( .A(B[45]), .B(A[45]), .Z(n109) );
  AND U130 ( .A(n110), .B(n111), .Z(n108) );
  NAND U131 ( .A(B[44]), .B(n112), .Z(n111) );
  NANDN U132 ( .A(A[44]), .B(n113), .Z(n112) );
  NANDN U133 ( .A(n113), .B(A[44]), .Z(n110) );
  XOR U134 ( .A(n113), .B(n114), .Z(SUM[44]) );
  XNOR U135 ( .A(B[44]), .B(A[44]), .Z(n114) );
  AND U136 ( .A(n115), .B(n116), .Z(n113) );
  NAND U137 ( .A(B[43]), .B(n117), .Z(n116) );
  NANDN U138 ( .A(A[43]), .B(n118), .Z(n117) );
  NANDN U139 ( .A(n118), .B(A[43]), .Z(n115) );
  XOR U140 ( .A(n118), .B(n119), .Z(SUM[43]) );
  XNOR U141 ( .A(B[43]), .B(A[43]), .Z(n119) );
  AND U142 ( .A(n120), .B(n121), .Z(n118) );
  NAND U143 ( .A(B[42]), .B(n122), .Z(n121) );
  NANDN U144 ( .A(A[42]), .B(n123), .Z(n122) );
  NANDN U145 ( .A(n123), .B(A[42]), .Z(n120) );
  XOR U146 ( .A(n123), .B(n124), .Z(SUM[42]) );
  XNOR U147 ( .A(B[42]), .B(A[42]), .Z(n124) );
  AND U148 ( .A(n125), .B(n126), .Z(n123) );
  NAND U149 ( .A(B[41]), .B(n127), .Z(n126) );
  NANDN U150 ( .A(A[41]), .B(n128), .Z(n127) );
  NANDN U151 ( .A(n128), .B(A[41]), .Z(n125) );
  XOR U152 ( .A(n128), .B(n129), .Z(SUM[41]) );
  XNOR U153 ( .A(B[41]), .B(A[41]), .Z(n129) );
  AND U154 ( .A(n130), .B(n131), .Z(n128) );
  NAND U155 ( .A(B[40]), .B(n132), .Z(n131) );
  NANDN U156 ( .A(A[40]), .B(n133), .Z(n132) );
  NANDN U157 ( .A(n133), .B(A[40]), .Z(n130) );
  XOR U158 ( .A(n133), .B(n134), .Z(SUM[40]) );
  XNOR U159 ( .A(B[40]), .B(A[40]), .Z(n134) );
  AND U160 ( .A(n135), .B(n136), .Z(n133) );
  NAND U161 ( .A(B[39]), .B(n137), .Z(n136) );
  NANDN U162 ( .A(A[39]), .B(n138), .Z(n137) );
  NANDN U163 ( .A(n138), .B(A[39]), .Z(n135) );
  XOR U164 ( .A(n139), .B(n140), .Z(SUM[3]) );
  XNOR U165 ( .A(B[3]), .B(A[3]), .Z(n140) );
  XOR U166 ( .A(n138), .B(n141), .Z(SUM[39]) );
  XNOR U167 ( .A(B[39]), .B(A[39]), .Z(n141) );
  AND U168 ( .A(n142), .B(n143), .Z(n138) );
  NAND U169 ( .A(B[38]), .B(n144), .Z(n143) );
  NANDN U170 ( .A(A[38]), .B(n145), .Z(n144) );
  NANDN U171 ( .A(n145), .B(A[38]), .Z(n142) );
  XOR U172 ( .A(n145), .B(n146), .Z(SUM[38]) );
  XNOR U173 ( .A(B[38]), .B(A[38]), .Z(n146) );
  AND U174 ( .A(n147), .B(n148), .Z(n145) );
  NAND U175 ( .A(B[37]), .B(n149), .Z(n148) );
  NANDN U176 ( .A(A[37]), .B(n150), .Z(n149) );
  NANDN U177 ( .A(n150), .B(A[37]), .Z(n147) );
  XOR U178 ( .A(n150), .B(n151), .Z(SUM[37]) );
  XNOR U179 ( .A(B[37]), .B(A[37]), .Z(n151) );
  AND U180 ( .A(n152), .B(n153), .Z(n150) );
  NAND U181 ( .A(B[36]), .B(n154), .Z(n153) );
  NANDN U182 ( .A(A[36]), .B(n155), .Z(n154) );
  NANDN U183 ( .A(n155), .B(A[36]), .Z(n152) );
  XOR U184 ( .A(n155), .B(n156), .Z(SUM[36]) );
  XNOR U185 ( .A(B[36]), .B(A[36]), .Z(n156) );
  AND U186 ( .A(n157), .B(n158), .Z(n155) );
  NAND U187 ( .A(B[35]), .B(n159), .Z(n158) );
  NANDN U188 ( .A(A[35]), .B(n160), .Z(n159) );
  NANDN U189 ( .A(n160), .B(A[35]), .Z(n157) );
  XOR U190 ( .A(n160), .B(n161), .Z(SUM[35]) );
  XNOR U191 ( .A(B[35]), .B(A[35]), .Z(n161) );
  AND U192 ( .A(n162), .B(n163), .Z(n160) );
  NAND U193 ( .A(B[34]), .B(n164), .Z(n163) );
  NANDN U194 ( .A(A[34]), .B(n165), .Z(n164) );
  NANDN U195 ( .A(n165), .B(A[34]), .Z(n162) );
  XOR U196 ( .A(n165), .B(n166), .Z(SUM[34]) );
  XNOR U197 ( .A(B[34]), .B(A[34]), .Z(n166) );
  AND U198 ( .A(n167), .B(n168), .Z(n165) );
  NAND U199 ( .A(B[33]), .B(n169), .Z(n168) );
  NANDN U200 ( .A(A[33]), .B(n170), .Z(n169) );
  NANDN U201 ( .A(n170), .B(A[33]), .Z(n167) );
  XOR U202 ( .A(n170), .B(n171), .Z(SUM[33]) );
  XNOR U203 ( .A(B[33]), .B(A[33]), .Z(n171) );
  AND U204 ( .A(n172), .B(n173), .Z(n170) );
  NAND U205 ( .A(B[32]), .B(n174), .Z(n173) );
  NANDN U206 ( .A(A[32]), .B(n175), .Z(n174) );
  NANDN U207 ( .A(n175), .B(A[32]), .Z(n172) );
  XOR U208 ( .A(n175), .B(n176), .Z(SUM[32]) );
  XNOR U209 ( .A(B[32]), .B(A[32]), .Z(n176) );
  AND U210 ( .A(n177), .B(n178), .Z(n175) );
  NAND U211 ( .A(B[31]), .B(n179), .Z(n178) );
  NANDN U212 ( .A(A[31]), .B(n180), .Z(n179) );
  NANDN U213 ( .A(n180), .B(A[31]), .Z(n177) );
  XOR U214 ( .A(n180), .B(n181), .Z(SUM[31]) );
  XNOR U215 ( .A(B[31]), .B(A[31]), .Z(n181) );
  AND U216 ( .A(n182), .B(n183), .Z(n180) );
  NAND U217 ( .A(B[30]), .B(n184), .Z(n183) );
  NANDN U218 ( .A(A[30]), .B(n185), .Z(n184) );
  NANDN U219 ( .A(n185), .B(A[30]), .Z(n182) );
  XOR U220 ( .A(n185), .B(n186), .Z(SUM[30]) );
  XNOR U221 ( .A(B[30]), .B(A[30]), .Z(n186) );
  AND U222 ( .A(n187), .B(n188), .Z(n185) );
  NAND U223 ( .A(B[29]), .B(n189), .Z(n188) );
  NANDN U224 ( .A(A[29]), .B(n190), .Z(n189) );
  NANDN U225 ( .A(n190), .B(A[29]), .Z(n187) );
  XOR U226 ( .A(n191), .B(n192), .Z(SUM[2]) );
  XOR U227 ( .A(B[2]), .B(A[2]), .Z(n192) );
  XOR U228 ( .A(n190), .B(n193), .Z(SUM[29]) );
  XNOR U229 ( .A(B[29]), .B(A[29]), .Z(n193) );
  AND U230 ( .A(n194), .B(n195), .Z(n190) );
  NAND U231 ( .A(B[28]), .B(n196), .Z(n195) );
  NANDN U232 ( .A(A[28]), .B(n197), .Z(n196) );
  NANDN U233 ( .A(n197), .B(A[28]), .Z(n194) );
  XOR U234 ( .A(n197), .B(n198), .Z(SUM[28]) );
  XNOR U235 ( .A(B[28]), .B(A[28]), .Z(n198) );
  AND U236 ( .A(n199), .B(n200), .Z(n197) );
  NAND U237 ( .A(B[27]), .B(n201), .Z(n200) );
  NANDN U238 ( .A(A[27]), .B(n202), .Z(n201) );
  NANDN U239 ( .A(n202), .B(A[27]), .Z(n199) );
  XOR U240 ( .A(n202), .B(n203), .Z(SUM[27]) );
  XNOR U241 ( .A(B[27]), .B(A[27]), .Z(n203) );
  AND U242 ( .A(n204), .B(n205), .Z(n202) );
  NAND U243 ( .A(B[26]), .B(n206), .Z(n205) );
  NANDN U244 ( .A(A[26]), .B(n207), .Z(n206) );
  NANDN U245 ( .A(n207), .B(A[26]), .Z(n204) );
  XOR U246 ( .A(n207), .B(n208), .Z(SUM[26]) );
  XNOR U247 ( .A(B[26]), .B(A[26]), .Z(n208) );
  AND U248 ( .A(n209), .B(n210), .Z(n207) );
  NAND U249 ( .A(B[25]), .B(n211), .Z(n210) );
  NANDN U250 ( .A(A[25]), .B(n212), .Z(n211) );
  NANDN U251 ( .A(n212), .B(A[25]), .Z(n209) );
  XOR U252 ( .A(n212), .B(n213), .Z(SUM[25]) );
  XNOR U253 ( .A(B[25]), .B(A[25]), .Z(n213) );
  AND U254 ( .A(n214), .B(n215), .Z(n212) );
  NAND U255 ( .A(B[24]), .B(n216), .Z(n215) );
  NANDN U256 ( .A(A[24]), .B(n217), .Z(n216) );
  NANDN U257 ( .A(n217), .B(A[24]), .Z(n214) );
  XOR U258 ( .A(n217), .B(n218), .Z(SUM[24]) );
  XNOR U259 ( .A(B[24]), .B(A[24]), .Z(n218) );
  AND U260 ( .A(n219), .B(n220), .Z(n217) );
  NAND U261 ( .A(B[23]), .B(n221), .Z(n220) );
  NANDN U262 ( .A(A[23]), .B(n222), .Z(n221) );
  NANDN U263 ( .A(n222), .B(A[23]), .Z(n219) );
  XOR U264 ( .A(n222), .B(n223), .Z(SUM[23]) );
  XNOR U265 ( .A(B[23]), .B(A[23]), .Z(n223) );
  AND U266 ( .A(n224), .B(n225), .Z(n222) );
  NAND U267 ( .A(B[22]), .B(n226), .Z(n225) );
  NANDN U268 ( .A(A[22]), .B(n227), .Z(n226) );
  NANDN U269 ( .A(n227), .B(A[22]), .Z(n224) );
  XOR U270 ( .A(n227), .B(n228), .Z(SUM[22]) );
  XNOR U271 ( .A(B[22]), .B(A[22]), .Z(n228) );
  AND U272 ( .A(n229), .B(n230), .Z(n227) );
  NAND U273 ( .A(B[21]), .B(n231), .Z(n230) );
  NANDN U274 ( .A(A[21]), .B(n232), .Z(n231) );
  NANDN U275 ( .A(n232), .B(A[21]), .Z(n229) );
  XOR U276 ( .A(n232), .B(n233), .Z(SUM[21]) );
  XNOR U277 ( .A(B[21]), .B(A[21]), .Z(n233) );
  AND U278 ( .A(n234), .B(n235), .Z(n232) );
  NAND U279 ( .A(B[20]), .B(n236), .Z(n235) );
  NANDN U280 ( .A(A[20]), .B(n237), .Z(n236) );
  NANDN U281 ( .A(n237), .B(A[20]), .Z(n234) );
  XOR U282 ( .A(n237), .B(n238), .Z(SUM[20]) );
  XNOR U283 ( .A(B[20]), .B(A[20]), .Z(n238) );
  AND U284 ( .A(n239), .B(n240), .Z(n237) );
  NAND U285 ( .A(B[19]), .B(n241), .Z(n240) );
  NANDN U286 ( .A(A[19]), .B(n242), .Z(n241) );
  NANDN U287 ( .A(n242), .B(A[19]), .Z(n239) );
  XOR U288 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U289 ( .A(n242), .B(n243), .Z(SUM[19]) );
  XNOR U290 ( .A(B[19]), .B(A[19]), .Z(n243) );
  AND U291 ( .A(n244), .B(n245), .Z(n242) );
  NAND U292 ( .A(B[18]), .B(n246), .Z(n245) );
  NANDN U293 ( .A(A[18]), .B(n247), .Z(n246) );
  NANDN U294 ( .A(n247), .B(A[18]), .Z(n244) );
  XOR U295 ( .A(n247), .B(n248), .Z(SUM[18]) );
  XNOR U296 ( .A(B[18]), .B(A[18]), .Z(n248) );
  AND U297 ( .A(n249), .B(n250), .Z(n247) );
  NAND U298 ( .A(B[17]), .B(n251), .Z(n250) );
  NANDN U299 ( .A(A[17]), .B(n252), .Z(n251) );
  NANDN U300 ( .A(n252), .B(A[17]), .Z(n249) );
  XOR U301 ( .A(n252), .B(n253), .Z(SUM[17]) );
  XNOR U302 ( .A(B[17]), .B(A[17]), .Z(n253) );
  AND U303 ( .A(n254), .B(n255), .Z(n252) );
  NAND U304 ( .A(B[16]), .B(n256), .Z(n255) );
  NANDN U305 ( .A(A[16]), .B(n257), .Z(n256) );
  NANDN U306 ( .A(n257), .B(A[16]), .Z(n254) );
  XOR U307 ( .A(n257), .B(n258), .Z(SUM[16]) );
  XNOR U308 ( .A(B[16]), .B(A[16]), .Z(n258) );
  AND U309 ( .A(n259), .B(n260), .Z(n257) );
  NAND U310 ( .A(B[15]), .B(n261), .Z(n260) );
  NANDN U311 ( .A(A[15]), .B(n262), .Z(n261) );
  NANDN U312 ( .A(n262), .B(A[15]), .Z(n259) );
  XOR U313 ( .A(n262), .B(n263), .Z(SUM[15]) );
  XNOR U314 ( .A(B[15]), .B(A[15]), .Z(n263) );
  AND U315 ( .A(n264), .B(n265), .Z(n262) );
  NAND U316 ( .A(B[14]), .B(n266), .Z(n265) );
  NANDN U317 ( .A(A[14]), .B(n267), .Z(n266) );
  NANDN U318 ( .A(n267), .B(A[14]), .Z(n264) );
  XOR U319 ( .A(n267), .B(n268), .Z(SUM[14]) );
  XNOR U320 ( .A(B[14]), .B(A[14]), .Z(n268) );
  AND U321 ( .A(n269), .B(n270), .Z(n267) );
  NAND U322 ( .A(B[13]), .B(n271), .Z(n270) );
  NANDN U323 ( .A(A[13]), .B(n272), .Z(n271) );
  NANDN U324 ( .A(n272), .B(A[13]), .Z(n269) );
  XOR U325 ( .A(n272), .B(n273), .Z(SUM[13]) );
  XNOR U326 ( .A(B[13]), .B(A[13]), .Z(n273) );
  AND U327 ( .A(n274), .B(n275), .Z(n272) );
  NAND U328 ( .A(B[12]), .B(n276), .Z(n275) );
  NANDN U329 ( .A(A[12]), .B(n277), .Z(n276) );
  NANDN U330 ( .A(n277), .B(A[12]), .Z(n274) );
  XOR U331 ( .A(n277), .B(n278), .Z(SUM[12]) );
  XNOR U332 ( .A(B[12]), .B(A[12]), .Z(n278) );
  AND U333 ( .A(n279), .B(n280), .Z(n277) );
  NAND U334 ( .A(B[11]), .B(n281), .Z(n280) );
  NANDN U335 ( .A(A[11]), .B(n282), .Z(n281) );
  NANDN U336 ( .A(n282), .B(A[11]), .Z(n279) );
  XOR U337 ( .A(n282), .B(n283), .Z(SUM[11]) );
  XNOR U338 ( .A(B[11]), .B(A[11]), .Z(n283) );
  AND U339 ( .A(n284), .B(n285), .Z(n282) );
  NAND U340 ( .A(B[10]), .B(n286), .Z(n285) );
  NANDN U341 ( .A(A[10]), .B(n287), .Z(n286) );
  NANDN U342 ( .A(n287), .B(A[10]), .Z(n284) );
  XOR U343 ( .A(n287), .B(n288), .Z(SUM[10]) );
  XNOR U344 ( .A(B[10]), .B(A[10]), .Z(n288) );
  AND U345 ( .A(n289), .B(n290), .Z(n287) );
  NAND U346 ( .A(B[9]), .B(n291), .Z(n290) );
  OR U347 ( .A(n1), .B(A[9]), .Z(n291) );
  NAND U348 ( .A(A[9]), .B(n1), .Z(n289) );
  NAND U349 ( .A(n292), .B(n293), .Z(n1) );
  NAND U350 ( .A(B[8]), .B(n294), .Z(n293) );
  NANDN U351 ( .A(A[8]), .B(n3), .Z(n294) );
  NANDN U352 ( .A(n3), .B(A[8]), .Z(n292) );
  AND U353 ( .A(n295), .B(n296), .Z(n3) );
  NAND U354 ( .A(B[7]), .B(n297), .Z(n296) );
  NANDN U355 ( .A(A[7]), .B(n5), .Z(n297) );
  NANDN U356 ( .A(n5), .B(A[7]), .Z(n295) );
  AND U357 ( .A(n298), .B(n299), .Z(n5) );
  NAND U358 ( .A(B[6]), .B(n300), .Z(n299) );
  NANDN U359 ( .A(A[6]), .B(n7), .Z(n300) );
  NANDN U360 ( .A(n7), .B(A[6]), .Z(n298) );
  AND U361 ( .A(n301), .B(n302), .Z(n7) );
  NAND U362 ( .A(B[5]), .B(n303), .Z(n302) );
  NANDN U363 ( .A(A[5]), .B(n35), .Z(n303) );
  NANDN U364 ( .A(n35), .B(A[5]), .Z(n301) );
  AND U365 ( .A(n304), .B(n305), .Z(n35) );
  NAND U366 ( .A(B[4]), .B(n306), .Z(n305) );
  NANDN U367 ( .A(A[4]), .B(n87), .Z(n306) );
  NANDN U368 ( .A(n87), .B(A[4]), .Z(n304) );
  AND U369 ( .A(n307), .B(n308), .Z(n87) );
  NAND U370 ( .A(B[3]), .B(n309), .Z(n308) );
  NANDN U371 ( .A(A[3]), .B(n139), .Z(n309) );
  NANDN U372 ( .A(n139), .B(A[3]), .Z(n307) );
  AND U373 ( .A(n310), .B(n311), .Z(n139) );
  NAND U374 ( .A(B[2]), .B(n312), .Z(n311) );
  OR U375 ( .A(n191), .B(A[2]), .Z(n312) );
  NAND U376 ( .A(A[2]), .B(n191), .Z(n310) );
  AND U377 ( .A(B[1]), .B(A[1]), .Z(n191) );
endmodule


module modmult_step_N64 ( xregN_1, y, n, zin, zout );
  input [63:0] y;
  input [63:0] n;
  input [65:0] zin;
  output [65:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N72, N73, N74, N75,
         N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N204, N203, N202, N201, N200, N199, N198, N197, N196,
         N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185,
         N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174,
         N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163,
         N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152,
         N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141,
         N138, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271;
  wire   [65:0] z2;
  wire   [65:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N64_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N204, N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, 
        N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, 
        N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, 
        N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, 
        N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, 
        N142, N141}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N64_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N138), .TC(1'b0), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__0, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141}) );
  modmult_step_N64_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N138) );
  modmult_step_N64_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(1'b0), 
        .DIFF({N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, 
        N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        N76, N75, N74, N73, N72}) );
  modmult_step_N64_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(1'b0), .TC(1'b0), .LT_LE(N70) );
  modmult_step_N64_DW01_add_0 add_119 ( .A({zin[64:0], 1'b0}), .B({1'b0, 1'b0, 
        y}), .CI(1'b0), .SUM({N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N70), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N81), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[8]) );
  NANDN U9 ( .A(N70), .B(z2[8]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N80), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[7]) );
  NANDN U17 ( .A(N70), .B(z2[7]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N79), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[6]) );
  NANDN U20 ( .A(N70), .B(z2[6]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N78), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[65]) );
  NANDN U23 ( .A(N70), .B(z2[65]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N137), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[64]) );
  NANDN U26 ( .A(N70), .B(z2[64]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N136), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[63]) );
  NANDN U29 ( .A(N70), .B(z2[63]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N135), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[62]) );
  NANDN U32 ( .A(N70), .B(z2[62]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N134), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[61]) );
  NANDN U35 ( .A(N70), .B(z2[61]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N133), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[60]) );
  NANDN U38 ( .A(N70), .B(z2[60]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N132), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[5]) );
  NANDN U41 ( .A(N70), .B(z2[5]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N77), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[59]) );
  NANDN U44 ( .A(N70), .B(z2[59]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N131), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[58]) );
  NANDN U47 ( .A(N70), .B(z2[58]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N130), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[57]) );
  NANDN U50 ( .A(N70), .B(z2[57]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N129), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[56]) );
  NANDN U53 ( .A(N70), .B(z2[56]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N128), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[55]) );
  NANDN U56 ( .A(N70), .B(z2[55]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N127), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[54]) );
  NANDN U59 ( .A(N70), .B(z2[54]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N126), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[53]) );
  NANDN U62 ( .A(N70), .B(z2[53]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N125), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[52]) );
  NANDN U65 ( .A(N70), .B(z2[52]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N124), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[51]) );
  NANDN U68 ( .A(N70), .B(z2[51]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N123), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[50]) );
  NANDN U71 ( .A(N70), .B(z2[50]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N122), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[4]) );
  NANDN U74 ( .A(N70), .B(z2[4]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N76), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[49]) );
  NANDN U77 ( .A(N70), .B(z2[49]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N121), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[48]) );
  NANDN U80 ( .A(N70), .B(z2[48]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N120), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[47]) );
  NANDN U83 ( .A(N70), .B(z2[47]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N119), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[46]) );
  NANDN U86 ( .A(N70), .B(z2[46]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N118), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[45]) );
  NANDN U89 ( .A(N70), .B(z2[45]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N117), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[44]) );
  NANDN U92 ( .A(N70), .B(z2[44]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N116), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[43]) );
  NANDN U95 ( .A(N70), .B(z2[43]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N115), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[42]) );
  NANDN U98 ( .A(N70), .B(z2[42]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N114), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[41]) );
  NANDN U101 ( .A(N70), .B(z2[41]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N113), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[40]) );
  NANDN U104 ( .A(N70), .B(z2[40]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N112), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[3]) );
  NANDN U107 ( .A(N70), .B(z2[3]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N75), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[39]) );
  NANDN U110 ( .A(N70), .B(z2[39]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N111), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[38]) );
  NANDN U113 ( .A(N70), .B(z2[38]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N110), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[37]) );
  NANDN U116 ( .A(N70), .B(z2[37]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N109), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[36]) );
  NANDN U119 ( .A(N70), .B(z2[36]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N108), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[35]) );
  NANDN U122 ( .A(N70), .B(z2[35]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N107), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[34]) );
  NANDN U125 ( .A(N70), .B(z2[34]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N106), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[33]) );
  NANDN U128 ( .A(N70), .B(z2[33]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N105), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[32]) );
  NANDN U131 ( .A(N70), .B(z2[32]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N104), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[31]) );
  NANDN U134 ( .A(N70), .B(z2[31]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N103), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[30]) );
  NANDN U137 ( .A(N70), .B(z2[30]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N102), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[2]) );
  NANDN U140 ( .A(N70), .B(z2[2]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N74), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[29]) );
  NANDN U143 ( .A(N70), .B(z2[29]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N101), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[28]) );
  NANDN U146 ( .A(N70), .B(z2[28]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N100), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[27]) );
  NANDN U149 ( .A(N70), .B(z2[27]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N99), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[26]) );
  NANDN U152 ( .A(N70), .B(z2[26]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N98), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[25]) );
  NANDN U155 ( .A(N70), .B(z2[25]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N97), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[24]) );
  NANDN U158 ( .A(N70), .B(z2[24]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N96), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[23]) );
  NANDN U161 ( .A(N70), .B(z2[23]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N95), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[22]) );
  NANDN U164 ( .A(N70), .B(z2[22]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N94), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[21]) );
  NANDN U167 ( .A(N70), .B(z2[21]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N93), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[20]) );
  NANDN U170 ( .A(N70), .B(z2[20]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N92), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[1]) );
  NANDN U173 ( .A(N70), .B(z2[1]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N73), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[19]) );
  NANDN U176 ( .A(N70), .B(z2[19]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N91), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[18]) );
  NANDN U179 ( .A(N70), .B(z2[18]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N90), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[17]) );
  NANDN U182 ( .A(N70), .B(z2[17]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N89), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[16]) );
  NANDN U185 ( .A(N70), .B(z2[16]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N88), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[15]) );
  NANDN U188 ( .A(N70), .B(z2[15]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N87), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[14]) );
  NANDN U191 ( .A(N70), .B(z2[14]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N86), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[13]) );
  NANDN U194 ( .A(N70), .B(z2[13]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N85), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[12]) );
  NANDN U197 ( .A(N70), .B(z2[12]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N84), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[11]) );
  NANDN U200 ( .A(N70), .B(z2[11]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N83), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[10]) );
  NANDN U203 ( .A(N70), .B(z2[10]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N82), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[0]) );
  NANDN U206 ( .A(N70), .B(z2[0]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N72), .Z(n140) );
  IV U208 ( .A(N70), .Z(n3) );
  NAND U209 ( .A(n142), .B(n143), .Z(z2[9]) );
  NANDN U210 ( .A(xregN_1), .B(zin[8]), .Z(n143) );
  NAND U211 ( .A(N13), .B(xregN_1), .Z(n142) );
  NAND U212 ( .A(n144), .B(n145), .Z(z2[8]) );
  NANDN U213 ( .A(xregN_1), .B(zin[7]), .Z(n145) );
  NAND U214 ( .A(N12), .B(xregN_1), .Z(n144) );
  NAND U215 ( .A(n146), .B(n147), .Z(z2[7]) );
  NANDN U216 ( .A(xregN_1), .B(zin[6]), .Z(n147) );
  NAND U217 ( .A(N11), .B(xregN_1), .Z(n146) );
  NAND U218 ( .A(n148), .B(n149), .Z(z2[6]) );
  NANDN U219 ( .A(xregN_1), .B(zin[5]), .Z(n149) );
  NAND U220 ( .A(N10), .B(xregN_1), .Z(n148) );
  NAND U221 ( .A(n150), .B(n151), .Z(z2[65]) );
  NANDN U222 ( .A(xregN_1), .B(zin[64]), .Z(n151) );
  NAND U223 ( .A(N69), .B(xregN_1), .Z(n150) );
  NAND U224 ( .A(n152), .B(n153), .Z(z2[64]) );
  NANDN U225 ( .A(xregN_1), .B(zin[63]), .Z(n153) );
  NAND U226 ( .A(N68), .B(xregN_1), .Z(n152) );
  NAND U227 ( .A(n154), .B(n155), .Z(z2[63]) );
  NANDN U228 ( .A(xregN_1), .B(zin[62]), .Z(n155) );
  NAND U229 ( .A(N67), .B(xregN_1), .Z(n154) );
  NAND U230 ( .A(n156), .B(n157), .Z(z2[62]) );
  NANDN U231 ( .A(xregN_1), .B(zin[61]), .Z(n157) );
  NAND U232 ( .A(N66), .B(xregN_1), .Z(n156) );
  NAND U233 ( .A(n158), .B(n159), .Z(z2[61]) );
  NANDN U234 ( .A(xregN_1), .B(zin[60]), .Z(n159) );
  NAND U235 ( .A(N65), .B(xregN_1), .Z(n158) );
  NAND U236 ( .A(n160), .B(n161), .Z(z2[60]) );
  NANDN U237 ( .A(xregN_1), .B(zin[59]), .Z(n161) );
  NAND U238 ( .A(N64), .B(xregN_1), .Z(n160) );
  NAND U239 ( .A(n162), .B(n163), .Z(z2[5]) );
  NANDN U240 ( .A(xregN_1), .B(zin[4]), .Z(n163) );
  NAND U241 ( .A(N9), .B(xregN_1), .Z(n162) );
  NAND U242 ( .A(n164), .B(n165), .Z(z2[59]) );
  NANDN U243 ( .A(xregN_1), .B(zin[58]), .Z(n165) );
  NAND U244 ( .A(N63), .B(xregN_1), .Z(n164) );
  NAND U245 ( .A(n166), .B(n167), .Z(z2[58]) );
  NANDN U246 ( .A(xregN_1), .B(zin[57]), .Z(n167) );
  NAND U247 ( .A(N62), .B(xregN_1), .Z(n166) );
  NAND U248 ( .A(n168), .B(n169), .Z(z2[57]) );
  NANDN U249 ( .A(xregN_1), .B(zin[56]), .Z(n169) );
  NAND U250 ( .A(N61), .B(xregN_1), .Z(n168) );
  NAND U251 ( .A(n170), .B(n171), .Z(z2[56]) );
  NANDN U252 ( .A(xregN_1), .B(zin[55]), .Z(n171) );
  NAND U253 ( .A(N60), .B(xregN_1), .Z(n170) );
  NAND U254 ( .A(n172), .B(n173), .Z(z2[55]) );
  NANDN U255 ( .A(xregN_1), .B(zin[54]), .Z(n173) );
  NAND U256 ( .A(N59), .B(xregN_1), .Z(n172) );
  NAND U257 ( .A(n174), .B(n175), .Z(z2[54]) );
  NANDN U258 ( .A(xregN_1), .B(zin[53]), .Z(n175) );
  NAND U259 ( .A(N58), .B(xregN_1), .Z(n174) );
  NAND U260 ( .A(n176), .B(n177), .Z(z2[53]) );
  NANDN U261 ( .A(xregN_1), .B(zin[52]), .Z(n177) );
  NAND U262 ( .A(N57), .B(xregN_1), .Z(n176) );
  NAND U263 ( .A(n178), .B(n179), .Z(z2[52]) );
  NANDN U264 ( .A(xregN_1), .B(zin[51]), .Z(n179) );
  NAND U265 ( .A(N56), .B(xregN_1), .Z(n178) );
  NAND U266 ( .A(n180), .B(n181), .Z(z2[51]) );
  NANDN U267 ( .A(xregN_1), .B(zin[50]), .Z(n181) );
  NAND U268 ( .A(N55), .B(xregN_1), .Z(n180) );
  NAND U269 ( .A(n182), .B(n183), .Z(z2[50]) );
  NANDN U270 ( .A(xregN_1), .B(zin[49]), .Z(n183) );
  NAND U271 ( .A(N54), .B(xregN_1), .Z(n182) );
  NAND U272 ( .A(n184), .B(n185), .Z(z2[4]) );
  NANDN U273 ( .A(xregN_1), .B(zin[3]), .Z(n185) );
  NAND U274 ( .A(N8), .B(xregN_1), .Z(n184) );
  NAND U275 ( .A(n186), .B(n187), .Z(z2[49]) );
  NANDN U276 ( .A(xregN_1), .B(zin[48]), .Z(n187) );
  NAND U277 ( .A(N53), .B(xregN_1), .Z(n186) );
  NAND U278 ( .A(n188), .B(n189), .Z(z2[48]) );
  NANDN U279 ( .A(xregN_1), .B(zin[47]), .Z(n189) );
  NAND U280 ( .A(N52), .B(xregN_1), .Z(n188) );
  NAND U281 ( .A(n190), .B(n191), .Z(z2[47]) );
  NANDN U282 ( .A(xregN_1), .B(zin[46]), .Z(n191) );
  NAND U283 ( .A(N51), .B(xregN_1), .Z(n190) );
  NAND U284 ( .A(n192), .B(n193), .Z(z2[46]) );
  NANDN U285 ( .A(xregN_1), .B(zin[45]), .Z(n193) );
  NAND U286 ( .A(N50), .B(xregN_1), .Z(n192) );
  NAND U287 ( .A(n194), .B(n195), .Z(z2[45]) );
  NANDN U288 ( .A(xregN_1), .B(zin[44]), .Z(n195) );
  NAND U289 ( .A(N49), .B(xregN_1), .Z(n194) );
  NAND U290 ( .A(n196), .B(n197), .Z(z2[44]) );
  NANDN U291 ( .A(xregN_1), .B(zin[43]), .Z(n197) );
  NAND U292 ( .A(N48), .B(xregN_1), .Z(n196) );
  NAND U293 ( .A(n198), .B(n199), .Z(z2[43]) );
  NANDN U294 ( .A(xregN_1), .B(zin[42]), .Z(n199) );
  NAND U295 ( .A(N47), .B(xregN_1), .Z(n198) );
  NAND U296 ( .A(n200), .B(n201), .Z(z2[42]) );
  NANDN U297 ( .A(xregN_1), .B(zin[41]), .Z(n201) );
  NAND U298 ( .A(N46), .B(xregN_1), .Z(n200) );
  NAND U299 ( .A(n202), .B(n203), .Z(z2[41]) );
  NANDN U300 ( .A(xregN_1), .B(zin[40]), .Z(n203) );
  NAND U301 ( .A(N45), .B(xregN_1), .Z(n202) );
  NAND U302 ( .A(n204), .B(n205), .Z(z2[40]) );
  NANDN U303 ( .A(xregN_1), .B(zin[39]), .Z(n205) );
  NAND U304 ( .A(N44), .B(xregN_1), .Z(n204) );
  NAND U305 ( .A(n206), .B(n207), .Z(z2[3]) );
  NANDN U306 ( .A(xregN_1), .B(zin[2]), .Z(n207) );
  NAND U307 ( .A(N7), .B(xregN_1), .Z(n206) );
  NAND U308 ( .A(n208), .B(n209), .Z(z2[39]) );
  NANDN U309 ( .A(xregN_1), .B(zin[38]), .Z(n209) );
  NAND U310 ( .A(N43), .B(xregN_1), .Z(n208) );
  NAND U311 ( .A(n210), .B(n211), .Z(z2[38]) );
  NANDN U312 ( .A(xregN_1), .B(zin[37]), .Z(n211) );
  NAND U313 ( .A(N42), .B(xregN_1), .Z(n210) );
  NAND U314 ( .A(n212), .B(n213), .Z(z2[37]) );
  NANDN U315 ( .A(xregN_1), .B(zin[36]), .Z(n213) );
  NAND U316 ( .A(N41), .B(xregN_1), .Z(n212) );
  NAND U317 ( .A(n214), .B(n215), .Z(z2[36]) );
  NANDN U318 ( .A(xregN_1), .B(zin[35]), .Z(n215) );
  NAND U319 ( .A(N40), .B(xregN_1), .Z(n214) );
  NAND U320 ( .A(n216), .B(n217), .Z(z2[35]) );
  NANDN U321 ( .A(xregN_1), .B(zin[34]), .Z(n217) );
  NAND U322 ( .A(N39), .B(xregN_1), .Z(n216) );
  NAND U323 ( .A(n218), .B(n219), .Z(z2[34]) );
  NANDN U324 ( .A(xregN_1), .B(zin[33]), .Z(n219) );
  NAND U325 ( .A(N38), .B(xregN_1), .Z(n218) );
  NAND U326 ( .A(n220), .B(n221), .Z(z2[33]) );
  NANDN U327 ( .A(xregN_1), .B(zin[32]), .Z(n221) );
  NAND U328 ( .A(N37), .B(xregN_1), .Z(n220) );
  NAND U329 ( .A(n222), .B(n223), .Z(z2[32]) );
  NANDN U330 ( .A(xregN_1), .B(zin[31]), .Z(n223) );
  NAND U331 ( .A(N36), .B(xregN_1), .Z(n222) );
  NAND U332 ( .A(n224), .B(n225), .Z(z2[31]) );
  NANDN U333 ( .A(xregN_1), .B(zin[30]), .Z(n225) );
  NAND U334 ( .A(N35), .B(xregN_1), .Z(n224) );
  NAND U335 ( .A(n226), .B(n227), .Z(z2[30]) );
  NANDN U336 ( .A(xregN_1), .B(zin[29]), .Z(n227) );
  NAND U337 ( .A(N34), .B(xregN_1), .Z(n226) );
  NAND U338 ( .A(n228), .B(n229), .Z(z2[2]) );
  NANDN U339 ( .A(xregN_1), .B(zin[1]), .Z(n229) );
  NAND U340 ( .A(N6), .B(xregN_1), .Z(n228) );
  NAND U341 ( .A(n230), .B(n231), .Z(z2[29]) );
  NANDN U342 ( .A(xregN_1), .B(zin[28]), .Z(n231) );
  NAND U343 ( .A(N33), .B(xregN_1), .Z(n230) );
  NAND U344 ( .A(n232), .B(n233), .Z(z2[28]) );
  NANDN U345 ( .A(xregN_1), .B(zin[27]), .Z(n233) );
  NAND U346 ( .A(N32), .B(xregN_1), .Z(n232) );
  NAND U347 ( .A(n234), .B(n235), .Z(z2[27]) );
  NANDN U348 ( .A(xregN_1), .B(zin[26]), .Z(n235) );
  NAND U349 ( .A(N31), .B(xregN_1), .Z(n234) );
  NAND U350 ( .A(n236), .B(n237), .Z(z2[26]) );
  NANDN U351 ( .A(xregN_1), .B(zin[25]), .Z(n237) );
  NAND U352 ( .A(N30), .B(xregN_1), .Z(n236) );
  NAND U353 ( .A(n238), .B(n239), .Z(z2[25]) );
  NANDN U354 ( .A(xregN_1), .B(zin[24]), .Z(n239) );
  NAND U355 ( .A(N29), .B(xregN_1), .Z(n238) );
  NAND U356 ( .A(n240), .B(n241), .Z(z2[24]) );
  NANDN U357 ( .A(xregN_1), .B(zin[23]), .Z(n241) );
  NAND U358 ( .A(N28), .B(xregN_1), .Z(n240) );
  NAND U359 ( .A(n242), .B(n243), .Z(z2[23]) );
  NANDN U360 ( .A(xregN_1), .B(zin[22]), .Z(n243) );
  NAND U361 ( .A(N27), .B(xregN_1), .Z(n242) );
  NAND U362 ( .A(n244), .B(n245), .Z(z2[22]) );
  NANDN U363 ( .A(xregN_1), .B(zin[21]), .Z(n245) );
  NAND U364 ( .A(N26), .B(xregN_1), .Z(n244) );
  NAND U365 ( .A(n246), .B(n247), .Z(z2[21]) );
  NANDN U366 ( .A(xregN_1), .B(zin[20]), .Z(n247) );
  NAND U367 ( .A(N25), .B(xregN_1), .Z(n246) );
  NAND U368 ( .A(n248), .B(n249), .Z(z2[20]) );
  NANDN U369 ( .A(xregN_1), .B(zin[19]), .Z(n249) );
  NAND U370 ( .A(N24), .B(xregN_1), .Z(n248) );
  NAND U371 ( .A(n250), .B(n251), .Z(z2[1]) );
  NANDN U372 ( .A(xregN_1), .B(zin[0]), .Z(n251) );
  NAND U373 ( .A(N5), .B(xregN_1), .Z(n250) );
  NAND U374 ( .A(n252), .B(n253), .Z(z2[19]) );
  NANDN U375 ( .A(xregN_1), .B(zin[18]), .Z(n253) );
  NAND U376 ( .A(N23), .B(xregN_1), .Z(n252) );
  NAND U377 ( .A(n254), .B(n255), .Z(z2[18]) );
  NANDN U378 ( .A(xregN_1), .B(zin[17]), .Z(n255) );
  NAND U379 ( .A(N22), .B(xregN_1), .Z(n254) );
  NAND U380 ( .A(n256), .B(n257), .Z(z2[17]) );
  NANDN U381 ( .A(xregN_1), .B(zin[16]), .Z(n257) );
  NAND U382 ( .A(N21), .B(xregN_1), .Z(n256) );
  NAND U383 ( .A(n258), .B(n259), .Z(z2[16]) );
  NANDN U384 ( .A(xregN_1), .B(zin[15]), .Z(n259) );
  NAND U385 ( .A(N20), .B(xregN_1), .Z(n258) );
  NAND U386 ( .A(n260), .B(n261), .Z(z2[15]) );
  NANDN U387 ( .A(xregN_1), .B(zin[14]), .Z(n261) );
  NAND U388 ( .A(N19), .B(xregN_1), .Z(n260) );
  NAND U389 ( .A(n262), .B(n263), .Z(z2[14]) );
  NANDN U390 ( .A(xregN_1), .B(zin[13]), .Z(n263) );
  NAND U391 ( .A(N18), .B(xregN_1), .Z(n262) );
  NAND U392 ( .A(n264), .B(n265), .Z(z2[13]) );
  NANDN U393 ( .A(xregN_1), .B(zin[12]), .Z(n265) );
  NAND U394 ( .A(N17), .B(xregN_1), .Z(n264) );
  NAND U395 ( .A(n266), .B(n267), .Z(z2[12]) );
  NANDN U396 ( .A(xregN_1), .B(zin[11]), .Z(n267) );
  NAND U397 ( .A(N16), .B(xregN_1), .Z(n266) );
  NAND U398 ( .A(n268), .B(n269), .Z(z2[11]) );
  NANDN U399 ( .A(xregN_1), .B(zin[10]), .Z(n269) );
  NAND U400 ( .A(N15), .B(xregN_1), .Z(n268) );
  NAND U401 ( .A(n270), .B(n271), .Z(z2[10]) );
  NANDN U402 ( .A(xregN_1), .B(zin[9]), .Z(n271) );
  NAND U403 ( .A(N14), .B(xregN_1), .Z(n270) );
  AND U404 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_N64_CC64 ( clk, rst, start, x, y, n, o );
  input [63:0] x;
  input [63:0] y;
  input [63:0] n;
  output [63:0] o;
  input clk, rst, start;
  wire   \zout[0][65] , \zout[0][64] , \zin[0][65] , \zin[0][64] ,
         \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] ,
         \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] ,
         \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] ,
         \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] ,
         \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] ,
         \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] ,
         \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] ,
         \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] ,
         \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] ,
         \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] ,
         \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] ,
         \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] ,
         \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127;
  wire   [65:0] zreg;
  wire   [63:0] xin;
  wire   [63:0] xreg;

  DFF \xreg_reg[1]  ( .D(n127), .CLK(clk), .RST(rst), .Q(xreg[1]) );
  DFF \xreg_reg[2]  ( .D(xin[1]), .CLK(clk), .RST(rst), .Q(xreg[2]) );
  DFF \xreg_reg[3]  ( .D(xin[2]), .CLK(clk), .RST(rst), .Q(xreg[3]) );
  DFF \xreg_reg[4]  ( .D(xin[3]), .CLK(clk), .RST(rst), .Q(xreg[4]) );
  DFF \xreg_reg[5]  ( .D(xin[4]), .CLK(clk), .RST(rst), .Q(xreg[5]) );
  DFF \xreg_reg[6]  ( .D(xin[5]), .CLK(clk), .RST(rst), .Q(xreg[6]) );
  DFF \xreg_reg[7]  ( .D(xin[6]), .CLK(clk), .RST(rst), .Q(xreg[7]) );
  DFF \xreg_reg[8]  ( .D(xin[7]), .CLK(clk), .RST(rst), .Q(xreg[8]) );
  DFF \xreg_reg[9]  ( .D(xin[8]), .CLK(clk), .RST(rst), .Q(xreg[9]) );
  DFF \xreg_reg[10]  ( .D(xin[9]), .CLK(clk), .RST(rst), .Q(xreg[10]) );
  DFF \xreg_reg[11]  ( .D(xin[10]), .CLK(clk), .RST(rst), .Q(xreg[11]) );
  DFF \xreg_reg[12]  ( .D(xin[11]), .CLK(clk), .RST(rst), .Q(xreg[12]) );
  DFF \xreg_reg[13]  ( .D(xin[12]), .CLK(clk), .RST(rst), .Q(xreg[13]) );
  DFF \xreg_reg[14]  ( .D(xin[13]), .CLK(clk), .RST(rst), .Q(xreg[14]) );
  DFF \xreg_reg[15]  ( .D(xin[14]), .CLK(clk), .RST(rst), .Q(xreg[15]) );
  DFF \xreg_reg[16]  ( .D(xin[15]), .CLK(clk), .RST(rst), .Q(xreg[16]) );
  DFF \xreg_reg[17]  ( .D(xin[16]), .CLK(clk), .RST(rst), .Q(xreg[17]) );
  DFF \xreg_reg[18]  ( .D(xin[17]), .CLK(clk), .RST(rst), .Q(xreg[18]) );
  DFF \xreg_reg[19]  ( .D(xin[18]), .CLK(clk), .RST(rst), .Q(xreg[19]) );
  DFF \xreg_reg[20]  ( .D(xin[19]), .CLK(clk), .RST(rst), .Q(xreg[20]) );
  DFF \xreg_reg[21]  ( .D(xin[20]), .CLK(clk), .RST(rst), .Q(xreg[21]) );
  DFF \xreg_reg[22]  ( .D(xin[21]), .CLK(clk), .RST(rst), .Q(xreg[22]) );
  DFF \xreg_reg[23]  ( .D(xin[22]), .CLK(clk), .RST(rst), .Q(xreg[23]) );
  DFF \xreg_reg[24]  ( .D(xin[23]), .CLK(clk), .RST(rst), .Q(xreg[24]) );
  DFF \xreg_reg[25]  ( .D(xin[24]), .CLK(clk), .RST(rst), .Q(xreg[25]) );
  DFF \xreg_reg[26]  ( .D(xin[25]), .CLK(clk), .RST(rst), .Q(xreg[26]) );
  DFF \xreg_reg[27]  ( .D(xin[26]), .CLK(clk), .RST(rst), .Q(xreg[27]) );
  DFF \xreg_reg[28]  ( .D(xin[27]), .CLK(clk), .RST(rst), .Q(xreg[28]) );
  DFF \xreg_reg[29]  ( .D(xin[28]), .CLK(clk), .RST(rst), .Q(xreg[29]) );
  DFF \xreg_reg[30]  ( .D(xin[29]), .CLK(clk), .RST(rst), .Q(xreg[30]) );
  DFF \xreg_reg[31]  ( .D(xin[30]), .CLK(clk), .RST(rst), .Q(xreg[31]) );
  DFF \xreg_reg[32]  ( .D(xin[31]), .CLK(clk), .RST(rst), .Q(xreg[32]) );
  DFF \xreg_reg[33]  ( .D(xin[32]), .CLK(clk), .RST(rst), .Q(xreg[33]) );
  DFF \xreg_reg[34]  ( .D(xin[33]), .CLK(clk), .RST(rst), .Q(xreg[34]) );
  DFF \xreg_reg[35]  ( .D(xin[34]), .CLK(clk), .RST(rst), .Q(xreg[35]) );
  DFF \xreg_reg[36]  ( .D(xin[35]), .CLK(clk), .RST(rst), .Q(xreg[36]) );
  DFF \xreg_reg[37]  ( .D(xin[36]), .CLK(clk), .RST(rst), .Q(xreg[37]) );
  DFF \xreg_reg[38]  ( .D(xin[37]), .CLK(clk), .RST(rst), .Q(xreg[38]) );
  DFF \xreg_reg[39]  ( .D(xin[38]), .CLK(clk), .RST(rst), .Q(xreg[39]) );
  DFF \xreg_reg[40]  ( .D(xin[39]), .CLK(clk), .RST(rst), .Q(xreg[40]) );
  DFF \xreg_reg[41]  ( .D(xin[40]), .CLK(clk), .RST(rst), .Q(xreg[41]) );
  DFF \xreg_reg[42]  ( .D(xin[41]), .CLK(clk), .RST(rst), .Q(xreg[42]) );
  DFF \xreg_reg[43]  ( .D(xin[42]), .CLK(clk), .RST(rst), .Q(xreg[43]) );
  DFF \xreg_reg[44]  ( .D(xin[43]), .CLK(clk), .RST(rst), .Q(xreg[44]) );
  DFF \xreg_reg[45]  ( .D(xin[44]), .CLK(clk), .RST(rst), .Q(xreg[45]) );
  DFF \xreg_reg[46]  ( .D(xin[45]), .CLK(clk), .RST(rst), .Q(xreg[46]) );
  DFF \xreg_reg[47]  ( .D(xin[46]), .CLK(clk), .RST(rst), .Q(xreg[47]) );
  DFF \xreg_reg[48]  ( .D(xin[47]), .CLK(clk), .RST(rst), .Q(xreg[48]) );
  DFF \xreg_reg[49]  ( .D(xin[48]), .CLK(clk), .RST(rst), .Q(xreg[49]) );
  DFF \xreg_reg[50]  ( .D(xin[49]), .CLK(clk), .RST(rst), .Q(xreg[50]) );
  DFF \xreg_reg[51]  ( .D(xin[50]), .CLK(clk), .RST(rst), .Q(xreg[51]) );
  DFF \xreg_reg[52]  ( .D(xin[51]), .CLK(clk), .RST(rst), .Q(xreg[52]) );
  DFF \xreg_reg[53]  ( .D(xin[52]), .CLK(clk), .RST(rst), .Q(xreg[53]) );
  DFF \xreg_reg[54]  ( .D(xin[53]), .CLK(clk), .RST(rst), .Q(xreg[54]) );
  DFF \xreg_reg[55]  ( .D(xin[54]), .CLK(clk), .RST(rst), .Q(xreg[55]) );
  DFF \xreg_reg[56]  ( .D(xin[55]), .CLK(clk), .RST(rst), .Q(xreg[56]) );
  DFF \xreg_reg[57]  ( .D(xin[56]), .CLK(clk), .RST(rst), .Q(xreg[57]) );
  DFF \xreg_reg[58]  ( .D(xin[57]), .CLK(clk), .RST(rst), .Q(xreg[58]) );
  DFF \xreg_reg[59]  ( .D(xin[58]), .CLK(clk), .RST(rst), .Q(xreg[59]) );
  DFF \xreg_reg[60]  ( .D(xin[59]), .CLK(clk), .RST(rst), .Q(xreg[60]) );
  DFF \xreg_reg[61]  ( .D(xin[60]), .CLK(clk), .RST(rst), .Q(xreg[61]) );
  DFF \xreg_reg[62]  ( .D(xin[61]), .CLK(clk), .RST(rst), .Q(xreg[62]) );
  DFF \xreg_reg[63]  ( .D(xin[62]), .CLK(clk), .RST(rst), .Q(xreg[63]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(zreg[0]) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(zreg[1]) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(zreg[2]) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(zreg[3]) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(zreg[4]) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(zreg[5]) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(zreg[6]) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(zreg[7]) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(zreg[8]) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(zreg[9]) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(zreg[10]) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(zreg[11]) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(zreg[12]) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(zreg[13]) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .Q(zreg[14]) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .Q(zreg[15]) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .Q(zreg[16]) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .Q(zreg[17]) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .Q(zreg[18]) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .Q(zreg[19]) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .Q(zreg[20]) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .Q(zreg[21]) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .Q(zreg[22]) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .Q(zreg[23]) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .Q(zreg[24]) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .Q(zreg[25]) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .Q(zreg[26]) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .Q(zreg[27]) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .Q(zreg[28]) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .Q(zreg[29]) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .Q(zreg[30]) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .Q(zreg[31]) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .Q(zreg[32]) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .Q(zreg[33]) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .Q(zreg[34]) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .Q(zreg[35]) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .Q(zreg[36]) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .Q(zreg[37]) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .Q(zreg[38]) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .Q(zreg[39]) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .Q(zreg[40]) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .Q(zreg[41]) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .Q(zreg[42]) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .Q(zreg[43]) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .Q(zreg[44]) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .Q(zreg[45]) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .Q(zreg[46]) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .Q(zreg[47]) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .Q(zreg[48]) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .Q(zreg[49]) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .Q(zreg[50]) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .Q(zreg[51]) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .Q(zreg[52]) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .Q(zreg[53]) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .Q(zreg[54]) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .Q(zreg[55]) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .Q(zreg[56]) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .Q(zreg[57]) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .Q(zreg[58]) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .Q(zreg[59]) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .Q(zreg[60]) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .Q(zreg[61]) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .Q(zreg[62]) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .Q(zreg[63]) );
  DFF \zreg_reg[64]  ( .D(\zout[0][64] ), .CLK(clk), .RST(rst), .Q(zreg[64])
         );
  DFF \zreg_reg[65]  ( .D(\zout[0][65] ), .CLK(clk), .RST(rst), .Q(zreg[65])
         );
  modmult_step_N64 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[63]), .y(y), 
        .n(n), .zin({\zin[0][65] , \zin[0][64] , \zin[0][63] , \zin[0][62] , 
        \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] , \zin[0][57] , 
        \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] , \zin[0][52] , 
        \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] , \zin[0][47] , 
        \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] , \zin[0][42] , 
        \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] , \zin[0][37] , 
        \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] , \zin[0][32] , 
        \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] , \zin[0][27] , 
        \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] , \zin[0][22] , 
        \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] , \zin[0][17] , 
        \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] , \zin[0][12] , 
        \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] , \zin[0][7] , 
        \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] , \zin[0][2] , 
        \zin[0][1] , \zin[0][0] }), .zout({\zout[0][65] , \zout[0][64] , o})
         );
  ANDN U3 ( .B(zreg[9]), .A(start), .Z(\zin[0][9] ) );
  ANDN U4 ( .B(zreg[8]), .A(start), .Z(\zin[0][8] ) );
  ANDN U5 ( .B(zreg[7]), .A(start), .Z(\zin[0][7] ) );
  ANDN U6 ( .B(zreg[6]), .A(start), .Z(\zin[0][6] ) );
  ANDN U7 ( .B(zreg[65]), .A(start), .Z(\zin[0][65] ) );
  ANDN U8 ( .B(zreg[64]), .A(start), .Z(\zin[0][64] ) );
  ANDN U9 ( .B(zreg[63]), .A(start), .Z(\zin[0][63] ) );
  ANDN U10 ( .B(zreg[62]), .A(start), .Z(\zin[0][62] ) );
  ANDN U11 ( .B(zreg[61]), .A(start), .Z(\zin[0][61] ) );
  ANDN U12 ( .B(zreg[60]), .A(start), .Z(\zin[0][60] ) );
  ANDN U13 ( .B(zreg[5]), .A(start), .Z(\zin[0][5] ) );
  ANDN U14 ( .B(zreg[59]), .A(start), .Z(\zin[0][59] ) );
  ANDN U15 ( .B(zreg[58]), .A(start), .Z(\zin[0][58] ) );
  ANDN U16 ( .B(zreg[57]), .A(start), .Z(\zin[0][57] ) );
  ANDN U17 ( .B(zreg[56]), .A(start), .Z(\zin[0][56] ) );
  ANDN U18 ( .B(zreg[55]), .A(start), .Z(\zin[0][55] ) );
  ANDN U19 ( .B(zreg[54]), .A(start), .Z(\zin[0][54] ) );
  ANDN U20 ( .B(zreg[53]), .A(start), .Z(\zin[0][53] ) );
  ANDN U21 ( .B(zreg[52]), .A(start), .Z(\zin[0][52] ) );
  ANDN U22 ( .B(zreg[51]), .A(start), .Z(\zin[0][51] ) );
  ANDN U23 ( .B(zreg[50]), .A(start), .Z(\zin[0][50] ) );
  ANDN U24 ( .B(zreg[4]), .A(start), .Z(\zin[0][4] ) );
  ANDN U25 ( .B(zreg[49]), .A(start), .Z(\zin[0][49] ) );
  ANDN U26 ( .B(zreg[48]), .A(start), .Z(\zin[0][48] ) );
  ANDN U27 ( .B(zreg[47]), .A(start), .Z(\zin[0][47] ) );
  ANDN U28 ( .B(zreg[46]), .A(start), .Z(\zin[0][46] ) );
  ANDN U29 ( .B(zreg[45]), .A(start), .Z(\zin[0][45] ) );
  ANDN U30 ( .B(zreg[44]), .A(start), .Z(\zin[0][44] ) );
  ANDN U31 ( .B(zreg[43]), .A(start), .Z(\zin[0][43] ) );
  ANDN U32 ( .B(zreg[42]), .A(start), .Z(\zin[0][42] ) );
  ANDN U33 ( .B(zreg[41]), .A(start), .Z(\zin[0][41] ) );
  ANDN U34 ( .B(zreg[40]), .A(start), .Z(\zin[0][40] ) );
  ANDN U35 ( .B(zreg[3]), .A(start), .Z(\zin[0][3] ) );
  ANDN U36 ( .B(zreg[39]), .A(start), .Z(\zin[0][39] ) );
  ANDN U37 ( .B(zreg[38]), .A(start), .Z(\zin[0][38] ) );
  ANDN U38 ( .B(zreg[37]), .A(start), .Z(\zin[0][37] ) );
  ANDN U39 ( .B(zreg[36]), .A(start), .Z(\zin[0][36] ) );
  ANDN U40 ( .B(zreg[35]), .A(start), .Z(\zin[0][35] ) );
  ANDN U41 ( .B(zreg[34]), .A(start), .Z(\zin[0][34] ) );
  ANDN U42 ( .B(zreg[33]), .A(start), .Z(\zin[0][33] ) );
  ANDN U43 ( .B(zreg[32]), .A(start), .Z(\zin[0][32] ) );
  ANDN U44 ( .B(zreg[31]), .A(start), .Z(\zin[0][31] ) );
  ANDN U45 ( .B(zreg[30]), .A(start), .Z(\zin[0][30] ) );
  ANDN U46 ( .B(zreg[2]), .A(start), .Z(\zin[0][2] ) );
  ANDN U47 ( .B(zreg[29]), .A(start), .Z(\zin[0][29] ) );
  ANDN U48 ( .B(zreg[28]), .A(start), .Z(\zin[0][28] ) );
  ANDN U49 ( .B(zreg[27]), .A(start), .Z(\zin[0][27] ) );
  ANDN U50 ( .B(zreg[26]), .A(start), .Z(\zin[0][26] ) );
  ANDN U51 ( .B(zreg[25]), .A(start), .Z(\zin[0][25] ) );
  ANDN U52 ( .B(zreg[24]), .A(start), .Z(\zin[0][24] ) );
  ANDN U53 ( .B(zreg[23]), .A(start), .Z(\zin[0][23] ) );
  ANDN U54 ( .B(zreg[22]), .A(start), .Z(\zin[0][22] ) );
  ANDN U55 ( .B(zreg[21]), .A(start), .Z(\zin[0][21] ) );
  ANDN U56 ( .B(zreg[20]), .A(start), .Z(\zin[0][20] ) );
  ANDN U57 ( .B(zreg[1]), .A(start), .Z(\zin[0][1] ) );
  ANDN U58 ( .B(zreg[19]), .A(start), .Z(\zin[0][19] ) );
  ANDN U59 ( .B(zreg[18]), .A(start), .Z(\zin[0][18] ) );
  ANDN U60 ( .B(zreg[17]), .A(start), .Z(\zin[0][17] ) );
  ANDN U61 ( .B(zreg[16]), .A(start), .Z(\zin[0][16] ) );
  ANDN U62 ( .B(zreg[15]), .A(start), .Z(\zin[0][15] ) );
  ANDN U63 ( .B(zreg[14]), .A(start), .Z(\zin[0][14] ) );
  ANDN U64 ( .B(zreg[13]), .A(start), .Z(\zin[0][13] ) );
  ANDN U65 ( .B(zreg[12]), .A(start), .Z(\zin[0][12] ) );
  ANDN U66 ( .B(zreg[11]), .A(start), .Z(\zin[0][11] ) );
  ANDN U67 ( .B(zreg[10]), .A(start), .Z(\zin[0][10] ) );
  ANDN U68 ( .B(zreg[0]), .A(start), .Z(\zin[0][0] ) );
  NAND U69 ( .A(n1), .B(n2), .Z(xin[9]) );
  NANDN U70 ( .A(start), .B(xreg[9]), .Z(n2) );
  NAND U71 ( .A(x[9]), .B(start), .Z(n1) );
  NAND U72 ( .A(n3), .B(n4), .Z(xin[8]) );
  NANDN U73 ( .A(start), .B(xreg[8]), .Z(n4) );
  NAND U74 ( .A(x[8]), .B(start), .Z(n3) );
  NAND U75 ( .A(n5), .B(n6), .Z(xin[7]) );
  NANDN U76 ( .A(start), .B(xreg[7]), .Z(n6) );
  NAND U77 ( .A(x[7]), .B(start), .Z(n5) );
  NAND U78 ( .A(n7), .B(n8), .Z(xin[6]) );
  NANDN U79 ( .A(start), .B(xreg[6]), .Z(n8) );
  NAND U80 ( .A(x[6]), .B(start), .Z(n7) );
  NAND U81 ( .A(n9), .B(n10), .Z(xin[63]) );
  NANDN U82 ( .A(start), .B(xreg[63]), .Z(n10) );
  NAND U83 ( .A(x[63]), .B(start), .Z(n9) );
  NAND U84 ( .A(n11), .B(n12), .Z(xin[62]) );
  NANDN U85 ( .A(start), .B(xreg[62]), .Z(n12) );
  NAND U86 ( .A(x[62]), .B(start), .Z(n11) );
  NAND U87 ( .A(n13), .B(n14), .Z(xin[61]) );
  NANDN U88 ( .A(start), .B(xreg[61]), .Z(n14) );
  NAND U89 ( .A(x[61]), .B(start), .Z(n13) );
  NAND U90 ( .A(n15), .B(n16), .Z(xin[60]) );
  NANDN U91 ( .A(start), .B(xreg[60]), .Z(n16) );
  NAND U92 ( .A(x[60]), .B(start), .Z(n15) );
  NAND U93 ( .A(n17), .B(n18), .Z(xin[5]) );
  NANDN U94 ( .A(start), .B(xreg[5]), .Z(n18) );
  NAND U95 ( .A(x[5]), .B(start), .Z(n17) );
  NAND U96 ( .A(n19), .B(n20), .Z(xin[59]) );
  NANDN U97 ( .A(start), .B(xreg[59]), .Z(n20) );
  NAND U98 ( .A(x[59]), .B(start), .Z(n19) );
  NAND U99 ( .A(n21), .B(n22), .Z(xin[58]) );
  NANDN U100 ( .A(start), .B(xreg[58]), .Z(n22) );
  NAND U101 ( .A(x[58]), .B(start), .Z(n21) );
  NAND U102 ( .A(n23), .B(n24), .Z(xin[57]) );
  NANDN U103 ( .A(start), .B(xreg[57]), .Z(n24) );
  NAND U104 ( .A(x[57]), .B(start), .Z(n23) );
  NAND U105 ( .A(n25), .B(n26), .Z(xin[56]) );
  NANDN U106 ( .A(start), .B(xreg[56]), .Z(n26) );
  NAND U107 ( .A(x[56]), .B(start), .Z(n25) );
  NAND U108 ( .A(n27), .B(n28), .Z(xin[55]) );
  NANDN U109 ( .A(start), .B(xreg[55]), .Z(n28) );
  NAND U110 ( .A(x[55]), .B(start), .Z(n27) );
  NAND U111 ( .A(n29), .B(n30), .Z(xin[54]) );
  NANDN U112 ( .A(start), .B(xreg[54]), .Z(n30) );
  NAND U113 ( .A(x[54]), .B(start), .Z(n29) );
  NAND U114 ( .A(n31), .B(n32), .Z(xin[53]) );
  NANDN U115 ( .A(start), .B(xreg[53]), .Z(n32) );
  NAND U116 ( .A(x[53]), .B(start), .Z(n31) );
  NAND U117 ( .A(n33), .B(n34), .Z(xin[52]) );
  NANDN U118 ( .A(start), .B(xreg[52]), .Z(n34) );
  NAND U119 ( .A(x[52]), .B(start), .Z(n33) );
  NAND U120 ( .A(n35), .B(n36), .Z(xin[51]) );
  NANDN U121 ( .A(start), .B(xreg[51]), .Z(n36) );
  NAND U122 ( .A(x[51]), .B(start), .Z(n35) );
  NAND U123 ( .A(n37), .B(n38), .Z(xin[50]) );
  NANDN U124 ( .A(start), .B(xreg[50]), .Z(n38) );
  NAND U125 ( .A(x[50]), .B(start), .Z(n37) );
  NAND U126 ( .A(n39), .B(n40), .Z(xin[4]) );
  NANDN U127 ( .A(start), .B(xreg[4]), .Z(n40) );
  NAND U128 ( .A(x[4]), .B(start), .Z(n39) );
  NAND U129 ( .A(n41), .B(n42), .Z(xin[49]) );
  NANDN U130 ( .A(start), .B(xreg[49]), .Z(n42) );
  NAND U131 ( .A(x[49]), .B(start), .Z(n41) );
  NAND U132 ( .A(n43), .B(n44), .Z(xin[48]) );
  NANDN U133 ( .A(start), .B(xreg[48]), .Z(n44) );
  NAND U134 ( .A(x[48]), .B(start), .Z(n43) );
  NAND U135 ( .A(n45), .B(n46), .Z(xin[47]) );
  NANDN U136 ( .A(start), .B(xreg[47]), .Z(n46) );
  NAND U137 ( .A(x[47]), .B(start), .Z(n45) );
  NAND U138 ( .A(n47), .B(n48), .Z(xin[46]) );
  NANDN U139 ( .A(start), .B(xreg[46]), .Z(n48) );
  NAND U140 ( .A(x[46]), .B(start), .Z(n47) );
  NAND U141 ( .A(n49), .B(n50), .Z(xin[45]) );
  NANDN U142 ( .A(start), .B(xreg[45]), .Z(n50) );
  NAND U143 ( .A(x[45]), .B(start), .Z(n49) );
  NAND U144 ( .A(n51), .B(n52), .Z(xin[44]) );
  NANDN U145 ( .A(start), .B(xreg[44]), .Z(n52) );
  NAND U146 ( .A(x[44]), .B(start), .Z(n51) );
  NAND U147 ( .A(n53), .B(n54), .Z(xin[43]) );
  NANDN U148 ( .A(start), .B(xreg[43]), .Z(n54) );
  NAND U149 ( .A(x[43]), .B(start), .Z(n53) );
  NAND U150 ( .A(n55), .B(n56), .Z(xin[42]) );
  NANDN U151 ( .A(start), .B(xreg[42]), .Z(n56) );
  NAND U152 ( .A(x[42]), .B(start), .Z(n55) );
  NAND U153 ( .A(n57), .B(n58), .Z(xin[41]) );
  NANDN U154 ( .A(start), .B(xreg[41]), .Z(n58) );
  NAND U155 ( .A(x[41]), .B(start), .Z(n57) );
  NAND U156 ( .A(n59), .B(n60), .Z(xin[40]) );
  NANDN U157 ( .A(start), .B(xreg[40]), .Z(n60) );
  NAND U158 ( .A(x[40]), .B(start), .Z(n59) );
  NAND U159 ( .A(n61), .B(n62), .Z(xin[3]) );
  NANDN U160 ( .A(start), .B(xreg[3]), .Z(n62) );
  NAND U161 ( .A(x[3]), .B(start), .Z(n61) );
  NAND U162 ( .A(n63), .B(n64), .Z(xin[39]) );
  NANDN U163 ( .A(start), .B(xreg[39]), .Z(n64) );
  NAND U164 ( .A(x[39]), .B(start), .Z(n63) );
  NAND U165 ( .A(n65), .B(n66), .Z(xin[38]) );
  NANDN U166 ( .A(start), .B(xreg[38]), .Z(n66) );
  NAND U167 ( .A(x[38]), .B(start), .Z(n65) );
  NAND U168 ( .A(n67), .B(n68), .Z(xin[37]) );
  NANDN U169 ( .A(start), .B(xreg[37]), .Z(n68) );
  NAND U170 ( .A(x[37]), .B(start), .Z(n67) );
  NAND U171 ( .A(n69), .B(n70), .Z(xin[36]) );
  NANDN U172 ( .A(start), .B(xreg[36]), .Z(n70) );
  NAND U173 ( .A(x[36]), .B(start), .Z(n69) );
  NAND U174 ( .A(n71), .B(n72), .Z(xin[35]) );
  NANDN U175 ( .A(start), .B(xreg[35]), .Z(n72) );
  NAND U176 ( .A(x[35]), .B(start), .Z(n71) );
  NAND U177 ( .A(n73), .B(n74), .Z(xin[34]) );
  NANDN U178 ( .A(start), .B(xreg[34]), .Z(n74) );
  NAND U179 ( .A(x[34]), .B(start), .Z(n73) );
  NAND U180 ( .A(n75), .B(n76), .Z(xin[33]) );
  NANDN U181 ( .A(start), .B(xreg[33]), .Z(n76) );
  NAND U182 ( .A(x[33]), .B(start), .Z(n75) );
  NAND U183 ( .A(n77), .B(n78), .Z(xin[32]) );
  NANDN U184 ( .A(start), .B(xreg[32]), .Z(n78) );
  NAND U185 ( .A(x[32]), .B(start), .Z(n77) );
  NAND U186 ( .A(n79), .B(n80), .Z(xin[31]) );
  NANDN U187 ( .A(start), .B(xreg[31]), .Z(n80) );
  NAND U188 ( .A(x[31]), .B(start), .Z(n79) );
  NAND U189 ( .A(n81), .B(n82), .Z(xin[30]) );
  NANDN U190 ( .A(start), .B(xreg[30]), .Z(n82) );
  NAND U191 ( .A(x[30]), .B(start), .Z(n81) );
  NAND U192 ( .A(n83), .B(n84), .Z(xin[2]) );
  NANDN U193 ( .A(start), .B(xreg[2]), .Z(n84) );
  NAND U194 ( .A(x[2]), .B(start), .Z(n83) );
  NAND U195 ( .A(n85), .B(n86), .Z(xin[29]) );
  NANDN U196 ( .A(start), .B(xreg[29]), .Z(n86) );
  NAND U197 ( .A(x[29]), .B(start), .Z(n85) );
  NAND U198 ( .A(n87), .B(n88), .Z(xin[28]) );
  NANDN U199 ( .A(start), .B(xreg[28]), .Z(n88) );
  NAND U200 ( .A(x[28]), .B(start), .Z(n87) );
  NAND U201 ( .A(n89), .B(n90), .Z(xin[27]) );
  NANDN U202 ( .A(start), .B(xreg[27]), .Z(n90) );
  NAND U203 ( .A(x[27]), .B(start), .Z(n89) );
  NAND U204 ( .A(n91), .B(n92), .Z(xin[26]) );
  NANDN U205 ( .A(start), .B(xreg[26]), .Z(n92) );
  NAND U206 ( .A(x[26]), .B(start), .Z(n91) );
  NAND U207 ( .A(n93), .B(n94), .Z(xin[25]) );
  NANDN U208 ( .A(start), .B(xreg[25]), .Z(n94) );
  NAND U209 ( .A(x[25]), .B(start), .Z(n93) );
  NAND U210 ( .A(n95), .B(n96), .Z(xin[24]) );
  NANDN U211 ( .A(start), .B(xreg[24]), .Z(n96) );
  NAND U212 ( .A(x[24]), .B(start), .Z(n95) );
  NAND U213 ( .A(n97), .B(n98), .Z(xin[23]) );
  NANDN U214 ( .A(start), .B(xreg[23]), .Z(n98) );
  NAND U215 ( .A(x[23]), .B(start), .Z(n97) );
  NAND U216 ( .A(n99), .B(n100), .Z(xin[22]) );
  NANDN U217 ( .A(start), .B(xreg[22]), .Z(n100) );
  NAND U218 ( .A(x[22]), .B(start), .Z(n99) );
  NAND U219 ( .A(n101), .B(n102), .Z(xin[21]) );
  NANDN U220 ( .A(start), .B(xreg[21]), .Z(n102) );
  NAND U221 ( .A(x[21]), .B(start), .Z(n101) );
  NAND U222 ( .A(n103), .B(n104), .Z(xin[20]) );
  NANDN U223 ( .A(start), .B(xreg[20]), .Z(n104) );
  NAND U224 ( .A(x[20]), .B(start), .Z(n103) );
  NAND U225 ( .A(n105), .B(n106), .Z(xin[1]) );
  NANDN U226 ( .A(start), .B(xreg[1]), .Z(n106) );
  NAND U227 ( .A(x[1]), .B(start), .Z(n105) );
  NAND U228 ( .A(n107), .B(n108), .Z(xin[19]) );
  NANDN U229 ( .A(start), .B(xreg[19]), .Z(n108) );
  NAND U230 ( .A(x[19]), .B(start), .Z(n107) );
  NAND U231 ( .A(n109), .B(n110), .Z(xin[18]) );
  NANDN U232 ( .A(start), .B(xreg[18]), .Z(n110) );
  NAND U233 ( .A(x[18]), .B(start), .Z(n109) );
  NAND U234 ( .A(n111), .B(n112), .Z(xin[17]) );
  NANDN U235 ( .A(start), .B(xreg[17]), .Z(n112) );
  NAND U236 ( .A(x[17]), .B(start), .Z(n111) );
  NAND U237 ( .A(n113), .B(n114), .Z(xin[16]) );
  NANDN U238 ( .A(start), .B(xreg[16]), .Z(n114) );
  NAND U239 ( .A(x[16]), .B(start), .Z(n113) );
  NAND U240 ( .A(n115), .B(n116), .Z(xin[15]) );
  NANDN U241 ( .A(start), .B(xreg[15]), .Z(n116) );
  NAND U242 ( .A(x[15]), .B(start), .Z(n115) );
  NAND U243 ( .A(n117), .B(n118), .Z(xin[14]) );
  NANDN U244 ( .A(start), .B(xreg[14]), .Z(n118) );
  NAND U245 ( .A(x[14]), .B(start), .Z(n117) );
  NAND U246 ( .A(n119), .B(n120), .Z(xin[13]) );
  NANDN U247 ( .A(start), .B(xreg[13]), .Z(n120) );
  NAND U248 ( .A(x[13]), .B(start), .Z(n119) );
  NAND U249 ( .A(n121), .B(n122), .Z(xin[12]) );
  NANDN U250 ( .A(start), .B(xreg[12]), .Z(n122) );
  NAND U251 ( .A(x[12]), .B(start), .Z(n121) );
  NAND U252 ( .A(n123), .B(n124), .Z(xin[11]) );
  NANDN U253 ( .A(start), .B(xreg[11]), .Z(n124) );
  NAND U254 ( .A(x[11]), .B(start), .Z(n123) );
  NAND U255 ( .A(n125), .B(n126), .Z(xin[10]) );
  NANDN U256 ( .A(start), .B(xreg[10]), .Z(n126) );
  NAND U257 ( .A(x[10]), .B(start), .Z(n125) );
  AND U258 ( .A(x[0]), .B(start), .Z(n127) );
endmodule


module modexp_2N_NN_N64_CC8192 ( clk, rst, m, e, n, c );
  input [63:0] m;
  input [63:0] e;
  input [63:0] n;
  output [63:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825;
  wire   [63:0] start_in;
  wire   [63:0] start_reg;
  wire   [63:0] ereg;
  wire   [63:0] o;
  wire   [63:0] creg;
  wire   [63:0] x;
  wire   [63:0] y;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(n1825), .CLK(clk), .RST(rst), .Q(start_reg[0])
         );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF mul_pow_reg ( .D(n977), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n976), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n975), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n974), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n973), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n972), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n971), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n970), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n969), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n968), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n967), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n966), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n965), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n964), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n963), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n962), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n961), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n960), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n959), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n958), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n957), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n956), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n955), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n954), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n953), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n952), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n951), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n950), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n949), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n948), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n947), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n946), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n945), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n944), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n943), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n942), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n941), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n940), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n939), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n938), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n937), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n936), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n935), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n934), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n933), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n932), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n931), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n930), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n929), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n928), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n927), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n926), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n925), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n924), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n923), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n922), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n921), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n920), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n919), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n918), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n917), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n916), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n915), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n914), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n913), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF first_one_reg ( .D(n848), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n911), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n910), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n909), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n908), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n907), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n906), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n905), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n904), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n903), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n902), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n901), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n900), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n899), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n898), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n897), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n896), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n895), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n894), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n893), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n892), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n891), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n890), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n889), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n888), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n887), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n886), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n885), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n884), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n883), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n882), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n881), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n880), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n879), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n878), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n877), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n876), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n875), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n874), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n873), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n872), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n871), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n870), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n869), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n868), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n867), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n866), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n865), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n864), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n863), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n862), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n861), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n860), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n859), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n858), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n857), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n856), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n855), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n854), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n853), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n852), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n851), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n850), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n849), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n912), .CLK(clk), .RST(rst), .Q(creg[63]) );
  modmult_N64_CC64 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), .x(x), .y(y), .n(n), .o(o) );
  NAND U1236 ( .A(n978), .B(n979), .Z(y[9]) );
  NAND U1237 ( .A(n980), .B(m[9]), .Z(n979) );
  NAND U1238 ( .A(n981), .B(creg[9]), .Z(n978) );
  NAND U1239 ( .A(n982), .B(n983), .Z(y[8]) );
  NAND U1240 ( .A(n980), .B(m[8]), .Z(n983) );
  NAND U1241 ( .A(n981), .B(creg[8]), .Z(n982) );
  NAND U1242 ( .A(n984), .B(n985), .Z(y[7]) );
  NAND U1243 ( .A(n980), .B(m[7]), .Z(n985) );
  NAND U1244 ( .A(n981), .B(creg[7]), .Z(n984) );
  NAND U1245 ( .A(n986), .B(n987), .Z(y[6]) );
  NAND U1246 ( .A(n980), .B(m[6]), .Z(n987) );
  NAND U1247 ( .A(n981), .B(creg[6]), .Z(n986) );
  NAND U1248 ( .A(n988), .B(n989), .Z(y[63]) );
  NAND U1249 ( .A(n980), .B(m[63]), .Z(n989) );
  NAND U1250 ( .A(n981), .B(creg[63]), .Z(n988) );
  NAND U1251 ( .A(n990), .B(n991), .Z(y[62]) );
  NAND U1252 ( .A(n980), .B(m[62]), .Z(n991) );
  NAND U1253 ( .A(n981), .B(creg[62]), .Z(n990) );
  NAND U1254 ( .A(n992), .B(n993), .Z(y[61]) );
  NAND U1255 ( .A(n980), .B(m[61]), .Z(n993) );
  NAND U1256 ( .A(n981), .B(creg[61]), .Z(n992) );
  NAND U1257 ( .A(n994), .B(n995), .Z(y[60]) );
  NAND U1258 ( .A(n980), .B(m[60]), .Z(n995) );
  NAND U1259 ( .A(n981), .B(creg[60]), .Z(n994) );
  NAND U1260 ( .A(n996), .B(n997), .Z(y[5]) );
  NAND U1261 ( .A(n980), .B(m[5]), .Z(n997) );
  NAND U1262 ( .A(n981), .B(creg[5]), .Z(n996) );
  NAND U1263 ( .A(n998), .B(n999), .Z(y[59]) );
  NAND U1264 ( .A(n980), .B(m[59]), .Z(n999) );
  NAND U1265 ( .A(n981), .B(creg[59]), .Z(n998) );
  NAND U1266 ( .A(n1000), .B(n1001), .Z(y[58]) );
  NAND U1267 ( .A(n980), .B(m[58]), .Z(n1001) );
  NAND U1268 ( .A(n981), .B(creg[58]), .Z(n1000) );
  NAND U1269 ( .A(n1002), .B(n1003), .Z(y[57]) );
  NAND U1270 ( .A(n980), .B(m[57]), .Z(n1003) );
  NAND U1271 ( .A(n981), .B(creg[57]), .Z(n1002) );
  NAND U1272 ( .A(n1004), .B(n1005), .Z(y[56]) );
  NAND U1273 ( .A(n980), .B(m[56]), .Z(n1005) );
  NAND U1274 ( .A(n981), .B(creg[56]), .Z(n1004) );
  NAND U1275 ( .A(n1006), .B(n1007), .Z(y[55]) );
  NAND U1276 ( .A(n980), .B(m[55]), .Z(n1007) );
  NAND U1277 ( .A(n981), .B(creg[55]), .Z(n1006) );
  NAND U1278 ( .A(n1008), .B(n1009), .Z(y[54]) );
  NAND U1279 ( .A(n980), .B(m[54]), .Z(n1009) );
  NAND U1280 ( .A(n981), .B(creg[54]), .Z(n1008) );
  NAND U1281 ( .A(n1010), .B(n1011), .Z(y[53]) );
  NAND U1282 ( .A(n980), .B(m[53]), .Z(n1011) );
  NAND U1283 ( .A(n981), .B(creg[53]), .Z(n1010) );
  NAND U1284 ( .A(n1012), .B(n1013), .Z(y[52]) );
  NAND U1285 ( .A(n980), .B(m[52]), .Z(n1013) );
  NAND U1286 ( .A(n981), .B(creg[52]), .Z(n1012) );
  NAND U1287 ( .A(n1014), .B(n1015), .Z(y[51]) );
  NAND U1288 ( .A(n980), .B(m[51]), .Z(n1015) );
  NAND U1289 ( .A(n981), .B(creg[51]), .Z(n1014) );
  NAND U1290 ( .A(n1016), .B(n1017), .Z(y[50]) );
  NAND U1291 ( .A(n980), .B(m[50]), .Z(n1017) );
  NAND U1292 ( .A(n981), .B(creg[50]), .Z(n1016) );
  NAND U1293 ( .A(n1018), .B(n1019), .Z(y[4]) );
  NAND U1294 ( .A(n980), .B(m[4]), .Z(n1019) );
  NAND U1295 ( .A(n981), .B(creg[4]), .Z(n1018) );
  NAND U1296 ( .A(n1020), .B(n1021), .Z(y[49]) );
  NAND U1297 ( .A(n980), .B(m[49]), .Z(n1021) );
  NAND U1298 ( .A(n981), .B(creg[49]), .Z(n1020) );
  NAND U1299 ( .A(n1022), .B(n1023), .Z(y[48]) );
  NAND U1300 ( .A(n980), .B(m[48]), .Z(n1023) );
  NAND U1301 ( .A(n981), .B(creg[48]), .Z(n1022) );
  NAND U1302 ( .A(n1024), .B(n1025), .Z(y[47]) );
  NAND U1303 ( .A(n980), .B(m[47]), .Z(n1025) );
  NAND U1304 ( .A(n981), .B(creg[47]), .Z(n1024) );
  NAND U1305 ( .A(n1026), .B(n1027), .Z(y[46]) );
  NAND U1306 ( .A(n980), .B(m[46]), .Z(n1027) );
  NAND U1307 ( .A(n981), .B(creg[46]), .Z(n1026) );
  NAND U1308 ( .A(n1028), .B(n1029), .Z(y[45]) );
  NAND U1309 ( .A(n980), .B(m[45]), .Z(n1029) );
  NAND U1310 ( .A(n981), .B(creg[45]), .Z(n1028) );
  NAND U1311 ( .A(n1030), .B(n1031), .Z(y[44]) );
  NAND U1312 ( .A(n980), .B(m[44]), .Z(n1031) );
  NAND U1313 ( .A(n981), .B(creg[44]), .Z(n1030) );
  NAND U1314 ( .A(n1032), .B(n1033), .Z(y[43]) );
  NAND U1315 ( .A(n980), .B(m[43]), .Z(n1033) );
  NAND U1316 ( .A(n981), .B(creg[43]), .Z(n1032) );
  NAND U1317 ( .A(n1034), .B(n1035), .Z(y[42]) );
  NAND U1318 ( .A(n980), .B(m[42]), .Z(n1035) );
  NAND U1319 ( .A(n981), .B(creg[42]), .Z(n1034) );
  NAND U1320 ( .A(n1036), .B(n1037), .Z(y[41]) );
  NAND U1321 ( .A(n980), .B(m[41]), .Z(n1037) );
  NAND U1322 ( .A(n981), .B(creg[41]), .Z(n1036) );
  NAND U1323 ( .A(n1038), .B(n1039), .Z(y[40]) );
  NAND U1324 ( .A(n980), .B(m[40]), .Z(n1039) );
  NAND U1325 ( .A(n981), .B(creg[40]), .Z(n1038) );
  NAND U1326 ( .A(n1040), .B(n1041), .Z(y[3]) );
  NAND U1327 ( .A(n980), .B(m[3]), .Z(n1041) );
  NAND U1328 ( .A(n981), .B(creg[3]), .Z(n1040) );
  NAND U1329 ( .A(n1042), .B(n1043), .Z(y[39]) );
  NAND U1330 ( .A(n980), .B(m[39]), .Z(n1043) );
  NAND U1331 ( .A(n981), .B(creg[39]), .Z(n1042) );
  NAND U1332 ( .A(n1044), .B(n1045), .Z(y[38]) );
  NAND U1333 ( .A(n980), .B(m[38]), .Z(n1045) );
  NAND U1334 ( .A(n981), .B(creg[38]), .Z(n1044) );
  NAND U1335 ( .A(n1046), .B(n1047), .Z(y[37]) );
  NAND U1336 ( .A(n980), .B(m[37]), .Z(n1047) );
  NAND U1337 ( .A(n981), .B(creg[37]), .Z(n1046) );
  NAND U1338 ( .A(n1048), .B(n1049), .Z(y[36]) );
  NAND U1339 ( .A(n980), .B(m[36]), .Z(n1049) );
  NAND U1340 ( .A(n981), .B(creg[36]), .Z(n1048) );
  NAND U1341 ( .A(n1050), .B(n1051), .Z(y[35]) );
  NAND U1342 ( .A(n980), .B(m[35]), .Z(n1051) );
  NAND U1343 ( .A(n981), .B(creg[35]), .Z(n1050) );
  NAND U1344 ( .A(n1052), .B(n1053), .Z(y[34]) );
  NAND U1345 ( .A(n980), .B(m[34]), .Z(n1053) );
  NAND U1346 ( .A(n981), .B(creg[34]), .Z(n1052) );
  NAND U1347 ( .A(n1054), .B(n1055), .Z(y[33]) );
  NAND U1348 ( .A(n980), .B(m[33]), .Z(n1055) );
  NAND U1349 ( .A(n981), .B(creg[33]), .Z(n1054) );
  NAND U1350 ( .A(n1056), .B(n1057), .Z(y[32]) );
  NAND U1351 ( .A(n980), .B(m[32]), .Z(n1057) );
  NAND U1352 ( .A(n981), .B(creg[32]), .Z(n1056) );
  NAND U1353 ( .A(n1058), .B(n1059), .Z(y[31]) );
  NAND U1354 ( .A(n980), .B(m[31]), .Z(n1059) );
  NAND U1355 ( .A(n981), .B(creg[31]), .Z(n1058) );
  NAND U1356 ( .A(n1060), .B(n1061), .Z(y[30]) );
  NAND U1357 ( .A(n980), .B(m[30]), .Z(n1061) );
  NAND U1358 ( .A(n981), .B(creg[30]), .Z(n1060) );
  NAND U1359 ( .A(n1062), .B(n1063), .Z(y[2]) );
  NAND U1360 ( .A(n980), .B(m[2]), .Z(n1063) );
  NAND U1361 ( .A(n981), .B(creg[2]), .Z(n1062) );
  NAND U1362 ( .A(n1064), .B(n1065), .Z(y[29]) );
  NAND U1363 ( .A(n980), .B(m[29]), .Z(n1065) );
  NAND U1364 ( .A(n981), .B(creg[29]), .Z(n1064) );
  NAND U1365 ( .A(n1066), .B(n1067), .Z(y[28]) );
  NAND U1366 ( .A(n980), .B(m[28]), .Z(n1067) );
  NAND U1367 ( .A(n981), .B(creg[28]), .Z(n1066) );
  NAND U1368 ( .A(n1068), .B(n1069), .Z(y[27]) );
  NAND U1369 ( .A(n980), .B(m[27]), .Z(n1069) );
  NAND U1370 ( .A(n981), .B(creg[27]), .Z(n1068) );
  NAND U1371 ( .A(n1070), .B(n1071), .Z(y[26]) );
  NAND U1372 ( .A(n980), .B(m[26]), .Z(n1071) );
  NAND U1373 ( .A(n981), .B(creg[26]), .Z(n1070) );
  NAND U1374 ( .A(n1072), .B(n1073), .Z(y[25]) );
  NAND U1375 ( .A(n980), .B(m[25]), .Z(n1073) );
  NAND U1376 ( .A(n981), .B(creg[25]), .Z(n1072) );
  NAND U1377 ( .A(n1074), .B(n1075), .Z(y[24]) );
  NAND U1378 ( .A(n980), .B(m[24]), .Z(n1075) );
  NAND U1379 ( .A(n981), .B(creg[24]), .Z(n1074) );
  NAND U1380 ( .A(n1076), .B(n1077), .Z(y[23]) );
  NAND U1381 ( .A(n980), .B(m[23]), .Z(n1077) );
  NAND U1382 ( .A(n981), .B(creg[23]), .Z(n1076) );
  NAND U1383 ( .A(n1078), .B(n1079), .Z(y[22]) );
  NAND U1384 ( .A(n980), .B(m[22]), .Z(n1079) );
  NAND U1385 ( .A(n981), .B(creg[22]), .Z(n1078) );
  NAND U1386 ( .A(n1080), .B(n1081), .Z(y[21]) );
  NAND U1387 ( .A(n980), .B(m[21]), .Z(n1081) );
  NAND U1388 ( .A(n981), .B(creg[21]), .Z(n1080) );
  NAND U1389 ( .A(n1082), .B(n1083), .Z(y[20]) );
  NAND U1390 ( .A(n980), .B(m[20]), .Z(n1083) );
  NAND U1391 ( .A(n981), .B(creg[20]), .Z(n1082) );
  NAND U1392 ( .A(n1084), .B(n1085), .Z(y[1]) );
  NAND U1393 ( .A(n980), .B(m[1]), .Z(n1085) );
  NAND U1394 ( .A(n981), .B(creg[1]), .Z(n1084) );
  NAND U1395 ( .A(n1086), .B(n1087), .Z(y[19]) );
  NAND U1396 ( .A(n980), .B(m[19]), .Z(n1087) );
  NAND U1397 ( .A(n981), .B(creg[19]), .Z(n1086) );
  NAND U1398 ( .A(n1088), .B(n1089), .Z(y[18]) );
  NAND U1399 ( .A(n980), .B(m[18]), .Z(n1089) );
  NAND U1400 ( .A(n981), .B(creg[18]), .Z(n1088) );
  NAND U1401 ( .A(n1090), .B(n1091), .Z(y[17]) );
  NAND U1402 ( .A(n980), .B(m[17]), .Z(n1091) );
  NAND U1403 ( .A(n981), .B(creg[17]), .Z(n1090) );
  NAND U1404 ( .A(n1092), .B(n1093), .Z(y[16]) );
  NAND U1405 ( .A(n980), .B(m[16]), .Z(n1093) );
  NAND U1406 ( .A(n981), .B(creg[16]), .Z(n1092) );
  NAND U1407 ( .A(n1094), .B(n1095), .Z(y[15]) );
  NAND U1408 ( .A(n980), .B(m[15]), .Z(n1095) );
  NAND U1409 ( .A(n981), .B(creg[15]), .Z(n1094) );
  NAND U1410 ( .A(n1096), .B(n1097), .Z(y[14]) );
  NAND U1411 ( .A(n980), .B(m[14]), .Z(n1097) );
  NAND U1412 ( .A(n981), .B(creg[14]), .Z(n1096) );
  NAND U1413 ( .A(n1098), .B(n1099), .Z(y[13]) );
  NAND U1414 ( .A(n980), .B(m[13]), .Z(n1099) );
  NAND U1415 ( .A(n981), .B(creg[13]), .Z(n1098) );
  NAND U1416 ( .A(n1100), .B(n1101), .Z(y[12]) );
  NAND U1417 ( .A(n980), .B(m[12]), .Z(n1101) );
  NAND U1418 ( .A(n981), .B(creg[12]), .Z(n1100) );
  NAND U1419 ( .A(n1102), .B(n1103), .Z(y[11]) );
  NAND U1420 ( .A(n980), .B(m[11]), .Z(n1103) );
  NAND U1421 ( .A(n981), .B(creg[11]), .Z(n1102) );
  NAND U1422 ( .A(n1104), .B(n1105), .Z(y[10]) );
  NAND U1423 ( .A(n980), .B(m[10]), .Z(n1105) );
  NAND U1424 ( .A(n981), .B(creg[10]), .Z(n1104) );
  NAND U1425 ( .A(n1106), .B(n1107), .Z(y[0]) );
  NAND U1426 ( .A(n980), .B(m[0]), .Z(n1107) );
  NAND U1427 ( .A(n981), .B(creg[0]), .Z(n1106) );
  IV U1428 ( .A(n980), .Z(n981) );
  NAND U1429 ( .A(n1108), .B(n1109), .Z(x[9]) );
  NAND U1430 ( .A(creg[9]), .B(init), .Z(n1108) );
  NAND U1431 ( .A(n1110), .B(n1111), .Z(x[8]) );
  NAND U1432 ( .A(creg[8]), .B(init), .Z(n1110) );
  NAND U1433 ( .A(n1112), .B(n1113), .Z(x[7]) );
  NAND U1434 ( .A(creg[7]), .B(init), .Z(n1112) );
  NAND U1435 ( .A(n1114), .B(n1115), .Z(x[6]) );
  NAND U1436 ( .A(creg[6]), .B(init), .Z(n1114) );
  NAND U1437 ( .A(n1116), .B(n1117), .Z(x[63]) );
  NAND U1438 ( .A(creg[63]), .B(init), .Z(n1116) );
  NAND U1439 ( .A(n1118), .B(n1119), .Z(x[62]) );
  NAND U1440 ( .A(creg[62]), .B(init), .Z(n1118) );
  NAND U1441 ( .A(n1120), .B(n1121), .Z(x[61]) );
  NAND U1442 ( .A(creg[61]), .B(init), .Z(n1120) );
  NAND U1443 ( .A(n1122), .B(n1123), .Z(x[60]) );
  NAND U1444 ( .A(creg[60]), .B(init), .Z(n1122) );
  NAND U1445 ( .A(n1124), .B(n1125), .Z(x[5]) );
  NAND U1446 ( .A(creg[5]), .B(init), .Z(n1124) );
  NAND U1447 ( .A(n1126), .B(n1127), .Z(x[59]) );
  NAND U1448 ( .A(creg[59]), .B(init), .Z(n1126) );
  NAND U1449 ( .A(n1128), .B(n1129), .Z(x[58]) );
  NAND U1450 ( .A(creg[58]), .B(init), .Z(n1128) );
  NAND U1451 ( .A(n1130), .B(n1131), .Z(x[57]) );
  NAND U1452 ( .A(creg[57]), .B(init), .Z(n1130) );
  NAND U1453 ( .A(n1132), .B(n1133), .Z(x[56]) );
  NAND U1454 ( .A(creg[56]), .B(init), .Z(n1132) );
  NAND U1455 ( .A(n1134), .B(n1135), .Z(x[55]) );
  NAND U1456 ( .A(creg[55]), .B(init), .Z(n1134) );
  NAND U1457 ( .A(n1136), .B(n1137), .Z(x[54]) );
  NAND U1458 ( .A(creg[54]), .B(init), .Z(n1136) );
  NAND U1459 ( .A(n1138), .B(n1139), .Z(x[53]) );
  NAND U1460 ( .A(creg[53]), .B(init), .Z(n1138) );
  NAND U1461 ( .A(n1140), .B(n1141), .Z(x[52]) );
  NAND U1462 ( .A(creg[52]), .B(init), .Z(n1140) );
  NAND U1463 ( .A(n1142), .B(n1143), .Z(x[51]) );
  NAND U1464 ( .A(creg[51]), .B(init), .Z(n1142) );
  NAND U1465 ( .A(n1144), .B(n1145), .Z(x[50]) );
  NAND U1466 ( .A(creg[50]), .B(init), .Z(n1144) );
  NAND U1467 ( .A(n1146), .B(n1147), .Z(x[4]) );
  NAND U1468 ( .A(creg[4]), .B(init), .Z(n1146) );
  NAND U1469 ( .A(n1148), .B(n1149), .Z(x[49]) );
  NAND U1470 ( .A(creg[49]), .B(init), .Z(n1148) );
  NAND U1471 ( .A(n1150), .B(n1151), .Z(x[48]) );
  NAND U1472 ( .A(creg[48]), .B(init), .Z(n1150) );
  NAND U1473 ( .A(n1152), .B(n1153), .Z(x[47]) );
  NAND U1474 ( .A(creg[47]), .B(init), .Z(n1152) );
  NAND U1475 ( .A(n1154), .B(n1155), .Z(x[46]) );
  NAND U1476 ( .A(creg[46]), .B(init), .Z(n1154) );
  NAND U1477 ( .A(n1156), .B(n1157), .Z(x[45]) );
  NAND U1478 ( .A(creg[45]), .B(init), .Z(n1156) );
  NAND U1479 ( .A(n1158), .B(n1159), .Z(x[44]) );
  NAND U1480 ( .A(creg[44]), .B(init), .Z(n1158) );
  NAND U1481 ( .A(n1160), .B(n1161), .Z(x[43]) );
  NAND U1482 ( .A(creg[43]), .B(init), .Z(n1160) );
  NAND U1483 ( .A(n1162), .B(n1163), .Z(x[42]) );
  NAND U1484 ( .A(creg[42]), .B(init), .Z(n1162) );
  NAND U1485 ( .A(n1164), .B(n1165), .Z(x[41]) );
  NAND U1486 ( .A(creg[41]), .B(init), .Z(n1164) );
  NAND U1487 ( .A(n1166), .B(n1167), .Z(x[40]) );
  NAND U1488 ( .A(creg[40]), .B(init), .Z(n1166) );
  NAND U1489 ( .A(n1168), .B(n1169), .Z(x[3]) );
  NAND U1490 ( .A(creg[3]), .B(init), .Z(n1168) );
  NAND U1491 ( .A(n1170), .B(n1171), .Z(x[39]) );
  NAND U1492 ( .A(creg[39]), .B(init), .Z(n1170) );
  NAND U1493 ( .A(n1172), .B(n1173), .Z(x[38]) );
  NAND U1494 ( .A(creg[38]), .B(init), .Z(n1172) );
  NAND U1495 ( .A(n1174), .B(n1175), .Z(x[37]) );
  NAND U1496 ( .A(creg[37]), .B(init), .Z(n1174) );
  NAND U1497 ( .A(n1176), .B(n1177), .Z(x[36]) );
  NAND U1498 ( .A(creg[36]), .B(init), .Z(n1176) );
  NAND U1499 ( .A(n1178), .B(n1179), .Z(x[35]) );
  NAND U1500 ( .A(creg[35]), .B(init), .Z(n1178) );
  NAND U1501 ( .A(n1180), .B(n1181), .Z(x[34]) );
  NAND U1502 ( .A(creg[34]), .B(init), .Z(n1180) );
  NAND U1503 ( .A(n1182), .B(n1183), .Z(x[33]) );
  NAND U1504 ( .A(creg[33]), .B(init), .Z(n1182) );
  NAND U1505 ( .A(n1184), .B(n1185), .Z(x[32]) );
  NAND U1506 ( .A(creg[32]), .B(init), .Z(n1184) );
  NAND U1507 ( .A(n1186), .B(n1187), .Z(x[31]) );
  NAND U1508 ( .A(creg[31]), .B(init), .Z(n1186) );
  NAND U1509 ( .A(n1188), .B(n1189), .Z(x[30]) );
  NAND U1510 ( .A(creg[30]), .B(init), .Z(n1188) );
  NAND U1511 ( .A(n1190), .B(n1191), .Z(x[2]) );
  NAND U1512 ( .A(creg[2]), .B(init), .Z(n1190) );
  NAND U1513 ( .A(n1192), .B(n1193), .Z(x[29]) );
  NAND U1514 ( .A(creg[29]), .B(init), .Z(n1192) );
  NAND U1515 ( .A(n1194), .B(n1195), .Z(x[28]) );
  NAND U1516 ( .A(creg[28]), .B(init), .Z(n1194) );
  NAND U1517 ( .A(n1196), .B(n1197), .Z(x[27]) );
  NAND U1518 ( .A(creg[27]), .B(init), .Z(n1196) );
  NAND U1519 ( .A(n1198), .B(n1199), .Z(x[26]) );
  NAND U1520 ( .A(creg[26]), .B(init), .Z(n1198) );
  NAND U1521 ( .A(n1200), .B(n1201), .Z(x[25]) );
  NAND U1522 ( .A(creg[25]), .B(init), .Z(n1200) );
  NAND U1523 ( .A(n1202), .B(n1203), .Z(x[24]) );
  NAND U1524 ( .A(creg[24]), .B(init), .Z(n1202) );
  NAND U1525 ( .A(n1204), .B(n1205), .Z(x[23]) );
  NAND U1526 ( .A(creg[23]), .B(init), .Z(n1204) );
  NAND U1527 ( .A(n1206), .B(n1207), .Z(x[22]) );
  NAND U1528 ( .A(creg[22]), .B(init), .Z(n1206) );
  NAND U1529 ( .A(n1208), .B(n1209), .Z(x[21]) );
  NAND U1530 ( .A(creg[21]), .B(init), .Z(n1208) );
  NAND U1531 ( .A(n1210), .B(n1211), .Z(x[20]) );
  NAND U1532 ( .A(creg[20]), .B(init), .Z(n1210) );
  NAND U1533 ( .A(n1212), .B(n1213), .Z(x[1]) );
  NAND U1534 ( .A(creg[1]), .B(init), .Z(n1212) );
  NAND U1535 ( .A(n1214), .B(n1215), .Z(x[19]) );
  NAND U1536 ( .A(creg[19]), .B(init), .Z(n1214) );
  NAND U1537 ( .A(n1216), .B(n1217), .Z(x[18]) );
  NAND U1538 ( .A(creg[18]), .B(init), .Z(n1216) );
  NAND U1539 ( .A(n1218), .B(n1219), .Z(x[17]) );
  NAND U1540 ( .A(creg[17]), .B(init), .Z(n1218) );
  NAND U1541 ( .A(n1220), .B(n1221), .Z(x[16]) );
  NAND U1542 ( .A(creg[16]), .B(init), .Z(n1220) );
  NAND U1543 ( .A(n1222), .B(n1223), .Z(x[15]) );
  NAND U1544 ( .A(creg[15]), .B(init), .Z(n1222) );
  NAND U1545 ( .A(n1224), .B(n1225), .Z(x[14]) );
  NAND U1546 ( .A(creg[14]), .B(init), .Z(n1224) );
  NAND U1547 ( .A(n1226), .B(n1227), .Z(x[13]) );
  NAND U1548 ( .A(creg[13]), .B(init), .Z(n1226) );
  NAND U1549 ( .A(n1228), .B(n1229), .Z(x[12]) );
  NAND U1550 ( .A(creg[12]), .B(init), .Z(n1228) );
  NAND U1551 ( .A(n1230), .B(n1231), .Z(x[11]) );
  NAND U1552 ( .A(creg[11]), .B(init), .Z(n1230) );
  NAND U1553 ( .A(n1232), .B(n1233), .Z(x[10]) );
  NAND U1554 ( .A(creg[10]), .B(init), .Z(n1232) );
  NAND U1555 ( .A(n1234), .B(n1235), .Z(x[0]) );
  NAND U1556 ( .A(creg[0]), .B(init), .Z(n1234) );
  AND U1557 ( .A(start_reg[9]), .B(init), .Z(start_in[9]) );
  AND U1558 ( .A(start_reg[8]), .B(init), .Z(start_in[8]) );
  AND U1559 ( .A(start_reg[7]), .B(init), .Z(start_in[7]) );
  AND U1560 ( .A(start_reg[6]), .B(init), .Z(start_in[6]) );
  AND U1561 ( .A(start_reg[62]), .B(init), .Z(start_in[62]) );
  AND U1562 ( .A(start_reg[61]), .B(init), .Z(start_in[61]) );
  AND U1563 ( .A(start_reg[60]), .B(init), .Z(start_in[60]) );
  AND U1564 ( .A(start_reg[5]), .B(init), .Z(start_in[5]) );
  AND U1565 ( .A(start_reg[59]), .B(init), .Z(start_in[59]) );
  AND U1566 ( .A(start_reg[58]), .B(init), .Z(start_in[58]) );
  AND U1567 ( .A(start_reg[57]), .B(init), .Z(start_in[57]) );
  AND U1568 ( .A(start_reg[56]), .B(init), .Z(start_in[56]) );
  AND U1569 ( .A(start_reg[55]), .B(init), .Z(start_in[55]) );
  AND U1570 ( .A(start_reg[54]), .B(init), .Z(start_in[54]) );
  AND U1571 ( .A(start_reg[53]), .B(init), .Z(start_in[53]) );
  AND U1572 ( .A(start_reg[52]), .B(init), .Z(start_in[52]) );
  AND U1573 ( .A(start_reg[51]), .B(init), .Z(start_in[51]) );
  AND U1574 ( .A(start_reg[50]), .B(init), .Z(start_in[50]) );
  AND U1575 ( .A(start_reg[4]), .B(init), .Z(start_in[4]) );
  AND U1576 ( .A(start_reg[49]), .B(init), .Z(start_in[49]) );
  AND U1577 ( .A(start_reg[48]), .B(init), .Z(start_in[48]) );
  AND U1578 ( .A(start_reg[47]), .B(init), .Z(start_in[47]) );
  AND U1579 ( .A(start_reg[46]), .B(init), .Z(start_in[46]) );
  AND U1580 ( .A(start_reg[45]), .B(init), .Z(start_in[45]) );
  AND U1581 ( .A(start_reg[44]), .B(init), .Z(start_in[44]) );
  AND U1582 ( .A(start_reg[43]), .B(init), .Z(start_in[43]) );
  AND U1583 ( .A(start_reg[42]), .B(init), .Z(start_in[42]) );
  AND U1584 ( .A(start_reg[41]), .B(init), .Z(start_in[41]) );
  AND U1585 ( .A(start_reg[40]), .B(init), .Z(start_in[40]) );
  AND U1586 ( .A(start_reg[3]), .B(init), .Z(start_in[3]) );
  AND U1587 ( .A(start_reg[39]), .B(init), .Z(start_in[39]) );
  AND U1588 ( .A(start_reg[38]), .B(init), .Z(start_in[38]) );
  AND U1589 ( .A(start_reg[37]), .B(init), .Z(start_in[37]) );
  AND U1590 ( .A(start_reg[36]), .B(init), .Z(start_in[36]) );
  AND U1591 ( .A(start_reg[35]), .B(init), .Z(start_in[35]) );
  AND U1592 ( .A(start_reg[34]), .B(init), .Z(start_in[34]) );
  AND U1593 ( .A(start_reg[33]), .B(init), .Z(start_in[33]) );
  AND U1594 ( .A(start_reg[32]), .B(init), .Z(start_in[32]) );
  AND U1595 ( .A(start_reg[31]), .B(init), .Z(start_in[31]) );
  AND U1596 ( .A(start_reg[30]), .B(init), .Z(start_in[30]) );
  AND U1597 ( .A(start_reg[2]), .B(init), .Z(start_in[2]) );
  AND U1598 ( .A(start_reg[29]), .B(init), .Z(start_in[29]) );
  AND U1599 ( .A(start_reg[28]), .B(init), .Z(start_in[28]) );
  AND U1600 ( .A(start_reg[27]), .B(init), .Z(start_in[27]) );
  AND U1601 ( .A(start_reg[26]), .B(init), .Z(start_in[26]) );
  AND U1602 ( .A(start_reg[25]), .B(init), .Z(start_in[25]) );
  AND U1603 ( .A(start_reg[24]), .B(init), .Z(start_in[24]) );
  AND U1604 ( .A(start_reg[23]), .B(init), .Z(start_in[23]) );
  AND U1605 ( .A(start_reg[22]), .B(init), .Z(start_in[22]) );
  AND U1606 ( .A(start_reg[21]), .B(init), .Z(start_in[21]) );
  AND U1607 ( .A(start_reg[20]), .B(init), .Z(start_in[20]) );
  AND U1608 ( .A(start_reg[1]), .B(init), .Z(start_in[1]) );
  AND U1609 ( .A(start_reg[19]), .B(init), .Z(start_in[19]) );
  AND U1610 ( .A(start_reg[18]), .B(init), .Z(start_in[18]) );
  AND U1611 ( .A(start_reg[17]), .B(init), .Z(start_in[17]) );
  AND U1612 ( .A(start_reg[16]), .B(init), .Z(start_in[16]) );
  AND U1613 ( .A(start_reg[15]), .B(init), .Z(start_in[15]) );
  AND U1614 ( .A(start_reg[14]), .B(init), .Z(start_in[14]) );
  AND U1615 ( .A(start_reg[13]), .B(init), .Z(start_in[13]) );
  AND U1616 ( .A(start_reg[12]), .B(init), .Z(start_in[12]) );
  AND U1617 ( .A(start_reg[11]), .B(init), .Z(start_in[11]) );
  AND U1618 ( .A(start_reg[10]), .B(init), .Z(start_in[10]) );
  NANDN U1619 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  XOR U1620 ( .A(mul_pow), .B(n1825), .Z(n977) );
  NAND U1621 ( .A(n1236), .B(n1237), .Z(n976) );
  NANDN U1622 ( .A(n1238), .B(ereg[0]), .Z(n1237) );
  NANDN U1623 ( .A(init), .B(e[0]), .Z(n1236) );
  NAND U1624 ( .A(n1239), .B(n1240), .Z(n975) );
  NANDN U1625 ( .A(init), .B(e[1]), .Z(n1240) );
  AND U1626 ( .A(n1241), .B(n1242), .Z(n1239) );
  NAND U1627 ( .A(n1243), .B(ereg[0]), .Z(n1242) );
  NANDN U1628 ( .A(n1238), .B(ereg[1]), .Z(n1241) );
  NAND U1629 ( .A(n1244), .B(n1245), .Z(n974) );
  NANDN U1630 ( .A(init), .B(e[2]), .Z(n1245) );
  AND U1631 ( .A(n1246), .B(n1247), .Z(n1244) );
  NAND U1632 ( .A(ereg[1]), .B(n1243), .Z(n1247) );
  NANDN U1633 ( .A(n1238), .B(ereg[2]), .Z(n1246) );
  NAND U1634 ( .A(n1248), .B(n1249), .Z(n973) );
  NANDN U1635 ( .A(init), .B(e[3]), .Z(n1249) );
  AND U1636 ( .A(n1250), .B(n1251), .Z(n1248) );
  NAND U1637 ( .A(ereg[2]), .B(n1243), .Z(n1251) );
  NANDN U1638 ( .A(n1238), .B(ereg[3]), .Z(n1250) );
  NAND U1639 ( .A(n1252), .B(n1253), .Z(n972) );
  NANDN U1640 ( .A(init), .B(e[4]), .Z(n1253) );
  AND U1641 ( .A(n1254), .B(n1255), .Z(n1252) );
  NAND U1642 ( .A(ereg[3]), .B(n1243), .Z(n1255) );
  NANDN U1643 ( .A(n1238), .B(ereg[4]), .Z(n1254) );
  NAND U1644 ( .A(n1256), .B(n1257), .Z(n971) );
  NANDN U1645 ( .A(init), .B(e[5]), .Z(n1257) );
  AND U1646 ( .A(n1258), .B(n1259), .Z(n1256) );
  NAND U1647 ( .A(ereg[4]), .B(n1243), .Z(n1259) );
  NANDN U1648 ( .A(n1238), .B(ereg[5]), .Z(n1258) );
  NAND U1649 ( .A(n1260), .B(n1261), .Z(n970) );
  NANDN U1650 ( .A(init), .B(e[6]), .Z(n1261) );
  AND U1651 ( .A(n1262), .B(n1263), .Z(n1260) );
  NAND U1652 ( .A(ereg[5]), .B(n1243), .Z(n1263) );
  NANDN U1653 ( .A(n1238), .B(ereg[6]), .Z(n1262) );
  NAND U1654 ( .A(n1264), .B(n1265), .Z(n969) );
  NANDN U1655 ( .A(init), .B(e[7]), .Z(n1265) );
  AND U1656 ( .A(n1266), .B(n1267), .Z(n1264) );
  NAND U1657 ( .A(ereg[6]), .B(n1243), .Z(n1267) );
  NANDN U1658 ( .A(n1238), .B(ereg[7]), .Z(n1266) );
  NAND U1659 ( .A(n1268), .B(n1269), .Z(n968) );
  NANDN U1660 ( .A(init), .B(e[8]), .Z(n1269) );
  AND U1661 ( .A(n1270), .B(n1271), .Z(n1268) );
  NAND U1662 ( .A(ereg[7]), .B(n1243), .Z(n1271) );
  NANDN U1663 ( .A(n1238), .B(ereg[8]), .Z(n1270) );
  NAND U1664 ( .A(n1272), .B(n1273), .Z(n967) );
  NANDN U1665 ( .A(init), .B(e[9]), .Z(n1273) );
  AND U1666 ( .A(n1274), .B(n1275), .Z(n1272) );
  NAND U1667 ( .A(ereg[8]), .B(n1243), .Z(n1275) );
  NANDN U1668 ( .A(n1238), .B(ereg[9]), .Z(n1274) );
  NAND U1669 ( .A(n1276), .B(n1277), .Z(n966) );
  NANDN U1670 ( .A(init), .B(e[10]), .Z(n1277) );
  AND U1671 ( .A(n1278), .B(n1279), .Z(n1276) );
  NAND U1672 ( .A(ereg[9]), .B(n1243), .Z(n1279) );
  NANDN U1673 ( .A(n1238), .B(ereg[10]), .Z(n1278) );
  NAND U1674 ( .A(n1280), .B(n1281), .Z(n965) );
  NANDN U1675 ( .A(init), .B(e[11]), .Z(n1281) );
  AND U1676 ( .A(n1282), .B(n1283), .Z(n1280) );
  NAND U1677 ( .A(ereg[10]), .B(n1243), .Z(n1283) );
  NANDN U1678 ( .A(n1238), .B(ereg[11]), .Z(n1282) );
  NAND U1679 ( .A(n1284), .B(n1285), .Z(n964) );
  NANDN U1680 ( .A(init), .B(e[12]), .Z(n1285) );
  AND U1681 ( .A(n1286), .B(n1287), .Z(n1284) );
  NAND U1682 ( .A(ereg[11]), .B(n1243), .Z(n1287) );
  NANDN U1683 ( .A(n1238), .B(ereg[12]), .Z(n1286) );
  NAND U1684 ( .A(n1288), .B(n1289), .Z(n963) );
  NANDN U1685 ( .A(init), .B(e[13]), .Z(n1289) );
  AND U1686 ( .A(n1290), .B(n1291), .Z(n1288) );
  NAND U1687 ( .A(ereg[12]), .B(n1243), .Z(n1291) );
  NANDN U1688 ( .A(n1238), .B(ereg[13]), .Z(n1290) );
  NAND U1689 ( .A(n1292), .B(n1293), .Z(n962) );
  NANDN U1690 ( .A(init), .B(e[14]), .Z(n1293) );
  AND U1691 ( .A(n1294), .B(n1295), .Z(n1292) );
  NAND U1692 ( .A(ereg[13]), .B(n1243), .Z(n1295) );
  NANDN U1693 ( .A(n1238), .B(ereg[14]), .Z(n1294) );
  NAND U1694 ( .A(n1296), .B(n1297), .Z(n961) );
  NANDN U1695 ( .A(init), .B(e[15]), .Z(n1297) );
  AND U1696 ( .A(n1298), .B(n1299), .Z(n1296) );
  NAND U1697 ( .A(ereg[14]), .B(n1243), .Z(n1299) );
  NANDN U1698 ( .A(n1238), .B(ereg[15]), .Z(n1298) );
  NAND U1699 ( .A(n1300), .B(n1301), .Z(n960) );
  NANDN U1700 ( .A(init), .B(e[16]), .Z(n1301) );
  AND U1701 ( .A(n1302), .B(n1303), .Z(n1300) );
  NAND U1702 ( .A(ereg[15]), .B(n1243), .Z(n1303) );
  NANDN U1703 ( .A(n1238), .B(ereg[16]), .Z(n1302) );
  NAND U1704 ( .A(n1304), .B(n1305), .Z(n959) );
  NANDN U1705 ( .A(init), .B(e[17]), .Z(n1305) );
  AND U1706 ( .A(n1306), .B(n1307), .Z(n1304) );
  NAND U1707 ( .A(ereg[16]), .B(n1243), .Z(n1307) );
  NANDN U1708 ( .A(n1238), .B(ereg[17]), .Z(n1306) );
  NAND U1709 ( .A(n1308), .B(n1309), .Z(n958) );
  NANDN U1710 ( .A(init), .B(e[18]), .Z(n1309) );
  AND U1711 ( .A(n1310), .B(n1311), .Z(n1308) );
  NAND U1712 ( .A(ereg[17]), .B(n1243), .Z(n1311) );
  NANDN U1713 ( .A(n1238), .B(ereg[18]), .Z(n1310) );
  NAND U1714 ( .A(n1312), .B(n1313), .Z(n957) );
  NANDN U1715 ( .A(init), .B(e[19]), .Z(n1313) );
  AND U1716 ( .A(n1314), .B(n1315), .Z(n1312) );
  NAND U1717 ( .A(ereg[18]), .B(n1243), .Z(n1315) );
  NANDN U1718 ( .A(n1238), .B(ereg[19]), .Z(n1314) );
  NAND U1719 ( .A(n1316), .B(n1317), .Z(n956) );
  NANDN U1720 ( .A(init), .B(e[20]), .Z(n1317) );
  AND U1721 ( .A(n1318), .B(n1319), .Z(n1316) );
  NAND U1722 ( .A(ereg[19]), .B(n1243), .Z(n1319) );
  NANDN U1723 ( .A(n1238), .B(ereg[20]), .Z(n1318) );
  NAND U1724 ( .A(n1320), .B(n1321), .Z(n955) );
  NANDN U1725 ( .A(init), .B(e[21]), .Z(n1321) );
  AND U1726 ( .A(n1322), .B(n1323), .Z(n1320) );
  NAND U1727 ( .A(ereg[20]), .B(n1243), .Z(n1323) );
  NANDN U1728 ( .A(n1238), .B(ereg[21]), .Z(n1322) );
  NAND U1729 ( .A(n1324), .B(n1325), .Z(n954) );
  NANDN U1730 ( .A(init), .B(e[22]), .Z(n1325) );
  AND U1731 ( .A(n1326), .B(n1327), .Z(n1324) );
  NAND U1732 ( .A(ereg[21]), .B(n1243), .Z(n1327) );
  NANDN U1733 ( .A(n1238), .B(ereg[22]), .Z(n1326) );
  NAND U1734 ( .A(n1328), .B(n1329), .Z(n953) );
  NANDN U1735 ( .A(init), .B(e[23]), .Z(n1329) );
  AND U1736 ( .A(n1330), .B(n1331), .Z(n1328) );
  NAND U1737 ( .A(ereg[22]), .B(n1243), .Z(n1331) );
  NANDN U1738 ( .A(n1238), .B(ereg[23]), .Z(n1330) );
  NAND U1739 ( .A(n1332), .B(n1333), .Z(n952) );
  NANDN U1740 ( .A(init), .B(e[24]), .Z(n1333) );
  AND U1741 ( .A(n1334), .B(n1335), .Z(n1332) );
  NAND U1742 ( .A(ereg[23]), .B(n1243), .Z(n1335) );
  NANDN U1743 ( .A(n1238), .B(ereg[24]), .Z(n1334) );
  NAND U1744 ( .A(n1336), .B(n1337), .Z(n951) );
  NANDN U1745 ( .A(init), .B(e[25]), .Z(n1337) );
  AND U1746 ( .A(n1338), .B(n1339), .Z(n1336) );
  NAND U1747 ( .A(ereg[24]), .B(n1243), .Z(n1339) );
  NANDN U1748 ( .A(n1238), .B(ereg[25]), .Z(n1338) );
  NAND U1749 ( .A(n1340), .B(n1341), .Z(n950) );
  NANDN U1750 ( .A(init), .B(e[26]), .Z(n1341) );
  AND U1751 ( .A(n1342), .B(n1343), .Z(n1340) );
  NAND U1752 ( .A(ereg[25]), .B(n1243), .Z(n1343) );
  NANDN U1753 ( .A(n1238), .B(ereg[26]), .Z(n1342) );
  NAND U1754 ( .A(n1344), .B(n1345), .Z(n949) );
  NANDN U1755 ( .A(init), .B(e[27]), .Z(n1345) );
  AND U1756 ( .A(n1346), .B(n1347), .Z(n1344) );
  NAND U1757 ( .A(ereg[26]), .B(n1243), .Z(n1347) );
  NANDN U1758 ( .A(n1238), .B(ereg[27]), .Z(n1346) );
  NAND U1759 ( .A(n1348), .B(n1349), .Z(n948) );
  NANDN U1760 ( .A(init), .B(e[28]), .Z(n1349) );
  AND U1761 ( .A(n1350), .B(n1351), .Z(n1348) );
  NAND U1762 ( .A(ereg[27]), .B(n1243), .Z(n1351) );
  NANDN U1763 ( .A(n1238), .B(ereg[28]), .Z(n1350) );
  NAND U1764 ( .A(n1352), .B(n1353), .Z(n947) );
  NANDN U1765 ( .A(init), .B(e[29]), .Z(n1353) );
  AND U1766 ( .A(n1354), .B(n1355), .Z(n1352) );
  NAND U1767 ( .A(ereg[28]), .B(n1243), .Z(n1355) );
  NANDN U1768 ( .A(n1238), .B(ereg[29]), .Z(n1354) );
  NAND U1769 ( .A(n1356), .B(n1357), .Z(n946) );
  NANDN U1770 ( .A(init), .B(e[30]), .Z(n1357) );
  AND U1771 ( .A(n1358), .B(n1359), .Z(n1356) );
  NAND U1772 ( .A(ereg[29]), .B(n1243), .Z(n1359) );
  NANDN U1773 ( .A(n1238), .B(ereg[30]), .Z(n1358) );
  NAND U1774 ( .A(n1360), .B(n1361), .Z(n945) );
  NANDN U1775 ( .A(init), .B(e[31]), .Z(n1361) );
  AND U1776 ( .A(n1362), .B(n1363), .Z(n1360) );
  NAND U1777 ( .A(ereg[30]), .B(n1243), .Z(n1363) );
  NANDN U1778 ( .A(n1238), .B(ereg[31]), .Z(n1362) );
  NAND U1779 ( .A(n1364), .B(n1365), .Z(n944) );
  NANDN U1780 ( .A(init), .B(e[32]), .Z(n1365) );
  AND U1781 ( .A(n1366), .B(n1367), .Z(n1364) );
  NAND U1782 ( .A(ereg[31]), .B(n1243), .Z(n1367) );
  NANDN U1783 ( .A(n1238), .B(ereg[32]), .Z(n1366) );
  NAND U1784 ( .A(n1368), .B(n1369), .Z(n943) );
  NANDN U1785 ( .A(init), .B(e[33]), .Z(n1369) );
  AND U1786 ( .A(n1370), .B(n1371), .Z(n1368) );
  NAND U1787 ( .A(ereg[32]), .B(n1243), .Z(n1371) );
  NANDN U1788 ( .A(n1238), .B(ereg[33]), .Z(n1370) );
  NAND U1789 ( .A(n1372), .B(n1373), .Z(n942) );
  NANDN U1790 ( .A(init), .B(e[34]), .Z(n1373) );
  AND U1791 ( .A(n1374), .B(n1375), .Z(n1372) );
  NAND U1792 ( .A(ereg[33]), .B(n1243), .Z(n1375) );
  NANDN U1793 ( .A(n1238), .B(ereg[34]), .Z(n1374) );
  NAND U1794 ( .A(n1376), .B(n1377), .Z(n941) );
  NANDN U1795 ( .A(init), .B(e[35]), .Z(n1377) );
  AND U1796 ( .A(n1378), .B(n1379), .Z(n1376) );
  NAND U1797 ( .A(ereg[34]), .B(n1243), .Z(n1379) );
  NANDN U1798 ( .A(n1238), .B(ereg[35]), .Z(n1378) );
  NAND U1799 ( .A(n1380), .B(n1381), .Z(n940) );
  NANDN U1800 ( .A(init), .B(e[36]), .Z(n1381) );
  AND U1801 ( .A(n1382), .B(n1383), .Z(n1380) );
  NAND U1802 ( .A(ereg[35]), .B(n1243), .Z(n1383) );
  NANDN U1803 ( .A(n1238), .B(ereg[36]), .Z(n1382) );
  NAND U1804 ( .A(n1384), .B(n1385), .Z(n939) );
  NANDN U1805 ( .A(init), .B(e[37]), .Z(n1385) );
  AND U1806 ( .A(n1386), .B(n1387), .Z(n1384) );
  NAND U1807 ( .A(ereg[36]), .B(n1243), .Z(n1387) );
  NANDN U1808 ( .A(n1238), .B(ereg[37]), .Z(n1386) );
  NAND U1809 ( .A(n1388), .B(n1389), .Z(n938) );
  NANDN U1810 ( .A(init), .B(e[38]), .Z(n1389) );
  AND U1811 ( .A(n1390), .B(n1391), .Z(n1388) );
  NAND U1812 ( .A(ereg[37]), .B(n1243), .Z(n1391) );
  NANDN U1813 ( .A(n1238), .B(ereg[38]), .Z(n1390) );
  NAND U1814 ( .A(n1392), .B(n1393), .Z(n937) );
  NANDN U1815 ( .A(init), .B(e[39]), .Z(n1393) );
  AND U1816 ( .A(n1394), .B(n1395), .Z(n1392) );
  NAND U1817 ( .A(ereg[38]), .B(n1243), .Z(n1395) );
  NANDN U1818 ( .A(n1238), .B(ereg[39]), .Z(n1394) );
  NAND U1819 ( .A(n1396), .B(n1397), .Z(n936) );
  NANDN U1820 ( .A(init), .B(e[40]), .Z(n1397) );
  AND U1821 ( .A(n1398), .B(n1399), .Z(n1396) );
  NAND U1822 ( .A(ereg[39]), .B(n1243), .Z(n1399) );
  NANDN U1823 ( .A(n1238), .B(ereg[40]), .Z(n1398) );
  NAND U1824 ( .A(n1400), .B(n1401), .Z(n935) );
  NANDN U1825 ( .A(init), .B(e[41]), .Z(n1401) );
  AND U1826 ( .A(n1402), .B(n1403), .Z(n1400) );
  NAND U1827 ( .A(ereg[40]), .B(n1243), .Z(n1403) );
  NANDN U1828 ( .A(n1238), .B(ereg[41]), .Z(n1402) );
  NAND U1829 ( .A(n1404), .B(n1405), .Z(n934) );
  NANDN U1830 ( .A(init), .B(e[42]), .Z(n1405) );
  AND U1831 ( .A(n1406), .B(n1407), .Z(n1404) );
  NAND U1832 ( .A(ereg[41]), .B(n1243), .Z(n1407) );
  NANDN U1833 ( .A(n1238), .B(ereg[42]), .Z(n1406) );
  NAND U1834 ( .A(n1408), .B(n1409), .Z(n933) );
  NANDN U1835 ( .A(init), .B(e[43]), .Z(n1409) );
  AND U1836 ( .A(n1410), .B(n1411), .Z(n1408) );
  NAND U1837 ( .A(ereg[42]), .B(n1243), .Z(n1411) );
  NANDN U1838 ( .A(n1238), .B(ereg[43]), .Z(n1410) );
  NAND U1839 ( .A(n1412), .B(n1413), .Z(n932) );
  NANDN U1840 ( .A(init), .B(e[44]), .Z(n1413) );
  AND U1841 ( .A(n1414), .B(n1415), .Z(n1412) );
  NAND U1842 ( .A(ereg[43]), .B(n1243), .Z(n1415) );
  NANDN U1843 ( .A(n1238), .B(ereg[44]), .Z(n1414) );
  NAND U1844 ( .A(n1416), .B(n1417), .Z(n931) );
  NANDN U1845 ( .A(init), .B(e[45]), .Z(n1417) );
  AND U1846 ( .A(n1418), .B(n1419), .Z(n1416) );
  NAND U1847 ( .A(ereg[44]), .B(n1243), .Z(n1419) );
  NANDN U1848 ( .A(n1238), .B(ereg[45]), .Z(n1418) );
  NAND U1849 ( .A(n1420), .B(n1421), .Z(n930) );
  NANDN U1850 ( .A(init), .B(e[46]), .Z(n1421) );
  AND U1851 ( .A(n1422), .B(n1423), .Z(n1420) );
  NAND U1852 ( .A(ereg[45]), .B(n1243), .Z(n1423) );
  NANDN U1853 ( .A(n1238), .B(ereg[46]), .Z(n1422) );
  NAND U1854 ( .A(n1424), .B(n1425), .Z(n929) );
  NANDN U1855 ( .A(init), .B(e[47]), .Z(n1425) );
  AND U1856 ( .A(n1426), .B(n1427), .Z(n1424) );
  NAND U1857 ( .A(ereg[46]), .B(n1243), .Z(n1427) );
  NANDN U1858 ( .A(n1238), .B(ereg[47]), .Z(n1426) );
  NAND U1859 ( .A(n1428), .B(n1429), .Z(n928) );
  NANDN U1860 ( .A(init), .B(e[48]), .Z(n1429) );
  AND U1861 ( .A(n1430), .B(n1431), .Z(n1428) );
  NAND U1862 ( .A(ereg[47]), .B(n1243), .Z(n1431) );
  NANDN U1863 ( .A(n1238), .B(ereg[48]), .Z(n1430) );
  NAND U1864 ( .A(n1432), .B(n1433), .Z(n927) );
  NANDN U1865 ( .A(init), .B(e[49]), .Z(n1433) );
  AND U1866 ( .A(n1434), .B(n1435), .Z(n1432) );
  NAND U1867 ( .A(ereg[48]), .B(n1243), .Z(n1435) );
  NANDN U1868 ( .A(n1238), .B(ereg[49]), .Z(n1434) );
  NAND U1869 ( .A(n1436), .B(n1437), .Z(n926) );
  NANDN U1870 ( .A(init), .B(e[50]), .Z(n1437) );
  AND U1871 ( .A(n1438), .B(n1439), .Z(n1436) );
  NAND U1872 ( .A(ereg[49]), .B(n1243), .Z(n1439) );
  NANDN U1873 ( .A(n1238), .B(ereg[50]), .Z(n1438) );
  NAND U1874 ( .A(n1440), .B(n1441), .Z(n925) );
  NANDN U1875 ( .A(init), .B(e[51]), .Z(n1441) );
  AND U1876 ( .A(n1442), .B(n1443), .Z(n1440) );
  NAND U1877 ( .A(ereg[50]), .B(n1243), .Z(n1443) );
  NANDN U1878 ( .A(n1238), .B(ereg[51]), .Z(n1442) );
  NAND U1879 ( .A(n1444), .B(n1445), .Z(n924) );
  NANDN U1880 ( .A(init), .B(e[52]), .Z(n1445) );
  AND U1881 ( .A(n1446), .B(n1447), .Z(n1444) );
  NAND U1882 ( .A(ereg[51]), .B(n1243), .Z(n1447) );
  NANDN U1883 ( .A(n1238), .B(ereg[52]), .Z(n1446) );
  NAND U1884 ( .A(n1448), .B(n1449), .Z(n923) );
  NANDN U1885 ( .A(init), .B(e[53]), .Z(n1449) );
  AND U1886 ( .A(n1450), .B(n1451), .Z(n1448) );
  NAND U1887 ( .A(ereg[52]), .B(n1243), .Z(n1451) );
  NANDN U1888 ( .A(n1238), .B(ereg[53]), .Z(n1450) );
  NAND U1889 ( .A(n1452), .B(n1453), .Z(n922) );
  NANDN U1890 ( .A(init), .B(e[54]), .Z(n1453) );
  AND U1891 ( .A(n1454), .B(n1455), .Z(n1452) );
  NAND U1892 ( .A(ereg[53]), .B(n1243), .Z(n1455) );
  NANDN U1893 ( .A(n1238), .B(ereg[54]), .Z(n1454) );
  NAND U1894 ( .A(n1456), .B(n1457), .Z(n921) );
  NANDN U1895 ( .A(init), .B(e[55]), .Z(n1457) );
  AND U1896 ( .A(n1458), .B(n1459), .Z(n1456) );
  NAND U1897 ( .A(ereg[54]), .B(n1243), .Z(n1459) );
  NANDN U1898 ( .A(n1238), .B(ereg[55]), .Z(n1458) );
  NAND U1899 ( .A(n1460), .B(n1461), .Z(n920) );
  NANDN U1900 ( .A(init), .B(e[56]), .Z(n1461) );
  AND U1901 ( .A(n1462), .B(n1463), .Z(n1460) );
  NAND U1902 ( .A(ereg[55]), .B(n1243), .Z(n1463) );
  NANDN U1903 ( .A(n1238), .B(ereg[56]), .Z(n1462) );
  NAND U1904 ( .A(n1464), .B(n1465), .Z(n919) );
  NANDN U1905 ( .A(init), .B(e[57]), .Z(n1465) );
  AND U1906 ( .A(n1466), .B(n1467), .Z(n1464) );
  NAND U1907 ( .A(ereg[56]), .B(n1243), .Z(n1467) );
  NANDN U1908 ( .A(n1238), .B(ereg[57]), .Z(n1466) );
  NAND U1909 ( .A(n1468), .B(n1469), .Z(n918) );
  NANDN U1910 ( .A(init), .B(e[58]), .Z(n1469) );
  AND U1911 ( .A(n1470), .B(n1471), .Z(n1468) );
  NAND U1912 ( .A(ereg[57]), .B(n1243), .Z(n1471) );
  NANDN U1913 ( .A(n1238), .B(ereg[58]), .Z(n1470) );
  NAND U1914 ( .A(n1472), .B(n1473), .Z(n917) );
  NANDN U1915 ( .A(init), .B(e[59]), .Z(n1473) );
  AND U1916 ( .A(n1474), .B(n1475), .Z(n1472) );
  NAND U1917 ( .A(ereg[58]), .B(n1243), .Z(n1475) );
  NANDN U1918 ( .A(n1238), .B(ereg[59]), .Z(n1474) );
  NAND U1919 ( .A(n1476), .B(n1477), .Z(n916) );
  NANDN U1920 ( .A(init), .B(e[60]), .Z(n1477) );
  AND U1921 ( .A(n1478), .B(n1479), .Z(n1476) );
  NAND U1922 ( .A(ereg[59]), .B(n1243), .Z(n1479) );
  NANDN U1923 ( .A(n1238), .B(ereg[60]), .Z(n1478) );
  NAND U1924 ( .A(n1480), .B(n1481), .Z(n915) );
  NANDN U1925 ( .A(init), .B(e[61]), .Z(n1481) );
  AND U1926 ( .A(n1482), .B(n1483), .Z(n1480) );
  NAND U1927 ( .A(ereg[60]), .B(n1243), .Z(n1483) );
  NANDN U1928 ( .A(n1238), .B(ereg[61]), .Z(n1482) );
  NAND U1929 ( .A(n1484), .B(n1485), .Z(n914) );
  NANDN U1930 ( .A(init), .B(e[62]), .Z(n1485) );
  AND U1931 ( .A(n1486), .B(n1487), .Z(n1484) );
  NAND U1932 ( .A(ereg[61]), .B(n1243), .Z(n1487) );
  NANDN U1933 ( .A(n1238), .B(ereg[62]), .Z(n1486) );
  NAND U1934 ( .A(n1488), .B(n1489), .Z(n913) );
  NANDN U1935 ( .A(init), .B(e[63]), .Z(n1489) );
  AND U1936 ( .A(n1490), .B(n1491), .Z(n1488) );
  NAND U1937 ( .A(ereg[62]), .B(n1243), .Z(n1491) );
  ANDN U1938 ( .B(n1238), .A(n1492), .Z(n1243) );
  NANDN U1939 ( .A(n1238), .B(ereg[63]), .Z(n1490) );
  AND U1940 ( .A(n1493), .B(n980), .Z(n1238) );
  NANDN U1941 ( .A(mul_pow), .B(init), .Z(n980) );
  NAND U1942 ( .A(n1492), .B(init), .Z(n1493) );
  NAND U1943 ( .A(n1494), .B(n1117), .Z(n912) );
  NANDN U1944 ( .A(init), .B(m[63]), .Z(n1117) );
  AND U1945 ( .A(n1495), .B(n1496), .Z(n1494) );
  NAND U1946 ( .A(o[63]), .B(n1497), .Z(n1496) );
  NANDN U1947 ( .A(n1498), .B(creg[63]), .Z(n1495) );
  NAND U1948 ( .A(n1499), .B(n1235), .Z(n911) );
  NANDN U1949 ( .A(init), .B(m[0]), .Z(n1235) );
  AND U1950 ( .A(n1500), .B(n1501), .Z(n1499) );
  NAND U1951 ( .A(o[0]), .B(n1497), .Z(n1501) );
  NANDN U1952 ( .A(n1498), .B(creg[0]), .Z(n1500) );
  NAND U1953 ( .A(n1502), .B(n1213), .Z(n910) );
  NANDN U1954 ( .A(init), .B(m[1]), .Z(n1213) );
  AND U1955 ( .A(n1503), .B(n1504), .Z(n1502) );
  NAND U1956 ( .A(o[1]), .B(n1497), .Z(n1504) );
  NANDN U1957 ( .A(n1498), .B(creg[1]), .Z(n1503) );
  NAND U1958 ( .A(n1505), .B(n1191), .Z(n909) );
  NANDN U1959 ( .A(init), .B(m[2]), .Z(n1191) );
  AND U1960 ( .A(n1506), .B(n1507), .Z(n1505) );
  NAND U1961 ( .A(o[2]), .B(n1497), .Z(n1507) );
  NANDN U1962 ( .A(n1498), .B(creg[2]), .Z(n1506) );
  NAND U1963 ( .A(n1508), .B(n1169), .Z(n908) );
  NANDN U1964 ( .A(init), .B(m[3]), .Z(n1169) );
  AND U1965 ( .A(n1509), .B(n1510), .Z(n1508) );
  NAND U1966 ( .A(o[3]), .B(n1497), .Z(n1510) );
  NANDN U1967 ( .A(n1498), .B(creg[3]), .Z(n1509) );
  NAND U1968 ( .A(n1511), .B(n1147), .Z(n907) );
  NANDN U1969 ( .A(init), .B(m[4]), .Z(n1147) );
  AND U1970 ( .A(n1512), .B(n1513), .Z(n1511) );
  NAND U1971 ( .A(o[4]), .B(n1497), .Z(n1513) );
  NANDN U1972 ( .A(n1498), .B(creg[4]), .Z(n1512) );
  NAND U1973 ( .A(n1514), .B(n1125), .Z(n906) );
  NANDN U1974 ( .A(init), .B(m[5]), .Z(n1125) );
  AND U1975 ( .A(n1515), .B(n1516), .Z(n1514) );
  NAND U1976 ( .A(o[5]), .B(n1497), .Z(n1516) );
  NANDN U1977 ( .A(n1498), .B(creg[5]), .Z(n1515) );
  NAND U1978 ( .A(n1517), .B(n1115), .Z(n905) );
  NANDN U1979 ( .A(init), .B(m[6]), .Z(n1115) );
  AND U1980 ( .A(n1518), .B(n1519), .Z(n1517) );
  NAND U1981 ( .A(o[6]), .B(n1497), .Z(n1519) );
  NANDN U1982 ( .A(n1498), .B(creg[6]), .Z(n1518) );
  NAND U1983 ( .A(n1520), .B(n1113), .Z(n904) );
  NANDN U1984 ( .A(init), .B(m[7]), .Z(n1113) );
  AND U1985 ( .A(n1521), .B(n1522), .Z(n1520) );
  NAND U1986 ( .A(o[7]), .B(n1497), .Z(n1522) );
  NANDN U1987 ( .A(n1498), .B(creg[7]), .Z(n1521) );
  NAND U1988 ( .A(n1523), .B(n1111), .Z(n903) );
  NANDN U1989 ( .A(init), .B(m[8]), .Z(n1111) );
  AND U1990 ( .A(n1524), .B(n1525), .Z(n1523) );
  NAND U1991 ( .A(o[8]), .B(n1497), .Z(n1525) );
  NANDN U1992 ( .A(n1498), .B(creg[8]), .Z(n1524) );
  NAND U1993 ( .A(n1526), .B(n1109), .Z(n902) );
  NANDN U1994 ( .A(init), .B(m[9]), .Z(n1109) );
  AND U1995 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1996 ( .A(o[9]), .B(n1497), .Z(n1528) );
  NANDN U1997 ( .A(n1498), .B(creg[9]), .Z(n1527) );
  NAND U1998 ( .A(n1529), .B(n1233), .Z(n901) );
  NANDN U1999 ( .A(init), .B(m[10]), .Z(n1233) );
  AND U2000 ( .A(n1530), .B(n1531), .Z(n1529) );
  NAND U2001 ( .A(o[10]), .B(n1497), .Z(n1531) );
  NANDN U2002 ( .A(n1498), .B(creg[10]), .Z(n1530) );
  NAND U2003 ( .A(n1532), .B(n1231), .Z(n900) );
  NANDN U2004 ( .A(init), .B(m[11]), .Z(n1231) );
  AND U2005 ( .A(n1533), .B(n1534), .Z(n1532) );
  NAND U2006 ( .A(o[11]), .B(n1497), .Z(n1534) );
  NANDN U2007 ( .A(n1498), .B(creg[11]), .Z(n1533) );
  NAND U2008 ( .A(n1535), .B(n1229), .Z(n899) );
  NANDN U2009 ( .A(init), .B(m[12]), .Z(n1229) );
  AND U2010 ( .A(n1536), .B(n1537), .Z(n1535) );
  NAND U2011 ( .A(o[12]), .B(n1497), .Z(n1537) );
  NANDN U2012 ( .A(n1498), .B(creg[12]), .Z(n1536) );
  NAND U2013 ( .A(n1538), .B(n1227), .Z(n898) );
  NANDN U2014 ( .A(init), .B(m[13]), .Z(n1227) );
  AND U2015 ( .A(n1539), .B(n1540), .Z(n1538) );
  NAND U2016 ( .A(o[13]), .B(n1497), .Z(n1540) );
  NANDN U2017 ( .A(n1498), .B(creg[13]), .Z(n1539) );
  NAND U2018 ( .A(n1541), .B(n1225), .Z(n897) );
  NANDN U2019 ( .A(init), .B(m[14]), .Z(n1225) );
  AND U2020 ( .A(n1542), .B(n1543), .Z(n1541) );
  NAND U2021 ( .A(o[14]), .B(n1497), .Z(n1543) );
  NANDN U2022 ( .A(n1498), .B(creg[14]), .Z(n1542) );
  NAND U2023 ( .A(n1544), .B(n1223), .Z(n896) );
  NANDN U2024 ( .A(init), .B(m[15]), .Z(n1223) );
  AND U2025 ( .A(n1545), .B(n1546), .Z(n1544) );
  NAND U2026 ( .A(o[15]), .B(n1497), .Z(n1546) );
  NANDN U2027 ( .A(n1498), .B(creg[15]), .Z(n1545) );
  NAND U2028 ( .A(n1547), .B(n1221), .Z(n895) );
  NANDN U2029 ( .A(init), .B(m[16]), .Z(n1221) );
  AND U2030 ( .A(n1548), .B(n1549), .Z(n1547) );
  NAND U2031 ( .A(o[16]), .B(n1497), .Z(n1549) );
  NANDN U2032 ( .A(n1498), .B(creg[16]), .Z(n1548) );
  NAND U2033 ( .A(n1550), .B(n1219), .Z(n894) );
  NANDN U2034 ( .A(init), .B(m[17]), .Z(n1219) );
  AND U2035 ( .A(n1551), .B(n1552), .Z(n1550) );
  NAND U2036 ( .A(o[17]), .B(n1497), .Z(n1552) );
  NANDN U2037 ( .A(n1498), .B(creg[17]), .Z(n1551) );
  NAND U2038 ( .A(n1553), .B(n1217), .Z(n893) );
  NANDN U2039 ( .A(init), .B(m[18]), .Z(n1217) );
  AND U2040 ( .A(n1554), .B(n1555), .Z(n1553) );
  NAND U2041 ( .A(o[18]), .B(n1497), .Z(n1555) );
  NANDN U2042 ( .A(n1498), .B(creg[18]), .Z(n1554) );
  NAND U2043 ( .A(n1556), .B(n1215), .Z(n892) );
  NANDN U2044 ( .A(init), .B(m[19]), .Z(n1215) );
  AND U2045 ( .A(n1557), .B(n1558), .Z(n1556) );
  NAND U2046 ( .A(o[19]), .B(n1497), .Z(n1558) );
  NANDN U2047 ( .A(n1498), .B(creg[19]), .Z(n1557) );
  NAND U2048 ( .A(n1559), .B(n1211), .Z(n891) );
  NANDN U2049 ( .A(init), .B(m[20]), .Z(n1211) );
  AND U2050 ( .A(n1560), .B(n1561), .Z(n1559) );
  NAND U2051 ( .A(o[20]), .B(n1497), .Z(n1561) );
  NANDN U2052 ( .A(n1498), .B(creg[20]), .Z(n1560) );
  NAND U2053 ( .A(n1562), .B(n1209), .Z(n890) );
  NANDN U2054 ( .A(init), .B(m[21]), .Z(n1209) );
  AND U2055 ( .A(n1563), .B(n1564), .Z(n1562) );
  NAND U2056 ( .A(o[21]), .B(n1497), .Z(n1564) );
  NANDN U2057 ( .A(n1498), .B(creg[21]), .Z(n1563) );
  NAND U2058 ( .A(n1565), .B(n1207), .Z(n889) );
  NANDN U2059 ( .A(init), .B(m[22]), .Z(n1207) );
  AND U2060 ( .A(n1566), .B(n1567), .Z(n1565) );
  NAND U2061 ( .A(o[22]), .B(n1497), .Z(n1567) );
  NANDN U2062 ( .A(n1498), .B(creg[22]), .Z(n1566) );
  NAND U2063 ( .A(n1568), .B(n1205), .Z(n888) );
  NANDN U2064 ( .A(init), .B(m[23]), .Z(n1205) );
  AND U2065 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U2066 ( .A(o[23]), .B(n1497), .Z(n1570) );
  NANDN U2067 ( .A(n1498), .B(creg[23]), .Z(n1569) );
  NAND U2068 ( .A(n1571), .B(n1203), .Z(n887) );
  NANDN U2069 ( .A(init), .B(m[24]), .Z(n1203) );
  AND U2070 ( .A(n1572), .B(n1573), .Z(n1571) );
  NAND U2071 ( .A(o[24]), .B(n1497), .Z(n1573) );
  NANDN U2072 ( .A(n1498), .B(creg[24]), .Z(n1572) );
  NAND U2073 ( .A(n1574), .B(n1201), .Z(n886) );
  NANDN U2074 ( .A(init), .B(m[25]), .Z(n1201) );
  AND U2075 ( .A(n1575), .B(n1576), .Z(n1574) );
  NAND U2076 ( .A(o[25]), .B(n1497), .Z(n1576) );
  NANDN U2077 ( .A(n1498), .B(creg[25]), .Z(n1575) );
  NAND U2078 ( .A(n1577), .B(n1199), .Z(n885) );
  NANDN U2079 ( .A(init), .B(m[26]), .Z(n1199) );
  AND U2080 ( .A(n1578), .B(n1579), .Z(n1577) );
  NAND U2081 ( .A(o[26]), .B(n1497), .Z(n1579) );
  NANDN U2082 ( .A(n1498), .B(creg[26]), .Z(n1578) );
  NAND U2083 ( .A(n1580), .B(n1197), .Z(n884) );
  NANDN U2084 ( .A(init), .B(m[27]), .Z(n1197) );
  AND U2085 ( .A(n1581), .B(n1582), .Z(n1580) );
  NAND U2086 ( .A(o[27]), .B(n1497), .Z(n1582) );
  NANDN U2087 ( .A(n1498), .B(creg[27]), .Z(n1581) );
  NAND U2088 ( .A(n1583), .B(n1195), .Z(n883) );
  NANDN U2089 ( .A(init), .B(m[28]), .Z(n1195) );
  AND U2090 ( .A(n1584), .B(n1585), .Z(n1583) );
  NAND U2091 ( .A(o[28]), .B(n1497), .Z(n1585) );
  NANDN U2092 ( .A(n1498), .B(creg[28]), .Z(n1584) );
  NAND U2093 ( .A(n1586), .B(n1193), .Z(n882) );
  NANDN U2094 ( .A(init), .B(m[29]), .Z(n1193) );
  AND U2095 ( .A(n1587), .B(n1588), .Z(n1586) );
  NAND U2096 ( .A(o[29]), .B(n1497), .Z(n1588) );
  NANDN U2097 ( .A(n1498), .B(creg[29]), .Z(n1587) );
  NAND U2098 ( .A(n1589), .B(n1189), .Z(n881) );
  NANDN U2099 ( .A(init), .B(m[30]), .Z(n1189) );
  AND U2100 ( .A(n1590), .B(n1591), .Z(n1589) );
  NAND U2101 ( .A(o[30]), .B(n1497), .Z(n1591) );
  NANDN U2102 ( .A(n1498), .B(creg[30]), .Z(n1590) );
  NAND U2103 ( .A(n1592), .B(n1187), .Z(n880) );
  NANDN U2104 ( .A(init), .B(m[31]), .Z(n1187) );
  AND U2105 ( .A(n1593), .B(n1594), .Z(n1592) );
  NAND U2106 ( .A(o[31]), .B(n1497), .Z(n1594) );
  NANDN U2107 ( .A(n1498), .B(creg[31]), .Z(n1593) );
  NAND U2108 ( .A(n1595), .B(n1185), .Z(n879) );
  NANDN U2109 ( .A(init), .B(m[32]), .Z(n1185) );
  AND U2110 ( .A(n1596), .B(n1597), .Z(n1595) );
  NAND U2111 ( .A(o[32]), .B(n1497), .Z(n1597) );
  NANDN U2112 ( .A(n1498), .B(creg[32]), .Z(n1596) );
  NAND U2113 ( .A(n1598), .B(n1183), .Z(n878) );
  NANDN U2114 ( .A(init), .B(m[33]), .Z(n1183) );
  AND U2115 ( .A(n1599), .B(n1600), .Z(n1598) );
  NAND U2116 ( .A(o[33]), .B(n1497), .Z(n1600) );
  NANDN U2117 ( .A(n1498), .B(creg[33]), .Z(n1599) );
  NAND U2118 ( .A(n1601), .B(n1181), .Z(n877) );
  NANDN U2119 ( .A(init), .B(m[34]), .Z(n1181) );
  AND U2120 ( .A(n1602), .B(n1603), .Z(n1601) );
  NAND U2121 ( .A(o[34]), .B(n1497), .Z(n1603) );
  NANDN U2122 ( .A(n1498), .B(creg[34]), .Z(n1602) );
  NAND U2123 ( .A(n1604), .B(n1179), .Z(n876) );
  NANDN U2124 ( .A(init), .B(m[35]), .Z(n1179) );
  AND U2125 ( .A(n1605), .B(n1606), .Z(n1604) );
  NAND U2126 ( .A(o[35]), .B(n1497), .Z(n1606) );
  NANDN U2127 ( .A(n1498), .B(creg[35]), .Z(n1605) );
  NAND U2128 ( .A(n1607), .B(n1177), .Z(n875) );
  NANDN U2129 ( .A(init), .B(m[36]), .Z(n1177) );
  AND U2130 ( .A(n1608), .B(n1609), .Z(n1607) );
  NAND U2131 ( .A(o[36]), .B(n1497), .Z(n1609) );
  NANDN U2132 ( .A(n1498), .B(creg[36]), .Z(n1608) );
  NAND U2133 ( .A(n1610), .B(n1175), .Z(n874) );
  NANDN U2134 ( .A(init), .B(m[37]), .Z(n1175) );
  AND U2135 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U2136 ( .A(o[37]), .B(n1497), .Z(n1612) );
  NANDN U2137 ( .A(n1498), .B(creg[37]), .Z(n1611) );
  NAND U2138 ( .A(n1613), .B(n1173), .Z(n873) );
  NANDN U2139 ( .A(init), .B(m[38]), .Z(n1173) );
  AND U2140 ( .A(n1614), .B(n1615), .Z(n1613) );
  NAND U2141 ( .A(o[38]), .B(n1497), .Z(n1615) );
  NANDN U2142 ( .A(n1498), .B(creg[38]), .Z(n1614) );
  NAND U2143 ( .A(n1616), .B(n1171), .Z(n872) );
  NANDN U2144 ( .A(init), .B(m[39]), .Z(n1171) );
  AND U2145 ( .A(n1617), .B(n1618), .Z(n1616) );
  NAND U2146 ( .A(o[39]), .B(n1497), .Z(n1618) );
  NANDN U2147 ( .A(n1498), .B(creg[39]), .Z(n1617) );
  NAND U2148 ( .A(n1619), .B(n1167), .Z(n871) );
  NANDN U2149 ( .A(init), .B(m[40]), .Z(n1167) );
  AND U2150 ( .A(n1620), .B(n1621), .Z(n1619) );
  NAND U2151 ( .A(o[40]), .B(n1497), .Z(n1621) );
  NANDN U2152 ( .A(n1498), .B(creg[40]), .Z(n1620) );
  NAND U2153 ( .A(n1622), .B(n1165), .Z(n870) );
  NANDN U2154 ( .A(init), .B(m[41]), .Z(n1165) );
  AND U2155 ( .A(n1623), .B(n1624), .Z(n1622) );
  NAND U2156 ( .A(o[41]), .B(n1497), .Z(n1624) );
  NANDN U2157 ( .A(n1498), .B(creg[41]), .Z(n1623) );
  NAND U2158 ( .A(n1625), .B(n1163), .Z(n869) );
  NANDN U2159 ( .A(init), .B(m[42]), .Z(n1163) );
  AND U2160 ( .A(n1626), .B(n1627), .Z(n1625) );
  NAND U2161 ( .A(o[42]), .B(n1497), .Z(n1627) );
  NANDN U2162 ( .A(n1498), .B(creg[42]), .Z(n1626) );
  NAND U2163 ( .A(n1628), .B(n1161), .Z(n868) );
  NANDN U2164 ( .A(init), .B(m[43]), .Z(n1161) );
  AND U2165 ( .A(n1629), .B(n1630), .Z(n1628) );
  NAND U2166 ( .A(o[43]), .B(n1497), .Z(n1630) );
  NANDN U2167 ( .A(n1498), .B(creg[43]), .Z(n1629) );
  NAND U2168 ( .A(n1631), .B(n1159), .Z(n867) );
  NANDN U2169 ( .A(init), .B(m[44]), .Z(n1159) );
  AND U2170 ( .A(n1632), .B(n1633), .Z(n1631) );
  NAND U2171 ( .A(o[44]), .B(n1497), .Z(n1633) );
  NANDN U2172 ( .A(n1498), .B(creg[44]), .Z(n1632) );
  NAND U2173 ( .A(n1634), .B(n1157), .Z(n866) );
  NANDN U2174 ( .A(init), .B(m[45]), .Z(n1157) );
  AND U2175 ( .A(n1635), .B(n1636), .Z(n1634) );
  NAND U2176 ( .A(o[45]), .B(n1497), .Z(n1636) );
  NANDN U2177 ( .A(n1498), .B(creg[45]), .Z(n1635) );
  NAND U2178 ( .A(n1637), .B(n1155), .Z(n865) );
  NANDN U2179 ( .A(init), .B(m[46]), .Z(n1155) );
  AND U2180 ( .A(n1638), .B(n1639), .Z(n1637) );
  NAND U2181 ( .A(o[46]), .B(n1497), .Z(n1639) );
  NANDN U2182 ( .A(n1498), .B(creg[46]), .Z(n1638) );
  NAND U2183 ( .A(n1640), .B(n1153), .Z(n864) );
  NANDN U2184 ( .A(init), .B(m[47]), .Z(n1153) );
  AND U2185 ( .A(n1641), .B(n1642), .Z(n1640) );
  NAND U2186 ( .A(o[47]), .B(n1497), .Z(n1642) );
  NANDN U2187 ( .A(n1498), .B(creg[47]), .Z(n1641) );
  NAND U2188 ( .A(n1643), .B(n1151), .Z(n863) );
  NANDN U2189 ( .A(init), .B(m[48]), .Z(n1151) );
  AND U2190 ( .A(n1644), .B(n1645), .Z(n1643) );
  NAND U2191 ( .A(o[48]), .B(n1497), .Z(n1645) );
  NANDN U2192 ( .A(n1498), .B(creg[48]), .Z(n1644) );
  NAND U2193 ( .A(n1646), .B(n1149), .Z(n862) );
  NANDN U2194 ( .A(init), .B(m[49]), .Z(n1149) );
  AND U2195 ( .A(n1647), .B(n1648), .Z(n1646) );
  NAND U2196 ( .A(o[49]), .B(n1497), .Z(n1648) );
  NANDN U2197 ( .A(n1498), .B(creg[49]), .Z(n1647) );
  NAND U2198 ( .A(n1649), .B(n1145), .Z(n861) );
  NANDN U2199 ( .A(init), .B(m[50]), .Z(n1145) );
  AND U2200 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U2201 ( .A(o[50]), .B(n1497), .Z(n1651) );
  NANDN U2202 ( .A(n1498), .B(creg[50]), .Z(n1650) );
  NAND U2203 ( .A(n1652), .B(n1143), .Z(n860) );
  NANDN U2204 ( .A(init), .B(m[51]), .Z(n1143) );
  AND U2205 ( .A(n1653), .B(n1654), .Z(n1652) );
  NAND U2206 ( .A(o[51]), .B(n1497), .Z(n1654) );
  NANDN U2207 ( .A(n1498), .B(creg[51]), .Z(n1653) );
  NAND U2208 ( .A(n1655), .B(n1141), .Z(n859) );
  NANDN U2209 ( .A(init), .B(m[52]), .Z(n1141) );
  AND U2210 ( .A(n1656), .B(n1657), .Z(n1655) );
  NAND U2211 ( .A(o[52]), .B(n1497), .Z(n1657) );
  NANDN U2212 ( .A(n1498), .B(creg[52]), .Z(n1656) );
  NAND U2213 ( .A(n1658), .B(n1139), .Z(n858) );
  NANDN U2214 ( .A(init), .B(m[53]), .Z(n1139) );
  AND U2215 ( .A(n1659), .B(n1660), .Z(n1658) );
  NAND U2216 ( .A(o[53]), .B(n1497), .Z(n1660) );
  NANDN U2217 ( .A(n1498), .B(creg[53]), .Z(n1659) );
  NAND U2218 ( .A(n1661), .B(n1137), .Z(n857) );
  NANDN U2219 ( .A(init), .B(m[54]), .Z(n1137) );
  AND U2220 ( .A(n1662), .B(n1663), .Z(n1661) );
  NAND U2221 ( .A(o[54]), .B(n1497), .Z(n1663) );
  NANDN U2222 ( .A(n1498), .B(creg[54]), .Z(n1662) );
  NAND U2223 ( .A(n1664), .B(n1135), .Z(n856) );
  NANDN U2224 ( .A(init), .B(m[55]), .Z(n1135) );
  AND U2225 ( .A(n1665), .B(n1666), .Z(n1664) );
  NAND U2226 ( .A(o[55]), .B(n1497), .Z(n1666) );
  NANDN U2227 ( .A(n1498), .B(creg[55]), .Z(n1665) );
  NAND U2228 ( .A(n1667), .B(n1133), .Z(n855) );
  NANDN U2229 ( .A(init), .B(m[56]), .Z(n1133) );
  AND U2230 ( .A(n1668), .B(n1669), .Z(n1667) );
  NAND U2231 ( .A(o[56]), .B(n1497), .Z(n1669) );
  NANDN U2232 ( .A(n1498), .B(creg[56]), .Z(n1668) );
  NAND U2233 ( .A(n1670), .B(n1131), .Z(n854) );
  NANDN U2234 ( .A(init), .B(m[57]), .Z(n1131) );
  AND U2235 ( .A(n1671), .B(n1672), .Z(n1670) );
  NAND U2236 ( .A(o[57]), .B(n1497), .Z(n1672) );
  NANDN U2237 ( .A(n1498), .B(creg[57]), .Z(n1671) );
  NAND U2238 ( .A(n1673), .B(n1129), .Z(n853) );
  NANDN U2239 ( .A(init), .B(m[58]), .Z(n1129) );
  AND U2240 ( .A(n1674), .B(n1675), .Z(n1673) );
  NAND U2241 ( .A(o[58]), .B(n1497), .Z(n1675) );
  NANDN U2242 ( .A(n1498), .B(creg[58]), .Z(n1674) );
  NAND U2243 ( .A(n1676), .B(n1127), .Z(n852) );
  NANDN U2244 ( .A(init), .B(m[59]), .Z(n1127) );
  AND U2245 ( .A(n1677), .B(n1678), .Z(n1676) );
  NAND U2246 ( .A(o[59]), .B(n1497), .Z(n1678) );
  NANDN U2247 ( .A(n1498), .B(creg[59]), .Z(n1677) );
  NAND U2248 ( .A(n1679), .B(n1123), .Z(n851) );
  NANDN U2249 ( .A(init), .B(m[60]), .Z(n1123) );
  AND U2250 ( .A(n1680), .B(n1681), .Z(n1679) );
  NAND U2251 ( .A(o[60]), .B(n1497), .Z(n1681) );
  NANDN U2252 ( .A(n1498), .B(creg[60]), .Z(n1680) );
  NAND U2253 ( .A(n1682), .B(n1121), .Z(n850) );
  NANDN U2254 ( .A(init), .B(m[61]), .Z(n1121) );
  AND U2255 ( .A(n1683), .B(n1684), .Z(n1682) );
  NAND U2256 ( .A(o[61]), .B(n1497), .Z(n1684) );
  NANDN U2257 ( .A(n1498), .B(creg[61]), .Z(n1683) );
  NAND U2258 ( .A(n1685), .B(n1119), .Z(n849) );
  NANDN U2259 ( .A(init), .B(m[62]), .Z(n1119) );
  AND U2260 ( .A(n1686), .B(n1687), .Z(n1685) );
  NAND U2261 ( .A(o[62]), .B(n1497), .Z(n1687) );
  ANDN U2262 ( .B(n1498), .A(n1492), .Z(n1497) );
  NANDN U2263 ( .A(n1498), .B(creg[62]), .Z(n1686) );
  NAND U2264 ( .A(init), .B(n1688), .Z(n1498) );
  NAND U2265 ( .A(first_one), .B(n1689), .Z(n1688) );
  AND U2266 ( .A(n1690), .B(n1825), .Z(n1689) );
  NAND U2267 ( .A(n1691), .B(mul_pow), .Z(n1690) );
  NANDN U2268 ( .A(first_one), .B(n1692), .Z(n848) );
  NAND U2269 ( .A(n1693), .B(ereg[63]), .Z(n1692) );
  AND U2270 ( .A(mul_pow), .B(n1825), .Z(n1693) );
  IV U2271 ( .A(n1492), .Z(n1825) );
  NAND U2272 ( .A(start_reg[63]), .B(init), .Z(n1492) );
  NAND U2273 ( .A(n1694), .B(n1695), .Z(c[9]) );
  NAND U2274 ( .A(n1696), .B(o[9]), .Z(n1695) );
  NAND U2275 ( .A(n1691), .B(creg[9]), .Z(n1694) );
  NAND U2276 ( .A(n1697), .B(n1698), .Z(c[8]) );
  NAND U2277 ( .A(n1696), .B(o[8]), .Z(n1698) );
  NAND U2278 ( .A(n1691), .B(creg[8]), .Z(n1697) );
  NAND U2279 ( .A(n1699), .B(n1700), .Z(c[7]) );
  NAND U2280 ( .A(n1696), .B(o[7]), .Z(n1700) );
  NAND U2281 ( .A(n1691), .B(creg[7]), .Z(n1699) );
  NAND U2282 ( .A(n1701), .B(n1702), .Z(c[6]) );
  NAND U2283 ( .A(n1696), .B(o[6]), .Z(n1702) );
  NAND U2284 ( .A(n1691), .B(creg[6]), .Z(n1701) );
  NAND U2285 ( .A(n1703), .B(n1704), .Z(c[63]) );
  NAND U2286 ( .A(n1696), .B(o[63]), .Z(n1704) );
  NAND U2287 ( .A(n1691), .B(creg[63]), .Z(n1703) );
  NAND U2288 ( .A(n1705), .B(n1706), .Z(c[62]) );
  NAND U2289 ( .A(n1696), .B(o[62]), .Z(n1706) );
  NAND U2290 ( .A(n1691), .B(creg[62]), .Z(n1705) );
  NAND U2291 ( .A(n1707), .B(n1708), .Z(c[61]) );
  NAND U2292 ( .A(n1696), .B(o[61]), .Z(n1708) );
  NAND U2293 ( .A(n1691), .B(creg[61]), .Z(n1707) );
  NAND U2294 ( .A(n1709), .B(n1710), .Z(c[60]) );
  NAND U2295 ( .A(n1696), .B(o[60]), .Z(n1710) );
  NAND U2296 ( .A(n1691), .B(creg[60]), .Z(n1709) );
  NAND U2297 ( .A(n1711), .B(n1712), .Z(c[5]) );
  NAND U2298 ( .A(n1696), .B(o[5]), .Z(n1712) );
  NAND U2299 ( .A(n1691), .B(creg[5]), .Z(n1711) );
  NAND U2300 ( .A(n1713), .B(n1714), .Z(c[59]) );
  NAND U2301 ( .A(n1696), .B(o[59]), .Z(n1714) );
  NAND U2302 ( .A(n1691), .B(creg[59]), .Z(n1713) );
  NAND U2303 ( .A(n1715), .B(n1716), .Z(c[58]) );
  NAND U2304 ( .A(n1696), .B(o[58]), .Z(n1716) );
  NAND U2305 ( .A(n1691), .B(creg[58]), .Z(n1715) );
  NAND U2306 ( .A(n1717), .B(n1718), .Z(c[57]) );
  NAND U2307 ( .A(n1696), .B(o[57]), .Z(n1718) );
  NAND U2308 ( .A(n1691), .B(creg[57]), .Z(n1717) );
  NAND U2309 ( .A(n1719), .B(n1720), .Z(c[56]) );
  NAND U2310 ( .A(n1696), .B(o[56]), .Z(n1720) );
  NAND U2311 ( .A(n1691), .B(creg[56]), .Z(n1719) );
  NAND U2312 ( .A(n1721), .B(n1722), .Z(c[55]) );
  NAND U2313 ( .A(n1696), .B(o[55]), .Z(n1722) );
  NAND U2314 ( .A(n1691), .B(creg[55]), .Z(n1721) );
  NAND U2315 ( .A(n1723), .B(n1724), .Z(c[54]) );
  NAND U2316 ( .A(n1696), .B(o[54]), .Z(n1724) );
  NAND U2317 ( .A(n1691), .B(creg[54]), .Z(n1723) );
  NAND U2318 ( .A(n1725), .B(n1726), .Z(c[53]) );
  NAND U2319 ( .A(n1696), .B(o[53]), .Z(n1726) );
  NAND U2320 ( .A(n1691), .B(creg[53]), .Z(n1725) );
  NAND U2321 ( .A(n1727), .B(n1728), .Z(c[52]) );
  NAND U2322 ( .A(n1696), .B(o[52]), .Z(n1728) );
  NAND U2323 ( .A(n1691), .B(creg[52]), .Z(n1727) );
  NAND U2324 ( .A(n1729), .B(n1730), .Z(c[51]) );
  NAND U2325 ( .A(n1696), .B(o[51]), .Z(n1730) );
  NAND U2326 ( .A(n1691), .B(creg[51]), .Z(n1729) );
  NAND U2327 ( .A(n1731), .B(n1732), .Z(c[50]) );
  NAND U2328 ( .A(n1696), .B(o[50]), .Z(n1732) );
  NAND U2329 ( .A(n1691), .B(creg[50]), .Z(n1731) );
  NAND U2330 ( .A(n1733), .B(n1734), .Z(c[4]) );
  NAND U2331 ( .A(n1696), .B(o[4]), .Z(n1734) );
  NAND U2332 ( .A(n1691), .B(creg[4]), .Z(n1733) );
  NAND U2333 ( .A(n1735), .B(n1736), .Z(c[49]) );
  NAND U2334 ( .A(n1696), .B(o[49]), .Z(n1736) );
  NAND U2335 ( .A(n1691), .B(creg[49]), .Z(n1735) );
  NAND U2336 ( .A(n1737), .B(n1738), .Z(c[48]) );
  NAND U2337 ( .A(n1696), .B(o[48]), .Z(n1738) );
  NAND U2338 ( .A(n1691), .B(creg[48]), .Z(n1737) );
  NAND U2339 ( .A(n1739), .B(n1740), .Z(c[47]) );
  NAND U2340 ( .A(n1696), .B(o[47]), .Z(n1740) );
  NAND U2341 ( .A(n1691), .B(creg[47]), .Z(n1739) );
  NAND U2342 ( .A(n1741), .B(n1742), .Z(c[46]) );
  NAND U2343 ( .A(n1696), .B(o[46]), .Z(n1742) );
  NAND U2344 ( .A(n1691), .B(creg[46]), .Z(n1741) );
  NAND U2345 ( .A(n1743), .B(n1744), .Z(c[45]) );
  NAND U2346 ( .A(n1696), .B(o[45]), .Z(n1744) );
  NAND U2347 ( .A(n1691), .B(creg[45]), .Z(n1743) );
  NAND U2348 ( .A(n1745), .B(n1746), .Z(c[44]) );
  NAND U2349 ( .A(n1696), .B(o[44]), .Z(n1746) );
  NAND U2350 ( .A(n1691), .B(creg[44]), .Z(n1745) );
  NAND U2351 ( .A(n1747), .B(n1748), .Z(c[43]) );
  NAND U2352 ( .A(n1696), .B(o[43]), .Z(n1748) );
  NAND U2353 ( .A(n1691), .B(creg[43]), .Z(n1747) );
  NAND U2354 ( .A(n1749), .B(n1750), .Z(c[42]) );
  NAND U2355 ( .A(n1696), .B(o[42]), .Z(n1750) );
  NAND U2356 ( .A(n1691), .B(creg[42]), .Z(n1749) );
  NAND U2357 ( .A(n1751), .B(n1752), .Z(c[41]) );
  NAND U2358 ( .A(n1696), .B(o[41]), .Z(n1752) );
  NAND U2359 ( .A(n1691), .B(creg[41]), .Z(n1751) );
  NAND U2360 ( .A(n1753), .B(n1754), .Z(c[40]) );
  NAND U2361 ( .A(n1696), .B(o[40]), .Z(n1754) );
  NAND U2362 ( .A(n1691), .B(creg[40]), .Z(n1753) );
  NAND U2363 ( .A(n1755), .B(n1756), .Z(c[3]) );
  NAND U2364 ( .A(n1696), .B(o[3]), .Z(n1756) );
  NAND U2365 ( .A(n1691), .B(creg[3]), .Z(n1755) );
  NAND U2366 ( .A(n1757), .B(n1758), .Z(c[39]) );
  NAND U2367 ( .A(n1696), .B(o[39]), .Z(n1758) );
  NAND U2368 ( .A(n1691), .B(creg[39]), .Z(n1757) );
  NAND U2369 ( .A(n1759), .B(n1760), .Z(c[38]) );
  NAND U2370 ( .A(n1696), .B(o[38]), .Z(n1760) );
  NAND U2371 ( .A(n1691), .B(creg[38]), .Z(n1759) );
  NAND U2372 ( .A(n1761), .B(n1762), .Z(c[37]) );
  NAND U2373 ( .A(n1696), .B(o[37]), .Z(n1762) );
  NAND U2374 ( .A(n1691), .B(creg[37]), .Z(n1761) );
  NAND U2375 ( .A(n1763), .B(n1764), .Z(c[36]) );
  NAND U2376 ( .A(n1696), .B(o[36]), .Z(n1764) );
  NAND U2377 ( .A(n1691), .B(creg[36]), .Z(n1763) );
  NAND U2378 ( .A(n1765), .B(n1766), .Z(c[35]) );
  NAND U2379 ( .A(n1696), .B(o[35]), .Z(n1766) );
  NAND U2380 ( .A(n1691), .B(creg[35]), .Z(n1765) );
  NAND U2381 ( .A(n1767), .B(n1768), .Z(c[34]) );
  NAND U2382 ( .A(n1696), .B(o[34]), .Z(n1768) );
  NAND U2383 ( .A(n1691), .B(creg[34]), .Z(n1767) );
  NAND U2384 ( .A(n1769), .B(n1770), .Z(c[33]) );
  NAND U2385 ( .A(n1696), .B(o[33]), .Z(n1770) );
  NAND U2386 ( .A(n1691), .B(creg[33]), .Z(n1769) );
  NAND U2387 ( .A(n1771), .B(n1772), .Z(c[32]) );
  NAND U2388 ( .A(n1696), .B(o[32]), .Z(n1772) );
  NAND U2389 ( .A(n1691), .B(creg[32]), .Z(n1771) );
  NAND U2390 ( .A(n1773), .B(n1774), .Z(c[31]) );
  NAND U2391 ( .A(n1696), .B(o[31]), .Z(n1774) );
  NAND U2392 ( .A(n1691), .B(creg[31]), .Z(n1773) );
  NAND U2393 ( .A(n1775), .B(n1776), .Z(c[30]) );
  NAND U2394 ( .A(n1696), .B(o[30]), .Z(n1776) );
  NAND U2395 ( .A(n1691), .B(creg[30]), .Z(n1775) );
  NAND U2396 ( .A(n1777), .B(n1778), .Z(c[2]) );
  NAND U2397 ( .A(n1696), .B(o[2]), .Z(n1778) );
  NAND U2398 ( .A(n1691), .B(creg[2]), .Z(n1777) );
  NAND U2399 ( .A(n1779), .B(n1780), .Z(c[29]) );
  NAND U2400 ( .A(n1696), .B(o[29]), .Z(n1780) );
  NAND U2401 ( .A(n1691), .B(creg[29]), .Z(n1779) );
  NAND U2402 ( .A(n1781), .B(n1782), .Z(c[28]) );
  NAND U2403 ( .A(n1696), .B(o[28]), .Z(n1782) );
  NAND U2404 ( .A(n1691), .B(creg[28]), .Z(n1781) );
  NAND U2405 ( .A(n1783), .B(n1784), .Z(c[27]) );
  NAND U2406 ( .A(n1696), .B(o[27]), .Z(n1784) );
  NAND U2407 ( .A(n1691), .B(creg[27]), .Z(n1783) );
  NAND U2408 ( .A(n1785), .B(n1786), .Z(c[26]) );
  NAND U2409 ( .A(n1696), .B(o[26]), .Z(n1786) );
  NAND U2410 ( .A(n1691), .B(creg[26]), .Z(n1785) );
  NAND U2411 ( .A(n1787), .B(n1788), .Z(c[25]) );
  NAND U2412 ( .A(n1696), .B(o[25]), .Z(n1788) );
  NAND U2413 ( .A(n1691), .B(creg[25]), .Z(n1787) );
  NAND U2414 ( .A(n1789), .B(n1790), .Z(c[24]) );
  NAND U2415 ( .A(n1696), .B(o[24]), .Z(n1790) );
  NAND U2416 ( .A(n1691), .B(creg[24]), .Z(n1789) );
  NAND U2417 ( .A(n1791), .B(n1792), .Z(c[23]) );
  NAND U2418 ( .A(n1696), .B(o[23]), .Z(n1792) );
  NAND U2419 ( .A(n1691), .B(creg[23]), .Z(n1791) );
  NAND U2420 ( .A(n1793), .B(n1794), .Z(c[22]) );
  NAND U2421 ( .A(n1696), .B(o[22]), .Z(n1794) );
  NAND U2422 ( .A(n1691), .B(creg[22]), .Z(n1793) );
  NAND U2423 ( .A(n1795), .B(n1796), .Z(c[21]) );
  NAND U2424 ( .A(n1696), .B(o[21]), .Z(n1796) );
  NAND U2425 ( .A(n1691), .B(creg[21]), .Z(n1795) );
  NAND U2426 ( .A(n1797), .B(n1798), .Z(c[20]) );
  NAND U2427 ( .A(n1696), .B(o[20]), .Z(n1798) );
  NAND U2428 ( .A(n1691), .B(creg[20]), .Z(n1797) );
  NAND U2429 ( .A(n1799), .B(n1800), .Z(c[1]) );
  NAND U2430 ( .A(n1696), .B(o[1]), .Z(n1800) );
  NAND U2431 ( .A(n1691), .B(creg[1]), .Z(n1799) );
  NAND U2432 ( .A(n1801), .B(n1802), .Z(c[19]) );
  NAND U2433 ( .A(n1696), .B(o[19]), .Z(n1802) );
  NAND U2434 ( .A(n1691), .B(creg[19]), .Z(n1801) );
  NAND U2435 ( .A(n1803), .B(n1804), .Z(c[18]) );
  NAND U2436 ( .A(n1696), .B(o[18]), .Z(n1804) );
  NAND U2437 ( .A(n1691), .B(creg[18]), .Z(n1803) );
  NAND U2438 ( .A(n1805), .B(n1806), .Z(c[17]) );
  NAND U2439 ( .A(n1696), .B(o[17]), .Z(n1806) );
  NAND U2440 ( .A(n1691), .B(creg[17]), .Z(n1805) );
  NAND U2441 ( .A(n1807), .B(n1808), .Z(c[16]) );
  NAND U2442 ( .A(n1696), .B(o[16]), .Z(n1808) );
  NAND U2443 ( .A(n1691), .B(creg[16]), .Z(n1807) );
  NAND U2444 ( .A(n1809), .B(n1810), .Z(c[15]) );
  NAND U2445 ( .A(n1696), .B(o[15]), .Z(n1810) );
  NAND U2446 ( .A(n1691), .B(creg[15]), .Z(n1809) );
  NAND U2447 ( .A(n1811), .B(n1812), .Z(c[14]) );
  NAND U2448 ( .A(n1696), .B(o[14]), .Z(n1812) );
  NAND U2449 ( .A(n1691), .B(creg[14]), .Z(n1811) );
  NAND U2450 ( .A(n1813), .B(n1814), .Z(c[13]) );
  NAND U2451 ( .A(n1696), .B(o[13]), .Z(n1814) );
  NAND U2452 ( .A(n1691), .B(creg[13]), .Z(n1813) );
  NAND U2453 ( .A(n1815), .B(n1816), .Z(c[12]) );
  NAND U2454 ( .A(n1696), .B(o[12]), .Z(n1816) );
  NAND U2455 ( .A(n1691), .B(creg[12]), .Z(n1815) );
  NAND U2456 ( .A(n1817), .B(n1818), .Z(c[11]) );
  NAND U2457 ( .A(n1696), .B(o[11]), .Z(n1818) );
  NAND U2458 ( .A(n1691), .B(creg[11]), .Z(n1817) );
  NAND U2459 ( .A(n1819), .B(n1820), .Z(c[10]) );
  NAND U2460 ( .A(n1696), .B(o[10]), .Z(n1820) );
  NAND U2461 ( .A(n1691), .B(creg[10]), .Z(n1819) );
  NAND U2462 ( .A(n1821), .B(n1822), .Z(c[0]) );
  NAND U2463 ( .A(n1696), .B(o[0]), .Z(n1822) );
  IV U2464 ( .A(n1691), .Z(n1696) );
  NAND U2465 ( .A(n1691), .B(creg[0]), .Z(n1821) );
  NAND U2466 ( .A(n1823), .B(n1824), .Z(n1691) );
  NANDN U2467 ( .A(ereg[63]), .B(init), .Z(n1824) );
  OR U2468 ( .A(init), .B(e[63]), .Z(n1823) );
endmodule

