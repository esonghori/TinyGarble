
module SubBytes_7 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n339), .B(n328), .Z(n341) );
  XOR U2963 ( .A(n493), .B(n494), .Z(n646) );
  XNOR U2964 ( .A(n170), .B(n162), .Z(n143) );
  IV U2965 ( .A(x[1]), .Z(n1447) );
  XOR U2966 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2967 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2968 ( .A(n1446), .Z(n3) );
  AND U2969 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2970 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2971 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2972 ( .A(n2), .B(n1), .Z(n66) );
  IV U2973 ( .A(n66), .Z(n12) );
  XNOR U2974 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2975 ( .A(x[7]), .Z(n4) );
  XNOR U2976 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2977 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2978 ( .A(n4), .B(n3), .Z(n11) );
  IV U2979 ( .A(n11), .Z(n1083) );
  XOR U2980 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2981 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2982 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2983 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2984 ( .A(n5), .Z(n790) );
  NANDN U2985 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2986 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2987 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2988 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2989 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2990 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2991 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2992 ( .A(n10), .B(n9), .Z(n46) );
  IV U2993 ( .A(n46), .Z(n52) );
  AND U2994 ( .A(n12), .B(n11), .Z(n17) );
  XOR U2995 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U2996 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U2997 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U2998 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U2999 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3000 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3001 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3002 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3003 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3004 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3005 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3006 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3007 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3008 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3009 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3010 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3011 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3012 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3013 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3014 ( .A(n52), .B(n25), .Z(n36) );
  IV U3015 ( .A(n42), .Z(n43) );
  IV U3016 ( .A(n44), .Z(n50) );
  XOR U3017 ( .A(n26), .B(n800), .Z(n29) );
  AND U3018 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3019 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3020 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3021 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3022 ( .A(n33), .B(n32), .Z(n54) );
  IV U3023 ( .A(n54), .Z(n49) );
  XOR U3024 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3025 ( .A(n43), .B(n34), .Z(n35) );
  AND U3026 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3027 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3028 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3029 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3030 ( .A(n44), .B(n38), .Z(n39) );
  AND U3031 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3032 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3033 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3034 ( .A(n52), .B(n42), .Z(n48) );
  AND U3035 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3036 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3037 ( .A(n46), .B(n45), .Z(n47) );
  AND U3038 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3039 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3040 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3041 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3042 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3043 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3044 ( .A(n806), .B(n791), .Z(n793) );
  OR U3045 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3046 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3047 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3048 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3049 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3050 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3051 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3052 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3053 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3054 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3055 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3056 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3057 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3058 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3059 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3060 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3061 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3062 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3063 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3064 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3065 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3066 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3067 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3068 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3069 ( .A(n70), .Z(n142) );
  NANDN U3070 ( .A(n128), .B(n142), .Z(n80) );
  IV U3071 ( .A(n135), .Z(n91) );
  XNOR U3072 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3073 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3074 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3075 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3076 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3077 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3078 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3079 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3080 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3081 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3082 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3083 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3084 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3085 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3086 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3087 ( .A(n78), .B(n77), .Z(n115) );
  IV U3088 ( .A(n115), .Z(n108) );
  XNOR U3089 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3090 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3091 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3092 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3093 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3094 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3095 ( .A(n81), .B(n171), .Z(n84) );
  AND U3096 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3097 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3098 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3099 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3100 ( .A(n94), .B(n86), .Z(n118) );
  AND U3101 ( .A(n129), .B(n161), .Z(n89) );
  IV U3102 ( .A(x[97]), .Z(n136) );
  XNOR U3103 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3104 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3105 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3106 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3107 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3108 ( .A(n108), .B(n90), .Z(n99) );
  IV U3109 ( .A(n118), .Z(n102) );
  NAND U3110 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3111 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3112 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3113 ( .A(n97), .B(n96), .Z(n114) );
  IV U3114 ( .A(n107), .Z(n116) );
  XOR U3115 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3116 ( .A(n102), .B(n111), .Z(n98) );
  AND U3117 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3118 ( .A(n118), .B(n108), .Z(n104) );
  AND U3119 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3120 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3121 ( .A(n102), .B(n101), .Z(n103) );
  AND U3122 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3123 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3124 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3125 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3126 ( .A(n131), .B(n106), .Z(n173) );
  IV U3127 ( .A(n114), .Z(n120) );
  NAND U3128 ( .A(n120), .B(n107), .Z(n113) );
  AND U3129 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3130 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3131 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3132 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3133 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3134 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3135 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3136 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3137 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3138 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3139 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3140 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3141 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3142 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3143 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3144 ( .B(n163), .A(n126), .Z(n184) );
  IV U3145 ( .A(n127), .Z(n162) );
  OR U3146 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3147 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3148 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3149 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3150 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3151 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3152 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3153 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3154 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3155 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3156 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3157 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3158 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3159 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3160 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3161 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3162 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3163 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3164 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3165 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3166 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3167 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3168 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3169 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3170 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3171 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3172 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3173 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3174 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3175 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3176 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3177 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3178 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3179 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3180 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3181 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3182 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3183 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3184 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3185 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3186 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3187 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3188 ( .A(x[105]), .Z(n292) );
  XOR U3189 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3190 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3191 ( .A(n291), .Z(n188) );
  AND U3192 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3193 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3194 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3195 ( .A(n187), .B(n186), .Z(n251) );
  IV U3196 ( .A(n251), .Z(n197) );
  XNOR U3197 ( .A(n197), .B(n291), .Z(n250) );
  IV U3198 ( .A(x[111]), .Z(n189) );
  XNOR U3199 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3200 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3201 ( .A(n189), .B(n188), .Z(n196) );
  IV U3202 ( .A(n196), .Z(n280) );
  XOR U3203 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3204 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3205 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3206 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3207 ( .A(n190), .Z(n255) );
  NANDN U3208 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3209 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3210 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3211 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3212 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3213 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3214 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3215 ( .A(n195), .B(n194), .Z(n231) );
  IV U3216 ( .A(n231), .Z(n237) );
  AND U3217 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3218 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3219 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3220 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3221 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3222 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3223 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3224 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3225 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3226 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3227 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3228 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3229 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3230 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3231 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3232 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3233 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3234 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3235 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3236 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3237 ( .A(n237), .B(n210), .Z(n221) );
  IV U3238 ( .A(n227), .Z(n228) );
  IV U3239 ( .A(n229), .Z(n235) );
  XOR U3240 ( .A(n211), .B(n265), .Z(n214) );
  AND U3241 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3242 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3243 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3244 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3245 ( .A(n218), .B(n217), .Z(n239) );
  IV U3246 ( .A(n239), .Z(n234) );
  XOR U3247 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3248 ( .A(n228), .B(n219), .Z(n220) );
  AND U3249 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3250 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3251 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3252 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3253 ( .A(n229), .B(n223), .Z(n224) );
  AND U3254 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3255 ( .A(n299), .B(n281), .Z(n256) );
  OR U3256 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3257 ( .A(n237), .B(n227), .Z(n233) );
  AND U3258 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3259 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3260 ( .A(n231), .B(n230), .Z(n232) );
  AND U3261 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3262 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3263 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3264 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3265 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3266 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3267 ( .A(n271), .B(n256), .Z(n258) );
  OR U3268 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3269 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3270 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3271 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3272 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3273 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3274 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3275 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3276 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3277 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3278 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3279 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3280 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3281 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3282 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3283 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3284 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3285 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3286 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3287 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3288 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3289 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3290 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3291 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3292 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3293 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3294 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3295 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3296 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3297 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3298 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3299 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3300 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3301 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3302 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3303 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3304 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3305 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3306 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3307 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3308 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3309 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3310 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3311 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3312 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3313 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3314 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3315 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3316 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3317 ( .A(x[15]), .Z(n311) );
  IV U3318 ( .A(x[10]), .Z(n315) );
  XOR U3319 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3320 ( .A(n315), .B(n307), .Z(n352) );
  IV U3321 ( .A(n352), .Z(n309) );
  XOR U3322 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3323 ( .A(x[9]), .Z(n655) );
  XNOR U3324 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3325 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3326 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3327 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3328 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3329 ( .A(n314), .B(n497), .Z(n318) );
  IV U3330 ( .A(x[13]), .Z(n353) );
  XOR U3331 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3332 ( .A(n353), .B(n310), .Z(n325) );
  IV U3333 ( .A(n325), .Z(n656) );
  XOR U3334 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3335 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3336 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3337 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3338 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3339 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3340 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3341 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3342 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3343 ( .A(n333), .B(n312), .Z(n328) );
  IV U3344 ( .A(n313), .Z(n647) );
  IV U3345 ( .A(n314), .Z(n507) );
  XNOR U3346 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3347 ( .A(n507), .B(n321), .Z(n501) );
  IV U3348 ( .A(n316), .Z(n344) );
  NANDN U3349 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3350 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3351 ( .A(n648), .B(n497), .Z(n498) );
  OR U3352 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3353 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3354 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3355 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3356 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3357 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3358 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3359 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3360 ( .A(n647), .B(n324), .Z(n356) );
  IV U3361 ( .A(n356), .Z(n359) );
  NAND U3362 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3363 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3364 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3365 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3366 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3367 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3368 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3369 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3370 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3371 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3372 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3373 ( .A(n348), .B(n358), .Z(n336) );
  AND U3374 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3375 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3376 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3377 ( .A(n342), .B(n340), .Z(n354) );
  OR U3378 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3379 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3380 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3381 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3382 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3383 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3384 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3385 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3386 ( .A(n347), .B(n346), .Z(n361) );
  OR U3387 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3388 ( .A(n496), .B(n349), .Z(n504) );
  AND U3389 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3390 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3391 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3392 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3393 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3394 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3395 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3396 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3397 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3398 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3399 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3400 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3401 ( .A(n670), .B(n519), .Z(n654) );
  IV U3402 ( .A(n654), .Z(z[10]) );
  XNOR U3403 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3404 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3405 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3406 ( .A(x[113]), .Z(n475) );
  XOR U3407 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3408 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3409 ( .A(n474), .Z(n371) );
  AND U3410 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3411 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3412 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3413 ( .A(n370), .B(n369), .Z(n434) );
  IV U3414 ( .A(n434), .Z(n380) );
  XNOR U3415 ( .A(n380), .B(n474), .Z(n433) );
  IV U3416 ( .A(x[119]), .Z(n372) );
  XNOR U3417 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3418 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3419 ( .A(n372), .B(n371), .Z(n379) );
  IV U3420 ( .A(n379), .Z(n463) );
  XOR U3421 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3422 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3423 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3424 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3425 ( .A(n373), .Z(n438) );
  NANDN U3426 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3427 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3428 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3429 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3430 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3431 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3432 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3433 ( .A(n378), .B(n377), .Z(n414) );
  IV U3434 ( .A(n414), .Z(n420) );
  AND U3435 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3436 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3437 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3438 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3439 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3440 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3441 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3442 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3443 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3444 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3445 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3446 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3447 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3448 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3449 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3450 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3451 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3452 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3453 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3454 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3455 ( .A(n420), .B(n393), .Z(n404) );
  IV U3456 ( .A(n410), .Z(n411) );
  IV U3457 ( .A(n412), .Z(n418) );
  XOR U3458 ( .A(n394), .B(n448), .Z(n397) );
  AND U3459 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3460 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3461 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3462 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3463 ( .A(n401), .B(n400), .Z(n422) );
  IV U3464 ( .A(n422), .Z(n417) );
  XOR U3465 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3466 ( .A(n411), .B(n402), .Z(n403) );
  AND U3467 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3468 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3469 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3470 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3471 ( .A(n412), .B(n406), .Z(n407) );
  AND U3472 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3473 ( .A(n482), .B(n464), .Z(n439) );
  OR U3474 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3475 ( .A(n420), .B(n410), .Z(n416) );
  AND U3476 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3477 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3478 ( .A(n414), .B(n413), .Z(n415) );
  AND U3479 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3480 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3481 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3482 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3483 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3484 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3485 ( .A(n454), .B(n439), .Z(n441) );
  OR U3486 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3487 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3488 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3489 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3490 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3491 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3492 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3493 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3494 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3495 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3496 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3497 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3498 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3499 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3500 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3501 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3502 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3503 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3504 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3505 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3506 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3507 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3508 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3509 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3510 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3511 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3512 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3513 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3514 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3515 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3516 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3517 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3518 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3519 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3520 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3521 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3522 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3523 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3524 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3525 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3526 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3527 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3528 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3529 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3530 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3531 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3532 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3533 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3534 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3535 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3536 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3537 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3538 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3539 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3540 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3541 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3542 ( .A(n506), .B(n672), .Z(n509) );
  OR U3543 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3544 ( .A(n650), .B(n499), .Z(n671) );
  OR U3545 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3546 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3547 ( .A(n511), .B(n503), .Z(n678) );
  AND U3548 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3549 ( .A(n507), .B(n506), .Z(n675) );
  OR U3550 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3551 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3552 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3553 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3554 ( .A(n515), .B(n514), .Z(n660) );
  OR U3555 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3556 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3557 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3558 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3559 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3560 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3561 ( .A(x[121]), .Z(n628) );
  XOR U3562 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3563 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3564 ( .A(n627), .Z(n524) );
  AND U3565 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3566 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3567 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3568 ( .A(n523), .B(n522), .Z(n587) );
  IV U3569 ( .A(n587), .Z(n533) );
  XNOR U3570 ( .A(n533), .B(n627), .Z(n586) );
  IV U3571 ( .A(x[127]), .Z(n525) );
  XNOR U3572 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3573 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3574 ( .A(n525), .B(n524), .Z(n532) );
  IV U3575 ( .A(n532), .Z(n616) );
  XOR U3576 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3577 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3578 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3579 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3580 ( .A(n526), .Z(n591) );
  NANDN U3581 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3582 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3583 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3584 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3585 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3586 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3587 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3588 ( .A(n531), .B(n530), .Z(n567) );
  IV U3589 ( .A(n567), .Z(n573) );
  AND U3590 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3591 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3592 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3593 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3594 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3595 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3596 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3597 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3598 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3599 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3600 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3601 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3602 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3603 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3604 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3605 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3606 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3607 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3608 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3609 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3610 ( .A(n573), .B(n546), .Z(n557) );
  IV U3611 ( .A(n563), .Z(n564) );
  IV U3612 ( .A(n565), .Z(n571) );
  XOR U3613 ( .A(n547), .B(n601), .Z(n550) );
  AND U3614 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3615 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3616 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3617 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3618 ( .A(n554), .B(n553), .Z(n575) );
  IV U3619 ( .A(n575), .Z(n570) );
  XOR U3620 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3621 ( .A(n564), .B(n555), .Z(n556) );
  AND U3622 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3623 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3624 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3625 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3626 ( .A(n565), .B(n559), .Z(n560) );
  AND U3627 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3628 ( .A(n635), .B(n617), .Z(n592) );
  OR U3629 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3630 ( .A(n573), .B(n563), .Z(n569) );
  AND U3631 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3632 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3633 ( .A(n567), .B(n566), .Z(n568) );
  AND U3634 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3635 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3636 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3637 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3638 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3639 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3640 ( .A(n607), .B(n592), .Z(n594) );
  OR U3641 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3642 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3643 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3644 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3645 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3646 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3647 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3648 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3649 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3650 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3651 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3652 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3653 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3654 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3655 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3656 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3657 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3658 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3659 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3660 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3661 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3662 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3663 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3664 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3665 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3666 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3667 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3668 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3669 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3670 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3671 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3672 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3673 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3674 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3675 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3676 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3677 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3678 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3679 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3680 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3681 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3682 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3683 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3684 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3685 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3686 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3687 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3688 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3689 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3690 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3691 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3692 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3693 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3694 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3695 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3696 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3697 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3698 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3699 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3700 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3701 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3702 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3703 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3704 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3705 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3706 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3707 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3708 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3709 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3710 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3711 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3712 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3713 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3714 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3715 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3716 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3717 ( .A(x[17]), .Z(n815) );
  XOR U3718 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U3719 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U3720 ( .A(n814), .Z(n686) );
  AND U3721 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3722 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3723 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3724 ( .A(n685), .B(n684), .Z(n749) );
  IV U3725 ( .A(n749), .Z(n695) );
  XNOR U3726 ( .A(n695), .B(n814), .Z(n748) );
  IV U3727 ( .A(x[23]), .Z(n687) );
  XNOR U3728 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3729 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3730 ( .A(n687), .B(n686), .Z(n694) );
  IV U3731 ( .A(n694), .Z(n778) );
  XOR U3732 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3733 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3734 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3735 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3736 ( .A(n688), .Z(n753) );
  NANDN U3737 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3738 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3739 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3740 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3741 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3742 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3743 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3744 ( .A(n693), .B(n692), .Z(n729) );
  IV U3745 ( .A(n729), .Z(n735) );
  AND U3746 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3747 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3748 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3749 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3750 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3751 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3752 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3753 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3754 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3755 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3756 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3757 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3758 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3759 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3760 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3761 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3762 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3763 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3764 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3765 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3766 ( .A(n735), .B(n708), .Z(n719) );
  IV U3767 ( .A(n725), .Z(n726) );
  IV U3768 ( .A(n727), .Z(n733) );
  XOR U3769 ( .A(n709), .B(n763), .Z(n712) );
  AND U3770 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3771 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3772 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3773 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3774 ( .A(n716), .B(n715), .Z(n737) );
  IV U3775 ( .A(n737), .Z(n732) );
  XOR U3776 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3777 ( .A(n726), .B(n717), .Z(n718) );
  AND U3778 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3779 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3780 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3781 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3782 ( .A(n727), .B(n721), .Z(n722) );
  AND U3783 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3784 ( .A(n822), .B(n779), .Z(n754) );
  OR U3785 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3786 ( .A(n735), .B(n725), .Z(n731) );
  AND U3787 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3788 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3789 ( .A(n729), .B(n728), .Z(n730) );
  AND U3790 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3791 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3792 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3793 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3794 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3795 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3796 ( .A(n769), .B(n754), .Z(n756) );
  OR U3797 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3798 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3799 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3800 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3801 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3802 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3803 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3804 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3805 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3806 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3807 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3808 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3809 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3810 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3811 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3812 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3813 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3814 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3815 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3816 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3817 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3818 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3819 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3820 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3821 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3822 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3823 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3824 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3825 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3826 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3827 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3828 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3829 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3830 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3831 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3832 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3833 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3834 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3835 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3836 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3837 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3838 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3839 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3840 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3841 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3842 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3843 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3844 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3845 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3846 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3847 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3848 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3849 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3850 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3851 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3852 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3853 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3854 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3855 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3856 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3857 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3858 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3859 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3860 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3861 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3862 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3863 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3864 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3865 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3866 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3867 ( .A(x[25]), .Z(n939) );
  XOR U3868 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3869 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3870 ( .A(n938), .Z(n835) );
  AND U3871 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3872 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3873 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3874 ( .A(n834), .B(n833), .Z(n898) );
  IV U3875 ( .A(n898), .Z(n844) );
  XNOR U3876 ( .A(n844), .B(n938), .Z(n897) );
  IV U3877 ( .A(x[31]), .Z(n836) );
  XNOR U3878 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3879 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3880 ( .A(n836), .B(n835), .Z(n843) );
  IV U3881 ( .A(n843), .Z(n927) );
  XOR U3882 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3883 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3884 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3885 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3886 ( .A(n837), .Z(n902) );
  NANDN U3887 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3888 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3889 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3890 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3891 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3892 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3893 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3894 ( .A(n842), .B(n841), .Z(n878) );
  IV U3895 ( .A(n878), .Z(n884) );
  AND U3896 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3897 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3898 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3899 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3900 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3901 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3902 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3903 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3904 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3905 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3906 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3907 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3908 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3909 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3910 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3911 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3912 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3913 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3914 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3915 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3916 ( .A(n884), .B(n857), .Z(n868) );
  IV U3917 ( .A(n874), .Z(n875) );
  IV U3918 ( .A(n876), .Z(n882) );
  XOR U3919 ( .A(n858), .B(n912), .Z(n861) );
  AND U3920 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3921 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3922 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3923 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3924 ( .A(n865), .B(n864), .Z(n886) );
  IV U3925 ( .A(n886), .Z(n881) );
  XOR U3926 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3927 ( .A(n875), .B(n866), .Z(n867) );
  AND U3928 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3929 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3930 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3931 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3932 ( .A(n876), .B(n870), .Z(n871) );
  AND U3933 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3934 ( .A(n946), .B(n928), .Z(n903) );
  OR U3935 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3936 ( .A(n884), .B(n874), .Z(n880) );
  AND U3937 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3938 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3939 ( .A(n878), .B(n877), .Z(n879) );
  AND U3940 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3941 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3942 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3943 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3944 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3945 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3946 ( .A(n918), .B(n903), .Z(n905) );
  OR U3947 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3948 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3949 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3950 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3951 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3952 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3953 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3954 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3955 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3956 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3957 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3958 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3959 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3960 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3961 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3962 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3963 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3964 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3965 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3966 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3967 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3968 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3969 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3970 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3971 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3972 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3973 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3974 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3975 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3976 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3977 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3978 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3979 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3980 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3981 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3982 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3983 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3984 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3985 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3986 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3987 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3988 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3989 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3990 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3991 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3992 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3993 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3994 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3995 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3996 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3997 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U3998 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U3999 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4000 ( .A(x[33]), .Z(n1065) );
  XOR U4001 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4002 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4003 ( .A(n1064), .Z(n961) );
  AND U4004 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4005 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4006 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4007 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4008 ( .A(n1024), .Z(n970) );
  XNOR U4009 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4010 ( .A(x[39]), .Z(n962) );
  XNOR U4011 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4012 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4013 ( .A(n962), .B(n961), .Z(n969) );
  IV U4014 ( .A(n969), .Z(n1053) );
  XOR U4015 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4016 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4017 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4018 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4019 ( .A(n963), .Z(n1028) );
  NANDN U4020 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4021 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4022 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4023 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4024 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4025 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4026 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4027 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4028 ( .A(n1004), .Z(n1010) );
  AND U4029 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4030 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4031 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4032 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4033 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4034 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4035 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4036 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4037 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4038 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4039 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4040 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4041 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4042 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4043 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4044 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4045 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4046 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4047 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4048 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4049 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4050 ( .A(n1000), .Z(n1001) );
  IV U4051 ( .A(n1002), .Z(n1008) );
  XOR U4052 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4053 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4054 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4055 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4056 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4057 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4058 ( .A(n1012), .Z(n1007) );
  XOR U4059 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4060 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4061 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4062 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4063 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4064 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4065 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4066 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4067 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4068 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4069 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4070 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4071 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4072 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4073 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4074 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4075 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4076 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4077 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4078 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4079 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4080 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4081 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4082 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4083 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4084 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4085 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4086 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4087 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4088 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4089 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4090 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4091 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4092 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4093 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4094 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4095 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4096 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4097 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4098 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4099 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4100 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4101 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4102 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4103 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4104 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4105 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4106 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4107 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4108 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4109 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4110 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4111 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4112 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4113 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4114 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4115 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4116 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4117 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4118 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4119 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4120 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4121 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4122 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4123 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4124 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4125 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4126 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4127 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4128 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4129 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4130 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4131 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4132 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4133 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4134 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4135 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4136 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4137 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4138 ( .A(x[41]), .Z(n1199) );
  XOR U4139 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4140 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4141 ( .A(n1198), .Z(n1095) );
  AND U4142 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4143 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4144 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4145 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4146 ( .A(n1158), .Z(n1104) );
  XNOR U4147 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4148 ( .A(x[47]), .Z(n1096) );
  XNOR U4149 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4150 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4151 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4152 ( .A(n1103), .Z(n1187) );
  XOR U4153 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4154 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4155 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4156 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4157 ( .A(n1097), .Z(n1162) );
  NANDN U4158 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4159 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4160 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4161 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4162 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4163 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4164 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4165 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4166 ( .A(n1138), .Z(n1144) );
  AND U4167 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4168 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4169 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4170 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4171 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4172 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4173 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4174 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4175 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4176 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4177 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4178 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4179 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4180 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4181 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4182 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4183 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4184 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4185 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4186 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4187 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4188 ( .A(n1134), .Z(n1135) );
  IV U4189 ( .A(n1136), .Z(n1142) );
  XOR U4190 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4191 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4192 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4193 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4194 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4195 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4196 ( .A(n1146), .Z(n1141) );
  XOR U4197 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4198 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4199 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4200 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4201 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4202 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4203 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4204 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4205 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4206 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4207 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4208 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4209 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4210 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4211 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4212 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4213 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4214 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4215 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4216 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4217 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4218 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4219 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4220 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4221 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4222 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4223 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4224 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4225 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4226 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4227 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4228 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4229 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4230 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4231 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4232 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4233 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4234 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4235 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4236 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4237 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4238 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4239 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4240 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4241 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4242 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4243 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4244 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4245 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4246 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4247 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4248 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4249 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4250 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4251 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4252 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4253 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4254 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4255 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4256 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4257 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4258 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4259 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4260 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4261 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4262 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4263 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4264 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4265 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4266 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4267 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4268 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4269 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4270 ( .A(x[49]), .Z(n1324) );
  XOR U4271 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4272 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4273 ( .A(n1323), .Z(n1219) );
  AND U4274 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4275 ( .A(x[51]), .B(n1324), .Z(n1222) );
  XNOR U4276 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4277 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4278 ( .A(n1282), .Z(n1228) );
  XNOR U4279 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4280 ( .A(x[55]), .Z(n1220) );
  XNOR U4281 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4282 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4283 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4284 ( .A(n1227), .Z(n1312) );
  XOR U4285 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4286 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4287 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4288 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4289 ( .A(n1221), .Z(n1286) );
  NANDN U4290 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4291 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4292 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4293 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4294 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4295 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4296 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4297 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4298 ( .A(n1262), .Z(n1268) );
  AND U4299 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4300 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4301 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4302 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4303 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4304 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4305 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4306 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4307 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4308 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4309 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4310 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4311 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4312 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4313 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4314 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4315 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4316 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4317 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4318 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4319 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4320 ( .A(n1258), .Z(n1259) );
  IV U4321 ( .A(n1260), .Z(n1266) );
  XOR U4322 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4323 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4324 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4325 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4326 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4327 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4328 ( .A(n1270), .Z(n1265) );
  XOR U4329 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4330 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4331 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4332 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4333 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4334 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4335 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4336 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4337 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4338 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4339 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4340 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4341 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4342 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4343 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4344 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4345 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4346 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4347 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4348 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4349 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4350 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4351 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4352 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4353 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4354 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4355 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4356 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4357 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4358 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4359 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4360 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4361 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4362 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4363 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4364 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4365 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4366 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4367 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4368 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4369 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4370 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4371 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4372 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4373 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4374 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4375 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4376 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4377 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4378 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4379 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4380 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4381 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4382 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4383 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4384 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4385 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4386 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4387 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4388 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4389 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4390 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4391 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4392 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4393 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4394 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4395 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4396 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4397 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4398 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4399 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4400 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4401 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4402 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4403 ( .A(x[57]), .Z(n1462) );
  XOR U4404 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4405 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4406 ( .A(n1461), .Z(n1344) );
  AND U4407 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4408 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4409 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4410 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4411 ( .A(n1407), .Z(n1353) );
  XNOR U4412 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4413 ( .A(x[63]), .Z(n1345) );
  XNOR U4414 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4415 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4416 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4417 ( .A(n1352), .Z(n1436) );
  XOR U4418 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4419 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4420 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4421 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4422 ( .A(n1346), .Z(n1411) );
  NANDN U4423 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4424 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4425 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4426 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4427 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4428 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4429 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4430 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4431 ( .A(n1387), .Z(n1393) );
  AND U4432 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4433 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4434 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4435 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4436 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4437 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4438 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4439 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4440 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4441 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4442 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4443 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4444 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4445 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4446 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4447 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4448 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4449 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4450 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4451 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4452 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4453 ( .A(n1383), .Z(n1384) );
  IV U4454 ( .A(n1385), .Z(n1391) );
  XOR U4455 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4456 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4457 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4458 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4459 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4460 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4461 ( .A(n1395), .Z(n1390) );
  XOR U4462 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4463 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4464 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4465 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4466 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4467 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4468 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4469 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4470 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4471 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4472 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4473 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4474 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4475 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4476 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4477 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4478 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4479 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4480 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4481 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4482 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4483 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4484 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4485 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4486 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4487 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4488 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4489 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4490 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4491 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4492 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4493 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4494 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4495 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4496 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4497 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4498 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4499 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4500 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4501 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4502 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4503 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4504 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4505 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4506 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4507 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4508 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4509 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4510 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4511 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4512 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4513 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4514 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4515 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4516 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4517 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4518 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4519 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4520 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4521 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4522 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4523 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4524 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4525 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4526 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4527 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4528 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4529 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4530 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4531 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4532 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4533 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4534 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4535 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4536 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4537 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4538 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4539 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4540 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4541 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4542 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4543 ( .A(x[65]), .Z(n1586) );
  XOR U4544 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4545 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4546 ( .A(n1585), .Z(n1482) );
  AND U4547 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4548 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4549 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4550 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4551 ( .A(n1545), .Z(n1491) );
  XNOR U4552 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4553 ( .A(x[71]), .Z(n1483) );
  XNOR U4554 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4555 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4556 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4557 ( .A(n1490), .Z(n1574) );
  XOR U4558 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4559 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4560 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4561 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4562 ( .A(n1484), .Z(n1549) );
  NANDN U4563 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4564 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4565 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4566 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4567 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4568 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4569 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4570 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4571 ( .A(n1525), .Z(n1531) );
  AND U4572 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4573 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4574 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4575 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4576 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4577 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4578 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4579 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4580 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4581 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4582 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4583 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4584 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4585 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4586 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4587 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4588 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4589 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4590 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4591 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4592 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4593 ( .A(n1521), .Z(n1522) );
  IV U4594 ( .A(n1523), .Z(n1529) );
  XOR U4595 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4596 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4597 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4598 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4599 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4600 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4601 ( .A(n1533), .Z(n1528) );
  XOR U4602 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4603 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4604 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4605 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4606 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4607 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4608 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4609 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4610 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4611 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4612 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4613 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4614 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4615 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4616 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4617 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4618 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4619 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4620 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4621 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4622 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4623 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4624 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4625 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4626 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4627 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4628 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4629 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4630 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4631 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4632 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4633 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4634 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4635 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4636 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4637 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4638 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4639 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4640 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4641 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4642 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4643 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4644 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4645 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4646 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4647 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4648 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4649 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4650 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4651 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4652 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4653 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4654 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4655 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4656 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4657 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4658 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4659 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4660 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4661 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4662 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4663 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4664 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4665 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4666 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4667 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4668 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4669 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4670 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4671 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4672 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4673 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4674 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4675 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4676 ( .A(x[73]), .Z(n1712) );
  XOR U4677 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4678 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4679 ( .A(n1711), .Z(n1608) );
  AND U4680 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4681 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4682 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4683 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4684 ( .A(n1671), .Z(n1617) );
  XNOR U4685 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4686 ( .A(x[79]), .Z(n1609) );
  XNOR U4687 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4688 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4689 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4690 ( .A(n1616), .Z(n1700) );
  XOR U4691 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4692 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4693 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4694 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4695 ( .A(n1610), .Z(n1675) );
  NANDN U4696 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4697 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4698 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4699 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4700 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4701 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4702 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4703 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4704 ( .A(n1651), .Z(n1657) );
  AND U4705 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4706 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4707 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4708 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4709 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4710 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4711 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4712 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4713 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4714 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4715 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4716 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4717 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4718 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4719 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4720 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4721 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4722 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4723 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4724 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4725 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4726 ( .A(n1647), .Z(n1648) );
  IV U4727 ( .A(n1649), .Z(n1655) );
  XOR U4728 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4729 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4730 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4731 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4732 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4733 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4734 ( .A(n1659), .Z(n1654) );
  XOR U4735 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4736 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4737 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4738 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4739 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4740 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4741 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4742 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4743 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4744 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4745 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4746 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4747 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4748 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4749 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4750 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4751 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4752 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4753 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4754 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4755 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4756 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4757 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4758 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4759 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4760 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4761 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4762 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4763 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4764 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4765 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4766 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4767 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4768 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4769 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4770 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4771 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4772 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4773 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4774 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4775 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4776 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4777 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4778 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4779 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4780 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4781 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4782 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4783 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4784 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4785 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4786 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4787 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4788 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4789 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4790 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4791 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4792 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4793 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4794 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4795 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4796 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4797 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4798 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4799 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4800 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4801 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4802 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4803 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4804 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4805 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4806 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4807 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4808 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4809 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4810 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4811 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4812 ( .A(n1838), .Z(n1735) );
  IV U4813 ( .A(x[81]), .Z(n1837) );
  NAND U4814 ( .A(n1735), .B(n1837), .Z(n1742) );
  XOR U4815 ( .A(x[83]), .B(x[81]), .Z(n1738) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_8 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n815), .B(x[19]), .Z(n689) );
  XOR U2963 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U2964 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2965 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2966 ( .A(n475), .B(x[115]), .Z(n374) );
  XNOR U2967 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2968 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2969 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2970 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2971 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2972 ( .A(x[1]), .Z(n1447) );
  XOR U2973 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2974 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2975 ( .A(n1446), .Z(n3) );
  AND U2976 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2977 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2978 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2979 ( .A(n2), .B(n1), .Z(n66) );
  IV U2980 ( .A(n66), .Z(n12) );
  XNOR U2981 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2982 ( .A(x[7]), .Z(n4) );
  XNOR U2983 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2984 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2985 ( .A(n4), .B(n3), .Z(n11) );
  IV U2986 ( .A(n11), .Z(n1083) );
  XOR U2987 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2988 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2989 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2990 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2991 ( .A(n5), .Z(n790) );
  NANDN U2992 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2993 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2994 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2995 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2996 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2997 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2998 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2999 ( .A(n10), .B(n9), .Z(n46) );
  IV U3000 ( .A(n46), .Z(n52) );
  AND U3001 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3002 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3003 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3004 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3005 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3006 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3007 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3008 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3009 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3010 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3011 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3012 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3013 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3014 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3015 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3016 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3017 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3018 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3019 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3020 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3021 ( .A(n52), .B(n25), .Z(n36) );
  IV U3022 ( .A(n42), .Z(n43) );
  IV U3023 ( .A(n44), .Z(n50) );
  XOR U3024 ( .A(n26), .B(n800), .Z(n29) );
  AND U3025 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3026 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3027 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3028 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3029 ( .A(n33), .B(n32), .Z(n54) );
  IV U3030 ( .A(n54), .Z(n49) );
  XOR U3031 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3032 ( .A(n43), .B(n34), .Z(n35) );
  AND U3033 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3034 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3035 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3036 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3037 ( .A(n44), .B(n38), .Z(n39) );
  AND U3038 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3039 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3040 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3041 ( .A(n52), .B(n42), .Z(n48) );
  AND U3042 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3043 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3044 ( .A(n46), .B(n45), .Z(n47) );
  AND U3045 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3046 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3047 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3048 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3049 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3050 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3051 ( .A(n806), .B(n791), .Z(n793) );
  OR U3052 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3053 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3054 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3055 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3056 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3057 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3058 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3059 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3060 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3061 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3062 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3063 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3064 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3065 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3066 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3067 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3068 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3069 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3070 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3071 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3072 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3073 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3074 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3075 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3076 ( .A(n70), .Z(n142) );
  NANDN U3077 ( .A(n128), .B(n142), .Z(n80) );
  IV U3078 ( .A(n135), .Z(n91) );
  XNOR U3079 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3080 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3081 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3082 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3083 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3084 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3085 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3086 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3087 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3088 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3089 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3090 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3091 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3092 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3093 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3094 ( .A(n78), .B(n77), .Z(n115) );
  IV U3095 ( .A(n115), .Z(n108) );
  XNOR U3096 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3097 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3098 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3099 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3100 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3101 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3102 ( .A(n81), .B(n171), .Z(n84) );
  AND U3103 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3104 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3105 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3106 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3107 ( .A(n94), .B(n86), .Z(n118) );
  AND U3108 ( .A(n129), .B(n161), .Z(n89) );
  IV U3109 ( .A(x[97]), .Z(n136) );
  XNOR U3110 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3111 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3112 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3113 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3114 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3115 ( .A(n108), .B(n90), .Z(n99) );
  IV U3116 ( .A(n118), .Z(n102) );
  NAND U3117 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3118 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3119 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3120 ( .A(n97), .B(n96), .Z(n114) );
  IV U3121 ( .A(n107), .Z(n116) );
  XOR U3122 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3123 ( .A(n102), .B(n111), .Z(n98) );
  AND U3124 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3125 ( .A(n118), .B(n108), .Z(n104) );
  AND U3126 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3127 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3128 ( .A(n102), .B(n101), .Z(n103) );
  AND U3129 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3130 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3131 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3132 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3133 ( .A(n131), .B(n106), .Z(n173) );
  IV U3134 ( .A(n114), .Z(n120) );
  NAND U3135 ( .A(n120), .B(n107), .Z(n113) );
  AND U3136 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3137 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3138 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3139 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3140 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3141 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3142 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3143 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3144 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3145 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3146 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3147 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3148 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3149 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3150 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3151 ( .B(n163), .A(n126), .Z(n184) );
  IV U3152 ( .A(n127), .Z(n162) );
  OR U3153 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3154 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3155 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3156 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3157 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3158 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3159 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3160 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3161 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3162 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3163 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3164 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3165 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3166 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3167 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3168 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3169 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3170 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3171 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3172 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3173 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3174 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3175 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3176 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3177 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3178 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3179 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3180 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3181 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3182 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3183 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3184 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3185 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3186 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3187 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3188 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3189 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3190 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3191 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3192 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3193 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3194 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3195 ( .A(x[105]), .Z(n292) );
  XOR U3196 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3197 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3198 ( .A(n291), .Z(n188) );
  AND U3199 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3200 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3201 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3202 ( .A(n187), .B(n186), .Z(n251) );
  IV U3203 ( .A(n251), .Z(n197) );
  XNOR U3204 ( .A(n197), .B(n291), .Z(n250) );
  IV U3205 ( .A(x[111]), .Z(n189) );
  XNOR U3206 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3207 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3208 ( .A(n189), .B(n188), .Z(n196) );
  IV U3209 ( .A(n196), .Z(n280) );
  XOR U3210 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3211 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3212 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3213 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3214 ( .A(n190), .Z(n255) );
  NANDN U3215 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3216 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3217 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3218 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3219 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3220 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3221 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3222 ( .A(n195), .B(n194), .Z(n231) );
  IV U3223 ( .A(n231), .Z(n237) );
  AND U3224 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3225 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3226 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3227 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3228 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3229 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3230 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3231 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3232 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3233 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3234 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3235 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3236 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3237 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3238 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3239 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3240 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3241 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3242 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3243 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3244 ( .A(n237), .B(n210), .Z(n221) );
  IV U3245 ( .A(n227), .Z(n228) );
  IV U3246 ( .A(n229), .Z(n235) );
  XOR U3247 ( .A(n211), .B(n265), .Z(n214) );
  AND U3248 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3249 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3250 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3251 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3252 ( .A(n218), .B(n217), .Z(n239) );
  IV U3253 ( .A(n239), .Z(n234) );
  XOR U3254 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3255 ( .A(n228), .B(n219), .Z(n220) );
  AND U3256 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3257 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3258 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3259 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3260 ( .A(n229), .B(n223), .Z(n224) );
  AND U3261 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3262 ( .A(n299), .B(n281), .Z(n256) );
  OR U3263 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3264 ( .A(n237), .B(n227), .Z(n233) );
  AND U3265 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3266 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3267 ( .A(n231), .B(n230), .Z(n232) );
  AND U3268 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3269 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3270 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3271 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3272 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3273 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3274 ( .A(n271), .B(n256), .Z(n258) );
  OR U3275 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3276 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3277 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3278 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3279 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3280 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3281 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3282 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3283 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3284 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3285 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3286 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3287 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3288 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3289 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3290 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3291 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3292 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3293 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3294 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3295 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3296 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3297 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3298 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3299 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3300 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3301 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3302 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3303 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3304 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3305 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3306 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3307 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3308 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3309 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3310 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3311 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3312 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3313 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3314 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3315 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3316 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3317 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3318 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3319 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3320 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3321 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3322 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3323 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3324 ( .A(x[15]), .Z(n311) );
  IV U3325 ( .A(x[10]), .Z(n315) );
  XOR U3326 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3327 ( .A(n315), .B(n307), .Z(n352) );
  IV U3328 ( .A(n352), .Z(n309) );
  XOR U3329 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3330 ( .A(x[9]), .Z(n655) );
  XNOR U3331 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3332 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3333 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3334 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3335 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3336 ( .A(n314), .B(n497), .Z(n318) );
  IV U3337 ( .A(x[13]), .Z(n353) );
  XOR U3338 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3339 ( .A(n353), .B(n310), .Z(n325) );
  IV U3340 ( .A(n325), .Z(n656) );
  XOR U3341 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3342 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3343 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3344 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3345 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3346 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3347 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3348 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3349 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3350 ( .A(n333), .B(n312), .Z(n328) );
  IV U3351 ( .A(n313), .Z(n647) );
  IV U3352 ( .A(n314), .Z(n507) );
  XNOR U3353 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3354 ( .A(n507), .B(n321), .Z(n501) );
  IV U3355 ( .A(n316), .Z(n344) );
  NANDN U3356 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3357 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3358 ( .A(n648), .B(n497), .Z(n498) );
  OR U3359 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3360 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3361 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3362 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3363 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3364 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3365 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3366 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3367 ( .A(n647), .B(n324), .Z(n356) );
  IV U3368 ( .A(n356), .Z(n359) );
  NAND U3369 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3370 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3371 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3372 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3373 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3374 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3375 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3376 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3377 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3378 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3379 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3380 ( .A(n348), .B(n358), .Z(n336) );
  AND U3381 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3382 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3383 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3384 ( .A(n342), .B(n340), .Z(n354) );
  OR U3385 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3386 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3387 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3388 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3389 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3390 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3391 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3392 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3393 ( .A(n347), .B(n346), .Z(n361) );
  OR U3394 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3395 ( .A(n496), .B(n349), .Z(n504) );
  AND U3396 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3397 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3398 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3399 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3400 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3401 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3402 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3403 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3404 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3405 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3406 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3407 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3408 ( .A(n670), .B(n519), .Z(n654) );
  IV U3409 ( .A(n654), .Z(z[10]) );
  XNOR U3410 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3411 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3412 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3413 ( .A(x[113]), .Z(n475) );
  XOR U3414 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3415 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3416 ( .A(n474), .Z(n371) );
  AND U3417 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3418 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3419 ( .A(n370), .B(n369), .Z(n434) );
  IV U3420 ( .A(n434), .Z(n380) );
  XNOR U3421 ( .A(n380), .B(n474), .Z(n433) );
  IV U3422 ( .A(x[119]), .Z(n372) );
  XNOR U3423 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3424 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3425 ( .A(n372), .B(n371), .Z(n379) );
  IV U3426 ( .A(n379), .Z(n463) );
  XOR U3427 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3428 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3429 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3430 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3431 ( .A(n373), .Z(n438) );
  NANDN U3432 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3433 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3434 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3435 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3436 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3437 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3438 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3439 ( .A(n378), .B(n377), .Z(n414) );
  IV U3440 ( .A(n414), .Z(n420) );
  AND U3441 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3442 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3443 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3444 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3445 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3446 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3447 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3448 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3449 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3450 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3451 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3452 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3453 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3454 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3455 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3456 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3457 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3458 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3459 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3460 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3461 ( .A(n420), .B(n393), .Z(n404) );
  IV U3462 ( .A(n410), .Z(n411) );
  IV U3463 ( .A(n412), .Z(n418) );
  XOR U3464 ( .A(n394), .B(n448), .Z(n397) );
  AND U3465 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3466 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3467 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3469 ( .A(n401), .B(n400), .Z(n422) );
  IV U3470 ( .A(n422), .Z(n417) );
  XOR U3471 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3472 ( .A(n411), .B(n402), .Z(n403) );
  AND U3473 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3474 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3475 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3476 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3477 ( .A(n412), .B(n406), .Z(n407) );
  AND U3478 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3479 ( .A(n482), .B(n464), .Z(n439) );
  OR U3480 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3481 ( .A(n420), .B(n410), .Z(n416) );
  AND U3482 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3483 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3484 ( .A(n414), .B(n413), .Z(n415) );
  AND U3485 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3486 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3487 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3488 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3489 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3490 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3491 ( .A(n454), .B(n439), .Z(n441) );
  OR U3492 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3493 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3494 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3495 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3496 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3497 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3498 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3499 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3500 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3501 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3502 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3503 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3504 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3505 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3506 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3507 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3508 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3509 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3510 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3511 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3512 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3513 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3514 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3515 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3516 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3517 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3518 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3519 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3520 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3521 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3522 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3523 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3524 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3525 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3526 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3527 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3528 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3529 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3530 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3531 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3532 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3533 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3534 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3536 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3537 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3538 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3539 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3540 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3541 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3542 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3543 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3544 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3545 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3546 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3547 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3548 ( .A(n506), .B(n672), .Z(n509) );
  OR U3549 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3550 ( .A(n650), .B(n499), .Z(n671) );
  OR U3551 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3552 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3553 ( .A(n511), .B(n503), .Z(n678) );
  AND U3554 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3555 ( .A(n507), .B(n506), .Z(n675) );
  OR U3556 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3557 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3558 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3559 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3560 ( .A(n515), .B(n514), .Z(n660) );
  OR U3561 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3562 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3563 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3564 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3565 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3566 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3567 ( .A(x[121]), .Z(n628) );
  XOR U3568 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3569 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3570 ( .A(n627), .Z(n524) );
  AND U3571 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3572 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3573 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3574 ( .A(n523), .B(n522), .Z(n587) );
  IV U3575 ( .A(n587), .Z(n533) );
  XNOR U3576 ( .A(n533), .B(n627), .Z(n586) );
  IV U3577 ( .A(x[127]), .Z(n525) );
  XNOR U3578 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3579 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3580 ( .A(n525), .B(n524), .Z(n532) );
  IV U3581 ( .A(n532), .Z(n616) );
  XOR U3582 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3583 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3584 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3585 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3586 ( .A(n526), .Z(n591) );
  NANDN U3587 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3588 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3589 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3590 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3591 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3592 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3593 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3594 ( .A(n531), .B(n530), .Z(n567) );
  IV U3595 ( .A(n567), .Z(n573) );
  AND U3596 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3597 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3598 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3599 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3600 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3601 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3602 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3603 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3604 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3605 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3606 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3607 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3608 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3609 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3610 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3611 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3612 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3613 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3614 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3615 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3616 ( .A(n573), .B(n546), .Z(n557) );
  IV U3617 ( .A(n563), .Z(n564) );
  IV U3618 ( .A(n565), .Z(n571) );
  XOR U3619 ( .A(n547), .B(n601), .Z(n550) );
  AND U3620 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3621 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3622 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3623 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3624 ( .A(n554), .B(n553), .Z(n575) );
  IV U3625 ( .A(n575), .Z(n570) );
  XOR U3626 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3627 ( .A(n564), .B(n555), .Z(n556) );
  AND U3628 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3629 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3630 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3631 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3632 ( .A(n565), .B(n559), .Z(n560) );
  AND U3633 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3634 ( .A(n635), .B(n617), .Z(n592) );
  OR U3635 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3636 ( .A(n573), .B(n563), .Z(n569) );
  AND U3637 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3638 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3639 ( .A(n567), .B(n566), .Z(n568) );
  AND U3640 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3641 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3642 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3643 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3644 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3645 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3646 ( .A(n607), .B(n592), .Z(n594) );
  OR U3647 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3648 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3649 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3650 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3651 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3652 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3653 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3654 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3655 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3656 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3657 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3658 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3659 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3660 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3661 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3662 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3663 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3664 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3665 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3666 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3667 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3668 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3669 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3670 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3671 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3672 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3673 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3674 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3675 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3676 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3677 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3678 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3679 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3680 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3681 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3682 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3683 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3684 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3685 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3686 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3687 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3688 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3689 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3690 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3691 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3692 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3693 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3694 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3695 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3696 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3697 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3698 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3699 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3700 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3701 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3702 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3703 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3704 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3705 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3706 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3707 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3708 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3709 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3710 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3711 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3712 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3713 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3714 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3715 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3716 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3717 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3718 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3719 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3720 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3721 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3722 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3723 ( .A(x[17]), .Z(n815) );
  IV U3724 ( .A(n814), .Z(n686) );
  AND U3725 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3726 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3727 ( .A(n685), .B(n684), .Z(n749) );
  IV U3728 ( .A(n749), .Z(n695) );
  XNOR U3729 ( .A(n695), .B(n814), .Z(n748) );
  IV U3730 ( .A(x[23]), .Z(n687) );
  XNOR U3731 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3732 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3733 ( .A(n687), .B(n686), .Z(n694) );
  IV U3734 ( .A(n694), .Z(n778) );
  XOR U3735 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3736 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3737 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3738 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3739 ( .A(n688), .Z(n753) );
  NANDN U3740 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3741 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3742 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3743 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3744 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3745 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3746 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3747 ( .A(n693), .B(n692), .Z(n729) );
  IV U3748 ( .A(n729), .Z(n735) );
  AND U3749 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3750 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3751 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3752 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3753 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3754 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3755 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3756 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3757 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3758 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3759 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3760 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3761 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3762 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3763 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3764 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3765 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3766 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3767 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3768 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3769 ( .A(n735), .B(n708), .Z(n719) );
  IV U3770 ( .A(n725), .Z(n726) );
  IV U3771 ( .A(n727), .Z(n733) );
  XOR U3772 ( .A(n709), .B(n763), .Z(n712) );
  AND U3773 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3774 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3775 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3776 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3777 ( .A(n716), .B(n715), .Z(n737) );
  IV U3778 ( .A(n737), .Z(n732) );
  XOR U3779 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3780 ( .A(n726), .B(n717), .Z(n718) );
  AND U3781 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3782 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3783 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3784 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3785 ( .A(n727), .B(n721), .Z(n722) );
  AND U3786 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3787 ( .A(n822), .B(n779), .Z(n754) );
  OR U3788 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3789 ( .A(n735), .B(n725), .Z(n731) );
  AND U3790 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3791 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3792 ( .A(n729), .B(n728), .Z(n730) );
  AND U3793 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3794 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3795 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3796 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3797 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3798 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3799 ( .A(n769), .B(n754), .Z(n756) );
  OR U3800 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3801 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3802 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3803 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3804 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3805 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3806 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3807 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3808 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3809 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3810 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3811 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3812 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3813 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3814 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3815 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3816 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3817 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3818 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3819 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3820 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3821 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3822 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3823 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3824 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3825 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3826 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3827 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3828 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3829 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3830 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3831 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3832 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3833 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3834 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3835 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3836 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3837 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3838 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3839 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3840 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3841 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3842 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3843 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3844 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3845 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3846 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3847 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3848 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3849 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3850 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3851 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3852 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3853 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3854 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3855 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3856 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3857 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3858 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3859 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3860 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3861 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3862 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3863 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3864 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3865 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3866 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3867 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3868 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3869 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3870 ( .A(x[25]), .Z(n939) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_9 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n815), .B(x[19]), .Z(n689) );
  XNOR U2963 ( .A(n628), .B(x[123]), .Z(n527) );
  XOR U2964 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2965 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2966 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2967 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2968 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2969 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2970 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3418 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3419 ( .A(n370), .B(n369), .Z(n434) );
  IV U3420 ( .A(n434), .Z(n380) );
  XNOR U3421 ( .A(n380), .B(n474), .Z(n433) );
  IV U3422 ( .A(x[119]), .Z(n372) );
  XNOR U3423 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3424 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3425 ( .A(n372), .B(n371), .Z(n379) );
  IV U3426 ( .A(n379), .Z(n463) );
  XOR U3427 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3428 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3429 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3430 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3431 ( .A(n373), .Z(n438) );
  NANDN U3432 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3433 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3434 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3435 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3436 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3437 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3438 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3439 ( .A(n378), .B(n377), .Z(n414) );
  IV U3440 ( .A(n414), .Z(n420) );
  AND U3441 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3442 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3443 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3444 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3445 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3446 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3447 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3448 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3449 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3450 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3451 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3452 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3453 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3454 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3455 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3456 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3457 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3458 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3459 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3460 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3461 ( .A(n420), .B(n393), .Z(n404) );
  IV U3462 ( .A(n410), .Z(n411) );
  IV U3463 ( .A(n412), .Z(n418) );
  XOR U3464 ( .A(n394), .B(n448), .Z(n397) );
  AND U3465 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3466 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3467 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3469 ( .A(n401), .B(n400), .Z(n422) );
  IV U3470 ( .A(n422), .Z(n417) );
  XOR U3471 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3472 ( .A(n411), .B(n402), .Z(n403) );
  AND U3473 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3474 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3475 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3476 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3477 ( .A(n412), .B(n406), .Z(n407) );
  AND U3478 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3479 ( .A(n482), .B(n464), .Z(n439) );
  OR U3480 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3481 ( .A(n420), .B(n410), .Z(n416) );
  AND U3482 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3483 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3484 ( .A(n414), .B(n413), .Z(n415) );
  AND U3485 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3486 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3487 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3488 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3489 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3490 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3491 ( .A(n454), .B(n439), .Z(n441) );
  OR U3492 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3493 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3494 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3495 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3496 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3497 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3498 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3499 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3500 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3501 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3502 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3503 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3504 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3505 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3506 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3507 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3508 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3509 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3510 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3511 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3512 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3513 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3514 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3515 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3516 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3517 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3518 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3519 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3520 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3521 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3522 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3523 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3524 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3525 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3526 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3527 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3528 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3529 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3530 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3531 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3532 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3533 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3534 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3536 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3537 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3538 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3539 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3540 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3541 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3542 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3543 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3544 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3545 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3546 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3547 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3548 ( .A(n506), .B(n672), .Z(n509) );
  OR U3549 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3550 ( .A(n650), .B(n499), .Z(n671) );
  OR U3551 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3552 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3553 ( .A(n511), .B(n503), .Z(n678) );
  AND U3554 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3555 ( .A(n507), .B(n506), .Z(n675) );
  OR U3556 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3557 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3558 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3559 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3560 ( .A(n515), .B(n514), .Z(n660) );
  OR U3561 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3562 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3563 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3564 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3565 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3566 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3567 ( .A(x[121]), .Z(n628) );
  XOR U3568 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3569 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3570 ( .A(n627), .Z(n524) );
  AND U3571 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3726 ( .A(n685), .B(n684), .Z(n749) );
  IV U3727 ( .A(n749), .Z(n695) );
  XNOR U3728 ( .A(n695), .B(n814), .Z(n748) );
  IV U3729 ( .A(x[23]), .Z(n687) );
  XNOR U3730 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3731 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3732 ( .A(n687), .B(n686), .Z(n694) );
  IV U3733 ( .A(n694), .Z(n778) );
  XOR U3734 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3735 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3736 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3737 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3738 ( .A(n688), .Z(n753) );
  NANDN U3739 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3740 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3741 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3742 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3743 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3744 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3745 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3746 ( .A(n693), .B(n692), .Z(n729) );
  IV U3747 ( .A(n729), .Z(n735) );
  AND U3748 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3749 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3750 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3751 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3752 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3753 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3754 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3755 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3756 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3757 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3758 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3759 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3760 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3761 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3762 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3763 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3764 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3765 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3766 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3767 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3768 ( .A(n735), .B(n708), .Z(n719) );
  IV U3769 ( .A(n725), .Z(n726) );
  IV U3770 ( .A(n727), .Z(n733) );
  XOR U3771 ( .A(n709), .B(n763), .Z(n712) );
  AND U3772 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3773 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3774 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3775 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3776 ( .A(n716), .B(n715), .Z(n737) );
  IV U3777 ( .A(n737), .Z(n732) );
  XOR U3778 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3779 ( .A(n726), .B(n717), .Z(n718) );
  AND U3780 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3781 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3782 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3783 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3784 ( .A(n727), .B(n721), .Z(n722) );
  AND U3785 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3786 ( .A(n822), .B(n779), .Z(n754) );
  OR U3787 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3788 ( .A(n735), .B(n725), .Z(n731) );
  AND U3789 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3790 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3791 ( .A(n729), .B(n728), .Z(n730) );
  AND U3792 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3793 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3794 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3795 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3796 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3797 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3798 ( .A(n769), .B(n754), .Z(n756) );
  OR U3799 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3800 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3801 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3802 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3803 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3804 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3805 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3806 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3807 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3808 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3809 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3810 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3811 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3812 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3813 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3814 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3815 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3816 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3817 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3818 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3819 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3820 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3821 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3822 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3823 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3824 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3825 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3826 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3827 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3828 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3829 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3830 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3831 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3832 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3833 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3834 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3835 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3836 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3837 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3838 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3839 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3840 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3841 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3842 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3843 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3844 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3845 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3846 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3847 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3848 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3849 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3850 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3851 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3852 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3853 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3854 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3855 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3856 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3857 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3858 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3859 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3860 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3861 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3862 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3863 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3864 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3865 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3866 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3867 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3868 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3869 ( .A(x[25]), .Z(n939) );
  XOR U3870 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_10 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U2963 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2964 ( .A(n339), .B(n328), .Z(n341) );
  XOR U2965 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2966 ( .A(n170), .B(n162), .Z(n143) );
  XNOR U2967 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2968 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2969 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2970 ( .A(x[1]), .Z(n1447) );
  XOR U2971 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2972 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2973 ( .A(n1446), .Z(n3) );
  AND U2974 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2975 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2976 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2977 ( .A(n2), .B(n1), .Z(n66) );
  IV U2978 ( .A(n66), .Z(n12) );
  XNOR U2979 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2980 ( .A(x[7]), .Z(n4) );
  XNOR U2981 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2982 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2983 ( .A(n4), .B(n3), .Z(n11) );
  IV U2984 ( .A(n11), .Z(n1083) );
  XOR U2985 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2986 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2987 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2988 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2989 ( .A(n5), .Z(n790) );
  NANDN U2990 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2991 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2992 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2993 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2994 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2995 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2996 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2997 ( .A(n10), .B(n9), .Z(n46) );
  IV U2998 ( .A(n46), .Z(n52) );
  AND U2999 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3000 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3001 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3002 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3003 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3004 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3005 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3006 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3007 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3008 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3009 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3010 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3011 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3012 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3013 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3014 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3015 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3016 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3017 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3018 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3019 ( .A(n52), .B(n25), .Z(n36) );
  IV U3020 ( .A(n42), .Z(n43) );
  IV U3021 ( .A(n44), .Z(n50) );
  XOR U3022 ( .A(n26), .B(n800), .Z(n29) );
  AND U3023 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3024 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3025 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3026 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3027 ( .A(n33), .B(n32), .Z(n54) );
  IV U3028 ( .A(n54), .Z(n49) );
  XOR U3029 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3030 ( .A(n43), .B(n34), .Z(n35) );
  AND U3031 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3032 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3033 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3034 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3035 ( .A(n44), .B(n38), .Z(n39) );
  AND U3036 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3037 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3038 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3039 ( .A(n52), .B(n42), .Z(n48) );
  AND U3040 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3041 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3042 ( .A(n46), .B(n45), .Z(n47) );
  AND U3043 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3044 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3045 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3046 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3047 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3048 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3049 ( .A(n806), .B(n791), .Z(n793) );
  OR U3050 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3051 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3052 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3053 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3054 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3055 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3056 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3057 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3058 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3059 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3060 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3061 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3062 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3063 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3064 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3065 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3066 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3067 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3068 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3069 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3070 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3071 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3072 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3073 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3074 ( .A(n70), .Z(n142) );
  NANDN U3075 ( .A(n128), .B(n142), .Z(n80) );
  IV U3076 ( .A(n135), .Z(n91) );
  XNOR U3077 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3078 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3079 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3080 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3081 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3082 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3083 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3084 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3085 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3086 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3087 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3088 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3089 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3090 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3091 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3092 ( .A(n78), .B(n77), .Z(n115) );
  IV U3093 ( .A(n115), .Z(n108) );
  XNOR U3094 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3095 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3096 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3097 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3098 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3099 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3100 ( .A(n81), .B(n171), .Z(n84) );
  AND U3101 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3102 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3103 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3104 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3105 ( .A(n94), .B(n86), .Z(n118) );
  AND U3106 ( .A(n129), .B(n161), .Z(n89) );
  IV U3107 ( .A(x[97]), .Z(n136) );
  XNOR U3108 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3109 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3110 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3111 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3112 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3113 ( .A(n108), .B(n90), .Z(n99) );
  IV U3114 ( .A(n118), .Z(n102) );
  NAND U3115 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3116 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3117 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3118 ( .A(n97), .B(n96), .Z(n114) );
  IV U3119 ( .A(n107), .Z(n116) );
  XOR U3120 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3121 ( .A(n102), .B(n111), .Z(n98) );
  AND U3122 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3123 ( .A(n118), .B(n108), .Z(n104) );
  AND U3124 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3125 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3126 ( .A(n102), .B(n101), .Z(n103) );
  AND U3127 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3128 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3129 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3130 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3131 ( .A(n131), .B(n106), .Z(n173) );
  IV U3132 ( .A(n114), .Z(n120) );
  NAND U3133 ( .A(n120), .B(n107), .Z(n113) );
  AND U3134 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3135 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3136 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3137 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3138 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3139 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3140 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3141 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3142 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3143 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3144 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3145 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3146 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3147 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3148 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3149 ( .B(n163), .A(n126), .Z(n184) );
  IV U3150 ( .A(n127), .Z(n162) );
  OR U3151 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3152 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3153 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3154 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3155 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3156 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3157 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3158 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3159 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3160 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3161 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3162 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3163 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3164 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3165 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3166 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3167 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3168 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3169 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3170 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3171 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3172 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3173 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3174 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3175 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3176 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3177 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3178 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3179 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3180 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3181 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3182 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3183 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3184 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3185 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3186 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3187 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3188 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3189 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3190 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3191 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3192 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3193 ( .A(x[105]), .Z(n292) );
  XOR U3194 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3195 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3196 ( .A(n291), .Z(n188) );
  AND U3197 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3198 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3199 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3200 ( .A(n187), .B(n186), .Z(n251) );
  IV U3201 ( .A(n251), .Z(n197) );
  XNOR U3202 ( .A(n197), .B(n291), .Z(n250) );
  IV U3203 ( .A(x[111]), .Z(n189) );
  XNOR U3204 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3205 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3206 ( .A(n189), .B(n188), .Z(n196) );
  IV U3207 ( .A(n196), .Z(n280) );
  XOR U3208 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3209 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3210 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3211 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3212 ( .A(n190), .Z(n255) );
  NANDN U3213 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3214 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3215 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3216 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3217 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3218 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3219 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3220 ( .A(n195), .B(n194), .Z(n231) );
  IV U3221 ( .A(n231), .Z(n237) );
  AND U3222 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3223 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3224 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3225 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3226 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3227 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3228 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3229 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3230 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3231 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3232 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3233 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3234 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3235 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3236 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3238 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3239 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3240 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3241 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3242 ( .A(n237), .B(n210), .Z(n221) );
  IV U3243 ( .A(n227), .Z(n228) );
  IV U3244 ( .A(n229), .Z(n235) );
  XOR U3245 ( .A(n211), .B(n265), .Z(n214) );
  AND U3246 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3247 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3248 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3249 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3250 ( .A(n218), .B(n217), .Z(n239) );
  IV U3251 ( .A(n239), .Z(n234) );
  XOR U3252 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3253 ( .A(n228), .B(n219), .Z(n220) );
  AND U3254 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3255 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3256 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3257 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3258 ( .A(n229), .B(n223), .Z(n224) );
  AND U3259 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3260 ( .A(n299), .B(n281), .Z(n256) );
  OR U3261 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3262 ( .A(n237), .B(n227), .Z(n233) );
  AND U3263 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3264 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3265 ( .A(n231), .B(n230), .Z(n232) );
  AND U3266 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3267 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3268 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3269 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3270 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3271 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3272 ( .A(n271), .B(n256), .Z(n258) );
  OR U3273 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3274 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3275 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3276 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3277 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3278 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3279 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3280 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3281 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3282 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3283 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3284 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3285 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3286 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3287 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3288 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3289 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3290 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3291 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3292 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3293 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3294 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3295 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3296 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3297 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3298 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3299 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3300 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3301 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3302 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3303 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3304 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3305 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3306 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3307 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3308 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3309 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3310 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3311 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3312 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3313 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3314 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3315 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3316 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3317 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3318 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3319 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3320 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3321 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3322 ( .A(x[15]), .Z(n311) );
  IV U3323 ( .A(x[10]), .Z(n315) );
  XOR U3324 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3325 ( .A(n315), .B(n307), .Z(n352) );
  IV U3326 ( .A(n352), .Z(n309) );
  XOR U3327 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3328 ( .A(x[9]), .Z(n655) );
  XNOR U3329 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3330 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3331 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3332 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3333 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3334 ( .A(n314), .B(n497), .Z(n318) );
  IV U3335 ( .A(x[13]), .Z(n353) );
  XOR U3336 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3337 ( .A(n353), .B(n310), .Z(n325) );
  IV U3338 ( .A(n325), .Z(n656) );
  XOR U3339 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3340 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3341 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3342 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3343 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3344 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3345 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3346 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3347 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3348 ( .A(n333), .B(n312), .Z(n328) );
  IV U3349 ( .A(n313), .Z(n647) );
  IV U3350 ( .A(n314), .Z(n507) );
  XNOR U3351 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3352 ( .A(n507), .B(n321), .Z(n501) );
  IV U3353 ( .A(n316), .Z(n344) );
  NANDN U3354 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3355 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3356 ( .A(n648), .B(n497), .Z(n498) );
  OR U3357 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3358 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3359 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3360 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3361 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3362 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3363 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3364 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3365 ( .A(n647), .B(n324), .Z(n356) );
  IV U3366 ( .A(n356), .Z(n359) );
  NAND U3367 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3368 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3369 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3370 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3371 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3372 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3373 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3374 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3375 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3376 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3377 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3378 ( .A(n348), .B(n358), .Z(n336) );
  AND U3379 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3380 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3381 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3382 ( .A(n342), .B(n340), .Z(n354) );
  OR U3383 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3384 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3385 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3386 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3387 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3388 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3389 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3390 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3391 ( .A(n347), .B(n346), .Z(n361) );
  OR U3392 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3393 ( .A(n496), .B(n349), .Z(n504) );
  AND U3394 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3395 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3396 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3397 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3398 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3399 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3400 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3401 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3402 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3403 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3404 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3405 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3406 ( .A(n670), .B(n519), .Z(n654) );
  IV U3407 ( .A(n654), .Z(z[10]) );
  XNOR U3408 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3409 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3410 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3411 ( .A(x[113]), .Z(n475) );
  XOR U3412 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3413 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3414 ( .A(n474), .Z(n371) );
  AND U3415 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3416 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3417 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3418 ( .A(n370), .B(n369), .Z(n434) );
  IV U3419 ( .A(n434), .Z(n380) );
  XNOR U3420 ( .A(n380), .B(n474), .Z(n433) );
  IV U3421 ( .A(x[119]), .Z(n372) );
  XNOR U3422 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3423 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3424 ( .A(n372), .B(n371), .Z(n379) );
  IV U3425 ( .A(n379), .Z(n463) );
  XOR U3426 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3427 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3428 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3429 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3430 ( .A(n373), .Z(n438) );
  NANDN U3431 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3432 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3433 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3434 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3435 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3436 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3437 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3438 ( .A(n378), .B(n377), .Z(n414) );
  IV U3439 ( .A(n414), .Z(n420) );
  AND U3440 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3441 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3442 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3443 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3444 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3445 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3446 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3447 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3448 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3449 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3450 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3451 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3452 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3453 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3454 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3455 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3456 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3457 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3458 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3459 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3460 ( .A(n420), .B(n393), .Z(n404) );
  IV U3461 ( .A(n410), .Z(n411) );
  IV U3462 ( .A(n412), .Z(n418) );
  XOR U3463 ( .A(n394), .B(n448), .Z(n397) );
  AND U3464 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3465 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3466 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3467 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3468 ( .A(n401), .B(n400), .Z(n422) );
  IV U3469 ( .A(n422), .Z(n417) );
  XOR U3470 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3471 ( .A(n411), .B(n402), .Z(n403) );
  AND U3472 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3473 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3474 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3475 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3476 ( .A(n412), .B(n406), .Z(n407) );
  AND U3477 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3478 ( .A(n482), .B(n464), .Z(n439) );
  OR U3479 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3480 ( .A(n420), .B(n410), .Z(n416) );
  AND U3481 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3482 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3483 ( .A(n414), .B(n413), .Z(n415) );
  AND U3484 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3485 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3486 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3487 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3488 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3489 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3490 ( .A(n454), .B(n439), .Z(n441) );
  OR U3491 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3492 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3493 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3494 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3495 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3496 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3497 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3498 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3499 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3500 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3501 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3502 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3503 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3504 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3505 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3506 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3507 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3508 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3509 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3510 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3511 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3512 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3513 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3514 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3515 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3516 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3517 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3518 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3519 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3520 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3521 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3522 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3523 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3524 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3525 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3526 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3527 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3528 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3529 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3530 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3531 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3532 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3533 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3534 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3535 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3536 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3537 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3538 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3539 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3540 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3541 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3542 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3543 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3544 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3545 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3546 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3547 ( .A(n506), .B(n672), .Z(n509) );
  OR U3548 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3549 ( .A(n650), .B(n499), .Z(n671) );
  OR U3550 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3551 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3552 ( .A(n511), .B(n503), .Z(n678) );
  AND U3553 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3554 ( .A(n507), .B(n506), .Z(n675) );
  OR U3555 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3556 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3557 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3558 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3559 ( .A(n515), .B(n514), .Z(n660) );
  OR U3560 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3561 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3562 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3563 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3564 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3565 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3566 ( .A(x[121]), .Z(n628) );
  XOR U3567 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3568 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3569 ( .A(n627), .Z(n524) );
  AND U3570 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3571 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3726 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3727 ( .A(n685), .B(n684), .Z(n749) );
  IV U3728 ( .A(n749), .Z(n695) );
  XNOR U3729 ( .A(n695), .B(n814), .Z(n748) );
  IV U3730 ( .A(x[23]), .Z(n687) );
  XNOR U3731 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3732 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3733 ( .A(n687), .B(n686), .Z(n694) );
  IV U3734 ( .A(n694), .Z(n778) );
  XOR U3735 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3736 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3737 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3738 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3739 ( .A(n688), .Z(n753) );
  NANDN U3740 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3741 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3742 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3743 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3744 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3745 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3746 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3747 ( .A(n693), .B(n692), .Z(n729) );
  IV U3748 ( .A(n729), .Z(n735) );
  AND U3749 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3750 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3751 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3752 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3753 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3754 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3755 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3756 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3757 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3758 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3759 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3760 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3761 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3762 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3763 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3764 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3765 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3766 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3767 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3768 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3769 ( .A(n735), .B(n708), .Z(n719) );
  IV U3770 ( .A(n725), .Z(n726) );
  IV U3771 ( .A(n727), .Z(n733) );
  XOR U3772 ( .A(n709), .B(n763), .Z(n712) );
  AND U3773 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3774 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3775 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3776 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3777 ( .A(n716), .B(n715), .Z(n737) );
  IV U3778 ( .A(n737), .Z(n732) );
  XOR U3779 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3780 ( .A(n726), .B(n717), .Z(n718) );
  AND U3781 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3782 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3783 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3784 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3785 ( .A(n727), .B(n721), .Z(n722) );
  AND U3786 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3787 ( .A(n822), .B(n779), .Z(n754) );
  OR U3788 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3789 ( .A(n735), .B(n725), .Z(n731) );
  AND U3790 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3791 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3792 ( .A(n729), .B(n728), .Z(n730) );
  AND U3793 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3794 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3795 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3796 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3797 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3798 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3799 ( .A(n769), .B(n754), .Z(n756) );
  OR U3800 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3801 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3802 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3803 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3804 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3805 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3806 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3807 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3808 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3809 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3810 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3811 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3812 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3813 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3814 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3815 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3816 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3817 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3818 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3819 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3820 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3821 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3822 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3823 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3824 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3825 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3826 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3827 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3828 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3829 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3830 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3831 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3832 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3833 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3834 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3835 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3836 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3837 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3838 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3839 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3840 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3841 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3842 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3843 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3844 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3845 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3846 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3847 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3848 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3849 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3850 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3851 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3852 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3853 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3854 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3855 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3856 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3857 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3858 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3859 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3860 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3861 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3862 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3863 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3864 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3865 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3866 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3867 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3868 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3869 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3870 ( .A(x[25]), .Z(n939) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_11 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U2963 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2964 ( .A(n475), .B(x[115]), .Z(n374) );
  XOR U2965 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2966 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2967 ( .A(n170), .B(n162), .Z(n143) );
  XNOR U2968 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2969 ( .A(x[21]), .B(n685), .Z(n814) );
  XOR U2970 ( .A(n493), .B(n494), .Z(n646) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3418 ( .A(n370), .B(n369), .Z(n434) );
  IV U3419 ( .A(n434), .Z(n380) );
  XNOR U3420 ( .A(n380), .B(n474), .Z(n433) );
  IV U3421 ( .A(x[119]), .Z(n372) );
  XNOR U3422 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3423 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3424 ( .A(n372), .B(n371), .Z(n379) );
  IV U3425 ( .A(n379), .Z(n463) );
  XOR U3426 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3427 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3428 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3429 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3430 ( .A(n373), .Z(n438) );
  NANDN U3431 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3432 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3433 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3434 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3435 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3436 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3437 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3438 ( .A(n378), .B(n377), .Z(n414) );
  IV U3439 ( .A(n414), .Z(n420) );
  AND U3440 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3441 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3442 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3443 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3444 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3445 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3446 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3447 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3448 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3449 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3450 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3451 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3452 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3453 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3454 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3455 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3456 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3457 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3458 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3459 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3460 ( .A(n420), .B(n393), .Z(n404) );
  IV U3461 ( .A(n410), .Z(n411) );
  IV U3462 ( .A(n412), .Z(n418) );
  XOR U3463 ( .A(n394), .B(n448), .Z(n397) );
  AND U3464 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3465 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3466 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3467 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3468 ( .A(n401), .B(n400), .Z(n422) );
  IV U3469 ( .A(n422), .Z(n417) );
  XOR U3470 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3471 ( .A(n411), .B(n402), .Z(n403) );
  AND U3472 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3473 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3474 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3475 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3476 ( .A(n412), .B(n406), .Z(n407) );
  AND U3477 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3478 ( .A(n482), .B(n464), .Z(n439) );
  OR U3479 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3480 ( .A(n420), .B(n410), .Z(n416) );
  AND U3481 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3482 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3483 ( .A(n414), .B(n413), .Z(n415) );
  AND U3484 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3485 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3486 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3487 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3488 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3489 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3490 ( .A(n454), .B(n439), .Z(n441) );
  OR U3491 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3492 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3493 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3494 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3495 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3496 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3497 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3498 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3499 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3500 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3501 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3502 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3503 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3504 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3505 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3506 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3507 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3508 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3509 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3510 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3511 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3512 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3513 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3514 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3515 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3516 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3517 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3518 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3519 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3520 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3521 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3522 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3523 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3524 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3525 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3526 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3527 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3528 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3529 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3530 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3531 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3532 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3533 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3534 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3535 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3536 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3537 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3538 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3539 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3540 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3541 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3542 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3543 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3544 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3545 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3546 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3547 ( .A(n506), .B(n672), .Z(n509) );
  OR U3548 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3549 ( .A(n650), .B(n499), .Z(n671) );
  OR U3550 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3551 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3552 ( .A(n511), .B(n503), .Z(n678) );
  AND U3553 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3554 ( .A(n507), .B(n506), .Z(n675) );
  OR U3555 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3556 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3557 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3558 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3559 ( .A(n515), .B(n514), .Z(n660) );
  OR U3560 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3561 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3562 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3563 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3564 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3565 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3566 ( .A(x[121]), .Z(n628) );
  XOR U3567 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3568 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3569 ( .A(n627), .Z(n524) );
  AND U3570 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3571 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3726 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3727 ( .A(n685), .B(n684), .Z(n749) );
  IV U3728 ( .A(n749), .Z(n695) );
  XNOR U3729 ( .A(n695), .B(n814), .Z(n748) );
  IV U3730 ( .A(x[23]), .Z(n687) );
  XNOR U3731 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3732 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3733 ( .A(n687), .B(n686), .Z(n694) );
  IV U3734 ( .A(n694), .Z(n778) );
  XOR U3735 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3736 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3737 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3738 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3739 ( .A(n688), .Z(n753) );
  NANDN U3740 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3741 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3742 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3743 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3744 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3745 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3746 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3747 ( .A(n693), .B(n692), .Z(n729) );
  IV U3748 ( .A(n729), .Z(n735) );
  AND U3749 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3750 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3751 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3752 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3753 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3754 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3755 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3756 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3757 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3758 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3759 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3760 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3761 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3762 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3763 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3764 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3765 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3766 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3767 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3768 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3769 ( .A(n735), .B(n708), .Z(n719) );
  IV U3770 ( .A(n725), .Z(n726) );
  IV U3771 ( .A(n727), .Z(n733) );
  XOR U3772 ( .A(n709), .B(n763), .Z(n712) );
  AND U3773 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3774 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3775 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3776 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3777 ( .A(n716), .B(n715), .Z(n737) );
  IV U3778 ( .A(n737), .Z(n732) );
  XOR U3779 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3780 ( .A(n726), .B(n717), .Z(n718) );
  AND U3781 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3782 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3783 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3784 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3785 ( .A(n727), .B(n721), .Z(n722) );
  AND U3786 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3787 ( .A(n822), .B(n779), .Z(n754) );
  OR U3788 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3789 ( .A(n735), .B(n725), .Z(n731) );
  AND U3790 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3791 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3792 ( .A(n729), .B(n728), .Z(n730) );
  AND U3793 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3794 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3795 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3796 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3797 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3798 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3799 ( .A(n769), .B(n754), .Z(n756) );
  OR U3800 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3801 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3802 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3803 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3804 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3805 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3806 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3807 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3808 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3809 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3810 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3811 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3812 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3813 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3814 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3815 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3816 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3817 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3818 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3819 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3820 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3821 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3822 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3823 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3824 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3825 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3826 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3827 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3828 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3829 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3830 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3831 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3832 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3833 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3834 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3835 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3836 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3837 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3838 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3839 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3840 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3841 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3842 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3843 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3844 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3845 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3846 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3847 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3848 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3849 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3850 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3851 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3852 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3853 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3854 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3855 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3856 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3857 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3858 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3859 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3860 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3861 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3862 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3863 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3864 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3865 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3866 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3867 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3868 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3869 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3870 ( .A(x[25]), .Z(n939) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_12 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U2963 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2964 ( .A(n475), .B(x[115]), .Z(n374) );
  XNOR U2965 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2966 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XNOR U2967 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2968 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2969 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2970 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3418 ( .A(n370), .B(n369), .Z(n434) );
  IV U3419 ( .A(n434), .Z(n380) );
  XNOR U3420 ( .A(n380), .B(n474), .Z(n433) );
  IV U3421 ( .A(x[119]), .Z(n372) );
  XNOR U3422 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3423 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3424 ( .A(n372), .B(n371), .Z(n379) );
  IV U3425 ( .A(n379), .Z(n463) );
  XOR U3426 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3427 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3428 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3429 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3430 ( .A(n373), .Z(n438) );
  NANDN U3431 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3432 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3433 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3434 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3435 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3436 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3437 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3438 ( .A(n378), .B(n377), .Z(n414) );
  IV U3439 ( .A(n414), .Z(n420) );
  AND U3440 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3441 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3442 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3443 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3444 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3445 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3446 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3447 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3448 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3449 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3450 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3451 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3452 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3453 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3454 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3455 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3456 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3457 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3458 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3459 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3460 ( .A(n420), .B(n393), .Z(n404) );
  IV U3461 ( .A(n410), .Z(n411) );
  IV U3462 ( .A(n412), .Z(n418) );
  XOR U3463 ( .A(n394), .B(n448), .Z(n397) );
  AND U3464 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3465 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3466 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3467 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3468 ( .A(n401), .B(n400), .Z(n422) );
  IV U3469 ( .A(n422), .Z(n417) );
  XOR U3470 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3471 ( .A(n411), .B(n402), .Z(n403) );
  AND U3472 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3473 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3474 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3475 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3476 ( .A(n412), .B(n406), .Z(n407) );
  AND U3477 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3478 ( .A(n482), .B(n464), .Z(n439) );
  OR U3479 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3480 ( .A(n420), .B(n410), .Z(n416) );
  AND U3481 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3482 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3483 ( .A(n414), .B(n413), .Z(n415) );
  AND U3484 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3485 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3486 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3487 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3488 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3489 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3490 ( .A(n454), .B(n439), .Z(n441) );
  OR U3491 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3492 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3493 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3494 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3495 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3496 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3497 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3498 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3499 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3500 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3501 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3502 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3503 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3504 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3505 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3506 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3507 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3508 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3509 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3510 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3511 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3512 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3513 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3514 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3515 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3516 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3517 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3518 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3519 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3520 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3521 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3522 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3523 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3524 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3525 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3526 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3527 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3528 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3529 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3530 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3531 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3532 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3533 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3534 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3535 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3536 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3537 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3538 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3539 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3540 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3541 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3542 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3543 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3544 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3545 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3546 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3547 ( .A(n506), .B(n672), .Z(n509) );
  OR U3548 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3549 ( .A(n650), .B(n499), .Z(n671) );
  OR U3550 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3551 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3552 ( .A(n511), .B(n503), .Z(n678) );
  AND U3553 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3554 ( .A(n507), .B(n506), .Z(n675) );
  OR U3555 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3556 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3557 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3558 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3559 ( .A(n515), .B(n514), .Z(n660) );
  OR U3560 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3561 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3562 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3563 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3564 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3565 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3566 ( .A(x[121]), .Z(n628) );
  XOR U3567 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3568 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3569 ( .A(n627), .Z(n524) );
  AND U3570 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3571 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3726 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3727 ( .A(n685), .B(n684), .Z(n749) );
  IV U3728 ( .A(n749), .Z(n695) );
  XNOR U3729 ( .A(n695), .B(n814), .Z(n748) );
  IV U3730 ( .A(x[23]), .Z(n687) );
  XNOR U3731 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3732 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3733 ( .A(n687), .B(n686), .Z(n694) );
  IV U3734 ( .A(n694), .Z(n778) );
  XOR U3735 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3736 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3737 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3738 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3739 ( .A(n688), .Z(n753) );
  NANDN U3740 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3741 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3742 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3743 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3744 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3745 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3746 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3747 ( .A(n693), .B(n692), .Z(n729) );
  IV U3748 ( .A(n729), .Z(n735) );
  AND U3749 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3750 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3751 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3752 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3753 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3754 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3755 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3756 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3757 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3758 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3759 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3760 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3761 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3762 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3763 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3764 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3765 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3766 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3767 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3768 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3769 ( .A(n735), .B(n708), .Z(n719) );
  IV U3770 ( .A(n725), .Z(n726) );
  IV U3771 ( .A(n727), .Z(n733) );
  XOR U3772 ( .A(n709), .B(n763), .Z(n712) );
  AND U3773 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3774 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3775 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3776 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3777 ( .A(n716), .B(n715), .Z(n737) );
  IV U3778 ( .A(n737), .Z(n732) );
  XOR U3779 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3780 ( .A(n726), .B(n717), .Z(n718) );
  AND U3781 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3782 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3783 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3784 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3785 ( .A(n727), .B(n721), .Z(n722) );
  AND U3786 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3787 ( .A(n822), .B(n779), .Z(n754) );
  OR U3788 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3789 ( .A(n735), .B(n725), .Z(n731) );
  AND U3790 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3791 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3792 ( .A(n729), .B(n728), .Z(n730) );
  AND U3793 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3794 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3795 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3796 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3797 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3798 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3799 ( .A(n769), .B(n754), .Z(n756) );
  OR U3800 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3801 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3802 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3803 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3804 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3805 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3806 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3807 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3808 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3809 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3810 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3811 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3812 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3813 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3814 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3815 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3816 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3817 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3818 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3819 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3820 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3821 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3822 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3823 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3824 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3825 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3826 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3827 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3828 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3829 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3830 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3831 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3832 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3833 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3834 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3835 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3836 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3837 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3838 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3839 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3840 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3841 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3842 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3843 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3844 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3845 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3846 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3847 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3848 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3849 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3850 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3851 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3852 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3853 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3854 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3855 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3856 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3857 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3858 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3859 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3860 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3861 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3862 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3863 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3864 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3865 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3866 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3867 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3868 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3869 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3870 ( .A(x[25]), .Z(n939) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_13 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U2963 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XOR U2964 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2965 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2966 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XNOR U2967 ( .A(n628), .B(x[123]), .Z(n527) );
  XNOR U2968 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2969 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2970 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3418 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3419 ( .A(n370), .B(n369), .Z(n434) );
  IV U3420 ( .A(n434), .Z(n380) );
  XNOR U3421 ( .A(n380), .B(n474), .Z(n433) );
  IV U3422 ( .A(x[119]), .Z(n372) );
  XNOR U3423 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3424 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3425 ( .A(n372), .B(n371), .Z(n379) );
  IV U3426 ( .A(n379), .Z(n463) );
  XOR U3427 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3428 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3429 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3430 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3431 ( .A(n373), .Z(n438) );
  NANDN U3432 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3433 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3434 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3435 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3436 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3437 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3438 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3439 ( .A(n378), .B(n377), .Z(n414) );
  IV U3440 ( .A(n414), .Z(n420) );
  AND U3441 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3442 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3443 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3444 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3445 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3446 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3447 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3448 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3449 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3450 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3451 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3452 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3453 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3454 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3455 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3456 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3457 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3458 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3459 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3460 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3461 ( .A(n420), .B(n393), .Z(n404) );
  IV U3462 ( .A(n410), .Z(n411) );
  IV U3463 ( .A(n412), .Z(n418) );
  XOR U3464 ( .A(n394), .B(n448), .Z(n397) );
  AND U3465 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3466 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3467 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3469 ( .A(n401), .B(n400), .Z(n422) );
  IV U3470 ( .A(n422), .Z(n417) );
  XOR U3471 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3472 ( .A(n411), .B(n402), .Z(n403) );
  AND U3473 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3474 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3475 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3476 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3477 ( .A(n412), .B(n406), .Z(n407) );
  AND U3478 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3479 ( .A(n482), .B(n464), .Z(n439) );
  OR U3480 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3481 ( .A(n420), .B(n410), .Z(n416) );
  AND U3482 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3483 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3484 ( .A(n414), .B(n413), .Z(n415) );
  AND U3485 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3486 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3487 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3488 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3489 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3490 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3491 ( .A(n454), .B(n439), .Z(n441) );
  OR U3492 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3493 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3494 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3495 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3496 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3497 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3498 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3499 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3500 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3501 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3502 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3503 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3504 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3505 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3506 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3507 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3508 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3509 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3510 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3511 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3512 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3513 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3514 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3515 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3516 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3517 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3518 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3519 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3520 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3521 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3522 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3523 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3524 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3525 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3526 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3527 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3528 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3529 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3530 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3531 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3532 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3533 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3534 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3536 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3537 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3538 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3539 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3540 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3541 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3542 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3543 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3544 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3545 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3546 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3547 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3548 ( .A(n506), .B(n672), .Z(n509) );
  OR U3549 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3550 ( .A(n650), .B(n499), .Z(n671) );
  OR U3551 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3552 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3553 ( .A(n511), .B(n503), .Z(n678) );
  AND U3554 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3555 ( .A(n507), .B(n506), .Z(n675) );
  OR U3556 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3557 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3558 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3559 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3560 ( .A(n515), .B(n514), .Z(n660) );
  OR U3561 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3562 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3563 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3564 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3565 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3566 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3567 ( .A(x[121]), .Z(n628) );
  XOR U3568 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3569 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3570 ( .A(n627), .Z(n524) );
  AND U3571 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3726 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3727 ( .A(n685), .B(n684), .Z(n749) );
  IV U3728 ( .A(n749), .Z(n695) );
  XNOR U3729 ( .A(n695), .B(n814), .Z(n748) );
  IV U3730 ( .A(x[23]), .Z(n687) );
  XNOR U3731 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3732 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3733 ( .A(n687), .B(n686), .Z(n694) );
  IV U3734 ( .A(n694), .Z(n778) );
  XOR U3735 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3736 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3737 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3738 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3739 ( .A(n688), .Z(n753) );
  NANDN U3740 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3741 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3742 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3743 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3744 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3745 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3746 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3747 ( .A(n693), .B(n692), .Z(n729) );
  IV U3748 ( .A(n729), .Z(n735) );
  AND U3749 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3750 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3751 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3752 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3753 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3754 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3755 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3756 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3757 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3758 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3759 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3760 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3761 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3762 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3763 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3764 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3765 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3766 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3767 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3768 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3769 ( .A(n735), .B(n708), .Z(n719) );
  IV U3770 ( .A(n725), .Z(n726) );
  IV U3771 ( .A(n727), .Z(n733) );
  XOR U3772 ( .A(n709), .B(n763), .Z(n712) );
  AND U3773 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3774 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3775 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3776 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3777 ( .A(n716), .B(n715), .Z(n737) );
  IV U3778 ( .A(n737), .Z(n732) );
  XOR U3779 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3780 ( .A(n726), .B(n717), .Z(n718) );
  AND U3781 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3782 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3783 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3784 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3785 ( .A(n727), .B(n721), .Z(n722) );
  AND U3786 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3787 ( .A(n822), .B(n779), .Z(n754) );
  OR U3788 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3789 ( .A(n735), .B(n725), .Z(n731) );
  AND U3790 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3791 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3792 ( .A(n729), .B(n728), .Z(n730) );
  AND U3793 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3794 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3795 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3796 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3797 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3798 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3799 ( .A(n769), .B(n754), .Z(n756) );
  OR U3800 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3801 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3802 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3803 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3804 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3805 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3806 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3807 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3808 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3809 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3810 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3811 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3812 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3813 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3814 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3815 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3816 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3817 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3818 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3819 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3820 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3821 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3822 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3823 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3824 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3825 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3826 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3827 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3828 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3829 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3830 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3831 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3832 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3833 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3834 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3835 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3836 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3837 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3838 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3839 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3840 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3841 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3842 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3843 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3844 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3845 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3846 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3847 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3848 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3849 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3850 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3851 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3852 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3853 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3854 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3855 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3856 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3857 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3858 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3859 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3860 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3861 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3862 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3863 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3864 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3865 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3866 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3867 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3868 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3869 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3870 ( .A(x[25]), .Z(n939) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_14 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n815), .B(x[19]), .Z(n689) );
  XOR U2963 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2964 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2965 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2966 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2967 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2968 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2969 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2970 ( .A(x[1]), .Z(n1447) );
  XOR U2971 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2972 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2973 ( .A(n1446), .Z(n3) );
  AND U2974 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2975 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2976 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2977 ( .A(n2), .B(n1), .Z(n66) );
  IV U2978 ( .A(n66), .Z(n12) );
  XNOR U2979 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2980 ( .A(x[7]), .Z(n4) );
  XNOR U2981 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2982 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2983 ( .A(n4), .B(n3), .Z(n11) );
  IV U2984 ( .A(n11), .Z(n1083) );
  XOR U2985 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2986 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2987 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2988 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2989 ( .A(n5), .Z(n790) );
  NANDN U2990 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2991 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2992 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2993 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2994 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2995 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2996 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2997 ( .A(n10), .B(n9), .Z(n46) );
  IV U2998 ( .A(n46), .Z(n52) );
  AND U2999 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3000 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3001 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3002 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3003 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3004 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3005 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3006 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3007 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3008 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3009 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3010 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3011 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3012 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3013 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3014 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3015 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3016 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3017 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3018 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3019 ( .A(n52), .B(n25), .Z(n36) );
  IV U3020 ( .A(n42), .Z(n43) );
  IV U3021 ( .A(n44), .Z(n50) );
  XOR U3022 ( .A(n26), .B(n800), .Z(n29) );
  AND U3023 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3024 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3025 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3026 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3027 ( .A(n33), .B(n32), .Z(n54) );
  IV U3028 ( .A(n54), .Z(n49) );
  XOR U3029 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3030 ( .A(n43), .B(n34), .Z(n35) );
  AND U3031 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3032 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3033 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3034 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3035 ( .A(n44), .B(n38), .Z(n39) );
  AND U3036 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3037 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3038 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3039 ( .A(n52), .B(n42), .Z(n48) );
  AND U3040 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3041 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3042 ( .A(n46), .B(n45), .Z(n47) );
  AND U3043 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3044 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3045 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3046 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3047 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3048 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3049 ( .A(n806), .B(n791), .Z(n793) );
  OR U3050 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3051 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3052 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3053 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3054 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3055 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3056 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3057 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3058 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3059 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3060 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3061 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3062 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3063 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3064 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3065 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3066 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3067 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3068 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3069 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3070 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3071 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3072 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3073 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3074 ( .A(n70), .Z(n142) );
  NANDN U3075 ( .A(n128), .B(n142), .Z(n80) );
  IV U3076 ( .A(n135), .Z(n91) );
  XNOR U3077 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3078 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3079 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3080 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3081 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3082 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3083 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3084 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3085 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3086 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3087 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3088 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3089 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3090 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3091 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3092 ( .A(n78), .B(n77), .Z(n115) );
  IV U3093 ( .A(n115), .Z(n108) );
  XNOR U3094 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3095 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3096 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3097 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3098 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3099 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3100 ( .A(n81), .B(n171), .Z(n84) );
  AND U3101 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3102 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3103 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3104 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3105 ( .A(n94), .B(n86), .Z(n118) );
  AND U3106 ( .A(n129), .B(n161), .Z(n89) );
  IV U3107 ( .A(x[97]), .Z(n136) );
  XNOR U3108 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3109 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3110 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3111 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3112 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3113 ( .A(n108), .B(n90), .Z(n99) );
  IV U3114 ( .A(n118), .Z(n102) );
  NAND U3115 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3116 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3117 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3118 ( .A(n97), .B(n96), .Z(n114) );
  IV U3119 ( .A(n107), .Z(n116) );
  XOR U3120 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3121 ( .A(n102), .B(n111), .Z(n98) );
  AND U3122 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3123 ( .A(n118), .B(n108), .Z(n104) );
  AND U3124 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3125 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3126 ( .A(n102), .B(n101), .Z(n103) );
  AND U3127 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3128 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3129 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3130 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3131 ( .A(n131), .B(n106), .Z(n173) );
  IV U3132 ( .A(n114), .Z(n120) );
  NAND U3133 ( .A(n120), .B(n107), .Z(n113) );
  AND U3134 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3135 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3136 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3137 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3138 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3139 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3140 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3141 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3142 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3143 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3144 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3145 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3146 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3147 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3148 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3149 ( .B(n163), .A(n126), .Z(n184) );
  IV U3150 ( .A(n127), .Z(n162) );
  OR U3151 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3152 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3153 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3154 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3155 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3156 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3157 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3158 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3159 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3160 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3161 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3162 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3163 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3164 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3165 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3166 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3167 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3168 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3169 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3170 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3171 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3172 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3173 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3174 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3175 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3176 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3177 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3178 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3179 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3180 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3181 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3182 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3183 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3184 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3185 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3186 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3187 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3188 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3189 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3190 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3191 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3192 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3193 ( .A(x[105]), .Z(n292) );
  XOR U3194 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3195 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3196 ( .A(n291), .Z(n188) );
  AND U3197 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3198 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3199 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3200 ( .A(n187), .B(n186), .Z(n251) );
  IV U3201 ( .A(n251), .Z(n197) );
  XNOR U3202 ( .A(n197), .B(n291), .Z(n250) );
  IV U3203 ( .A(x[111]), .Z(n189) );
  XNOR U3204 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3205 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3206 ( .A(n189), .B(n188), .Z(n196) );
  IV U3207 ( .A(n196), .Z(n280) );
  XOR U3208 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3209 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3210 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3211 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3212 ( .A(n190), .Z(n255) );
  NANDN U3213 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3214 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3215 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3216 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3217 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3218 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3219 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3220 ( .A(n195), .B(n194), .Z(n231) );
  IV U3221 ( .A(n231), .Z(n237) );
  AND U3222 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3223 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3224 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3225 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3226 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3227 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3228 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3229 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3230 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3231 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3232 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3233 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3234 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3235 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3236 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3238 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3239 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3240 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3241 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3242 ( .A(n237), .B(n210), .Z(n221) );
  IV U3243 ( .A(n227), .Z(n228) );
  IV U3244 ( .A(n229), .Z(n235) );
  XOR U3245 ( .A(n211), .B(n265), .Z(n214) );
  AND U3246 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3247 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3248 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3249 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3250 ( .A(n218), .B(n217), .Z(n239) );
  IV U3251 ( .A(n239), .Z(n234) );
  XOR U3252 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3253 ( .A(n228), .B(n219), .Z(n220) );
  AND U3254 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3255 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3256 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3257 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3258 ( .A(n229), .B(n223), .Z(n224) );
  AND U3259 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3260 ( .A(n299), .B(n281), .Z(n256) );
  OR U3261 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3262 ( .A(n237), .B(n227), .Z(n233) );
  AND U3263 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3264 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3265 ( .A(n231), .B(n230), .Z(n232) );
  AND U3266 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3267 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3268 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3269 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3270 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3271 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3272 ( .A(n271), .B(n256), .Z(n258) );
  OR U3273 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3274 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3275 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3276 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3277 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3278 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3279 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3280 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3281 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3282 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3283 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3284 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3285 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3286 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3287 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3288 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3289 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3290 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3291 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3292 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3293 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3294 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3295 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3296 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3297 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3298 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3299 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3300 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3301 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3302 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3303 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3304 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3305 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3306 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3307 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3308 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3309 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3310 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3311 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3312 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3313 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3314 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3315 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3316 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3317 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3318 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3319 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3320 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3321 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3322 ( .A(x[15]), .Z(n311) );
  IV U3323 ( .A(x[10]), .Z(n315) );
  XOR U3324 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3325 ( .A(n315), .B(n307), .Z(n352) );
  IV U3326 ( .A(n352), .Z(n309) );
  XOR U3327 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3328 ( .A(x[9]), .Z(n655) );
  XNOR U3329 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3330 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3331 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3332 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3333 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3334 ( .A(n314), .B(n497), .Z(n318) );
  IV U3335 ( .A(x[13]), .Z(n353) );
  XOR U3336 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3337 ( .A(n353), .B(n310), .Z(n325) );
  IV U3338 ( .A(n325), .Z(n656) );
  XOR U3339 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3340 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3341 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3342 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3343 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3344 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3345 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3346 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3347 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3348 ( .A(n333), .B(n312), .Z(n328) );
  IV U3349 ( .A(n313), .Z(n647) );
  IV U3350 ( .A(n314), .Z(n507) );
  XNOR U3351 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3352 ( .A(n507), .B(n321), .Z(n501) );
  IV U3353 ( .A(n316), .Z(n344) );
  NANDN U3354 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3355 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3356 ( .A(n648), .B(n497), .Z(n498) );
  OR U3357 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3358 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3359 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3360 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3361 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3362 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3363 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3364 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3365 ( .A(n647), .B(n324), .Z(n356) );
  IV U3366 ( .A(n356), .Z(n359) );
  NAND U3367 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3368 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3369 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3370 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3371 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3372 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3373 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3374 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3375 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3376 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3377 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3378 ( .A(n348), .B(n358), .Z(n336) );
  AND U3379 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3380 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3381 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3382 ( .A(n342), .B(n340), .Z(n354) );
  OR U3383 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3384 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3385 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3386 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3387 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3388 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3389 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3390 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3391 ( .A(n347), .B(n346), .Z(n361) );
  OR U3392 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3393 ( .A(n496), .B(n349), .Z(n504) );
  AND U3394 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3395 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3396 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3397 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3398 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3399 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3400 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3401 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3402 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3403 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3404 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3405 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3406 ( .A(n670), .B(n519), .Z(n654) );
  IV U3407 ( .A(n654), .Z(z[10]) );
  XNOR U3408 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3409 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3410 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3411 ( .A(x[113]), .Z(n475) );
  XOR U3412 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3413 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3414 ( .A(n474), .Z(n371) );
  AND U3415 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3416 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3417 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3418 ( .A(n370), .B(n369), .Z(n434) );
  IV U3419 ( .A(n434), .Z(n380) );
  XNOR U3420 ( .A(n380), .B(n474), .Z(n433) );
  IV U3421 ( .A(x[119]), .Z(n372) );
  XNOR U3422 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3423 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3424 ( .A(n372), .B(n371), .Z(n379) );
  IV U3425 ( .A(n379), .Z(n463) );
  XOR U3426 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3427 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3428 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3429 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3430 ( .A(n373), .Z(n438) );
  NANDN U3431 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3432 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3433 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3434 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3435 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3436 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3437 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3438 ( .A(n378), .B(n377), .Z(n414) );
  IV U3439 ( .A(n414), .Z(n420) );
  AND U3440 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3441 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3442 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3443 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3444 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3445 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3446 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3447 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3448 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3449 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3450 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3451 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3452 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3453 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3454 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3455 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3456 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3457 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3458 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3459 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3460 ( .A(n420), .B(n393), .Z(n404) );
  IV U3461 ( .A(n410), .Z(n411) );
  IV U3462 ( .A(n412), .Z(n418) );
  XOR U3463 ( .A(n394), .B(n448), .Z(n397) );
  AND U3464 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3465 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3466 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3467 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3468 ( .A(n401), .B(n400), .Z(n422) );
  IV U3469 ( .A(n422), .Z(n417) );
  XOR U3470 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3471 ( .A(n411), .B(n402), .Z(n403) );
  AND U3472 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3473 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3474 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3475 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3476 ( .A(n412), .B(n406), .Z(n407) );
  AND U3477 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3478 ( .A(n482), .B(n464), .Z(n439) );
  OR U3479 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3480 ( .A(n420), .B(n410), .Z(n416) );
  AND U3481 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3482 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3483 ( .A(n414), .B(n413), .Z(n415) );
  AND U3484 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3485 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3486 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3487 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3488 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3489 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3490 ( .A(n454), .B(n439), .Z(n441) );
  OR U3491 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3492 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3493 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3494 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3495 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3496 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3497 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3498 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3499 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3500 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3501 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3502 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3503 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3504 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3505 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3506 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3507 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3508 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3509 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3510 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3511 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3512 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3513 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3514 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3515 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3516 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3517 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3518 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3519 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3520 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3521 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3522 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3523 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3524 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3525 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3526 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3527 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3528 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3529 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3530 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3531 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3532 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3533 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3534 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3535 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3536 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3537 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3538 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3539 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3540 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3541 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3542 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3543 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3544 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3545 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3546 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3547 ( .A(n506), .B(n672), .Z(n509) );
  OR U3548 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3549 ( .A(n650), .B(n499), .Z(n671) );
  OR U3550 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3551 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3552 ( .A(n511), .B(n503), .Z(n678) );
  AND U3553 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3554 ( .A(n507), .B(n506), .Z(n675) );
  OR U3555 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3556 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3557 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3558 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3559 ( .A(n515), .B(n514), .Z(n660) );
  OR U3560 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3561 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3562 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3563 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3564 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3565 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3566 ( .A(x[121]), .Z(n628) );
  XOR U3567 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3568 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3569 ( .A(n627), .Z(n524) );
  AND U3570 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3571 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3726 ( .A(n685), .B(n684), .Z(n749) );
  IV U3727 ( .A(n749), .Z(n695) );
  XNOR U3728 ( .A(n695), .B(n814), .Z(n748) );
  IV U3729 ( .A(x[23]), .Z(n687) );
  XNOR U3730 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3731 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3732 ( .A(n687), .B(n686), .Z(n694) );
  IV U3733 ( .A(n694), .Z(n778) );
  XOR U3734 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3735 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3736 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3737 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3738 ( .A(n688), .Z(n753) );
  NANDN U3739 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3740 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3741 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3742 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3743 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3744 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3745 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3746 ( .A(n693), .B(n692), .Z(n729) );
  IV U3747 ( .A(n729), .Z(n735) );
  AND U3748 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3749 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3750 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3751 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3752 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3753 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3754 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3755 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3756 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3757 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3758 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3759 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3760 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3761 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3762 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3763 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3764 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3765 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3766 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3767 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3768 ( .A(n735), .B(n708), .Z(n719) );
  IV U3769 ( .A(n725), .Z(n726) );
  IV U3770 ( .A(n727), .Z(n733) );
  XOR U3771 ( .A(n709), .B(n763), .Z(n712) );
  AND U3772 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3773 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3774 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3775 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3776 ( .A(n716), .B(n715), .Z(n737) );
  IV U3777 ( .A(n737), .Z(n732) );
  XOR U3778 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3779 ( .A(n726), .B(n717), .Z(n718) );
  AND U3780 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3781 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3782 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3783 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3784 ( .A(n727), .B(n721), .Z(n722) );
  AND U3785 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3786 ( .A(n822), .B(n779), .Z(n754) );
  OR U3787 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3788 ( .A(n735), .B(n725), .Z(n731) );
  AND U3789 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3790 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3791 ( .A(n729), .B(n728), .Z(n730) );
  AND U3792 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3793 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3794 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3795 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3796 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3797 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3798 ( .A(n769), .B(n754), .Z(n756) );
  OR U3799 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3800 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3801 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3802 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3803 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3804 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3805 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3806 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3807 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3808 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3809 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3810 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3811 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3812 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3813 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3814 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3815 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3816 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3817 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3818 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3819 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3820 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3821 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3822 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3823 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3824 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3825 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3826 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3827 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3828 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3829 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3830 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3831 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3832 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3833 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3834 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3835 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3836 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3837 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3838 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3839 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3840 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3841 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3842 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3843 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3844 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3845 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3846 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3847 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3848 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3849 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3850 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3851 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3852 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3853 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3854 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3855 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3856 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3857 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3858 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3859 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3860 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3861 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3862 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3863 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3864 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3865 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3866 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3867 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3868 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3869 ( .A(x[25]), .Z(n939) );
  XOR U3870 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_15 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n475), .B(x[115]), .Z(n374) );
  XNOR U2963 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2964 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2965 ( .A(n339), .B(n328), .Z(n341) );
  XOR U2966 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XOR U2967 ( .A(n493), .B(n494), .Z(n646) );
  XNOR U2968 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2969 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2970 ( .A(x[1]), .Z(n1447) );
  XOR U2971 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2972 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2973 ( .A(n1446), .Z(n3) );
  AND U2974 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2975 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2976 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2977 ( .A(n2), .B(n1), .Z(n66) );
  IV U2978 ( .A(n66), .Z(n12) );
  XNOR U2979 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2980 ( .A(x[7]), .Z(n4) );
  XNOR U2981 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2982 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2983 ( .A(n4), .B(n3), .Z(n11) );
  IV U2984 ( .A(n11), .Z(n1083) );
  XOR U2985 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2986 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2987 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2988 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2989 ( .A(n5), .Z(n790) );
  NANDN U2990 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2991 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2992 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2993 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2994 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2995 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2996 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2997 ( .A(n10), .B(n9), .Z(n46) );
  IV U2998 ( .A(n46), .Z(n52) );
  AND U2999 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3000 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3001 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3002 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3003 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3004 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3005 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3006 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3007 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3008 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3009 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3010 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3011 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3012 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3013 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3014 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3015 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3016 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3017 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3018 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3019 ( .A(n52), .B(n25), .Z(n36) );
  IV U3020 ( .A(n42), .Z(n43) );
  IV U3021 ( .A(n44), .Z(n50) );
  XOR U3022 ( .A(n26), .B(n800), .Z(n29) );
  AND U3023 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3024 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3025 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3026 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3027 ( .A(n33), .B(n32), .Z(n54) );
  IV U3028 ( .A(n54), .Z(n49) );
  XOR U3029 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3030 ( .A(n43), .B(n34), .Z(n35) );
  AND U3031 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3032 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3033 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3034 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3035 ( .A(n44), .B(n38), .Z(n39) );
  AND U3036 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3037 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3038 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3039 ( .A(n52), .B(n42), .Z(n48) );
  AND U3040 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3041 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3042 ( .A(n46), .B(n45), .Z(n47) );
  AND U3043 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3044 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3045 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3046 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3047 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3048 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3049 ( .A(n806), .B(n791), .Z(n793) );
  OR U3050 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3051 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3052 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3053 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3054 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3055 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3056 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3057 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3058 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3059 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3060 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3061 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3062 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3063 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3064 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3065 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3066 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3067 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3068 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3069 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3070 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3071 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3072 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3073 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3074 ( .A(n70), .Z(n142) );
  NANDN U3075 ( .A(n128), .B(n142), .Z(n80) );
  IV U3076 ( .A(n135), .Z(n91) );
  XNOR U3077 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3078 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3079 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3080 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3081 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3082 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3083 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3084 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3085 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3086 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3087 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3088 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3089 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3090 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3091 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3092 ( .A(n78), .B(n77), .Z(n115) );
  IV U3093 ( .A(n115), .Z(n108) );
  XNOR U3094 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3095 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3096 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3097 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3098 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3099 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3100 ( .A(n81), .B(n171), .Z(n84) );
  AND U3101 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3102 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3103 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3104 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3105 ( .A(n94), .B(n86), .Z(n118) );
  AND U3106 ( .A(n129), .B(n161), .Z(n89) );
  IV U3107 ( .A(x[97]), .Z(n136) );
  XNOR U3108 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3109 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3110 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3111 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3112 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3113 ( .A(n108), .B(n90), .Z(n99) );
  IV U3114 ( .A(n118), .Z(n102) );
  NAND U3115 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3116 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3117 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3118 ( .A(n97), .B(n96), .Z(n114) );
  IV U3119 ( .A(n107), .Z(n116) );
  XOR U3120 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3121 ( .A(n102), .B(n111), .Z(n98) );
  AND U3122 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3123 ( .A(n118), .B(n108), .Z(n104) );
  AND U3124 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3125 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3126 ( .A(n102), .B(n101), .Z(n103) );
  AND U3127 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3128 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3129 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3130 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3131 ( .A(n131), .B(n106), .Z(n173) );
  IV U3132 ( .A(n114), .Z(n120) );
  NAND U3133 ( .A(n120), .B(n107), .Z(n113) );
  AND U3134 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3135 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3136 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3137 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3138 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3139 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3140 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3141 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3142 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3143 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3144 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3145 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3146 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3147 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3148 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3149 ( .B(n163), .A(n126), .Z(n184) );
  IV U3150 ( .A(n127), .Z(n162) );
  OR U3151 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3152 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3153 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3154 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3155 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3156 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3157 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3158 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3159 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3160 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3161 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3162 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3163 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3164 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3165 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3166 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3167 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3168 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3169 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3170 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3171 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3172 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3173 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3174 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3175 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3176 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3177 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3178 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3179 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3180 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3181 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3182 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3183 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3184 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3185 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3186 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3187 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3188 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3189 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3190 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3191 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3192 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3193 ( .A(x[105]), .Z(n292) );
  XOR U3194 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3195 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3196 ( .A(n291), .Z(n188) );
  AND U3197 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3198 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3199 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3200 ( .A(n187), .B(n186), .Z(n251) );
  IV U3201 ( .A(n251), .Z(n197) );
  XNOR U3202 ( .A(n197), .B(n291), .Z(n250) );
  IV U3203 ( .A(x[111]), .Z(n189) );
  XNOR U3204 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3205 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3206 ( .A(n189), .B(n188), .Z(n196) );
  IV U3207 ( .A(n196), .Z(n280) );
  XOR U3208 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3209 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3210 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3211 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3212 ( .A(n190), .Z(n255) );
  NANDN U3213 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3214 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3215 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3216 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3217 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3218 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3219 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3220 ( .A(n195), .B(n194), .Z(n231) );
  IV U3221 ( .A(n231), .Z(n237) );
  AND U3222 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3223 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3224 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3225 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3226 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3227 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3228 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3229 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3230 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3231 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3232 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3233 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3234 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3235 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3236 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3238 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3239 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3240 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3241 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3242 ( .A(n237), .B(n210), .Z(n221) );
  IV U3243 ( .A(n227), .Z(n228) );
  IV U3244 ( .A(n229), .Z(n235) );
  XOR U3245 ( .A(n211), .B(n265), .Z(n214) );
  AND U3246 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3247 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3248 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3249 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3250 ( .A(n218), .B(n217), .Z(n239) );
  IV U3251 ( .A(n239), .Z(n234) );
  XOR U3252 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3253 ( .A(n228), .B(n219), .Z(n220) );
  AND U3254 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3255 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3256 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3257 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3258 ( .A(n229), .B(n223), .Z(n224) );
  AND U3259 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3260 ( .A(n299), .B(n281), .Z(n256) );
  OR U3261 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3262 ( .A(n237), .B(n227), .Z(n233) );
  AND U3263 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3264 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3265 ( .A(n231), .B(n230), .Z(n232) );
  AND U3266 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3267 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3268 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3269 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3270 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3271 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3272 ( .A(n271), .B(n256), .Z(n258) );
  OR U3273 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3274 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3275 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3276 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3277 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3278 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3279 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3280 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3281 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3282 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3283 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3284 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3285 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3286 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3287 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3288 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3289 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3290 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3291 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3292 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3293 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3294 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3295 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3296 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3297 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3298 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3299 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3300 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3301 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3302 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3303 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3304 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3305 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3306 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3307 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3308 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3309 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3310 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3311 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3312 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3313 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3314 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3315 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3316 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3317 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3318 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3319 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3320 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3321 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3322 ( .A(x[15]), .Z(n311) );
  IV U3323 ( .A(x[10]), .Z(n315) );
  XOR U3324 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3325 ( .A(n315), .B(n307), .Z(n352) );
  IV U3326 ( .A(n352), .Z(n309) );
  XOR U3327 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3328 ( .A(x[9]), .Z(n655) );
  XNOR U3329 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3330 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3331 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3332 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3333 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3334 ( .A(n314), .B(n497), .Z(n318) );
  IV U3335 ( .A(x[13]), .Z(n353) );
  XOR U3336 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3337 ( .A(n353), .B(n310), .Z(n325) );
  IV U3338 ( .A(n325), .Z(n656) );
  XOR U3339 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3340 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3341 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3342 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3343 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3344 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3345 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3346 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3347 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3348 ( .A(n333), .B(n312), .Z(n328) );
  IV U3349 ( .A(n313), .Z(n647) );
  IV U3350 ( .A(n314), .Z(n507) );
  XNOR U3351 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3352 ( .A(n507), .B(n321), .Z(n501) );
  IV U3353 ( .A(n316), .Z(n344) );
  NANDN U3354 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3355 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3356 ( .A(n648), .B(n497), .Z(n498) );
  OR U3357 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3358 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3359 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3360 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3361 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3362 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3363 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3364 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3365 ( .A(n647), .B(n324), .Z(n356) );
  IV U3366 ( .A(n356), .Z(n359) );
  NAND U3367 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3368 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3369 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3370 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3371 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3372 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3373 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3374 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3375 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3376 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3377 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3378 ( .A(n348), .B(n358), .Z(n336) );
  AND U3379 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3380 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3381 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3382 ( .A(n342), .B(n340), .Z(n354) );
  OR U3383 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3384 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3385 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3386 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3387 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3388 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3389 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3390 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3391 ( .A(n347), .B(n346), .Z(n361) );
  OR U3392 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3393 ( .A(n496), .B(n349), .Z(n504) );
  AND U3394 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3395 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3396 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3397 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3398 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3399 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3400 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3401 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3402 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3403 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3404 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3405 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3406 ( .A(n670), .B(n519), .Z(n654) );
  IV U3407 ( .A(n654), .Z(z[10]) );
  XNOR U3408 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3409 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3410 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3411 ( .A(x[113]), .Z(n475) );
  XOR U3412 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3413 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3414 ( .A(n474), .Z(n371) );
  AND U3415 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3416 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3417 ( .A(n370), .B(n369), .Z(n434) );
  IV U3418 ( .A(n434), .Z(n380) );
  XNOR U3419 ( .A(n380), .B(n474), .Z(n433) );
  IV U3420 ( .A(x[119]), .Z(n372) );
  XNOR U3421 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3422 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3423 ( .A(n372), .B(n371), .Z(n379) );
  IV U3424 ( .A(n379), .Z(n463) );
  XOR U3425 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3426 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3427 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3428 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3429 ( .A(n373), .Z(n438) );
  NANDN U3430 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3431 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3432 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3433 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3434 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3435 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3436 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3437 ( .A(n378), .B(n377), .Z(n414) );
  IV U3438 ( .A(n414), .Z(n420) );
  AND U3439 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3440 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3441 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3442 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3443 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3444 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3445 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3446 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3447 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3448 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3449 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3450 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3451 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3452 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3453 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3454 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3455 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3456 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3457 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3458 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3459 ( .A(n420), .B(n393), .Z(n404) );
  IV U3460 ( .A(n410), .Z(n411) );
  IV U3461 ( .A(n412), .Z(n418) );
  XOR U3462 ( .A(n394), .B(n448), .Z(n397) );
  AND U3463 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3464 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3465 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3466 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3467 ( .A(n401), .B(n400), .Z(n422) );
  IV U3468 ( .A(n422), .Z(n417) );
  XOR U3469 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3470 ( .A(n411), .B(n402), .Z(n403) );
  AND U3471 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3472 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3473 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3474 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3475 ( .A(n412), .B(n406), .Z(n407) );
  AND U3476 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3477 ( .A(n482), .B(n464), .Z(n439) );
  OR U3478 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3479 ( .A(n420), .B(n410), .Z(n416) );
  AND U3480 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3481 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3482 ( .A(n414), .B(n413), .Z(n415) );
  AND U3483 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3484 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3485 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3486 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3487 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3488 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3489 ( .A(n454), .B(n439), .Z(n441) );
  OR U3490 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3491 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3492 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3493 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3494 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3495 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3496 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3497 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3498 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3499 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3500 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3501 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3502 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3503 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3504 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3505 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3506 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3507 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3508 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3509 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3510 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3511 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3512 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3513 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3514 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3515 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3516 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3517 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3518 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3519 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3520 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3521 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3522 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3523 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3524 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3525 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3526 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3527 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3528 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3529 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3530 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3531 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3532 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3533 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3534 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3535 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3536 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3537 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3538 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3539 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3540 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3541 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3542 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3543 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3544 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3545 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3546 ( .A(n506), .B(n672), .Z(n509) );
  OR U3547 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3548 ( .A(n650), .B(n499), .Z(n671) );
  OR U3549 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3550 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3551 ( .A(n511), .B(n503), .Z(n678) );
  AND U3552 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3553 ( .A(n507), .B(n506), .Z(n675) );
  OR U3554 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3555 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3556 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3557 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3558 ( .A(n515), .B(n514), .Z(n660) );
  OR U3559 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3560 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3561 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3562 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3563 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3564 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3565 ( .A(x[121]), .Z(n628) );
  XOR U3566 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3567 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3568 ( .A(n627), .Z(n524) );
  AND U3569 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3570 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3571 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3572 ( .A(n523), .B(n522), .Z(n587) );
  IV U3573 ( .A(n587), .Z(n533) );
  XNOR U3574 ( .A(n533), .B(n627), .Z(n586) );
  IV U3575 ( .A(x[127]), .Z(n525) );
  XNOR U3576 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3577 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3578 ( .A(n525), .B(n524), .Z(n532) );
  IV U3579 ( .A(n532), .Z(n616) );
  XOR U3580 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3581 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3582 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3583 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3584 ( .A(n526), .Z(n591) );
  NANDN U3585 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3586 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3587 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3588 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3589 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3590 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3591 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3592 ( .A(n531), .B(n530), .Z(n567) );
  IV U3593 ( .A(n567), .Z(n573) );
  AND U3594 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3595 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3596 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3597 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3598 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3599 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3600 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3601 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3602 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3603 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3604 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3605 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3606 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3607 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3608 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3609 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3610 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3611 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3612 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3613 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3614 ( .A(n573), .B(n546), .Z(n557) );
  IV U3615 ( .A(n563), .Z(n564) );
  IV U3616 ( .A(n565), .Z(n571) );
  XOR U3617 ( .A(n547), .B(n601), .Z(n550) );
  AND U3618 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3619 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3620 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3621 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3622 ( .A(n554), .B(n553), .Z(n575) );
  IV U3623 ( .A(n575), .Z(n570) );
  XOR U3624 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3625 ( .A(n564), .B(n555), .Z(n556) );
  AND U3626 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3627 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3628 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3629 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3630 ( .A(n565), .B(n559), .Z(n560) );
  AND U3631 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3632 ( .A(n635), .B(n617), .Z(n592) );
  OR U3633 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3634 ( .A(n573), .B(n563), .Z(n569) );
  AND U3635 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3636 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3637 ( .A(n567), .B(n566), .Z(n568) );
  AND U3638 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3639 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3640 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3641 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3642 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3643 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3644 ( .A(n607), .B(n592), .Z(n594) );
  OR U3645 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3646 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3647 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3648 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3649 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3650 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3651 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3652 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3653 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3654 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3655 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3656 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3657 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3658 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3659 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3660 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3661 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3662 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3663 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3664 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3665 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3666 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3667 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3668 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3669 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3670 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3671 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3672 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3673 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3674 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3675 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3676 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3677 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3678 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3679 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3680 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3681 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3682 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3683 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3684 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3685 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3686 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3687 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3688 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3689 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3690 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3691 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3692 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3693 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3694 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3695 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3696 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3697 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3698 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3699 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3700 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3701 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3702 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3703 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3704 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3705 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3706 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3707 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3708 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3709 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3710 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3711 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3712 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3713 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3714 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3715 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3716 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3717 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3718 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3719 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3720 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3721 ( .A(x[17]), .Z(n815) );
  IV U3722 ( .A(n814), .Z(n686) );
  AND U3723 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3724 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3725 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3726 ( .A(n685), .B(n684), .Z(n749) );
  IV U3727 ( .A(n749), .Z(n695) );
  XNOR U3728 ( .A(n695), .B(n814), .Z(n748) );
  IV U3729 ( .A(x[23]), .Z(n687) );
  XNOR U3730 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3731 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3732 ( .A(n687), .B(n686), .Z(n694) );
  IV U3733 ( .A(n694), .Z(n778) );
  XOR U3734 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3735 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3736 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3737 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3738 ( .A(n688), .Z(n753) );
  NANDN U3739 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3740 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3741 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3742 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3743 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3744 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3745 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3746 ( .A(n693), .B(n692), .Z(n729) );
  IV U3747 ( .A(n729), .Z(n735) );
  AND U3748 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3749 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3750 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3751 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3752 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3753 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3754 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3755 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3756 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3757 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3758 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3759 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3760 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3761 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3762 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3763 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3764 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3765 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3766 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3767 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3768 ( .A(n735), .B(n708), .Z(n719) );
  IV U3769 ( .A(n725), .Z(n726) );
  IV U3770 ( .A(n727), .Z(n733) );
  XOR U3771 ( .A(n709), .B(n763), .Z(n712) );
  AND U3772 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3773 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3774 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3775 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3776 ( .A(n716), .B(n715), .Z(n737) );
  IV U3777 ( .A(n737), .Z(n732) );
  XOR U3778 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3779 ( .A(n726), .B(n717), .Z(n718) );
  AND U3780 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3781 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3782 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3783 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3784 ( .A(n727), .B(n721), .Z(n722) );
  AND U3785 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3786 ( .A(n822), .B(n779), .Z(n754) );
  OR U3787 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3788 ( .A(n735), .B(n725), .Z(n731) );
  AND U3789 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3790 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3791 ( .A(n729), .B(n728), .Z(n730) );
  AND U3792 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3793 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3794 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3795 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3796 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3797 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3798 ( .A(n769), .B(n754), .Z(n756) );
  OR U3799 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3800 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3801 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3802 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3803 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3804 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3805 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3806 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3807 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3808 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3809 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3810 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3811 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3812 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3813 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3814 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3815 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3816 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3817 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3818 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3819 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3820 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3821 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3822 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3823 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3824 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3825 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3826 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3827 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3828 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3829 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3830 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3831 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3832 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3833 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3834 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3835 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3836 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3837 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3838 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3839 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3840 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3841 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3842 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3843 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3844 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3845 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3846 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3847 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3848 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3849 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3850 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3851 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3852 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3853 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3854 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3855 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3856 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3857 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3858 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3859 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3860 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3861 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3862 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3863 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3864 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3865 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3866 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3867 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3868 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3869 ( .A(x[25]), .Z(n939) );
  XOR U3870 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_16 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U2963 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2964 ( .A(n339), .B(n328), .Z(n341) );
  XNOR U2965 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2966 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2967 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2968 ( .A(n493), .B(n494), .Z(n646) );
  XNOR U2969 ( .A(n628), .B(x[123]), .Z(n527) );
  XOR U2970 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3418 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3419 ( .A(n370), .B(n369), .Z(n434) );
  IV U3420 ( .A(n434), .Z(n380) );
  XNOR U3421 ( .A(n380), .B(n474), .Z(n433) );
  IV U3422 ( .A(x[119]), .Z(n372) );
  XNOR U3423 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3424 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3425 ( .A(n372), .B(n371), .Z(n379) );
  IV U3426 ( .A(n379), .Z(n463) );
  XOR U3427 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3428 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3429 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3430 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3431 ( .A(n373), .Z(n438) );
  NANDN U3432 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3433 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3434 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3435 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3436 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3437 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3438 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3439 ( .A(n378), .B(n377), .Z(n414) );
  IV U3440 ( .A(n414), .Z(n420) );
  AND U3441 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3442 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3443 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3444 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3445 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3446 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3447 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3448 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3449 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3450 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3451 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3452 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3453 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3454 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3455 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3456 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3457 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3458 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3459 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3460 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3461 ( .A(n420), .B(n393), .Z(n404) );
  IV U3462 ( .A(n410), .Z(n411) );
  IV U3463 ( .A(n412), .Z(n418) );
  XOR U3464 ( .A(n394), .B(n448), .Z(n397) );
  AND U3465 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3466 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3467 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3469 ( .A(n401), .B(n400), .Z(n422) );
  IV U3470 ( .A(n422), .Z(n417) );
  XOR U3471 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3472 ( .A(n411), .B(n402), .Z(n403) );
  AND U3473 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3474 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3475 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3476 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3477 ( .A(n412), .B(n406), .Z(n407) );
  AND U3478 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3479 ( .A(n482), .B(n464), .Z(n439) );
  OR U3480 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3481 ( .A(n420), .B(n410), .Z(n416) );
  AND U3482 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3483 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3484 ( .A(n414), .B(n413), .Z(n415) );
  AND U3485 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3486 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3487 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3488 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3489 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3490 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3491 ( .A(n454), .B(n439), .Z(n441) );
  OR U3492 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3493 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3494 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3495 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3496 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3497 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3498 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3499 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3500 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3501 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3502 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3503 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3504 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3505 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3506 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3507 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3508 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3509 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3510 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3511 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3512 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3513 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3514 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3515 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3516 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3517 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3518 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3519 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3520 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3521 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3522 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3523 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3524 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3525 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3526 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3527 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3528 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3529 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3530 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3531 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3532 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3533 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3534 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3536 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3537 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3538 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3539 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3540 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3541 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3542 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3543 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3544 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3545 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3546 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3547 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3548 ( .A(n506), .B(n672), .Z(n509) );
  OR U3549 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3550 ( .A(n650), .B(n499), .Z(n671) );
  OR U3551 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3552 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3553 ( .A(n511), .B(n503), .Z(n678) );
  AND U3554 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3555 ( .A(n507), .B(n506), .Z(n675) );
  OR U3556 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3557 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3558 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3559 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3560 ( .A(n515), .B(n514), .Z(n660) );
  OR U3561 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3562 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3563 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3564 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3565 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3566 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3567 ( .A(x[121]), .Z(n628) );
  XOR U3568 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3569 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3570 ( .A(n627), .Z(n524) );
  AND U3571 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3572 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3573 ( .A(n523), .B(n522), .Z(n587) );
  IV U3574 ( .A(n587), .Z(n533) );
  XNOR U3575 ( .A(n533), .B(n627), .Z(n586) );
  IV U3576 ( .A(x[127]), .Z(n525) );
  XNOR U3577 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3578 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3579 ( .A(n525), .B(n524), .Z(n532) );
  IV U3580 ( .A(n532), .Z(n616) );
  XOR U3581 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3582 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3583 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3584 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3585 ( .A(n526), .Z(n591) );
  NANDN U3586 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3587 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3588 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3589 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3590 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3591 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3592 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3593 ( .A(n531), .B(n530), .Z(n567) );
  IV U3594 ( .A(n567), .Z(n573) );
  AND U3595 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3596 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3597 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3598 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3599 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3600 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3601 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3602 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3603 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3604 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3605 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3606 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3607 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3608 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3609 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3610 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3611 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3612 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3613 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3614 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3615 ( .A(n573), .B(n546), .Z(n557) );
  IV U3616 ( .A(n563), .Z(n564) );
  IV U3617 ( .A(n565), .Z(n571) );
  XOR U3618 ( .A(n547), .B(n601), .Z(n550) );
  AND U3619 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3620 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3621 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3622 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3623 ( .A(n554), .B(n553), .Z(n575) );
  IV U3624 ( .A(n575), .Z(n570) );
  XOR U3625 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3626 ( .A(n564), .B(n555), .Z(n556) );
  AND U3627 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3628 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3629 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3630 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3631 ( .A(n565), .B(n559), .Z(n560) );
  AND U3632 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3633 ( .A(n635), .B(n617), .Z(n592) );
  OR U3634 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3635 ( .A(n573), .B(n563), .Z(n569) );
  AND U3636 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3637 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3638 ( .A(n567), .B(n566), .Z(n568) );
  AND U3639 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3640 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3641 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3642 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3643 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3644 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3645 ( .A(n607), .B(n592), .Z(n594) );
  OR U3646 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3647 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3648 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3649 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3650 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3651 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3652 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3653 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3654 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3655 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3656 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3657 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3658 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3659 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3660 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3661 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3662 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3663 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3664 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3665 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3666 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3667 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3668 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3669 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3670 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3671 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3672 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3673 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3674 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3675 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3676 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3677 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3678 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3679 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3680 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3681 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3682 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3683 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3684 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3685 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3686 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3687 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3688 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3689 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3690 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3691 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3692 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3693 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3694 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3695 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3696 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3697 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3698 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3699 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3700 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3701 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3702 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3703 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3704 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3705 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3706 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3707 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3708 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3709 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3710 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3711 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3712 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3713 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3714 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3715 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3716 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3717 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3718 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3719 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3720 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3721 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3722 ( .A(x[17]), .Z(n815) );
  IV U3723 ( .A(n814), .Z(n686) );
  AND U3724 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3725 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3726 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3727 ( .A(n685), .B(n684), .Z(n749) );
  IV U3728 ( .A(n749), .Z(n695) );
  XNOR U3729 ( .A(n695), .B(n814), .Z(n748) );
  IV U3730 ( .A(x[23]), .Z(n687) );
  XNOR U3731 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3732 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3733 ( .A(n687), .B(n686), .Z(n694) );
  IV U3734 ( .A(n694), .Z(n778) );
  XOR U3735 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3736 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3737 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3738 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3739 ( .A(n688), .Z(n753) );
  NANDN U3740 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3741 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3742 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3743 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3744 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3745 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3746 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3747 ( .A(n693), .B(n692), .Z(n729) );
  IV U3748 ( .A(n729), .Z(n735) );
  AND U3749 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3750 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3751 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3752 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3753 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3754 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3755 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3756 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3757 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3758 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3759 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3760 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3761 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3762 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3763 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3764 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3765 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3766 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3767 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3768 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3769 ( .A(n735), .B(n708), .Z(n719) );
  IV U3770 ( .A(n725), .Z(n726) );
  IV U3771 ( .A(n727), .Z(n733) );
  XOR U3772 ( .A(n709), .B(n763), .Z(n712) );
  AND U3773 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3774 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3775 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3776 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3777 ( .A(n716), .B(n715), .Z(n737) );
  IV U3778 ( .A(n737), .Z(n732) );
  XOR U3779 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3780 ( .A(n726), .B(n717), .Z(n718) );
  AND U3781 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3782 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3783 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3784 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3785 ( .A(n727), .B(n721), .Z(n722) );
  AND U3786 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3787 ( .A(n822), .B(n779), .Z(n754) );
  OR U3788 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3789 ( .A(n735), .B(n725), .Z(n731) );
  AND U3790 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3791 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3792 ( .A(n729), .B(n728), .Z(n730) );
  AND U3793 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3794 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3795 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3796 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3797 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3798 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3799 ( .A(n769), .B(n754), .Z(n756) );
  OR U3800 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3801 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3802 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3803 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3804 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3805 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3806 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3807 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3808 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3809 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3810 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3811 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3812 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3813 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3814 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3815 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3816 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3817 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3818 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3819 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3820 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3821 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3822 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3823 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3824 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3825 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3826 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3827 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3828 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3829 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3830 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3831 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3832 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3833 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3834 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3835 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3836 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3837 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3838 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3839 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3840 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3841 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3842 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3843 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3844 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3845 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3846 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3847 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3848 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3849 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3850 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3851 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3852 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3853 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3854 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3855 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3856 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3857 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3858 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3859 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3860 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3861 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3862 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3863 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3864 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3865 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3866 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3867 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3868 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3869 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3870 ( .A(x[25]), .Z(n939) );
  XOR U3871 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3872 ( .A(n938), .Z(n835) );
  AND U3873 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3874 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3875 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3876 ( .A(n834), .B(n833), .Z(n898) );
  IV U3877 ( .A(n898), .Z(n844) );
  XNOR U3878 ( .A(n844), .B(n938), .Z(n897) );
  IV U3879 ( .A(x[31]), .Z(n836) );
  XNOR U3880 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3881 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3882 ( .A(n836), .B(n835), .Z(n843) );
  IV U3883 ( .A(n843), .Z(n927) );
  XOR U3884 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3885 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3886 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3887 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3888 ( .A(n837), .Z(n902) );
  NANDN U3889 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3890 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3891 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3892 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3893 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3894 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3895 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3896 ( .A(n842), .B(n841), .Z(n878) );
  IV U3897 ( .A(n878), .Z(n884) );
  AND U3898 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3899 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3900 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3901 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3902 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3903 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3904 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3905 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3906 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3907 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3908 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3909 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3910 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3911 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3912 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3913 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3914 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3915 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3916 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3917 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3918 ( .A(n884), .B(n857), .Z(n868) );
  IV U3919 ( .A(n874), .Z(n875) );
  IV U3920 ( .A(n876), .Z(n882) );
  XOR U3921 ( .A(n858), .B(n912), .Z(n861) );
  AND U3922 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3923 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3924 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3925 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3926 ( .A(n865), .B(n864), .Z(n886) );
  IV U3927 ( .A(n886), .Z(n881) );
  XOR U3928 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3929 ( .A(n875), .B(n866), .Z(n867) );
  AND U3930 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3931 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3932 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3933 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3934 ( .A(n876), .B(n870), .Z(n871) );
  AND U3935 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3936 ( .A(n946), .B(n928), .Z(n903) );
  OR U3937 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3938 ( .A(n884), .B(n874), .Z(n880) );
  AND U3939 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3940 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3941 ( .A(n878), .B(n877), .Z(n879) );
  AND U3942 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3943 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3944 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3945 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3946 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3947 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3948 ( .A(n918), .B(n903), .Z(n905) );
  OR U3949 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3950 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3951 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3952 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3953 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3954 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3955 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3956 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3957 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3958 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3959 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3960 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3961 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3962 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3963 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3964 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3965 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3966 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3967 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3968 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3969 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3970 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3971 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3972 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3973 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3974 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3975 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3976 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3977 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3978 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3979 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3980 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3981 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3982 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3983 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3984 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3985 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3986 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3987 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3988 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3989 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3990 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3991 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3992 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3993 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3994 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3995 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3996 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3997 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3998 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3999 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4000 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4001 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4002 ( .A(x[33]), .Z(n1065) );
  XOR U4003 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4004 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4005 ( .A(n1064), .Z(n961) );
  AND U4006 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4007 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4008 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4009 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4010 ( .A(n1024), .Z(n970) );
  XNOR U4011 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4012 ( .A(x[39]), .Z(n962) );
  XNOR U4013 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4014 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4015 ( .A(n962), .B(n961), .Z(n969) );
  IV U4016 ( .A(n969), .Z(n1053) );
  XOR U4017 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4018 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4019 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4020 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4021 ( .A(n963), .Z(n1028) );
  NANDN U4022 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4023 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4024 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4025 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4026 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4027 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4028 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4029 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4030 ( .A(n1004), .Z(n1010) );
  AND U4031 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4032 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4033 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4035 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4036 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4037 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4038 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4039 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4040 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4041 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4042 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4043 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4044 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4045 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4046 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4047 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4048 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4049 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4050 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4051 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4052 ( .A(n1000), .Z(n1001) );
  IV U4053 ( .A(n1002), .Z(n1008) );
  XOR U4054 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4055 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4056 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4057 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4058 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4059 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4060 ( .A(n1012), .Z(n1007) );
  XOR U4061 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4062 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4063 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4064 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4065 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4066 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4067 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4068 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4069 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4070 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4071 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4072 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4073 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4074 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4075 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4076 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4077 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4078 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4079 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4080 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4081 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4082 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4083 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4084 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4085 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4086 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4087 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4088 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4089 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4090 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4091 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4092 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4093 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4094 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4095 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4096 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4097 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4098 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4099 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4100 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4101 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4102 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4103 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4104 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4105 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4106 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4107 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4108 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4109 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4110 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4111 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4112 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4113 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4114 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4115 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4116 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4117 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4118 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4119 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4120 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4121 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4122 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4123 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4124 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4125 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4126 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4127 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4128 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4129 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4130 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4131 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4132 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4133 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4134 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4135 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4136 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4137 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4138 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4139 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4140 ( .A(x[41]), .Z(n1199) );
  XOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4142 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4143 ( .A(n1198), .Z(n1095) );
  AND U4144 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4145 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4146 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4147 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4148 ( .A(n1158), .Z(n1104) );
  XNOR U4149 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4150 ( .A(x[47]), .Z(n1096) );
  XNOR U4151 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4152 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4153 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4154 ( .A(n1103), .Z(n1187) );
  XOR U4155 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4156 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4157 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4158 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4159 ( .A(n1097), .Z(n1162) );
  NANDN U4160 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4161 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4162 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4164 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4165 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4166 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4167 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4168 ( .A(n1138), .Z(n1144) );
  AND U4169 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4170 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4171 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4172 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4173 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4174 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4175 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4176 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4177 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4178 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4179 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4180 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4181 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4182 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4183 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4184 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4185 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4186 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4187 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4188 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4189 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4190 ( .A(n1134), .Z(n1135) );
  IV U4191 ( .A(n1136), .Z(n1142) );
  XOR U4192 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4193 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4194 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4195 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4196 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4197 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4198 ( .A(n1146), .Z(n1141) );
  XOR U4199 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4200 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4201 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4202 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4203 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4204 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4205 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4206 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4207 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4208 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4209 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4210 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4211 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4212 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4213 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4214 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4215 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4216 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4217 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4218 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4219 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4220 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4221 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4222 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4223 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4224 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4225 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4226 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4227 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4228 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4229 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4230 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4231 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4232 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4233 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4234 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4235 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4236 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4237 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4238 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4239 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4240 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4241 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4242 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4243 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4244 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4245 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4246 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4247 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4248 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4249 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4250 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4251 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4252 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4253 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4254 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4255 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4256 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4257 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4258 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4259 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4260 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4261 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4262 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4263 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4264 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4265 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4266 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4267 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4268 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4269 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4270 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4271 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4272 ( .A(x[49]), .Z(n1324) );
  XOR U4273 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4274 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4275 ( .A(n1323), .Z(n1219) );
  AND U4276 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4277 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4278 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4279 ( .A(n1282), .Z(n1228) );
  XNOR U4280 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4281 ( .A(x[55]), .Z(n1220) );
  XNOR U4282 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4283 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4284 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4285 ( .A(n1227), .Z(n1312) );
  XOR U4286 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4287 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4288 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4289 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4290 ( .A(n1221), .Z(n1286) );
  NANDN U4291 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4292 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4293 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4294 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4295 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4296 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4297 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4298 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4299 ( .A(n1262), .Z(n1268) );
  AND U4300 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4301 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4302 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4303 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4304 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4305 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4306 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4307 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4308 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4309 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4310 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4311 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4312 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4313 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4314 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4315 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4316 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4317 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4318 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4319 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4320 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4321 ( .A(n1258), .Z(n1259) );
  IV U4322 ( .A(n1260), .Z(n1266) );
  XOR U4323 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4324 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4325 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4326 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4327 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4328 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4329 ( .A(n1270), .Z(n1265) );
  XOR U4330 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4331 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4332 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4333 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4334 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4335 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4336 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4337 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4338 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4339 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4340 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4341 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4342 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4343 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4344 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4345 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4346 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4347 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4348 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4349 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4350 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4351 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4352 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4353 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4354 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4355 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4356 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4357 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4358 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4359 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4360 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4361 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4362 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4363 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4364 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4365 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4366 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4367 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4368 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4369 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4370 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4371 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4372 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4373 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4374 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4375 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4376 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4377 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4378 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4379 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4380 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4381 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4382 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4383 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4384 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4385 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4386 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4387 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4388 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4389 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4390 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4391 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4392 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4393 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4394 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4395 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4396 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4397 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4398 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4399 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4400 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4401 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4402 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4403 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4404 ( .A(x[57]), .Z(n1462) );
  XOR U4405 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4406 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4407 ( .A(n1461), .Z(n1344) );
  AND U4408 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4409 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4410 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4411 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4412 ( .A(n1407), .Z(n1353) );
  XNOR U4413 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4414 ( .A(x[63]), .Z(n1345) );
  XNOR U4415 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4416 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4417 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4418 ( .A(n1352), .Z(n1436) );
  XOR U4419 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4420 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4421 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4422 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4423 ( .A(n1346), .Z(n1411) );
  NANDN U4424 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4425 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4426 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4427 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4428 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4429 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4430 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4431 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4432 ( .A(n1387), .Z(n1393) );
  AND U4433 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4434 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4435 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4436 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4437 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4438 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4439 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4440 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4441 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4442 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4443 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4444 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4445 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4446 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4447 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4448 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4449 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4450 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4451 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4452 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4453 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4454 ( .A(n1383), .Z(n1384) );
  IV U4455 ( .A(n1385), .Z(n1391) );
  XOR U4456 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4457 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4458 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4459 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4460 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4461 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4462 ( .A(n1395), .Z(n1390) );
  XOR U4463 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4464 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4465 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4466 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4467 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4468 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4469 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4470 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4471 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4472 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4473 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4474 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4475 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4476 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4477 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4478 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4479 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4480 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4481 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4482 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4483 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4484 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4485 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4486 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4487 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4488 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4489 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4490 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4491 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4492 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4493 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4494 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4495 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4496 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4497 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4498 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4499 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4500 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4501 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4502 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4503 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4504 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4505 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4506 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4507 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4508 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4509 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4510 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4511 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4512 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4513 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4514 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4515 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4516 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4517 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4518 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4519 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4520 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4521 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4522 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4523 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4524 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4525 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4526 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4527 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4528 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4529 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4530 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4531 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4532 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4533 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4534 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4535 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4536 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4537 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4538 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4539 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4540 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4541 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4542 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4543 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4544 ( .A(x[65]), .Z(n1586) );
  XOR U4545 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4546 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4547 ( .A(n1585), .Z(n1482) );
  AND U4548 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4549 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4550 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4551 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4552 ( .A(n1545), .Z(n1491) );
  XNOR U4553 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4554 ( .A(x[71]), .Z(n1483) );
  XNOR U4555 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4556 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4557 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4558 ( .A(n1490), .Z(n1574) );
  XOR U4559 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4560 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4561 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4562 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4563 ( .A(n1484), .Z(n1549) );
  NANDN U4564 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4565 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4566 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4567 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4568 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4569 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4570 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4571 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4572 ( .A(n1525), .Z(n1531) );
  AND U4573 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4574 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4575 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4576 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4577 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4578 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4579 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4580 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4581 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4582 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4583 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4584 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4585 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4586 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4587 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4588 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4589 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4590 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4591 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4592 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4593 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4594 ( .A(n1521), .Z(n1522) );
  IV U4595 ( .A(n1523), .Z(n1529) );
  XOR U4596 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4597 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4598 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4599 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4600 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4601 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4602 ( .A(n1533), .Z(n1528) );
  XOR U4603 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4604 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4605 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4606 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4607 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4608 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4609 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4610 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4611 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4612 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4613 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4614 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4615 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4616 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4617 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4618 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4619 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4620 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4621 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4622 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4623 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4624 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4625 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4626 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4627 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4628 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4629 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4630 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4631 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4632 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4633 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4634 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4635 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4636 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4637 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4638 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4639 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4640 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4641 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4642 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4643 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4644 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4645 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4646 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4647 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4648 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4649 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4650 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4651 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4652 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4653 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4654 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4655 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4656 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4657 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4658 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4659 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4660 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4661 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4662 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4663 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4664 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4665 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4666 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4667 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4668 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4669 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4670 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4671 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4672 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4673 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4674 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4675 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4676 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4677 ( .A(x[73]), .Z(n1712) );
  XOR U4678 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4679 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4680 ( .A(n1711), .Z(n1608) );
  AND U4681 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4682 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4683 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4684 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4685 ( .A(n1671), .Z(n1617) );
  XNOR U4686 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4687 ( .A(x[79]), .Z(n1609) );
  XNOR U4688 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4689 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4690 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4691 ( .A(n1616), .Z(n1700) );
  XOR U4692 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4693 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4694 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4695 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4696 ( .A(n1610), .Z(n1675) );
  NANDN U4697 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4698 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4699 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4700 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4701 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4702 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4703 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4704 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4705 ( .A(n1651), .Z(n1657) );
  AND U4706 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4707 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4708 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4709 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4710 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4711 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4712 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4713 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4714 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4715 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4716 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4717 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4718 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4719 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4720 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4721 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4722 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4723 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4724 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4725 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4726 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4727 ( .A(n1647), .Z(n1648) );
  IV U4728 ( .A(n1649), .Z(n1655) );
  XOR U4729 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4730 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4731 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4732 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4733 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4734 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4735 ( .A(n1659), .Z(n1654) );
  XOR U4736 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4737 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4738 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4739 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4740 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4741 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4742 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4743 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4744 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4745 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4746 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4747 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4748 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4749 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4750 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4751 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4752 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4753 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4754 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4755 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4756 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4757 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4758 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4759 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4760 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4761 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4762 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4763 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4764 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4765 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4766 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4767 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4768 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4769 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4770 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4771 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4772 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4773 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4774 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4775 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4776 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4777 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4778 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4779 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4780 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4781 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4782 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4783 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4784 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4785 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4786 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4787 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4788 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4789 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4790 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4791 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4792 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4793 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4794 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4795 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4796 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4797 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4798 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4799 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4800 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4801 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4802 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4803 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4804 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4805 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4806 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4807 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4808 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4809 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4810 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4811 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4812 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module aes_comb ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [1279:0] key;
  output [127:0] out;
  input clk, rst;
  wire   \w1[9][127] , \w1[9][126] , \w1[9][125] , \w1[9][124] , \w1[9][123] ,
         \w1[9][122] , \w1[9][121] , \w1[9][120] , \w1[9][119] , \w1[9][118] ,
         \w1[9][117] , \w1[9][116] , \w1[9][115] , \w1[9][114] , \w1[9][113] ,
         \w1[9][112] , \w1[9][111] , \w1[9][110] , \w1[9][109] , \w1[9][108] ,
         \w1[9][107] , \w1[9][106] , \w1[9][105] , \w1[9][104] , \w1[9][103] ,
         \w1[9][102] , \w1[9][101] , \w1[9][100] , \w1[9][99] , \w1[9][98] ,
         \w1[9][97] , \w1[9][96] , \w1[9][95] , \w1[9][94] , \w1[9][93] ,
         \w1[9][92] , \w1[9][91] , \w1[9][90] , \w1[9][89] , \w1[9][88] ,
         \w1[9][87] , \w1[9][86] , \w1[9][85] , \w1[9][84] , \w1[9][83] ,
         \w1[9][82] , \w1[9][81] , \w1[9][80] , \w1[9][79] , \w1[9][78] ,
         \w1[9][77] , \w1[9][76] , \w1[9][75] , \w1[9][74] , \w1[9][73] ,
         \w1[9][72] , \w1[9][71] , \w1[9][70] , \w1[9][69] , \w1[9][68] ,
         \w1[9][67] , \w1[9][66] , \w1[9][65] , \w1[9][64] , \w1[9][63] ,
         \w1[9][62] , \w1[9][61] , \w1[9][60] , \w1[9][59] , \w1[9][58] ,
         \w1[9][57] , \w1[9][56] , \w1[9][55] , \w1[9][54] , \w1[9][53] ,
         \w1[9][52] , \w1[9][51] , \w1[9][50] , \w1[9][49] , \w1[9][48] ,
         \w1[9][47] , \w1[9][46] , \w1[9][45] , \w1[9][44] , \w1[9][43] ,
         \w1[9][42] , \w1[9][41] , \w1[9][40] , \w1[9][39] , \w1[9][38] ,
         \w1[9][37] , \w1[9][36] , \w1[9][35] , \w1[9][34] , \w1[9][33] ,
         \w1[9][32] , \w1[9][31] , \w1[9][30] , \w1[9][29] , \w1[9][28] ,
         \w1[9][27] , \w1[9][26] , \w1[9][25] , \w1[9][24] , \w1[9][23] ,
         \w1[9][22] , \w1[9][21] , \w1[9][20] , \w1[9][19] , \w1[9][18] ,
         \w1[9][17] , \w1[9][16] , \w1[9][15] , \w1[9][14] , \w1[9][13] ,
         \w1[9][12] , \w1[9][11] , \w1[9][10] , \w1[9][9] , \w1[9][8] ,
         \w1[9][7] , \w1[9][6] , \w1[9][5] , \w1[9][4] , \w1[9][3] ,
         \w1[9][2] , \w1[9][1] , \w1[9][0] , \w1[8][127] , \w1[8][126] ,
         \w1[8][125] , \w1[8][124] , \w1[8][123] , \w1[8][122] , \w1[8][121] ,
         \w1[8][120] , \w1[8][119] , \w1[8][118] , \w1[8][117] , \w1[8][116] ,
         \w1[8][115] , \w1[8][114] , \w1[8][113] , \w1[8][112] , \w1[8][111] ,
         \w1[8][110] , \w1[8][109] , \w1[8][108] , \w1[8][107] , \w1[8][106] ,
         \w1[8][105] , \w1[8][104] , \w1[8][103] , \w1[8][102] , \w1[8][101] ,
         \w1[8][100] , \w1[8][99] , \w1[8][98] , \w1[8][97] , \w1[8][96] ,
         \w1[8][95] , \w1[8][94] , \w1[8][93] , \w1[8][92] , \w1[8][91] ,
         \w1[8][90] , \w1[8][89] , \w1[8][88] , \w1[8][87] , \w1[8][86] ,
         \w1[8][85] , \w1[8][84] , \w1[8][83] , \w1[8][82] , \w1[8][81] ,
         \w1[8][80] , \w1[8][79] , \w1[8][78] , \w1[8][77] , \w1[8][76] ,
         \w1[8][75] , \w1[8][74] , \w1[8][73] , \w1[8][72] , \w1[8][71] ,
         \w1[8][70] , \w1[8][69] , \w1[8][68] , \w1[8][67] , \w1[8][66] ,
         \w1[8][65] , \w1[8][64] , \w1[8][63] , \w1[8][62] , \w1[8][61] ,
         \w1[8][60] , \w1[8][59] , \w1[8][58] , \w1[8][57] , \w1[8][56] ,
         \w1[8][55] , \w1[8][54] , \w1[8][53] , \w1[8][52] , \w1[8][51] ,
         \w1[8][50] , \w1[8][49] , \w1[8][48] , \w1[8][47] , \w1[8][46] ,
         \w1[8][45] , \w1[8][44] , \w1[8][43] , \w1[8][42] , \w1[8][41] ,
         \w1[8][40] , \w1[8][39] , \w1[8][38] , \w1[8][37] , \w1[8][36] ,
         \w1[8][35] , \w1[8][34] , \w1[8][33] , \w1[8][32] , \w1[8][31] ,
         \w1[8][30] , \w1[8][29] , \w1[8][28] , \w1[8][27] , \w1[8][26] ,
         \w1[8][25] , \w1[8][24] , \w1[8][23] , \w1[8][22] , \w1[8][21] ,
         \w1[8][20] , \w1[8][19] , \w1[8][18] , \w1[8][17] , \w1[8][16] ,
         \w1[8][15] , \w1[8][14] , \w1[8][13] , \w1[8][12] , \w1[8][11] ,
         \w1[8][10] , \w1[8][9] , \w1[8][8] , \w1[8][7] , \w1[8][6] ,
         \w1[8][5] , \w1[8][4] , \w1[8][3] , \w1[8][2] , \w1[8][1] ,
         \w1[8][0] , \w1[7][127] , \w1[7][126] , \w1[7][125] , \w1[7][124] ,
         \w1[7][123] , \w1[7][122] , \w1[7][121] , \w1[7][120] , \w1[7][119] ,
         \w1[7][118] , \w1[7][117] , \w1[7][116] , \w1[7][115] , \w1[7][114] ,
         \w1[7][113] , \w1[7][112] , \w1[7][111] , \w1[7][110] , \w1[7][109] ,
         \w1[7][108] , \w1[7][107] , \w1[7][106] , \w1[7][105] , \w1[7][104] ,
         \w1[7][103] , \w1[7][102] , \w1[7][101] , \w1[7][100] , \w1[7][99] ,
         \w1[7][98] , \w1[7][97] , \w1[7][96] , \w1[7][95] , \w1[7][94] ,
         \w1[7][93] , \w1[7][92] , \w1[7][91] , \w1[7][90] , \w1[7][89] ,
         \w1[7][88] , \w1[7][87] , \w1[7][86] , \w1[7][85] , \w1[7][84] ,
         \w1[7][83] , \w1[7][82] , \w1[7][81] , \w1[7][80] , \w1[7][79] ,
         \w1[7][78] , \w1[7][77] , \w1[7][76] , \w1[7][75] , \w1[7][74] ,
         \w1[7][73] , \w1[7][72] , \w1[7][71] , \w1[7][70] , \w1[7][69] ,
         \w1[7][68] , \w1[7][67] , \w1[7][66] , \w1[7][65] , \w1[7][64] ,
         \w1[7][63] , \w1[7][62] , \w1[7][61] , \w1[7][60] , \w1[7][59] ,
         \w1[7][58] , \w1[7][57] , \w1[7][56] , \w1[7][55] , \w1[7][54] ,
         \w1[7][53] , \w1[7][52] , \w1[7][51] , \w1[7][50] , \w1[7][49] ,
         \w1[7][48] , \w1[7][47] , \w1[7][46] , \w1[7][45] , \w1[7][44] ,
         \w1[7][43] , \w1[7][42] , \w1[7][41] , \w1[7][40] , \w1[7][39] ,
         \w1[7][38] , \w1[7][37] , \w1[7][36] , \w1[7][35] , \w1[7][34] ,
         \w1[7][33] , \w1[7][32] , \w1[7][31] , \w1[7][30] , \w1[7][29] ,
         \w1[7][28] , \w1[7][27] , \w1[7][26] , \w1[7][25] , \w1[7][24] ,
         \w1[7][23] , \w1[7][22] , \w1[7][21] , \w1[7][20] , \w1[7][19] ,
         \w1[7][18] , \w1[7][17] , \w1[7][16] , \w1[7][15] , \w1[7][14] ,
         \w1[7][13] , \w1[7][12] , \w1[7][11] , \w1[7][10] , \w1[7][9] ,
         \w1[7][8] , \w1[7][7] , \w1[7][6] , \w1[7][5] , \w1[7][4] ,
         \w1[7][3] , \w1[7][2] , \w1[7][1] , \w1[7][0] , \w1[6][127] ,
         \w1[6][126] , \w1[6][125] , \w1[6][124] , \w1[6][123] , \w1[6][122] ,
         \w1[6][121] , \w1[6][120] , \w1[6][119] , \w1[6][118] , \w1[6][117] ,
         \w1[6][116] , \w1[6][115] , \w1[6][114] , \w1[6][113] , \w1[6][112] ,
         \w1[6][111] , \w1[6][110] , \w1[6][109] , \w1[6][108] , \w1[6][107] ,
         \w1[6][106] , \w1[6][105] , \w1[6][104] , \w1[6][103] , \w1[6][102] ,
         \w1[6][101] , \w1[6][100] , \w1[6][99] , \w1[6][98] , \w1[6][97] ,
         \w1[6][96] , \w1[6][95] , \w1[6][94] , \w1[6][93] , \w1[6][92] ,
         \w1[6][91] , \w1[6][90] , \w1[6][89] , \w1[6][88] , \w1[6][87] ,
         \w1[6][86] , \w1[6][85] , \w1[6][84] , \w1[6][83] , \w1[6][82] ,
         \w1[6][81] , \w1[6][80] , \w1[6][79] , \w1[6][78] , \w1[6][77] ,
         \w1[6][76] , \w1[6][75] , \w1[6][74] , \w1[6][73] , \w1[6][72] ,
         \w1[6][71] , \w1[6][70] , \w1[6][69] , \w1[6][68] , \w1[6][67] ,
         \w1[6][66] , \w1[6][65] , \w1[6][64] , \w1[6][63] , \w1[6][62] ,
         \w1[6][61] , \w1[6][60] , \w1[6][59] , \w1[6][58] , \w1[6][57] ,
         \w1[6][56] , \w1[6][55] , \w1[6][54] , \w1[6][53] , \w1[6][52] ,
         \w1[6][51] , \w1[6][50] , \w1[6][49] , \w1[6][48] , \w1[6][47] ,
         \w1[6][46] , \w1[6][45] , \w1[6][44] , \w1[6][43] , \w1[6][42] ,
         \w1[6][41] , \w1[6][40] , \w1[6][39] , \w1[6][38] , \w1[6][37] ,
         \w1[6][36] , \w1[6][35] , \w1[6][34] , \w1[6][33] , \w1[6][32] ,
         \w1[6][31] , \w1[6][30] , \w1[6][29] , \w1[6][28] , \w1[6][27] ,
         \w1[6][26] , \w1[6][25] , \w1[6][24] , \w1[6][23] , \w1[6][22] ,
         \w1[6][21] , \w1[6][20] , \w1[6][19] , \w1[6][18] , \w1[6][17] ,
         \w1[6][16] , \w1[6][15] , \w1[6][14] , \w1[6][13] , \w1[6][12] ,
         \w1[6][11] , \w1[6][10] , \w1[6][9] , \w1[6][8] , \w1[6][7] ,
         \w1[6][6] , \w1[6][5] , \w1[6][4] , \w1[6][3] , \w1[6][2] ,
         \w1[6][1] , \w1[6][0] , \w1[5][127] , \w1[5][126] , \w1[5][125] ,
         \w1[5][124] , \w1[5][123] , \w1[5][122] , \w1[5][121] , \w1[5][120] ,
         \w1[5][119] , \w1[5][118] , \w1[5][117] , \w1[5][116] , \w1[5][115] ,
         \w1[5][114] , \w1[5][113] , \w1[5][112] , \w1[5][111] , \w1[5][110] ,
         \w1[5][109] , \w1[5][108] , \w1[5][107] , \w1[5][106] , \w1[5][105] ,
         \w1[5][104] , \w1[5][103] , \w1[5][102] , \w1[5][101] , \w1[5][100] ,
         \w1[5][99] , \w1[5][98] , \w1[5][97] , \w1[5][96] , \w1[5][95] ,
         \w1[5][94] , \w1[5][93] , \w1[5][92] , \w1[5][91] , \w1[5][90] ,
         \w1[5][89] , \w1[5][88] , \w1[5][87] , \w1[5][86] , \w1[5][85] ,
         \w1[5][84] , \w1[5][83] , \w1[5][82] , \w1[5][81] , \w1[5][80] ,
         \w1[5][79] , \w1[5][78] , \w1[5][77] , \w1[5][76] , \w1[5][75] ,
         \w1[5][74] , \w1[5][73] , \w1[5][72] , \w1[5][71] , \w1[5][70] ,
         \w1[5][69] , \w1[5][68] , \w1[5][67] , \w1[5][66] , \w1[5][65] ,
         \w1[5][64] , \w1[5][63] , \w1[5][62] , \w1[5][61] , \w1[5][60] ,
         \w1[5][59] , \w1[5][58] , \w1[5][57] , \w1[5][56] , \w1[5][55] ,
         \w1[5][54] , \w1[5][53] , \w1[5][52] , \w1[5][51] , \w1[5][50] ,
         \w1[5][49] , \w1[5][48] , \w1[5][47] , \w1[5][46] , \w1[5][45] ,
         \w1[5][44] , \w1[5][43] , \w1[5][42] , \w1[5][41] , \w1[5][40] ,
         \w1[5][39] , \w1[5][38] , \w1[5][37] , \w1[5][36] , \w1[5][35] ,
         \w1[5][34] , \w1[5][33] , \w1[5][32] , \w1[5][31] , \w1[5][30] ,
         \w1[5][29] , \w1[5][28] , \w1[5][27] , \w1[5][26] , \w1[5][25] ,
         \w1[5][24] , \w1[5][23] , \w1[5][22] , \w1[5][21] , \w1[5][20] ,
         \w1[5][19] , \w1[5][18] , \w1[5][17] , \w1[5][16] , \w1[5][15] ,
         \w1[5][14] , \w1[5][13] , \w1[5][12] , \w1[5][11] , \w1[5][10] ,
         \w1[5][9] , \w1[5][8] , \w1[5][7] , \w1[5][6] , \w1[5][5] ,
         \w1[5][4] , \w1[5][3] , \w1[5][2] , \w1[5][1] , \w1[5][0] ,
         \w1[4][127] , \w1[4][126] , \w1[4][125] , \w1[4][124] , \w1[4][123] ,
         \w1[4][122] , \w1[4][121] , \w1[4][120] , \w1[4][119] , \w1[4][118] ,
         \w1[4][117] , \w1[4][116] , \w1[4][115] , \w1[4][114] , \w1[4][113] ,
         \w1[4][112] , \w1[4][111] , \w1[4][110] , \w1[4][109] , \w1[4][108] ,
         \w1[4][107] , \w1[4][106] , \w1[4][105] , \w1[4][104] , \w1[4][103] ,
         \w1[4][102] , \w1[4][101] , \w1[4][100] , \w1[4][99] , \w1[4][98] ,
         \w1[4][97] , \w1[4][96] , \w1[4][95] , \w1[4][94] , \w1[4][93] ,
         \w1[4][92] , \w1[4][91] , \w1[4][90] , \w1[4][89] , \w1[4][88] ,
         \w1[4][87] , \w1[4][86] , \w1[4][85] , \w1[4][84] , \w1[4][83] ,
         \w1[4][82] , \w1[4][81] , \w1[4][80] , \w1[4][79] , \w1[4][78] ,
         \w1[4][77] , \w1[4][76] , \w1[4][75] , \w1[4][74] , \w1[4][73] ,
         \w1[4][72] , \w1[4][71] , \w1[4][70] , \w1[4][69] , \w1[4][68] ,
         \w1[4][67] , \w1[4][66] , \w1[4][65] , \w1[4][64] , \w1[4][63] ,
         \w1[4][62] , \w1[4][61] , \w1[4][60] , \w1[4][59] , \w1[4][58] ,
         \w1[4][57] , \w1[4][56] , \w1[4][55] , \w1[4][54] , \w1[4][53] ,
         \w1[4][52] , \w1[4][51] , \w1[4][50] , \w1[4][49] , \w1[4][48] ,
         \w1[4][47] , \w1[4][46] , \w1[4][45] , \w1[4][44] , \w1[4][43] ,
         \w1[4][42] , \w1[4][41] , \w1[4][40] , \w1[4][39] , \w1[4][38] ,
         \w1[4][37] , \w1[4][36] , \w1[4][35] , \w1[4][34] , \w1[4][33] ,
         \w1[4][32] , \w1[4][31] , \w1[4][30] , \w1[4][29] , \w1[4][28] ,
         \w1[4][27] , \w1[4][26] , \w1[4][25] , \w1[4][24] , \w1[4][23] ,
         \w1[4][22] , \w1[4][21] , \w1[4][20] , \w1[4][19] , \w1[4][18] ,
         \w1[4][17] , \w1[4][16] , \w1[4][15] , \w1[4][14] , \w1[4][13] ,
         \w1[4][12] , \w1[4][11] , \w1[4][10] , \w1[4][9] , \w1[4][8] ,
         \w1[4][7] , \w1[4][6] , \w1[4][5] , \w1[4][4] , \w1[4][3] ,
         \w1[4][2] , \w1[4][1] , \w1[4][0] , \w1[3][127] , \w1[3][126] ,
         \w1[3][125] , \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] ,
         \w1[3][120] , \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] ,
         \w1[3][115] , \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] ,
         \w1[3][110] , \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] ,
         \w1[3][105] , \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] ,
         \w1[3][100] , \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] ,
         \w1[3][95] , \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] ,
         \w1[3][90] , \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] ,
         \w1[3][85] , \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] ,
         \w1[3][80] , \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] ,
         \w1[3][75] , \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] ,
         \w1[3][70] , \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] ,
         \w1[3][65] , \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] ,
         \w1[3][60] , \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] ,
         \w1[3][55] , \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] ,
         \w1[3][50] , \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] ,
         \w1[3][45] , \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] ,
         \w1[3][40] , \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] ,
         \w1[3][35] , \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] ,
         \w1[3][30] , \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] ,
         \w1[3][25] , \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] ,
         \w1[3][20] , \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] ,
         \w1[3][15] , \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] ,
         \w1[3][10] , \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] ,
         \w1[3][5] , \w1[3][4] , \w1[3][3] , \w1[3][2] , \w1[3][1] ,
         \w1[3][0] , \w1[2][127] , \w1[2][126] , \w1[2][125] , \w1[2][124] ,
         \w1[2][123] , \w1[2][122] , \w1[2][121] , \w1[2][120] , \w1[2][119] ,
         \w1[2][118] , \w1[2][117] , \w1[2][116] , \w1[2][115] , \w1[2][114] ,
         \w1[2][113] , \w1[2][112] , \w1[2][111] , \w1[2][110] , \w1[2][109] ,
         \w1[2][108] , \w1[2][107] , \w1[2][106] , \w1[2][105] , \w1[2][104] ,
         \w1[2][103] , \w1[2][102] , \w1[2][101] , \w1[2][100] , \w1[2][99] ,
         \w1[2][98] , \w1[2][97] , \w1[2][96] , \w1[2][95] , \w1[2][94] ,
         \w1[2][93] , \w1[2][92] , \w1[2][91] , \w1[2][90] , \w1[2][89] ,
         \w1[2][88] , \w1[2][87] , \w1[2][86] , \w1[2][85] , \w1[2][84] ,
         \w1[2][83] , \w1[2][82] , \w1[2][81] , \w1[2][80] , \w1[2][79] ,
         \w1[2][78] , \w1[2][77] , \w1[2][76] , \w1[2][75] , \w1[2][74] ,
         \w1[2][73] , \w1[2][72] , \w1[2][71] , \w1[2][70] , \w1[2][69] ,
         \w1[2][68] , \w1[2][67] , \w1[2][66] , \w1[2][65] , \w1[2][64] ,
         \w1[2][63] , \w1[2][62] , \w1[2][61] , \w1[2][60] , \w1[2][59] ,
         \w1[2][58] , \w1[2][57] , \w1[2][56] , \w1[2][55] , \w1[2][54] ,
         \w1[2][53] , \w1[2][52] , \w1[2][51] , \w1[2][50] , \w1[2][49] ,
         \w1[2][48] , \w1[2][47] , \w1[2][46] , \w1[2][45] , \w1[2][44] ,
         \w1[2][43] , \w1[2][42] , \w1[2][41] , \w1[2][40] , \w1[2][39] ,
         \w1[2][38] , \w1[2][37] , \w1[2][36] , \w1[2][35] , \w1[2][34] ,
         \w1[2][33] , \w1[2][32] , \w1[2][31] , \w1[2][30] , \w1[2][29] ,
         \w1[2][28] , \w1[2][27] , \w1[2][26] , \w1[2][25] , \w1[2][24] ,
         \w1[2][23] , \w1[2][22] , \w1[2][21] , \w1[2][20] , \w1[2][19] ,
         \w1[2][18] , \w1[2][17] , \w1[2][16] , \w1[2][15] , \w1[2][14] ,
         \w1[2][13] , \w1[2][12] , \w1[2][11] , \w1[2][10] , \w1[2][9] ,
         \w1[2][8] , \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] ,
         \w1[2][3] , \w1[2][2] , \w1[2][1] , \w1[2][0] , \w1[1][127] ,
         \w1[1][126] , \w1[1][125] , \w1[1][124] , \w1[1][123] , \w1[1][122] ,
         \w1[1][121] , \w1[1][120] , \w1[1][119] , \w1[1][118] , \w1[1][117] ,
         \w1[1][116] , \w1[1][115] , \w1[1][114] , \w1[1][113] , \w1[1][112] ,
         \w1[1][111] , \w1[1][110] , \w1[1][109] , \w1[1][108] , \w1[1][107] ,
         \w1[1][106] , \w1[1][105] , \w1[1][104] , \w1[1][103] , \w1[1][102] ,
         \w1[1][101] , \w1[1][100] , \w1[1][99] , \w1[1][98] , \w1[1][97] ,
         \w1[1][96] , \w1[1][95] , \w1[1][94] , \w1[1][93] , \w1[1][92] ,
         \w1[1][91] , \w1[1][90] , \w1[1][89] , \w1[1][88] , \w1[1][87] ,
         \w1[1][86] , \w1[1][85] , \w1[1][84] , \w1[1][83] , \w1[1][82] ,
         \w1[1][81] , \w1[1][80] , \w1[1][79] , \w1[1][78] , \w1[1][77] ,
         \w1[1][76] , \w1[1][75] , \w1[1][74] , \w1[1][73] , \w1[1][72] ,
         \w1[1][71] , \w1[1][70] , \w1[1][69] , \w1[1][68] , \w1[1][67] ,
         \w1[1][66] , \w1[1][65] , \w1[1][64] , \w1[1][63] , \w1[1][62] ,
         \w1[1][61] , \w1[1][60] , \w1[1][59] , \w1[1][58] , \w1[1][57] ,
         \w1[1][56] , \w1[1][55] , \w1[1][54] , \w1[1][53] , \w1[1][52] ,
         \w1[1][51] , \w1[1][50] , \w1[1][49] , \w1[1][48] , \w1[1][47] ,
         \w1[1][46] , \w1[1][45] , \w1[1][44] , \w1[1][43] , \w1[1][42] ,
         \w1[1][41] , \w1[1][40] , \w1[1][39] , \w1[1][38] , \w1[1][37] ,
         \w1[1][36] , \w1[1][35] , \w1[1][34] , \w1[1][33] , \w1[1][32] ,
         \w1[1][31] , \w1[1][30] , \w1[1][29] , \w1[1][28] , \w1[1][27] ,
         \w1[1][26] , \w1[1][25] , \w1[1][24] , \w1[1][23] , \w1[1][22] ,
         \w1[1][21] , \w1[1][20] , \w1[1][19] , \w1[1][18] , \w1[1][17] ,
         \w1[1][16] , \w1[1][15] , \w1[1][14] , \w1[1][13] , \w1[1][12] ,
         \w1[1][11] , \w1[1][10] , \w1[1][9] , \w1[1][8] , \w1[1][7] ,
         \w1[1][6] , \w1[1][5] , \w1[1][4] , \w1[1][3] , \w1[1][2] ,
         \w1[1][1] , \w1[1][0] , \w1[0][127] , \w1[0][126] , \w1[0][125] ,
         \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] ,
         \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] ,
         \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] ,
         \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] ,
         \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] ,
         \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] ,
         \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] ,
         \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] ,
         \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] ,
         \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] ,
         \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] ,
         \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] ,
         \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] ,
         \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] ,
         \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] ,
         \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] ,
         \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] ,
         \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] ,
         \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] ,
         \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] ,
         \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] ,
         \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] ,
         \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] ,
         \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] ,
         \w1[0][4] , \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] ,
         \w3[9][127] , \w3[9][126] , \w3[9][125] , \w3[9][124] , \w3[9][123] ,
         \w3[9][122] , \w3[9][121] , \w3[9][120] , \w3[9][119] , \w3[9][118] ,
         \w3[9][117] , \w3[9][116] , \w3[9][115] , \w3[9][114] , \w3[9][113] ,
         \w3[9][112] , \w3[9][111] , \w3[9][110] , \w3[9][109] , \w3[9][108] ,
         \w3[9][107] , \w3[9][106] , \w3[9][105] , \w3[9][104] , \w3[9][103] ,
         \w3[9][102] , \w3[9][101] , \w3[9][100] , \w3[9][99] , \w3[9][98] ,
         \w3[9][97] , \w3[9][96] , \w3[9][95] , \w3[9][94] , \w3[9][93] ,
         \w3[9][92] , \w3[9][91] , \w3[9][90] , \w3[9][89] , \w3[9][88] ,
         \w3[9][87] , \w3[9][86] , \w3[9][85] , \w3[9][84] , \w3[9][83] ,
         \w3[9][82] , \w3[9][81] , \w3[9][80] , \w3[9][79] , \w3[9][78] ,
         \w3[9][77] , \w3[9][76] , \w3[9][75] , \w3[9][74] , \w3[9][73] ,
         \w3[9][72] , \w3[9][71] , \w3[9][70] , \w3[9][69] , \w3[9][68] ,
         \w3[9][67] , \w3[9][66] , \w3[9][65] , \w3[9][64] , \w3[9][63] ,
         \w3[9][62] , \w3[9][61] , \w3[9][60] , \w3[9][59] , \w3[9][58] ,
         \w3[9][57] , \w3[9][56] , \w3[9][55] , \w3[9][54] , \w3[9][53] ,
         \w3[9][52] , \w3[9][51] , \w3[9][50] , \w3[9][49] , \w3[9][48] ,
         \w3[9][47] , \w3[9][46] , \w3[9][45] , \w3[9][44] , \w3[9][43] ,
         \w3[9][42] , \w3[9][41] , \w3[9][40] , \w3[9][39] , \w3[9][38] ,
         \w3[9][37] , \w3[9][36] , \w3[9][35] , \w3[9][34] , \w3[9][33] ,
         \w3[9][32] , \w3[9][31] , \w3[9][30] , \w3[9][29] , \w3[9][28] ,
         \w3[9][27] , \w3[9][26] , \w3[9][25] , \w3[9][24] , \w3[9][23] ,
         \w3[9][22] , \w3[9][21] , \w3[9][20] , \w3[9][19] , \w3[9][18] ,
         \w3[9][17] , \w3[9][16] , \w3[9][15] , \w3[9][14] , \w3[9][13] ,
         \w3[9][12] , \w3[9][11] , \w3[9][10] , \w3[9][9] , \w3[9][8] ,
         \w3[9][7] , \w3[9][6] , \w3[9][5] , \w3[9][4] , \w3[9][3] ,
         \w3[9][2] , \w3[9][1] , \w3[9][0] , \w3[8][127] , \w3[8][126] ,
         \w3[8][125] , \w3[8][124] , \w3[8][123] , \w3[8][122] , \w3[8][121] ,
         \w3[8][120] , \w3[8][119] , \w3[8][118] , \w3[8][117] , \w3[8][116] ,
         \w3[8][115] , \w3[8][114] , \w3[8][113] , \w3[8][112] , \w3[8][111] ,
         \w3[8][110] , \w3[8][109] , \w3[8][108] , \w3[8][107] , \w3[8][106] ,
         \w3[8][105] , \w3[8][104] , \w3[8][103] , \w3[8][102] , \w3[8][101] ,
         \w3[8][100] , \w3[8][99] , \w3[8][98] , \w3[8][97] , \w3[8][96] ,
         \w3[8][95] , \w3[8][94] , \w3[8][93] , \w3[8][92] , \w3[8][91] ,
         \w3[8][90] , \w3[8][89] , \w3[8][88] , \w3[8][87] , \w3[8][86] ,
         \w3[8][85] , \w3[8][84] , \w3[8][83] , \w3[8][82] , \w3[8][81] ,
         \w3[8][80] , \w3[8][79] , \w3[8][78] , \w3[8][77] , \w3[8][76] ,
         \w3[8][75] , \w3[8][74] , \w3[8][73] , \w3[8][72] , \w3[8][71] ,
         \w3[8][70] , \w3[8][69] , \w3[8][68] , \w3[8][67] , \w3[8][66] ,
         \w3[8][65] , \w3[8][64] , \w3[8][63] , \w3[8][62] , \w3[8][61] ,
         \w3[8][60] , \w3[8][59] , \w3[8][58] , \w3[8][57] , \w3[8][56] ,
         \w3[8][55] , \w3[8][54] , \w3[8][53] , \w3[8][52] , \w3[8][51] ,
         \w3[8][50] , \w3[8][49] , \w3[8][48] , \w3[8][47] , \w3[8][46] ,
         \w3[8][45] , \w3[8][44] , \w3[8][43] , \w3[8][42] , \w3[8][41] ,
         \w3[8][40] , \w3[8][39] , \w3[8][38] , \w3[8][37] , \w3[8][36] ,
         \w3[8][35] , \w3[8][34] , \w3[8][33] , \w3[8][32] , \w3[8][31] ,
         \w3[8][30] , \w3[8][29] , \w3[8][28] , \w3[8][27] , \w3[8][26] ,
         \w3[8][25] , \w3[8][24] , \w3[8][23] , \w3[8][22] , \w3[8][21] ,
         \w3[8][20] , \w3[8][19] , \w3[8][18] , \w3[8][17] , \w3[8][16] ,
         \w3[8][15] , \w3[8][14] , \w3[8][13] , \w3[8][12] , \w3[8][11] ,
         \w3[8][10] , \w3[8][9] , \w3[8][8] , \w3[8][7] , \w3[8][6] ,
         \w3[8][5] , \w3[8][4] , \w3[8][3] , \w3[8][2] , \w3[8][1] ,
         \w3[8][0] , \w3[7][127] , \w3[7][126] , \w3[7][125] , \w3[7][124] ,
         \w3[7][123] , \w3[7][122] , \w3[7][121] , \w3[7][120] , \w3[7][119] ,
         \w3[7][118] , \w3[7][117] , \w3[7][116] , \w3[7][115] , \w3[7][114] ,
         \w3[7][113] , \w3[7][112] , \w3[7][111] , \w3[7][110] , \w3[7][109] ,
         \w3[7][108] , \w3[7][107] , \w3[7][106] , \w3[7][105] , \w3[7][104] ,
         \w3[7][103] , \w3[7][102] , \w3[7][101] , \w3[7][100] , \w3[7][99] ,
         \w3[7][98] , \w3[7][97] , \w3[7][96] , \w3[7][95] , \w3[7][94] ,
         \w3[7][93] , \w3[7][92] , \w3[7][91] , \w3[7][90] , \w3[7][89] ,
         \w3[7][88] , \w3[7][87] , \w3[7][86] , \w3[7][85] , \w3[7][84] ,
         \w3[7][83] , \w3[7][82] , \w3[7][81] , \w3[7][80] , \w3[7][79] ,
         \w3[7][78] , \w3[7][77] , \w3[7][76] , \w3[7][75] , \w3[7][74] ,
         \w3[7][73] , \w3[7][72] , \w3[7][71] , \w3[7][70] , \w3[7][69] ,
         \w3[7][68] , \w3[7][67] , \w3[7][66] , \w3[7][65] , \w3[7][64] ,
         \w3[7][63] , \w3[7][62] , \w3[7][61] , \w3[7][60] , \w3[7][59] ,
         \w3[7][58] , \w3[7][57] , \w3[7][56] , \w3[7][55] , \w3[7][54] ,
         \w3[7][53] , \w3[7][52] , \w3[7][51] , \w3[7][50] , \w3[7][49] ,
         \w3[7][48] , \w3[7][47] , \w3[7][46] , \w3[7][45] , \w3[7][44] ,
         \w3[7][43] , \w3[7][42] , \w3[7][41] , \w3[7][40] , \w3[7][39] ,
         \w3[7][38] , \w3[7][37] , \w3[7][36] , \w3[7][35] , \w3[7][34] ,
         \w3[7][33] , \w3[7][32] , \w3[7][31] , \w3[7][30] , \w3[7][29] ,
         \w3[7][28] , \w3[7][27] , \w3[7][26] , \w3[7][25] , \w3[7][24] ,
         \w3[7][23] , \w3[7][22] , \w3[7][21] , \w3[7][20] , \w3[7][19] ,
         \w3[7][18] , \w3[7][17] , \w3[7][16] , \w3[7][15] , \w3[7][14] ,
         \w3[7][13] , \w3[7][12] , \w3[7][11] , \w3[7][10] , \w3[7][9] ,
         \w3[7][8] , \w3[7][7] , \w3[7][6] , \w3[7][5] , \w3[7][4] ,
         \w3[7][3] , \w3[7][2] , \w3[7][1] , \w3[7][0] , \w3[6][127] ,
         \w3[6][126] , \w3[6][125] , \w3[6][124] , \w3[6][123] , \w3[6][122] ,
         \w3[6][121] , \w3[6][120] , \w3[6][119] , \w3[6][118] , \w3[6][117] ,
         \w3[6][116] , \w3[6][115] , \w3[6][114] , \w3[6][113] , \w3[6][112] ,
         \w3[6][111] , \w3[6][110] , \w3[6][109] , \w3[6][108] , \w3[6][107] ,
         \w3[6][106] , \w3[6][105] , \w3[6][104] , \w3[6][103] , \w3[6][102] ,
         \w3[6][101] , \w3[6][100] , \w3[6][99] , \w3[6][98] , \w3[6][97] ,
         \w3[6][96] , \w3[6][95] , \w3[6][94] , \w3[6][93] , \w3[6][92] ,
         \w3[6][91] , \w3[6][90] , \w3[6][89] , \w3[6][88] , \w3[6][87] ,
         \w3[6][86] , \w3[6][85] , \w3[6][84] , \w3[6][83] , \w3[6][82] ,
         \w3[6][81] , \w3[6][80] , \w3[6][79] , \w3[6][78] , \w3[6][77] ,
         \w3[6][76] , \w3[6][75] , \w3[6][74] , \w3[6][73] , \w3[6][72] ,
         \w3[6][71] , \w3[6][70] , \w3[6][69] , \w3[6][68] , \w3[6][67] ,
         \w3[6][66] , \w3[6][65] , \w3[6][64] , \w3[6][63] , \w3[6][62] ,
         \w3[6][61] , \w3[6][60] , \w3[6][59] , \w3[6][58] , \w3[6][57] ,
         \w3[6][56] , \w3[6][55] , \w3[6][54] , \w3[6][53] , \w3[6][52] ,
         \w3[6][51] , \w3[6][50] , \w3[6][49] , \w3[6][48] , \w3[6][47] ,
         \w3[6][46] , \w3[6][45] , \w3[6][44] , \w3[6][43] , \w3[6][42] ,
         \w3[6][41] , \w3[6][40] , \w3[6][39] , \w3[6][38] , \w3[6][37] ,
         \w3[6][36] , \w3[6][35] , \w3[6][34] , \w3[6][33] , \w3[6][32] ,
         \w3[6][31] , \w3[6][30] , \w3[6][29] , \w3[6][28] , \w3[6][27] ,
         \w3[6][26] , \w3[6][25] , \w3[6][24] , \w3[6][23] , \w3[6][22] ,
         \w3[6][21] , \w3[6][20] , \w3[6][19] , \w3[6][18] , \w3[6][17] ,
         \w3[6][16] , \w3[6][15] , \w3[6][14] , \w3[6][13] , \w3[6][12] ,
         \w3[6][11] , \w3[6][10] , \w3[6][9] , \w3[6][8] , \w3[6][7] ,
         \w3[6][6] , \w3[6][5] , \w3[6][4] , \w3[6][3] , \w3[6][2] ,
         \w3[6][1] , \w3[6][0] , \w3[5][127] , \w3[5][126] , \w3[5][125] ,
         \w3[5][124] , \w3[5][123] , \w3[5][122] , \w3[5][121] , \w3[5][120] ,
         \w3[5][119] , \w3[5][118] , \w3[5][117] , \w3[5][116] , \w3[5][115] ,
         \w3[5][114] , \w3[5][113] , \w3[5][112] , \w3[5][111] , \w3[5][110] ,
         \w3[5][109] , \w3[5][108] , \w3[5][107] , \w3[5][106] , \w3[5][105] ,
         \w3[5][104] , \w3[5][103] , \w3[5][102] , \w3[5][101] , \w3[5][100] ,
         \w3[5][99] , \w3[5][98] , \w3[5][97] , \w3[5][96] , \w3[5][95] ,
         \w3[5][94] , \w3[5][93] , \w3[5][92] , \w3[5][91] , \w3[5][90] ,
         \w3[5][89] , \w3[5][88] , \w3[5][87] , \w3[5][86] , \w3[5][85] ,
         \w3[5][84] , \w3[5][83] , \w3[5][82] , \w3[5][81] , \w3[5][80] ,
         \w3[5][79] , \w3[5][78] , \w3[5][77] , \w3[5][76] , \w3[5][75] ,
         \w3[5][74] , \w3[5][73] , \w3[5][72] , \w3[5][71] , \w3[5][70] ,
         \w3[5][69] , \w3[5][68] , \w3[5][67] , \w3[5][66] , \w3[5][65] ,
         \w3[5][64] , \w3[5][63] , \w3[5][62] , \w3[5][61] , \w3[5][60] ,
         \w3[5][59] , \w3[5][58] , \w3[5][57] , \w3[5][56] , \w3[5][55] ,
         \w3[5][54] , \w3[5][53] , \w3[5][52] , \w3[5][51] , \w3[5][50] ,
         \w3[5][49] , \w3[5][48] , \w3[5][47] , \w3[5][46] , \w3[5][45] ,
         \w3[5][44] , \w3[5][43] , \w3[5][42] , \w3[5][41] , \w3[5][40] ,
         \w3[5][39] , \w3[5][38] , \w3[5][37] , \w3[5][36] , \w3[5][35] ,
         \w3[5][34] , \w3[5][33] , \w3[5][32] , \w3[5][31] , \w3[5][30] ,
         \w3[5][29] , \w3[5][28] , \w3[5][27] , \w3[5][26] , \w3[5][25] ,
         \w3[5][24] , \w3[5][23] , \w3[5][22] , \w3[5][21] , \w3[5][20] ,
         \w3[5][19] , \w3[5][18] , \w3[5][17] , \w3[5][16] , \w3[5][15] ,
         \w3[5][14] , \w3[5][13] , \w3[5][12] , \w3[5][11] , \w3[5][10] ,
         \w3[5][9] , \w3[5][8] , \w3[5][7] , \w3[5][6] , \w3[5][5] ,
         \w3[5][4] , \w3[5][3] , \w3[5][2] , \w3[5][1] , \w3[5][0] ,
         \w3[4][127] , \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] ,
         \w3[4][122] , \w3[4][121] , \w3[4][120] , \w3[4][119] , \w3[4][118] ,
         \w3[4][117] , \w3[4][116] , \w3[4][115] , \w3[4][114] , \w3[4][113] ,
         \w3[4][112] , \w3[4][111] , \w3[4][110] , \w3[4][109] , \w3[4][108] ,
         \w3[4][107] , \w3[4][106] , \w3[4][105] , \w3[4][104] , \w3[4][103] ,
         \w3[4][102] , \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] ,
         \w3[4][97] , \w3[4][96] , \w3[4][95] , \w3[4][94] , \w3[4][93] ,
         \w3[4][92] , \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] ,
         \w3[4][87] , \w3[4][86] , \w3[4][85] , \w3[4][84] , \w3[4][83] ,
         \w3[4][82] , \w3[4][81] , \w3[4][80] , \w3[4][79] , \w3[4][78] ,
         \w3[4][77] , \w3[4][76] , \w3[4][75] , \w3[4][74] , \w3[4][73] ,
         \w3[4][72] , \w3[4][71] , \w3[4][70] , \w3[4][69] , \w3[4][68] ,
         \w3[4][67] , \w3[4][66] , \w3[4][65] , \w3[4][64] , \w3[4][63] ,
         \w3[4][62] , \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] ,
         \w3[4][57] , \w3[4][56] , \w3[4][55] , \w3[4][54] , \w3[4][53] ,
         \w3[4][52] , \w3[4][51] , \w3[4][50] , \w3[4][49] , \w3[4][48] ,
         \w3[4][47] , \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] ,
         \w3[4][42] , \w3[4][41] , \w3[4][40] , \w3[4][39] , \w3[4][38] ,
         \w3[4][37] , \w3[4][36] , \w3[4][35] , \w3[4][34] , \w3[4][33] ,
         \w3[4][32] , \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] ,
         \w3[4][27] , \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][23] ,
         \w3[4][22] , \w3[4][21] , \w3[4][20] , \w3[4][19] , \w3[4][18] ,
         \w3[4][17] , \w3[4][16] , \w3[4][15] , \w3[4][14] , \w3[4][13] ,
         \w3[4][12] , \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] ,
         \w3[4][7] , \w3[4][6] , \w3[4][5] , \w3[4][4] , \w3[4][3] ,
         \w3[4][2] , \w3[4][1] , \w3[4][0] , \w3[3][127] , \w3[3][126] ,
         \w3[3][125] , \w3[3][124] , \w3[3][123] , \w3[3][122] , \w3[3][121] ,
         \w3[3][120] , \w3[3][119] , \w3[3][118] , \w3[3][117] , \w3[3][116] ,
         \w3[3][115] , \w3[3][114] , \w3[3][113] , \w3[3][112] , \w3[3][111] ,
         \w3[3][110] , \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] ,
         \w3[3][105] , \w3[3][104] , \w3[3][103] , \w3[3][102] , \w3[3][101] ,
         \w3[3][100] , \w3[3][99] , \w3[3][98] , \w3[3][97] , \w3[3][96] ,
         \w3[3][95] , \w3[3][94] , \w3[3][93] , \w3[3][92] , \w3[3][91] ,
         \w3[3][90] , \w3[3][89] , \w3[3][88] , \w3[3][87] , \w3[3][86] ,
         \w3[3][85] , \w3[3][84] , \w3[3][83] , \w3[3][82] , \w3[3][81] ,
         \w3[3][80] , \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] ,
         \w3[3][75] , \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][71] ,
         \w3[3][70] , \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] ,
         \w3[3][65] , \w3[3][64] , \w3[3][63] , \w3[3][62] , \w3[3][61] ,
         \w3[3][60] , \w3[3][59] , \w3[3][58] , \w3[3][57] , \w3[3][56] ,
         \w3[3][55] , \w3[3][54] , \w3[3][53] , \w3[3][52] , \w3[3][51] ,
         \w3[3][50] , \w3[3][49] , \w3[3][48] , \w3[3][47] , \w3[3][46] ,
         \w3[3][45] , \w3[3][44] , \w3[3][43] , \w3[3][42] , \w3[3][41] ,
         \w3[3][40] , \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] ,
         \w3[3][35] , \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][31] ,
         \w3[3][30] , \w3[3][29] , \w3[3][28] , \w3[3][27] , \w3[3][26] ,
         \w3[3][25] , \w3[3][24] , \w3[3][23] , \w3[3][22] , \w3[3][21] ,
         \w3[3][20] , \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] ,
         \w3[3][15] , \w3[3][14] , \w3[3][13] , \w3[3][12] , \w3[3][11] ,
         \w3[3][10] , \w3[3][9] , \w3[3][8] , \w3[3][7] , \w3[3][6] ,
         \w3[3][5] , \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] ,
         \w3[3][0] , \w3[2][127] , \w3[2][126] , \w3[2][125] , \w3[2][124] ,
         \w3[2][123] , \w3[2][122] , \w3[2][121] , \w3[2][120] , \w3[2][119] ,
         \w3[2][118] , \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] ,
         \w3[2][113] , \w3[2][112] , \w3[2][111] , \w3[2][110] , \w3[2][109] ,
         \w3[2][108] , \w3[2][107] , \w3[2][106] , \w3[2][105] , \w3[2][104] ,
         \w3[2][103] , \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] ,
         \w3[2][98] , \w3[2][97] , \w3[2][96] , \w3[2][95] , \w3[2][94] ,
         \w3[2][93] , \w3[2][92] , \w3[2][91] , \w3[2][90] , \w3[2][89] ,
         \w3[2][88] , \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] ,
         \w3[2][83] , \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][79] ,
         \w3[2][78] , \w3[2][77] , \w3[2][76] , \w3[2][75] , \w3[2][74] ,
         \w3[2][73] , \w3[2][72] , \w3[2][71] , \w3[2][70] , \w3[2][69] ,
         \w3[2][68] , \w3[2][67] , \w3[2][66] , \w3[2][65] , \w3[2][64] ,
         \w3[2][63] , \w3[2][62] , \w3[2][61] , \w3[2][60] , \w3[2][59] ,
         \w3[2][58] , \w3[2][57] , \w3[2][56] , \w3[2][55] , \w3[2][54] ,
         \w3[2][53] , \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] ,
         \w3[2][48] , \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] ,
         \w3[2][43] , \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][39] ,
         \w3[2][38] , \w3[2][37] , \w3[2][36] , \w3[2][35] , \w3[2][34] ,
         \w3[2][33] , \w3[2][32] , \w3[2][31] , \w3[2][30] , \w3[2][29] ,
         \w3[2][28] , \w3[2][27] , \w3[2][26] , \w3[2][25] , \w3[2][24] ,
         \w3[2][23] , \w3[2][22] , \w3[2][21] , \w3[2][20] , \w3[2][19] ,
         \w3[2][18] , \w3[2][17] , \w3[2][16] , \w3[2][15] , \w3[2][14] ,
         \w3[2][13] , \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] ,
         \w3[2][8] , \w3[2][7] , \w3[2][6] , \w3[2][5] , \w3[2][4] ,
         \w3[2][3] , \w3[2][2] , \w3[2][1] , \w3[2][0] , \w3[1][127] ,
         \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] ,
         \w3[1][121] , \w3[1][120] , \w3[1][119] , \w3[1][118] , \w3[1][117] ,
         \w3[1][116] , \w3[1][115] , \w3[1][114] , \w3[1][113] , \w3[1][112] ,
         \w3[1][111] , \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] ,
         \w3[1][106] , \w3[1][105] , \w3[1][104] , \w3[1][103] , \w3[1][102] ,
         \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , \w3[1][97] ,
         \w3[1][96] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] ,
         \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][87] ,
         \w3[1][86] , \w3[1][85] , \w3[1][84] , \w3[1][83] , \w3[1][82] ,
         \w3[1][81] , \w3[1][80] , \w3[1][79] , \w3[1][78] , \w3[1][77] ,
         \w3[1][76] , \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] ,
         \w3[1][71] , \w3[1][70] , \w3[1][69] , \w3[1][68] , \w3[1][67] ,
         \w3[1][66] , \w3[1][65] , \w3[1][64] , \w3[1][63] , \w3[1][62] ,
         \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] ,
         \w3[1][56] , \w3[1][55] , \w3[1][54] , \w3[1][53] , \w3[1][52] ,
         \w3[1][51] , \w3[1][50] , \w3[1][49] , \w3[1][48] , \w3[1][47] ,
         \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , \w3[1][42] ,
         \w3[1][41] , \w3[1][40] , \w3[1][39] , \w3[1][38] , \w3[1][37] ,
         \w3[1][36] , \w3[1][35] , \w3[1][34] , \w3[1][33] , \w3[1][32] ,
         \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] ,
         \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][23] , \w3[1][22] ,
         \w3[1][21] , \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] ,
         \w3[1][16] , \w3[1][15] , \w3[1][14] , \w3[1][13] , \w3[1][12] ,
         \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , \w3[1][7] ,
         \w3[1][6] , \w3[1][5] , \w3[1][4] , \w3[1][3] , \w3[1][2] ,
         \w3[1][1] , \w3[1][0] , \w3[0][127] , \w3[0][126] , \w3[0][125] ,
         \w3[0][124] , \w3[0][123] , \w3[0][122] , \w3[0][121] , \w3[0][120] ,
         \w3[0][119] , \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] ,
         \w3[0][114] , \w3[0][113] , \w3[0][112] , \w3[0][111] , \w3[0][110] ,
         \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , \w3[0][105] ,
         \w3[0][104] , \w3[0][103] , \w3[0][102] , \w3[0][101] , \w3[0][100] ,
         \w3[0][99] , \w3[0][98] , \w3[0][97] , \w3[0][96] , \w3[0][95] ,
         \w3[0][94] , \w3[0][93] , \w3[0][92] , \w3[0][91] , \w3[0][90] ,
         \w3[0][89] , \w3[0][88] , \w3[0][87] , \w3[0][86] , \w3[0][85] ,
         \w3[0][84] , \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] ,
         \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , \w3[0][75] ,
         \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][71] , \w3[0][70] ,
         \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] ,
         \w3[0][64] , \w3[0][63] , \w3[0][62] , \w3[0][61] , \w3[0][60] ,
         \w3[0][59] , \w3[0][58] , \w3[0][57] , \w3[0][56] , \w3[0][55] ,
         \w3[0][54] , \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] ,
         \w3[0][49] , \w3[0][48] , \w3[0][47] , \w3[0][46] , \w3[0][45] ,
         \w3[0][44] , \w3[0][43] , \w3[0][42] , \w3[0][41] , \w3[0][40] ,
         \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] ,
         \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][31] , \w3[0][30] ,
         \w3[0][29] , \w3[0][28] , \w3[0][27] , \w3[0][26] , \w3[0][25] ,
         \w3[0][24] , \w3[0][23] , \w3[0][22] , \w3[0][21] , \w3[0][20] ,
         \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , \w3[0][15] ,
         \w3[0][14] , \w3[0][13] , \w3[0][12] , \w3[0][11] , \w3[0][10] ,
         \w3[0][9] , \w3[0][8] , \w3[0][7] , \w3[0][6] , \w3[0][5] ,
         \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202;

  SubBytes_7 \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  SubBytes_16 \SUBBYTES[1].a  ( .x({\w1[1][127] , \w1[1][126] , \w1[1][125] , 
        \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] , \w1[1][120] , 
        \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] , \w1[1][115] , 
        \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] , \w1[1][110] , 
        \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] , \w1[1][105] , 
        \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] , \w1[1][100] , 
        \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] , \w1[1][95] , 
        \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] , \w1[1][90] , 
        \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] , \w1[1][85] , 
        \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] , \w1[1][80] , 
        \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] , \w1[1][75] , 
        \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] , \w1[1][70] , 
        \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] , \w1[1][65] , 
        \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] , \w1[1][60] , 
        \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] , \w1[1][55] , 
        \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] , \w1[1][50] , 
        \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] , \w1[1][45] , 
        \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] , \w1[1][40] , 
        \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] , \w1[1][35] , 
        \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] , \w1[1][30] , 
        \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] , \w1[1][25] , 
        \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] , \w1[1][20] , 
        \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] , \w1[1][15] , 
        \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] , \w1[1][10] , 
        \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] , \w1[1][5] , \w1[1][4] , 
        \w1[1][3] , \w1[1][2] , \w1[1][1] , \w1[1][0] }), .z({\w3[1][127] , 
        \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , 
        \w3[1][121] , \w3[1][120] , \w3[1][23] , \w3[1][22] , \w3[1][21] , 
        \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] , 
        \w3[1][47] , \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , 
        \w3[1][42] , \w3[1][41] , \w3[1][40] , \w3[1][71] , \w3[1][70] , 
        \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] , \w3[1][65] , 
        \w3[1][64] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , 
        \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][119] , 
        \w3[1][118] , \w3[1][117] , \w3[1][116] , \w3[1][115] , \w3[1][114] , 
        \w3[1][113] , \w3[1][112] , \w3[1][15] , \w3[1][14] , \w3[1][13] , 
        \w3[1][12] , \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , 
        \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] , \w3[1][35] , 
        \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][63] , \w3[1][62] , 
        \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , 
        \w3[1][56] , \w3[1][87] , \w3[1][86] , \w3[1][85] , \w3[1][84] , 
        \w3[1][83] , \w3[1][82] , \w3[1][81] , \w3[1][80] , \w3[1][111] , 
        \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] , 
        \w3[1][105] , \w3[1][104] , \w3[1][7] , \w3[1][6] , \w3[1][5] , 
        \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] , \w3[1][0] , 
        \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , 
        \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][55] , \w3[1][54] , 
        \w3[1][53] , \w3[1][52] , \w3[1][51] , \w3[1][50] , \w3[1][49] , 
        \w3[1][48] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] , 
        \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][103] , 
        \w3[1][102] , \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , 
        \w3[1][97] , \w3[1][96] }) );
  SubBytes_15 \SUBBYTES[2].a  ( .x({\w1[2][127] , \w1[2][126] , \w1[2][125] , 
        \w1[2][124] , \w1[2][123] , \w1[2][122] , \w1[2][121] , \w1[2][120] , 
        \w1[2][119] , \w1[2][118] , \w1[2][117] , \w1[2][116] , \w1[2][115] , 
        \w1[2][114] , \w1[2][113] , \w1[2][112] , \w1[2][111] , \w1[2][110] , 
        \w1[2][109] , \w1[2][108] , \w1[2][107] , \w1[2][106] , \w1[2][105] , 
        \w1[2][104] , \w1[2][103] , \w1[2][102] , \w1[2][101] , \w1[2][100] , 
        \w1[2][99] , \w1[2][98] , \w1[2][97] , \w1[2][96] , \w1[2][95] , 
        \w1[2][94] , \w1[2][93] , \w1[2][92] , \w1[2][91] , \w1[2][90] , 
        \w1[2][89] , \w1[2][88] , \w1[2][87] , \w1[2][86] , \w1[2][85] , 
        \w1[2][84] , \w1[2][83] , \w1[2][82] , \w1[2][81] , \w1[2][80] , 
        \w1[2][79] , \w1[2][78] , \w1[2][77] , \w1[2][76] , \w1[2][75] , 
        \w1[2][74] , \w1[2][73] , \w1[2][72] , \w1[2][71] , \w1[2][70] , 
        \w1[2][69] , \w1[2][68] , \w1[2][67] , \w1[2][66] , \w1[2][65] , 
        \w1[2][64] , \w1[2][63] , \w1[2][62] , \w1[2][61] , \w1[2][60] , 
        \w1[2][59] , \w1[2][58] , \w1[2][57] , \w1[2][56] , \w1[2][55] , 
        \w1[2][54] , \w1[2][53] , \w1[2][52] , \w1[2][51] , \w1[2][50] , 
        \w1[2][49] , \w1[2][48] , \w1[2][47] , \w1[2][46] , \w1[2][45] , 
        \w1[2][44] , \w1[2][43] , \w1[2][42] , \w1[2][41] , \w1[2][40] , 
        \w1[2][39] , \w1[2][38] , \w1[2][37] , \w1[2][36] , \w1[2][35] , 
        \w1[2][34] , \w1[2][33] , \w1[2][32] , \w1[2][31] , \w1[2][30] , 
        \w1[2][29] , \w1[2][28] , \w1[2][27] , \w1[2][26] , \w1[2][25] , 
        \w1[2][24] , \w1[2][23] , \w1[2][22] , \w1[2][21] , \w1[2][20] , 
        \w1[2][19] , \w1[2][18] , \w1[2][17] , \w1[2][16] , \w1[2][15] , 
        \w1[2][14] , \w1[2][13] , \w1[2][12] , \w1[2][11] , \w1[2][10] , 
        \w1[2][9] , \w1[2][8] , \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] , 
        \w1[2][3] , \w1[2][2] , \w1[2][1] , \w1[2][0] }), .z({\w3[2][127] , 
        \w3[2][126] , \w3[2][125] , \w3[2][124] , \w3[2][123] , \w3[2][122] , 
        \w3[2][121] , \w3[2][120] , \w3[2][23] , \w3[2][22] , \w3[2][21] , 
        \w3[2][20] , \w3[2][19] , \w3[2][18] , \w3[2][17] , \w3[2][16] , 
        \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] , \w3[2][43] , 
        \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][71] , \w3[2][70] , 
        \w3[2][69] , \w3[2][68] , \w3[2][67] , \w3[2][66] , \w3[2][65] , 
        \w3[2][64] , \w3[2][95] , \w3[2][94] , \w3[2][93] , \w3[2][92] , 
        \w3[2][91] , \w3[2][90] , \w3[2][89] , \w3[2][88] , \w3[2][119] , 
        \w3[2][118] , \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] , 
        \w3[2][113] , \w3[2][112] , \w3[2][15] , \w3[2][14] , \w3[2][13] , 
        \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] , \w3[2][8] , 
        \w3[2][39] , \w3[2][38] , \w3[2][37] , \w3[2][36] , \w3[2][35] , 
        \w3[2][34] , \w3[2][33] , \w3[2][32] , \w3[2][63] , \w3[2][62] , 
        \w3[2][61] , \w3[2][60] , \w3[2][59] , \w3[2][58] , \w3[2][57] , 
        \w3[2][56] , \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] , 
        \w3[2][83] , \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][111] , 
        \w3[2][110] , \w3[2][109] , \w3[2][108] , \w3[2][107] , \w3[2][106] , 
        \w3[2][105] , \w3[2][104] , \w3[2][7] , \w3[2][6] , \w3[2][5] , 
        \w3[2][4] , \w3[2][3] , \w3[2][2] , \w3[2][1] , \w3[2][0] , 
        \w3[2][31] , \w3[2][30] , \w3[2][29] , \w3[2][28] , \w3[2][27] , 
        \w3[2][26] , \w3[2][25] , \w3[2][24] , \w3[2][55] , \w3[2][54] , 
        \w3[2][53] , \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] , 
        \w3[2][48] , \w3[2][79] , \w3[2][78] , \w3[2][77] , \w3[2][76] , 
        \w3[2][75] , \w3[2][74] , \w3[2][73] , \w3[2][72] , \w3[2][103] , 
        \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] , \w3[2][98] , 
        \w3[2][97] , \w3[2][96] }) );
  SubBytes_14 \SUBBYTES[3].a  ( .x({\w1[3][127] , \w1[3][126] , \w1[3][125] , 
        \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] , \w1[3][120] , 
        \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] , \w1[3][115] , 
        \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] , \w1[3][110] , 
        \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] , \w1[3][105] , 
        \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] , \w1[3][100] , 
        \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] , \w1[3][95] , 
        \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] , \w1[3][90] , 
        \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] , \w1[3][85] , 
        \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] , \w1[3][80] , 
        \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] , \w1[3][75] , 
        \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] , \w1[3][70] , 
        \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] , \w1[3][65] , 
        \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] , \w1[3][60] , 
        \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] , \w1[3][55] , 
        \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] , \w1[3][50] , 
        \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] , \w1[3][45] , 
        \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] , \w1[3][40] , 
        \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] , \w1[3][35] , 
        \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] , \w1[3][30] , 
        \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] , \w1[3][25] , 
        \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] , \w1[3][20] , 
        \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] , \w1[3][15] , 
        \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] , \w1[3][10] , 
        \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] , \w1[3][5] , \w1[3][4] , 
        \w1[3][3] , \w1[3][2] , \w1[3][1] , \w1[3][0] }), .z({\w3[3][127] , 
        \w3[3][126] , \w3[3][125] , \w3[3][124] , \w3[3][123] , \w3[3][122] , 
        \w3[3][121] , \w3[3][120] , \w3[3][23] , \w3[3][22] , \w3[3][21] , 
        \w3[3][20] , \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] , 
        \w3[3][47] , \w3[3][46] , \w3[3][45] , \w3[3][44] , \w3[3][43] , 
        \w3[3][42] , \w3[3][41] , \w3[3][40] , \w3[3][71] , \w3[3][70] , 
        \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] , \w3[3][65] , 
        \w3[3][64] , \w3[3][95] , \w3[3][94] , \w3[3][93] , \w3[3][92] , 
        \w3[3][91] , \w3[3][90] , \w3[3][89] , \w3[3][88] , \w3[3][119] , 
        \w3[3][118] , \w3[3][117] , \w3[3][116] , \w3[3][115] , \w3[3][114] , 
        \w3[3][113] , \w3[3][112] , \w3[3][15] , \w3[3][14] , \w3[3][13] , 
        \w3[3][12] , \w3[3][11] , \w3[3][10] , \w3[3][9] , \w3[3][8] , 
        \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] , \w3[3][35] , 
        \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][63] , \w3[3][62] , 
        \w3[3][61] , \w3[3][60] , \w3[3][59] , \w3[3][58] , \w3[3][57] , 
        \w3[3][56] , \w3[3][87] , \w3[3][86] , \w3[3][85] , \w3[3][84] , 
        \w3[3][83] , \w3[3][82] , \w3[3][81] , \w3[3][80] , \w3[3][111] , 
        \w3[3][110] , \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] , 
        \w3[3][105] , \w3[3][104] , \w3[3][7] , \w3[3][6] , \w3[3][5] , 
        \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] , \w3[3][0] , 
        \w3[3][31] , \w3[3][30] , \w3[3][29] , \w3[3][28] , \w3[3][27] , 
        \w3[3][26] , \w3[3][25] , \w3[3][24] , \w3[3][55] , \w3[3][54] , 
        \w3[3][53] , \w3[3][52] , \w3[3][51] , \w3[3][50] , \w3[3][49] , 
        \w3[3][48] , \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] , 
        \w3[3][75] , \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][103] , 
        \w3[3][102] , \w3[3][101] , \w3[3][100] , \w3[3][99] , \w3[3][98] , 
        \w3[3][97] , \w3[3][96] }) );
  SubBytes_13 \SUBBYTES[4].a  ( .x({\w1[4][127] , \w1[4][126] , \w1[4][125] , 
        \w1[4][124] , \w1[4][123] , \w1[4][122] , \w1[4][121] , \w1[4][120] , 
        \w1[4][119] , \w1[4][118] , \w1[4][117] , \w1[4][116] , \w1[4][115] , 
        \w1[4][114] , \w1[4][113] , \w1[4][112] , \w1[4][111] , \w1[4][110] , 
        \w1[4][109] , \w1[4][108] , \w1[4][107] , \w1[4][106] , \w1[4][105] , 
        \w1[4][104] , \w1[4][103] , \w1[4][102] , \w1[4][101] , \w1[4][100] , 
        \w1[4][99] , \w1[4][98] , \w1[4][97] , \w1[4][96] , \w1[4][95] , 
        \w1[4][94] , \w1[4][93] , \w1[4][92] , \w1[4][91] , \w1[4][90] , 
        \w1[4][89] , \w1[4][88] , \w1[4][87] , \w1[4][86] , \w1[4][85] , 
        \w1[4][84] , \w1[4][83] , \w1[4][82] , \w1[4][81] , \w1[4][80] , 
        \w1[4][79] , \w1[4][78] , \w1[4][77] , \w1[4][76] , \w1[4][75] , 
        \w1[4][74] , \w1[4][73] , \w1[4][72] , \w1[4][71] , \w1[4][70] , 
        \w1[4][69] , \w1[4][68] , \w1[4][67] , \w1[4][66] , \w1[4][65] , 
        \w1[4][64] , \w1[4][63] , \w1[4][62] , \w1[4][61] , \w1[4][60] , 
        \w1[4][59] , \w1[4][58] , \w1[4][57] , \w1[4][56] , \w1[4][55] , 
        \w1[4][54] , \w1[4][53] , \w1[4][52] , \w1[4][51] , \w1[4][50] , 
        \w1[4][49] , \w1[4][48] , \w1[4][47] , \w1[4][46] , \w1[4][45] , 
        \w1[4][44] , \w1[4][43] , \w1[4][42] , \w1[4][41] , \w1[4][40] , 
        \w1[4][39] , \w1[4][38] , \w1[4][37] , \w1[4][36] , \w1[4][35] , 
        \w1[4][34] , \w1[4][33] , \w1[4][32] , \w1[4][31] , \w1[4][30] , 
        \w1[4][29] , \w1[4][28] , \w1[4][27] , \w1[4][26] , \w1[4][25] , 
        \w1[4][24] , \w1[4][23] , \w1[4][22] , \w1[4][21] , \w1[4][20] , 
        \w1[4][19] , \w1[4][18] , \w1[4][17] , \w1[4][16] , \w1[4][15] , 
        \w1[4][14] , \w1[4][13] , \w1[4][12] , \w1[4][11] , \w1[4][10] , 
        \w1[4][9] , \w1[4][8] , \w1[4][7] , \w1[4][6] , \w1[4][5] , \w1[4][4] , 
        \w1[4][3] , \w1[4][2] , \w1[4][1] , \w1[4][0] }), .z({\w3[4][127] , 
        \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] , \w3[4][122] , 
        \w3[4][121] , \w3[4][120] , \w3[4][23] , \w3[4][22] , \w3[4][21] , 
        \w3[4][20] , \w3[4][19] , \w3[4][18] , \w3[4][17] , \w3[4][16] , 
        \w3[4][47] , \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] , 
        \w3[4][42] , \w3[4][41] , \w3[4][40] , \w3[4][71] , \w3[4][70] , 
        \w3[4][69] , \w3[4][68] , \w3[4][67] , \w3[4][66] , \w3[4][65] , 
        \w3[4][64] , \w3[4][95] , \w3[4][94] , \w3[4][93] , \w3[4][92] , 
        \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] , \w3[4][119] , 
        \w3[4][118] , \w3[4][117] , \w3[4][116] , \w3[4][115] , \w3[4][114] , 
        \w3[4][113] , \w3[4][112] , \w3[4][15] , \w3[4][14] , \w3[4][13] , 
        \w3[4][12] , \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] , 
        \w3[4][39] , \w3[4][38] , \w3[4][37] , \w3[4][36] , \w3[4][35] , 
        \w3[4][34] , \w3[4][33] , \w3[4][32] , \w3[4][63] , \w3[4][62] , 
        \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] , \w3[4][57] , 
        \w3[4][56] , \w3[4][87] , \w3[4][86] , \w3[4][85] , \w3[4][84] , 
        \w3[4][83] , \w3[4][82] , \w3[4][81] , \w3[4][80] , \w3[4][111] , 
        \w3[4][110] , \w3[4][109] , \w3[4][108] , \w3[4][107] , \w3[4][106] , 
        \w3[4][105] , \w3[4][104] , \w3[4][7] , \w3[4][6] , \w3[4][5] , 
        \w3[4][4] , \w3[4][3] , \w3[4][2] , \w3[4][1] , \w3[4][0] , 
        \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] , \w3[4][27] , 
        \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][55] , \w3[4][54] , 
        \w3[4][53] , \w3[4][52] , \w3[4][51] , \w3[4][50] , \w3[4][49] , 
        \w3[4][48] , \w3[4][79] , \w3[4][78] , \w3[4][77] , \w3[4][76] , 
        \w3[4][75] , \w3[4][74] , \w3[4][73] , \w3[4][72] , \w3[4][103] , 
        \w3[4][102] , \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] , 
        \w3[4][97] , \w3[4][96] }) );
  SubBytes_12 \SUBBYTES[5].a  ( .x({\w1[5][127] , \w1[5][126] , \w1[5][125] , 
        \w1[5][124] , \w1[5][123] , \w1[5][122] , \w1[5][121] , \w1[5][120] , 
        \w1[5][119] , \w1[5][118] , \w1[5][117] , \w1[5][116] , \w1[5][115] , 
        \w1[5][114] , \w1[5][113] , \w1[5][112] , \w1[5][111] , \w1[5][110] , 
        \w1[5][109] , \w1[5][108] , \w1[5][107] , \w1[5][106] , \w1[5][105] , 
        \w1[5][104] , \w1[5][103] , \w1[5][102] , \w1[5][101] , \w1[5][100] , 
        \w1[5][99] , \w1[5][98] , \w1[5][97] , \w1[5][96] , \w1[5][95] , 
        \w1[5][94] , \w1[5][93] , \w1[5][92] , \w1[5][91] , \w1[5][90] , 
        \w1[5][89] , \w1[5][88] , \w1[5][87] , \w1[5][86] , \w1[5][85] , 
        \w1[5][84] , \w1[5][83] , \w1[5][82] , \w1[5][81] , \w1[5][80] , 
        \w1[5][79] , \w1[5][78] , \w1[5][77] , \w1[5][76] , \w1[5][75] , 
        \w1[5][74] , \w1[5][73] , \w1[5][72] , \w1[5][71] , \w1[5][70] , 
        \w1[5][69] , \w1[5][68] , \w1[5][67] , \w1[5][66] , \w1[5][65] , 
        \w1[5][64] , \w1[5][63] , \w1[5][62] , \w1[5][61] , \w1[5][60] , 
        \w1[5][59] , \w1[5][58] , \w1[5][57] , \w1[5][56] , \w1[5][55] , 
        \w1[5][54] , \w1[5][53] , \w1[5][52] , \w1[5][51] , \w1[5][50] , 
        \w1[5][49] , \w1[5][48] , \w1[5][47] , \w1[5][46] , \w1[5][45] , 
        \w1[5][44] , \w1[5][43] , \w1[5][42] , \w1[5][41] , \w1[5][40] , 
        \w1[5][39] , \w1[5][38] , \w1[5][37] , \w1[5][36] , \w1[5][35] , 
        \w1[5][34] , \w1[5][33] , \w1[5][32] , \w1[5][31] , \w1[5][30] , 
        \w1[5][29] , \w1[5][28] , \w1[5][27] , \w1[5][26] , \w1[5][25] , 
        \w1[5][24] , \w1[5][23] , \w1[5][22] , \w1[5][21] , \w1[5][20] , 
        \w1[5][19] , \w1[5][18] , \w1[5][17] , \w1[5][16] , \w1[5][15] , 
        \w1[5][14] , \w1[5][13] , \w1[5][12] , \w1[5][11] , \w1[5][10] , 
        \w1[5][9] , \w1[5][8] , \w1[5][7] , \w1[5][6] , \w1[5][5] , \w1[5][4] , 
        \w1[5][3] , \w1[5][2] , \w1[5][1] , \w1[5][0] }), .z({\w3[5][127] , 
        \w3[5][126] , \w3[5][125] , \w3[5][124] , \w3[5][123] , \w3[5][122] , 
        \w3[5][121] , \w3[5][120] , \w3[5][23] , \w3[5][22] , \w3[5][21] , 
        \w3[5][20] , \w3[5][19] , \w3[5][18] , \w3[5][17] , \w3[5][16] , 
        \w3[5][47] , \w3[5][46] , \w3[5][45] , \w3[5][44] , \w3[5][43] , 
        \w3[5][42] , \w3[5][41] , \w3[5][40] , \w3[5][71] , \w3[5][70] , 
        \w3[5][69] , \w3[5][68] , \w3[5][67] , \w3[5][66] , \w3[5][65] , 
        \w3[5][64] , \w3[5][95] , \w3[5][94] , \w3[5][93] , \w3[5][92] , 
        \w3[5][91] , \w3[5][90] , \w3[5][89] , \w3[5][88] , \w3[5][119] , 
        \w3[5][118] , \w3[5][117] , \w3[5][116] , \w3[5][115] , \w3[5][114] , 
        \w3[5][113] , \w3[5][112] , \w3[5][15] , \w3[5][14] , \w3[5][13] , 
        \w3[5][12] , \w3[5][11] , \w3[5][10] , \w3[5][9] , \w3[5][8] , 
        \w3[5][39] , \w3[5][38] , \w3[5][37] , \w3[5][36] , \w3[5][35] , 
        \w3[5][34] , \w3[5][33] , \w3[5][32] , \w3[5][63] , \w3[5][62] , 
        \w3[5][61] , \w3[5][60] , \w3[5][59] , \w3[5][58] , \w3[5][57] , 
        \w3[5][56] , \w3[5][87] , \w3[5][86] , \w3[5][85] , \w3[5][84] , 
        \w3[5][83] , \w3[5][82] , \w3[5][81] , \w3[5][80] , \w3[5][111] , 
        \w3[5][110] , \w3[5][109] , \w3[5][108] , \w3[5][107] , \w3[5][106] , 
        \w3[5][105] , \w3[5][104] , \w3[5][7] , \w3[5][6] , \w3[5][5] , 
        \w3[5][4] , \w3[5][3] , \w3[5][2] , \w3[5][1] , \w3[5][0] , 
        \w3[5][31] , \w3[5][30] , \w3[5][29] , \w3[5][28] , \w3[5][27] , 
        \w3[5][26] , \w3[5][25] , \w3[5][24] , \w3[5][55] , \w3[5][54] , 
        \w3[5][53] , \w3[5][52] , \w3[5][51] , \w3[5][50] , \w3[5][49] , 
        \w3[5][48] , \w3[5][79] , \w3[5][78] , \w3[5][77] , \w3[5][76] , 
        \w3[5][75] , \w3[5][74] , \w3[5][73] , \w3[5][72] , \w3[5][103] , 
        \w3[5][102] , \w3[5][101] , \w3[5][100] , \w3[5][99] , \w3[5][98] , 
        \w3[5][97] , \w3[5][96] }) );
  SubBytes_11 \SUBBYTES[6].a  ( .x({\w1[6][127] , \w1[6][126] , \w1[6][125] , 
        \w1[6][124] , \w1[6][123] , \w1[6][122] , \w1[6][121] , \w1[6][120] , 
        \w1[6][119] , \w1[6][118] , \w1[6][117] , \w1[6][116] , \w1[6][115] , 
        \w1[6][114] , \w1[6][113] , \w1[6][112] , \w1[6][111] , \w1[6][110] , 
        \w1[6][109] , \w1[6][108] , \w1[6][107] , \w1[6][106] , \w1[6][105] , 
        \w1[6][104] , \w1[6][103] , \w1[6][102] , \w1[6][101] , \w1[6][100] , 
        \w1[6][99] , \w1[6][98] , \w1[6][97] , \w1[6][96] , \w1[6][95] , 
        \w1[6][94] , \w1[6][93] , \w1[6][92] , \w1[6][91] , \w1[6][90] , 
        \w1[6][89] , \w1[6][88] , \w1[6][87] , \w1[6][86] , \w1[6][85] , 
        \w1[6][84] , \w1[6][83] , \w1[6][82] , \w1[6][81] , \w1[6][80] , 
        \w1[6][79] , \w1[6][78] , \w1[6][77] , \w1[6][76] , \w1[6][75] , 
        \w1[6][74] , \w1[6][73] , \w1[6][72] , \w1[6][71] , \w1[6][70] , 
        \w1[6][69] , \w1[6][68] , \w1[6][67] , \w1[6][66] , \w1[6][65] , 
        \w1[6][64] , \w1[6][63] , \w1[6][62] , \w1[6][61] , \w1[6][60] , 
        \w1[6][59] , \w1[6][58] , \w1[6][57] , \w1[6][56] , \w1[6][55] , 
        \w1[6][54] , \w1[6][53] , \w1[6][52] , \w1[6][51] , \w1[6][50] , 
        \w1[6][49] , \w1[6][48] , \w1[6][47] , \w1[6][46] , \w1[6][45] , 
        \w1[6][44] , \w1[6][43] , \w1[6][42] , \w1[6][41] , \w1[6][40] , 
        \w1[6][39] , \w1[6][38] , \w1[6][37] , \w1[6][36] , \w1[6][35] , 
        \w1[6][34] , \w1[6][33] , \w1[6][32] , \w1[6][31] , \w1[6][30] , 
        \w1[6][29] , \w1[6][28] , \w1[6][27] , \w1[6][26] , \w1[6][25] , 
        \w1[6][24] , \w1[6][23] , \w1[6][22] , \w1[6][21] , \w1[6][20] , 
        \w1[6][19] , \w1[6][18] , \w1[6][17] , \w1[6][16] , \w1[6][15] , 
        \w1[6][14] , \w1[6][13] , \w1[6][12] , \w1[6][11] , \w1[6][10] , 
        \w1[6][9] , \w1[6][8] , \w1[6][7] , \w1[6][6] , \w1[6][5] , \w1[6][4] , 
        \w1[6][3] , \w1[6][2] , \w1[6][1] , \w1[6][0] }), .z({\w3[6][127] , 
        \w3[6][126] , \w3[6][125] , \w3[6][124] , \w3[6][123] , \w3[6][122] , 
        \w3[6][121] , \w3[6][120] , \w3[6][23] , \w3[6][22] , \w3[6][21] , 
        \w3[6][20] , \w3[6][19] , \w3[6][18] , \w3[6][17] , \w3[6][16] , 
        \w3[6][47] , \w3[6][46] , \w3[6][45] , \w3[6][44] , \w3[6][43] , 
        \w3[6][42] , \w3[6][41] , \w3[6][40] , \w3[6][71] , \w3[6][70] , 
        \w3[6][69] , \w3[6][68] , \w3[6][67] , \w3[6][66] , \w3[6][65] , 
        \w3[6][64] , \w3[6][95] , \w3[6][94] , \w3[6][93] , \w3[6][92] , 
        \w3[6][91] , \w3[6][90] , \w3[6][89] , \w3[6][88] , \w3[6][119] , 
        \w3[6][118] , \w3[6][117] , \w3[6][116] , \w3[6][115] , \w3[6][114] , 
        \w3[6][113] , \w3[6][112] , \w3[6][15] , \w3[6][14] , \w3[6][13] , 
        \w3[6][12] , \w3[6][11] , \w3[6][10] , \w3[6][9] , \w3[6][8] , 
        \w3[6][39] , \w3[6][38] , \w3[6][37] , \w3[6][36] , \w3[6][35] , 
        \w3[6][34] , \w3[6][33] , \w3[6][32] , \w3[6][63] , \w3[6][62] , 
        \w3[6][61] , \w3[6][60] , \w3[6][59] , \w3[6][58] , \w3[6][57] , 
        \w3[6][56] , \w3[6][87] , \w3[6][86] , \w3[6][85] , \w3[6][84] , 
        \w3[6][83] , \w3[6][82] , \w3[6][81] , \w3[6][80] , \w3[6][111] , 
        \w3[6][110] , \w3[6][109] , \w3[6][108] , \w3[6][107] , \w3[6][106] , 
        \w3[6][105] , \w3[6][104] , \w3[6][7] , \w3[6][6] , \w3[6][5] , 
        \w3[6][4] , \w3[6][3] , \w3[6][2] , \w3[6][1] , \w3[6][0] , 
        \w3[6][31] , \w3[6][30] , \w3[6][29] , \w3[6][28] , \w3[6][27] , 
        \w3[6][26] , \w3[6][25] , \w3[6][24] , \w3[6][55] , \w3[6][54] , 
        \w3[6][53] , \w3[6][52] , \w3[6][51] , \w3[6][50] , \w3[6][49] , 
        \w3[6][48] , \w3[6][79] , \w3[6][78] , \w3[6][77] , \w3[6][76] , 
        \w3[6][75] , \w3[6][74] , \w3[6][73] , \w3[6][72] , \w3[6][103] , 
        \w3[6][102] , \w3[6][101] , \w3[6][100] , \w3[6][99] , \w3[6][98] , 
        \w3[6][97] , \w3[6][96] }) );
  SubBytes_10 \SUBBYTES[7].a  ( .x({\w1[7][127] , \w1[7][126] , \w1[7][125] , 
        \w1[7][124] , \w1[7][123] , \w1[7][122] , \w1[7][121] , \w1[7][120] , 
        \w1[7][119] , \w1[7][118] , \w1[7][117] , \w1[7][116] , \w1[7][115] , 
        \w1[7][114] , \w1[7][113] , \w1[7][112] , \w1[7][111] , \w1[7][110] , 
        \w1[7][109] , \w1[7][108] , \w1[7][107] , \w1[7][106] , \w1[7][105] , 
        \w1[7][104] , \w1[7][103] , \w1[7][102] , \w1[7][101] , \w1[7][100] , 
        \w1[7][99] , \w1[7][98] , \w1[7][97] , \w1[7][96] , \w1[7][95] , 
        \w1[7][94] , \w1[7][93] , \w1[7][92] , \w1[7][91] , \w1[7][90] , 
        \w1[7][89] , \w1[7][88] , \w1[7][87] , \w1[7][86] , \w1[7][85] , 
        \w1[7][84] , \w1[7][83] , \w1[7][82] , \w1[7][81] , \w1[7][80] , 
        \w1[7][79] , \w1[7][78] , \w1[7][77] , \w1[7][76] , \w1[7][75] , 
        \w1[7][74] , \w1[7][73] , \w1[7][72] , \w1[7][71] , \w1[7][70] , 
        \w1[7][69] , \w1[7][68] , \w1[7][67] , \w1[7][66] , \w1[7][65] , 
        \w1[7][64] , \w1[7][63] , \w1[7][62] , \w1[7][61] , \w1[7][60] , 
        \w1[7][59] , \w1[7][58] , \w1[7][57] , \w1[7][56] , \w1[7][55] , 
        \w1[7][54] , \w1[7][53] , \w1[7][52] , \w1[7][51] , \w1[7][50] , 
        \w1[7][49] , \w1[7][48] , \w1[7][47] , \w1[7][46] , \w1[7][45] , 
        \w1[7][44] , \w1[7][43] , \w1[7][42] , \w1[7][41] , \w1[7][40] , 
        \w1[7][39] , \w1[7][38] , \w1[7][37] , \w1[7][36] , \w1[7][35] , 
        \w1[7][34] , \w1[7][33] , \w1[7][32] , \w1[7][31] , \w1[7][30] , 
        \w1[7][29] , \w1[7][28] , \w1[7][27] , \w1[7][26] , \w1[7][25] , 
        \w1[7][24] , \w1[7][23] , \w1[7][22] , \w1[7][21] , \w1[7][20] , 
        \w1[7][19] , \w1[7][18] , \w1[7][17] , \w1[7][16] , \w1[7][15] , 
        \w1[7][14] , \w1[7][13] , \w1[7][12] , \w1[7][11] , \w1[7][10] , 
        \w1[7][9] , \w1[7][8] , \w1[7][7] , \w1[7][6] , \w1[7][5] , \w1[7][4] , 
        \w1[7][3] , \w1[7][2] , \w1[7][1] , \w1[7][0] }), .z({\w3[7][127] , 
        \w3[7][126] , \w3[7][125] , \w3[7][124] , \w3[7][123] , \w3[7][122] , 
        \w3[7][121] , \w3[7][120] , \w3[7][23] , \w3[7][22] , \w3[7][21] , 
        \w3[7][20] , \w3[7][19] , \w3[7][18] , \w3[7][17] , \w3[7][16] , 
        \w3[7][47] , \w3[7][46] , \w3[7][45] , \w3[7][44] , \w3[7][43] , 
        \w3[7][42] , \w3[7][41] , \w3[7][40] , \w3[7][71] , \w3[7][70] , 
        \w3[7][69] , \w3[7][68] , \w3[7][67] , \w3[7][66] , \w3[7][65] , 
        \w3[7][64] , \w3[7][95] , \w3[7][94] , \w3[7][93] , \w3[7][92] , 
        \w3[7][91] , \w3[7][90] , \w3[7][89] , \w3[7][88] , \w3[7][119] , 
        \w3[7][118] , \w3[7][117] , \w3[7][116] , \w3[7][115] , \w3[7][114] , 
        \w3[7][113] , \w3[7][112] , \w3[7][15] , \w3[7][14] , \w3[7][13] , 
        \w3[7][12] , \w3[7][11] , \w3[7][10] , \w3[7][9] , \w3[7][8] , 
        \w3[7][39] , \w3[7][38] , \w3[7][37] , \w3[7][36] , \w3[7][35] , 
        \w3[7][34] , \w3[7][33] , \w3[7][32] , \w3[7][63] , \w3[7][62] , 
        \w3[7][61] , \w3[7][60] , \w3[7][59] , \w3[7][58] , \w3[7][57] , 
        \w3[7][56] , \w3[7][87] , \w3[7][86] , \w3[7][85] , \w3[7][84] , 
        \w3[7][83] , \w3[7][82] , \w3[7][81] , \w3[7][80] , \w3[7][111] , 
        \w3[7][110] , \w3[7][109] , \w3[7][108] , \w3[7][107] , \w3[7][106] , 
        \w3[7][105] , \w3[7][104] , \w3[7][7] , \w3[7][6] , \w3[7][5] , 
        \w3[7][4] , \w3[7][3] , \w3[7][2] , \w3[7][1] , \w3[7][0] , 
        \w3[7][31] , \w3[7][30] , \w3[7][29] , \w3[7][28] , \w3[7][27] , 
        \w3[7][26] , \w3[7][25] , \w3[7][24] , \w3[7][55] , \w3[7][54] , 
        \w3[7][53] , \w3[7][52] , \w3[7][51] , \w3[7][50] , \w3[7][49] , 
        \w3[7][48] , \w3[7][79] , \w3[7][78] , \w3[7][77] , \w3[7][76] , 
        \w3[7][75] , \w3[7][74] , \w3[7][73] , \w3[7][72] , \w3[7][103] , 
        \w3[7][102] , \w3[7][101] , \w3[7][100] , \w3[7][99] , \w3[7][98] , 
        \w3[7][97] , \w3[7][96] }) );
  SubBytes_9 \SUBBYTES[8].a  ( .x({\w1[8][127] , \w1[8][126] , \w1[8][125] , 
        \w1[8][124] , \w1[8][123] , \w1[8][122] , \w1[8][121] , \w1[8][120] , 
        \w1[8][119] , \w1[8][118] , \w1[8][117] , \w1[8][116] , \w1[8][115] , 
        \w1[8][114] , \w1[8][113] , \w1[8][112] , \w1[8][111] , \w1[8][110] , 
        \w1[8][109] , \w1[8][108] , \w1[8][107] , \w1[8][106] , \w1[8][105] , 
        \w1[8][104] , \w1[8][103] , \w1[8][102] , \w1[8][101] , \w1[8][100] , 
        \w1[8][99] , \w1[8][98] , \w1[8][97] , \w1[8][96] , \w1[8][95] , 
        \w1[8][94] , \w1[8][93] , \w1[8][92] , \w1[8][91] , \w1[8][90] , 
        \w1[8][89] , \w1[8][88] , \w1[8][87] , \w1[8][86] , \w1[8][85] , 
        \w1[8][84] , \w1[8][83] , \w1[8][82] , \w1[8][81] , \w1[8][80] , 
        \w1[8][79] , \w1[8][78] , \w1[8][77] , \w1[8][76] , \w1[8][75] , 
        \w1[8][74] , \w1[8][73] , \w1[8][72] , \w1[8][71] , \w1[8][70] , 
        \w1[8][69] , \w1[8][68] , \w1[8][67] , \w1[8][66] , \w1[8][65] , 
        \w1[8][64] , \w1[8][63] , \w1[8][62] , \w1[8][61] , \w1[8][60] , 
        \w1[8][59] , \w1[8][58] , \w1[8][57] , \w1[8][56] , \w1[8][55] , 
        \w1[8][54] , \w1[8][53] , \w1[8][52] , \w1[8][51] , \w1[8][50] , 
        \w1[8][49] , \w1[8][48] , \w1[8][47] , \w1[8][46] , \w1[8][45] , 
        \w1[8][44] , \w1[8][43] , \w1[8][42] , \w1[8][41] , \w1[8][40] , 
        \w1[8][39] , \w1[8][38] , \w1[8][37] , \w1[8][36] , \w1[8][35] , 
        \w1[8][34] , \w1[8][33] , \w1[8][32] , \w1[8][31] , \w1[8][30] , 
        \w1[8][29] , \w1[8][28] , \w1[8][27] , \w1[8][26] , \w1[8][25] , 
        \w1[8][24] , \w1[8][23] , \w1[8][22] , \w1[8][21] , \w1[8][20] , 
        \w1[8][19] , \w1[8][18] , \w1[8][17] , \w1[8][16] , \w1[8][15] , 
        \w1[8][14] , \w1[8][13] , \w1[8][12] , \w1[8][11] , \w1[8][10] , 
        \w1[8][9] , \w1[8][8] , \w1[8][7] , \w1[8][6] , \w1[8][5] , \w1[8][4] , 
        \w1[8][3] , \w1[8][2] , \w1[8][1] , \w1[8][0] }), .z({\w3[8][127] , 
        \w3[8][126] , \w3[8][125] , \w3[8][124] , \w3[8][123] , \w3[8][122] , 
        \w3[8][121] , \w3[8][120] , \w3[8][23] , \w3[8][22] , \w3[8][21] , 
        \w3[8][20] , \w3[8][19] , \w3[8][18] , \w3[8][17] , \w3[8][16] , 
        \w3[8][47] , \w3[8][46] , \w3[8][45] , \w3[8][44] , \w3[8][43] , 
        \w3[8][42] , \w3[8][41] , \w3[8][40] , \w3[8][71] , \w3[8][70] , 
        \w3[8][69] , \w3[8][68] , \w3[8][67] , \w3[8][66] , \w3[8][65] , 
        \w3[8][64] , \w3[8][95] , \w3[8][94] , \w3[8][93] , \w3[8][92] , 
        \w3[8][91] , \w3[8][90] , \w3[8][89] , \w3[8][88] , \w3[8][119] , 
        \w3[8][118] , \w3[8][117] , \w3[8][116] , \w3[8][115] , \w3[8][114] , 
        \w3[8][113] , \w3[8][112] , \w3[8][15] , \w3[8][14] , \w3[8][13] , 
        \w3[8][12] , \w3[8][11] , \w3[8][10] , \w3[8][9] , \w3[8][8] , 
        \w3[8][39] , \w3[8][38] , \w3[8][37] , \w3[8][36] , \w3[8][35] , 
        \w3[8][34] , \w3[8][33] , \w3[8][32] , \w3[8][63] , \w3[8][62] , 
        \w3[8][61] , \w3[8][60] , \w3[8][59] , \w3[8][58] , \w3[8][57] , 
        \w3[8][56] , \w3[8][87] , \w3[8][86] , \w3[8][85] , \w3[8][84] , 
        \w3[8][83] , \w3[8][82] , \w3[8][81] , \w3[8][80] , \w3[8][111] , 
        \w3[8][110] , \w3[8][109] , \w3[8][108] , \w3[8][107] , \w3[8][106] , 
        \w3[8][105] , \w3[8][104] , \w3[8][7] , \w3[8][6] , \w3[8][5] , 
        \w3[8][4] , \w3[8][3] , \w3[8][2] , \w3[8][1] , \w3[8][0] , 
        \w3[8][31] , \w3[8][30] , \w3[8][29] , \w3[8][28] , \w3[8][27] , 
        \w3[8][26] , \w3[8][25] , \w3[8][24] , \w3[8][55] , \w3[8][54] , 
        \w3[8][53] , \w3[8][52] , \w3[8][51] , \w3[8][50] , \w3[8][49] , 
        \w3[8][48] , \w3[8][79] , \w3[8][78] , \w3[8][77] , \w3[8][76] , 
        \w3[8][75] , \w3[8][74] , \w3[8][73] , \w3[8][72] , \w3[8][103] , 
        \w3[8][102] , \w3[8][101] , \w3[8][100] , \w3[8][99] , \w3[8][98] , 
        \w3[8][97] , \w3[8][96] }) );
  SubBytes_8 \SUBBYTES[9].a  ( .x({\w1[9][127] , \w1[9][126] , \w1[9][125] , 
        \w1[9][124] , \w1[9][123] , \w1[9][122] , \w1[9][121] , \w1[9][120] , 
        \w1[9][119] , \w1[9][118] , \w1[9][117] , \w1[9][116] , \w1[9][115] , 
        \w1[9][114] , \w1[9][113] , \w1[9][112] , \w1[9][111] , \w1[9][110] , 
        \w1[9][109] , \w1[9][108] , \w1[9][107] , \w1[9][106] , \w1[9][105] , 
        \w1[9][104] , \w1[9][103] , \w1[9][102] , \w1[9][101] , \w1[9][100] , 
        \w1[9][99] , \w1[9][98] , \w1[9][97] , \w1[9][96] , \w1[9][95] , 
        \w1[9][94] , \w1[9][93] , \w1[9][92] , \w1[9][91] , \w1[9][90] , 
        \w1[9][89] , \w1[9][88] , \w1[9][87] , \w1[9][86] , \w1[9][85] , 
        \w1[9][84] , \w1[9][83] , \w1[9][82] , \w1[9][81] , \w1[9][80] , 
        \w1[9][79] , \w1[9][78] , \w1[9][77] , \w1[9][76] , \w1[9][75] , 
        \w1[9][74] , \w1[9][73] , \w1[9][72] , \w1[9][71] , \w1[9][70] , 
        \w1[9][69] , \w1[9][68] , \w1[9][67] , \w1[9][66] , \w1[9][65] , 
        \w1[9][64] , \w1[9][63] , \w1[9][62] , \w1[9][61] , \w1[9][60] , 
        \w1[9][59] , \w1[9][58] , \w1[9][57] , \w1[9][56] , \w1[9][55] , 
        \w1[9][54] , \w1[9][53] , \w1[9][52] , \w1[9][51] , \w1[9][50] , 
        \w1[9][49] , \w1[9][48] , \w1[9][47] , \w1[9][46] , \w1[9][45] , 
        \w1[9][44] , \w1[9][43] , \w1[9][42] , \w1[9][41] , \w1[9][40] , 
        \w1[9][39] , \w1[9][38] , \w1[9][37] , \w1[9][36] , \w1[9][35] , 
        \w1[9][34] , \w1[9][33] , \w1[9][32] , \w1[9][31] , \w1[9][30] , 
        \w1[9][29] , \w1[9][28] , \w1[9][27] , \w1[9][26] , \w1[9][25] , 
        \w1[9][24] , \w1[9][23] , \w1[9][22] , \w1[9][21] , \w1[9][20] , 
        \w1[9][19] , \w1[9][18] , \w1[9][17] , \w1[9][16] , \w1[9][15] , 
        \w1[9][14] , \w1[9][13] , \w1[9][12] , \w1[9][11] , \w1[9][10] , 
        \w1[9][9] , \w1[9][8] , \w1[9][7] , \w1[9][6] , \w1[9][5] , \w1[9][4] , 
        \w1[9][3] , \w1[9][2] , \w1[9][1] , \w1[9][0] }), .z({\w3[9][127] , 
        \w3[9][126] , \w3[9][125] , \w3[9][124] , \w3[9][123] , \w3[9][122] , 
        \w3[9][121] , \w3[9][120] , \w3[9][23] , \w3[9][22] , \w3[9][21] , 
        \w3[9][20] , \w3[9][19] , \w3[9][18] , \w3[9][17] , \w3[9][16] , 
        \w3[9][47] , \w3[9][46] , \w3[9][45] , \w3[9][44] , \w3[9][43] , 
        \w3[9][42] , \w3[9][41] , \w3[9][40] , \w3[9][71] , \w3[9][70] , 
        \w3[9][69] , \w3[9][68] , \w3[9][67] , \w3[9][66] , \w3[9][65] , 
        \w3[9][64] , \w3[9][95] , \w3[9][94] , \w3[9][93] , \w3[9][92] , 
        \w3[9][91] , \w3[9][90] , \w3[9][89] , \w3[9][88] , \w3[9][119] , 
        \w3[9][118] , \w3[9][117] , \w3[9][116] , \w3[9][115] , \w3[9][114] , 
        \w3[9][113] , \w3[9][112] , \w3[9][15] , \w3[9][14] , \w3[9][13] , 
        \w3[9][12] , \w3[9][11] , \w3[9][10] , \w3[9][9] , \w3[9][8] , 
        \w3[9][39] , \w3[9][38] , \w3[9][37] , \w3[9][36] , \w3[9][35] , 
        \w3[9][34] , \w3[9][33] , \w3[9][32] , \w3[9][63] , \w3[9][62] , 
        \w3[9][61] , \w3[9][60] , \w3[9][59] , \w3[9][58] , \w3[9][57] , 
        \w3[9][56] , \w3[9][87] , \w3[9][86] , \w3[9][85] , \w3[9][84] , 
        \w3[9][83] , \w3[9][82] , \w3[9][81] , \w3[9][80] , \w3[9][111] , 
        \w3[9][110] , \w3[9][109] , \w3[9][108] , \w3[9][107] , \w3[9][106] , 
        \w3[9][105] , \w3[9][104] , \w3[9][7] , \w3[9][6] , \w3[9][5] , 
        \w3[9][4] , \w3[9][3] , \w3[9][2] , \w3[9][1] , \w3[9][0] , 
        \w3[9][31] , \w3[9][30] , \w3[9][29] , \w3[9][28] , \w3[9][27] , 
        \w3[9][26] , \w3[9][25] , \w3[9][24] , \w3[9][55] , \w3[9][54] , 
        \w3[9][53] , \w3[9][52] , \w3[9][51] , \w3[9][50] , \w3[9][49] , 
        \w3[9][48] , \w3[9][79] , \w3[9][78] , \w3[9][77] , \w3[9][76] , 
        \w3[9][75] , \w3[9][74] , \w3[9][73] , \w3[9][72] , \w3[9][103] , 
        \w3[9][102] , \w3[9][101] , \w3[9][100] , \w3[9][99] , \w3[9][98] , 
        \w3[9][97] , \w3[9][96] }) );
  XOR U5567 ( .A(key[1171]), .B(n7892), .Z(n4159) );
  XNOR U5568 ( .A(\w3[8][11] ), .B(n7918), .Z(n4160) );
  XNOR U5569 ( .A(n4159), .B(n4160), .Z(\w1[9][19] ) );
  XOR U5570 ( .A(key[158]), .B(n4581), .Z(n4161) );
  XNOR U5571 ( .A(\w3[0][6] ), .B(n4720), .Z(n4162) );
  XNOR U5572 ( .A(n4161), .B(n4162), .Z(\w1[1][30] ) );
  XOR U5573 ( .A(key[403]), .B(n5380), .Z(n4163) );
  XNOR U5574 ( .A(\w3[2][11] ), .B(n5406), .Z(n4164) );
  XNOR U5575 ( .A(n4163), .B(n4164), .Z(\w1[3][19] ) );
  XOR U5576 ( .A(key[542]), .B(n5838), .Z(n4165) );
  XNOR U5577 ( .A(\w3[3][6] ), .B(n5976), .Z(n4166) );
  XNOR U5578 ( .A(n4165), .B(n4166), .Z(\w1[4][30] ) );
  XOR U5579 ( .A(key[662]), .B(n6226), .Z(n4167) );
  XNOR U5580 ( .A(\w3[4][14] ), .B(n6258), .Z(n4168) );
  XOR U5581 ( .A(n4167), .B(n4168), .Z(\w1[5][22] ) );
  XOR U5582 ( .A(\w3[4][1] ), .B(\w3[4][26] ), .Z(n4169) );
  XNOR U5583 ( .A(n6233), .B(key[665]), .Z(n4170) );
  XNOR U5584 ( .A(n4169), .B(n4170), .Z(n4171) );
  XNOR U5585 ( .A(n4171), .B(\w3[4][18] ), .Z(\w1[5][25] ) );
  XOR U5586 ( .A(key[798]), .B(n6680), .Z(n4172) );
  XNOR U5587 ( .A(\w3[5][6] ), .B(n6815), .Z(n4173) );
  XNOR U5588 ( .A(n4172), .B(n4173), .Z(\w1[6][30] ) );
  XOR U5589 ( .A(key[926]), .B(n7094), .Z(n4174) );
  XNOR U5590 ( .A(\w3[6][6] ), .B(n7229), .Z(n4175) );
  XNOR U5591 ( .A(n4174), .B(n4175), .Z(\w1[7][30] ) );
  XOR U5592 ( .A(key[1043]), .B(n7466), .Z(n4176) );
  XNOR U5593 ( .A(\w3[7][11] ), .B(n7492), .Z(n4177) );
  XNOR U5594 ( .A(n4176), .B(n4177), .Z(\w1[8][19] ) );
  XOR U5595 ( .A(key[1182]), .B(n7937), .Z(n4178) );
  XNOR U5596 ( .A(\w3[8][6] ), .B(n8073), .Z(n4179) );
  XNOR U5597 ( .A(n4178), .B(n4179), .Z(\w1[9][30] ) );
  XNOR U5598 ( .A(\w3[0][8] ), .B(\w3[0][12] ), .Z(n4180) );
  XNOR U5599 ( .A(n4576), .B(n4180), .Z(n4539) );
  XNOR U5600 ( .A(\w3[0][35] ), .B(\w3[0][59] ), .Z(n4615) );
  XNOR U5601 ( .A(\w3[0][67] ), .B(\w3[0][91] ), .Z(n4736) );
  XNOR U5602 ( .A(\w3[0][80] ), .B(\w3[0][85] ), .Z(n4808) );
  XOR U5603 ( .A(n4766), .B(\w3[0][74] ), .Z(n4181) );
  XNOR U5604 ( .A(n4765), .B(key[210]), .Z(n4182) );
  XNOR U5605 ( .A(n4181), .B(n4182), .Z(\w1[1][82] ) );
  XOR U5606 ( .A(\w3[0][96] ), .B(n4498), .Z(n4183) );
  XNOR U5607 ( .A(key[232]), .B(\w3[0][105] ), .Z(n4184) );
  XNOR U5608 ( .A(n4183), .B(n4184), .Z(n4185) );
  XOR U5609 ( .A(n4185), .B(n4825), .Z(\w1[1][104] ) );
  XOR U5610 ( .A(key[371]), .B(n4890), .Z(n4186) );
  XNOR U5611 ( .A(\w3[1][107] ), .B(n4923), .Z(n4187) );
  XNOR U5612 ( .A(n4186), .B(n4187), .Z(\w1[2][115] ) );
  XNOR U5613 ( .A(\w3[1][8] ), .B(\w3[1][12] ), .Z(n4188) );
  XNOR U5614 ( .A(n4997), .B(n4188), .Z(n4960) );
  XOR U5615 ( .A(key[150]), .B(n4549), .Z(n4189) );
  XNOR U5616 ( .A(\w3[0][14] ), .B(n4581), .Z(n4190) );
  XOR U5617 ( .A(n4189), .B(n4190), .Z(\w1[1][22] ) );
  XOR U5618 ( .A(\w3[0][1] ), .B(\w3[0][26] ), .Z(n4191) );
  XNOR U5619 ( .A(n4556), .B(key[153]), .Z(n4192) );
  XNOR U5620 ( .A(n4191), .B(n4192), .Z(n4193) );
  XNOR U5621 ( .A(n4193), .B(\w3[0][18] ), .Z(\w1[1][25] ) );
  XNOR U5622 ( .A(\w3[1][48] ), .B(\w3[1][53] ), .Z(n5109) );
  XNOR U5623 ( .A(\w3[1][80] ), .B(\w3[1][85] ), .Z(n5228) );
  XNOR U5624 ( .A(\w3[1][67] ), .B(\w3[1][91] ), .Z(n5156) );
  XOR U5625 ( .A(n5186), .B(\w3[1][74] ), .Z(n4194) );
  XNOR U5626 ( .A(n5185), .B(key[338]), .Z(n4195) );
  XNOR U5627 ( .A(n4194), .B(n4195), .Z(\w1[2][82] ) );
  XOR U5628 ( .A(key[307]), .B(n5069), .Z(n4196) );
  XNOR U5629 ( .A(\w3[1][43] ), .B(n5100), .Z(n4197) );
  XNOR U5630 ( .A(n4196), .B(n4197), .Z(\w1[2][51] ) );
  XOR U5631 ( .A(key[278]), .B(n4970), .Z(n4198) );
  XNOR U5632 ( .A(\w3[1][14] ), .B(n5002), .Z(n4199) );
  XOR U5633 ( .A(n4198), .B(n4199), .Z(\w1[2][22] ) );
  XNOR U5634 ( .A(\w3[2][8] ), .B(\w3[2][12] ), .Z(n4200) );
  XNOR U5635 ( .A(n5420), .B(n4200), .Z(n5380) );
  XOR U5636 ( .A(\w3[1][1] ), .B(\w3[1][26] ), .Z(n4201) );
  XNOR U5637 ( .A(n4977), .B(key[281]), .Z(n4202) );
  XNOR U5638 ( .A(n4201), .B(n4202), .Z(n4203) );
  XNOR U5639 ( .A(n4203), .B(\w3[1][18] ), .Z(\w1[2][25] ) );
  XOR U5640 ( .A(key[467]), .B(n5610), .Z(n4204) );
  XNOR U5641 ( .A(\w3[2][75] ), .B(n5646), .Z(n4205) );
  XNOR U5642 ( .A(n4204), .B(n4205), .Z(\w1[3][83] ) );
  XNOR U5643 ( .A(\w3[2][48] ), .B(\w3[2][53] ), .Z(n5532) );
  XNOR U5644 ( .A(\w3[2][80] ), .B(\w3[2][85] ), .Z(n5651) );
  XOR U5645 ( .A(key[435]), .B(n5492), .Z(n4206) );
  XNOR U5646 ( .A(\w3[2][43] ), .B(n5523), .Z(n4207) );
  XNOR U5647 ( .A(n4206), .B(n4207), .Z(\w1[3][51] ) );
  XOR U5648 ( .A(key[406]), .B(n5388), .Z(n4208) );
  XNOR U5649 ( .A(\w3[2][14] ), .B(n5425), .Z(n4209) );
  XOR U5650 ( .A(n4208), .B(n4209), .Z(\w1[3][22] ) );
  XNOR U5651 ( .A(\w3[3][8] ), .B(\w3[3][12] ), .Z(n4210) );
  XNOR U5652 ( .A(n5833), .B(n4210), .Z(n5796) );
  XNOR U5653 ( .A(\w3[3][48] ), .B(\w3[3][53] ), .Z(n5945) );
  XNOR U5654 ( .A(\w3[3][35] ), .B(\w3[3][59] ), .Z(n5870) );
  XNOR U5655 ( .A(\w3[3][80] ), .B(\w3[3][85] ), .Z(n6064) );
  XOR U5656 ( .A(key[595]), .B(n6023), .Z(n4211) );
  XNOR U5657 ( .A(\w3[3][75] ), .B(n6059), .Z(n4212) );
  XNOR U5658 ( .A(n4211), .B(n4212), .Z(\w1[4][83] ) );
  XOR U5659 ( .A(\w3[3][96] ), .B(n6081), .Z(n4213) );
  XNOR U5660 ( .A(key[616]), .B(\w3[3][105] ), .Z(n4214) );
  XNOR U5661 ( .A(n4213), .B(n4214), .Z(n4215) );
  XNOR U5662 ( .A(\w3[3][97] ), .B(n4215), .Z(\w1[4][104] ) );
  XNOR U5663 ( .A(\w3[4][8] ), .B(\w3[4][12] ), .Z(n4216) );
  XNOR U5664 ( .A(n6253), .B(n4216), .Z(n6216) );
  XOR U5665 ( .A(key[534]), .B(n5806), .Z(n4217) );
  XNOR U5666 ( .A(\w3[3][14] ), .B(n5838), .Z(n4218) );
  XOR U5667 ( .A(n4217), .B(n4218), .Z(\w1[4][22] ) );
  XOR U5668 ( .A(\w3[3][1] ), .B(\w3[3][26] ), .Z(n4219) );
  XNOR U5669 ( .A(n5813), .B(key[537]), .Z(n4220) );
  XNOR U5670 ( .A(n4219), .B(n4220), .Z(n4221) );
  XNOR U5671 ( .A(n4221), .B(\w3[3][18] ), .Z(\w1[4][25] ) );
  XOR U5672 ( .A(key[723]), .B(n6443), .Z(n4222) );
  XNOR U5673 ( .A(\w3[4][75] ), .B(n6480), .Z(n4223) );
  XNOR U5674 ( .A(n4222), .B(n4223), .Z(\w1[5][83] ) );
  XOR U5675 ( .A(key[755]), .B(n6146), .Z(n4224) );
  XNOR U5676 ( .A(\w3[4][107] ), .B(n6179), .Z(n4225) );
  XNOR U5677 ( .A(n4224), .B(n4225), .Z(\w1[5][115] ) );
  XNOR U5678 ( .A(\w3[4][48] ), .B(\w3[4][53] ), .Z(n6362) );
  XOR U5679 ( .A(key[691]), .B(n6322), .Z(n4226) );
  XNOR U5680 ( .A(\w3[4][43] ), .B(n6353), .Z(n4227) );
  XNOR U5681 ( .A(n4226), .B(n4227), .Z(\w1[5][51] ) );
  XNOR U5682 ( .A(\w3[5][8] ), .B(\w3[5][12] ), .Z(n4228) );
  XNOR U5683 ( .A(n6675), .B(n4228), .Z(n6638) );
  XNOR U5684 ( .A(\w3[5][80] ), .B(\w3[5][85] ), .Z(n6903) );
  XOR U5685 ( .A(key[670]), .B(n6258), .Z(n4229) );
  XNOR U5686 ( .A(\w3[4][6] ), .B(n6394), .Z(n4230) );
  XNOR U5687 ( .A(n4229), .B(n4230), .Z(\w1[5][30] ) );
  XOR U5688 ( .A(key[851]), .B(n6862), .Z(n4231) );
  XNOR U5689 ( .A(\w3[5][75] ), .B(n6898), .Z(n4232) );
  XNOR U5690 ( .A(n4231), .B(n4232), .Z(\w1[6][83] ) );
  XNOR U5691 ( .A(\w3[5][48] ), .B(\w3[5][53] ), .Z(n6784) );
  XOR U5692 ( .A(key[883]), .B(n6567), .Z(n4233) );
  XNOR U5693 ( .A(\w3[5][107] ), .B(n6601), .Z(n4234) );
  XNOR U5694 ( .A(n4233), .B(n4234), .Z(\w1[6][115] ) );
  XNOR U5695 ( .A(\w3[5][35] ), .B(\w3[5][59] ), .Z(n6713) );
  XOR U5696 ( .A(key[790]), .B(n6648), .Z(n4235) );
  XNOR U5697 ( .A(\w3[5][14] ), .B(n6680), .Z(n4236) );
  XOR U5698 ( .A(n4235), .B(n4236), .Z(\w1[6][22] ) );
  XOR U5699 ( .A(n6743), .B(\w3[5][42] ), .Z(n4237) );
  XNOR U5700 ( .A(n6742), .B(key[818]), .Z(n4238) );
  XNOR U5701 ( .A(n4237), .B(n4238), .Z(\w1[6][50] ) );
  XNOR U5702 ( .A(\w3[6][67] ), .B(\w3[6][91] ), .Z(n7245) );
  XNOR U5703 ( .A(\w3[6][8] ), .B(\w3[6][12] ), .Z(n4239) );
  XNOR U5704 ( .A(n7089), .B(n4239), .Z(n7052) );
  XNOR U5705 ( .A(\w3[6][48] ), .B(\w3[6][53] ), .Z(n7198) );
  XNOR U5706 ( .A(\w3[6][80] ), .B(\w3[6][85] ), .Z(n7317) );
  XOR U5707 ( .A(\w3[5][1] ), .B(\w3[5][26] ), .Z(n4240) );
  XNOR U5708 ( .A(n6655), .B(key[793]), .Z(n4241) );
  XNOR U5709 ( .A(n4240), .B(n4241), .Z(n4242) );
  XNOR U5710 ( .A(n4242), .B(\w3[5][18] ), .Z(\w1[6][25] ) );
  XOR U5711 ( .A(n7275), .B(\w3[6][74] ), .Z(n4243) );
  XNOR U5712 ( .A(n7274), .B(key[978]), .Z(n4244) );
  XNOR U5713 ( .A(n4243), .B(n4244), .Z(\w1[7][82] ) );
  XNOR U5714 ( .A(\w3[6][35] ), .B(\w3[6][59] ), .Z(n7127) );
  XOR U5715 ( .A(\w3[6][105] ), .B(n7333), .Z(n4245) );
  XNOR U5716 ( .A(n7341), .B(key[1009]), .Z(n4246) );
  XOR U5717 ( .A(n4245), .B(n4246), .Z(\w1[7][113] ) );
  XOR U5718 ( .A(n7157), .B(\w3[6][42] ), .Z(n4247) );
  XNOR U5719 ( .A(n7156), .B(key[946]), .Z(n4248) );
  XNOR U5720 ( .A(n4247), .B(n4248), .Z(\w1[7][50] ) );
  XNOR U5721 ( .A(\w3[7][48] ), .B(\w3[7][53] ), .Z(n7623) );
  XOR U5722 ( .A(key[918]), .B(n7062), .Z(n4249) );
  XNOR U5723 ( .A(\w3[6][14] ), .B(n7094), .Z(n4250) );
  XOR U5724 ( .A(n4249), .B(n4250), .Z(\w1[7][22] ) );
  XNOR U5725 ( .A(\w3[7][35] ), .B(\w3[7][59] ), .Z(n7549) );
  XNOR U5726 ( .A(\w3[7][80] ), .B(\w3[7][85] ), .Z(n7742) );
  XNOR U5727 ( .A(\w3[7][67] ), .B(\w3[7][91] ), .Z(n7670) );
  XNOR U5728 ( .A(\w3[7][8] ), .B(\w3[7][12] ), .Z(n4251) );
  XNOR U5729 ( .A(n7506), .B(n4251), .Z(n7466) );
  XOR U5730 ( .A(\w3[6][1] ), .B(\w3[6][26] ), .Z(n4252) );
  XNOR U5731 ( .A(n7069), .B(key[921]), .Z(n4253) );
  XNOR U5732 ( .A(n4252), .B(n4253), .Z(n4254) );
  XNOR U5733 ( .A(n4254), .B(\w3[6][18] ), .Z(\w1[7][25] ) );
  XOR U5734 ( .A(n7700), .B(\w3[7][74] ), .Z(n4255) );
  XNOR U5735 ( .A(n7699), .B(key[1106]), .Z(n4256) );
  XNOR U5736 ( .A(n4255), .B(n4256), .Z(\w1[8][82] ) );
  XOR U5737 ( .A(key[1147]), .B(n7432), .Z(n4257) );
  XNOR U5738 ( .A(\w3[7][99] ), .B(n7770), .Z(n4258) );
  XOR U5739 ( .A(n4257), .B(n4258), .Z(\w1[8][123] ) );
  XNOR U5740 ( .A(\w3[8][35] ), .B(\w3[8][59] ), .Z(n7970) );
  XNOR U5741 ( .A(\w3[8][67] ), .B(\w3[8][91] ), .Z(n8092) );
  XNOR U5742 ( .A(\w3[8][8] ), .B(\w3[8][12] ), .Z(n4259) );
  XNOR U5743 ( .A(n7932), .B(n4259), .Z(n7892) );
  XNOR U5744 ( .A(\w3[8][48] ), .B(\w3[8][53] ), .Z(n8042) );
  XOR U5745 ( .A(key[1046]), .B(n7474), .Z(n4260) );
  XNOR U5746 ( .A(\w3[7][14] ), .B(n7511), .Z(n4261) );
  XOR U5747 ( .A(n4260), .B(n4261), .Z(\w1[8][22] ) );
  XOR U5748 ( .A(key[1174]), .B(n7900), .Z(n4262) );
  XNOR U5749 ( .A(\w3[8][14] ), .B(n7937), .Z(n4263) );
  XOR U5750 ( .A(n4262), .B(n4263), .Z(\w1[9][22] ) );
  XOR U5751 ( .A(n8025), .B(\w3[8][58] ), .Z(n4264) );
  XNOR U5752 ( .A(\w3[8][50] ), .B(key[1209]), .Z(n4265) );
  XNOR U5753 ( .A(n4264), .B(n4265), .Z(n4266) );
  XOR U5754 ( .A(n8026), .B(n4266), .Z(\w1[9][57] ) );
  XNOR U5755 ( .A(\w3[0][48] ), .B(\w3[0][53] ), .Z(n4689) );
  XOR U5756 ( .A(key[179]), .B(n4648), .Z(n4267) );
  XNOR U5757 ( .A(\w3[0][43] ), .B(n4680), .Z(n4268) );
  XNOR U5758 ( .A(n4267), .B(n4268), .Z(\w1[1][51] ) );
  XOR U5759 ( .A(key[211]), .B(n4767), .Z(n4269) );
  XNOR U5760 ( .A(\w3[0][75] ), .B(n4803), .Z(n4270) );
  XNOR U5761 ( .A(n4269), .B(n4270), .Z(\w1[1][83] ) );
  XOR U5762 ( .A(\w3[0][65] ), .B(\w3[0][73] ), .Z(n4271) );
  XNOR U5763 ( .A(\w3[0][64] ), .B(key[200]), .Z(n4272) );
  XNOR U5764 ( .A(n4271), .B(n4272), .Z(n4273) );
  XNOR U5765 ( .A(n4821), .B(n4273), .Z(\w1[1][72] ) );
  XOR U5766 ( .A(n4665), .B(n4679), .Z(n4274) );
  XNOR U5767 ( .A(\w3[0][42] ), .B(key[169]), .Z(n4275) );
  XNOR U5768 ( .A(n4274), .B(n4275), .Z(n4276) );
  XNOR U5769 ( .A(\w3[0][33] ), .B(n4276), .Z(\w1[1][41] ) );
  XOR U5770 ( .A(key[251]), .B(n4505), .Z(n4277) );
  XNOR U5771 ( .A(\w3[0][99] ), .B(n4836), .Z(n4278) );
  XOR U5772 ( .A(n4277), .B(n4278), .Z(\w1[1][123] ) );
  XOR U5773 ( .A(\w3[0][25] ), .B(n4554), .Z(n4279) );
  XNOR U5774 ( .A(\w3[0][17] ), .B(key[152]), .Z(n4280) );
  XNOR U5775 ( .A(n4279), .B(n4280), .Z(n4281) );
  XNOR U5776 ( .A(n4555), .B(n4281), .Z(\w1[1][24] ) );
  XNOR U5777 ( .A(\w3[1][35] ), .B(\w3[1][59] ), .Z(n5038) );
  XOR U5778 ( .A(key[339]), .B(n5187), .Z(n4282) );
  XNOR U5779 ( .A(\w3[1][75] ), .B(n5223), .Z(n4283) );
  XNOR U5780 ( .A(n4282), .B(n4283), .Z(\w1[2][83] ) );
  XOR U5781 ( .A(key[149]), .B(n4548), .Z(n4284) );
  XNOR U5782 ( .A(\w3[0][13] ), .B(n4580), .Z(n4285) );
  XNOR U5783 ( .A(n4284), .B(n4285), .Z(\w1[1][21] ) );
  XOR U5784 ( .A(n5068), .B(\w3[1][42] ), .Z(n4286) );
  XNOR U5785 ( .A(n5067), .B(key[306]), .Z(n4287) );
  XNOR U5786 ( .A(n4286), .B(n4287), .Z(\w1[2][50] ) );
  XOR U5787 ( .A(\w3[1][96] ), .B(n4915), .Z(n4288) );
  XNOR U5788 ( .A(key[360]), .B(\w3[1][105] ), .Z(n4289) );
  XNOR U5789 ( .A(n4288), .B(n4289), .Z(n4290) );
  XOR U5790 ( .A(n4290), .B(n5245), .Z(\w1[2][104] ) );
  XOR U5791 ( .A(\w3[1][65] ), .B(\w3[1][73] ), .Z(n4291) );
  XNOR U5792 ( .A(\w3[1][64] ), .B(key[328]), .Z(n4292) );
  XNOR U5793 ( .A(n4291), .B(n4292), .Z(n4293) );
  XNOR U5794 ( .A(n5241), .B(n4293), .Z(\w1[2][72] ) );
  XOR U5795 ( .A(\w3[1][33] ), .B(\w3[1][41] ), .Z(n4294) );
  XNOR U5796 ( .A(\w3[1][32] ), .B(key[296]), .Z(n4295) );
  XNOR U5797 ( .A(n4294), .B(n4295), .Z(n4296) );
  XNOR U5798 ( .A(n5122), .B(n4296), .Z(\w1[2][40] ) );
  XOR U5799 ( .A(\w3[1][25] ), .B(n4975), .Z(n4297) );
  XNOR U5800 ( .A(\w3[1][17] ), .B(key[280]), .Z(n4298) );
  XNOR U5801 ( .A(n4297), .B(n4298), .Z(n4299) );
  XNOR U5802 ( .A(n4976), .B(n4299), .Z(\w1[2][24] ) );
  XOR U5803 ( .A(n5609), .B(\w3[2][74] ), .Z(n4300) );
  XNOR U5804 ( .A(n5608), .B(key[466]), .Z(n4301) );
  XNOR U5805 ( .A(n4300), .B(n4301), .Z(\w1[3][82] ) );
  XNOR U5806 ( .A(\w3[2][35] ), .B(\w3[2][59] ), .Z(n5461) );
  XNOR U5807 ( .A(\w3[2][67] ), .B(\w3[2][91] ), .Z(n5579) );
  XOR U5808 ( .A(key[277]), .B(n4969), .Z(n4302) );
  XNOR U5809 ( .A(\w3[1][13] ), .B(n5001), .Z(n4303) );
  XNOR U5810 ( .A(n4302), .B(n4303), .Z(\w1[2][21] ) );
  XOR U5811 ( .A(\w3[2][96] ), .B(n5336), .Z(n4304) );
  XNOR U5812 ( .A(key[488]), .B(\w3[2][105] ), .Z(n4305) );
  XNOR U5813 ( .A(n4304), .B(n4305), .Z(n4306) );
  XOR U5814 ( .A(n4306), .B(n5668), .Z(\w1[3][104] ) );
  XOR U5815 ( .A(n5491), .B(\w3[2][42] ), .Z(n4307) );
  XNOR U5816 ( .A(n5490), .B(key[434]), .Z(n4308) );
  XNOR U5817 ( .A(n4307), .B(n4308), .Z(\w1[3][50] ) );
  XOR U5818 ( .A(\w3[2][33] ), .B(\w3[2][41] ), .Z(n4309) );
  XNOR U5819 ( .A(\w3[2][32] ), .B(key[424]), .Z(n4310) );
  XNOR U5820 ( .A(n4309), .B(n4310), .Z(n4311) );
  XNOR U5821 ( .A(n5545), .B(n4311), .Z(\w1[3][40] ) );
  XOR U5822 ( .A(\w3[2][65] ), .B(\w3[2][73] ), .Z(n4312) );
  XNOR U5823 ( .A(\w3[2][64] ), .B(key[456]), .Z(n4313) );
  XNOR U5824 ( .A(n4312), .B(n4313), .Z(n4314) );
  XNOR U5825 ( .A(n5664), .B(n4314), .Z(\w1[3][72] ) );
  XOR U5826 ( .A(\w3[2][25] ), .B(n5393), .Z(n4315) );
  XNOR U5827 ( .A(\w3[2][17] ), .B(key[408]), .Z(n4316) );
  XNOR U5828 ( .A(n4315), .B(n4316), .Z(n4317) );
  XNOR U5829 ( .A(n5394), .B(n4317), .Z(\w1[3][24] ) );
  XOR U5830 ( .A(key[405]), .B(n5387), .Z(n4318) );
  XNOR U5831 ( .A(\w3[2][13] ), .B(n5424), .Z(n4319) );
  XNOR U5832 ( .A(n4318), .B(n4319), .Z(\w1[3][21] ) );
  XOR U5833 ( .A(key[563]), .B(n5904), .Z(n4320) );
  XNOR U5834 ( .A(\w3[3][43] ), .B(n5936), .Z(n4321) );
  XNOR U5835 ( .A(n4320), .B(n4321), .Z(\w1[4][51] ) );
  XOR U5836 ( .A(n6022), .B(\w3[3][74] ), .Z(n4322) );
  XNOR U5837 ( .A(n6021), .B(key[594]), .Z(n4323) );
  XNOR U5838 ( .A(n4322), .B(n4323), .Z(\w1[4][82] ) );
  XNOR U5839 ( .A(\w3[3][67] ), .B(\w3[3][91] ), .Z(n5992) );
  XOR U5840 ( .A(key[635]), .B(n5762), .Z(n4324) );
  XNOR U5841 ( .A(\w3[3][99] ), .B(n6092), .Z(n4325) );
  XOR U5842 ( .A(n4324), .B(n4325), .Z(\w1[4][123] ) );
  XOR U5843 ( .A(n5921), .B(n5935), .Z(n4326) );
  XNOR U5844 ( .A(\w3[3][42] ), .B(key[553]), .Z(n4327) );
  XNOR U5845 ( .A(n4326), .B(n4327), .Z(n4328) );
  XNOR U5846 ( .A(\w3[3][33] ), .B(n4328), .Z(\w1[4][41] ) );
  XOR U5847 ( .A(\w3[3][105] ), .B(n6080), .Z(n4329) );
  XNOR U5848 ( .A(n6088), .B(key[625]), .Z(n4330) );
  XOR U5849 ( .A(n4329), .B(n4330), .Z(\w1[4][113] ) );
  XOR U5850 ( .A(\w3[3][65] ), .B(\w3[3][73] ), .Z(n4331) );
  XNOR U5851 ( .A(\w3[3][64] ), .B(key[584]), .Z(n4332) );
  XNOR U5852 ( .A(n4331), .B(n4332), .Z(n4333) );
  XNOR U5853 ( .A(n6077), .B(n4333), .Z(\w1[4][72] ) );
  XNOR U5854 ( .A(\w3[4][80] ), .B(\w3[4][85] ), .Z(n6485) );
  XOR U5855 ( .A(\w3[3][25] ), .B(n5811), .Z(n4334) );
  XNOR U5856 ( .A(\w3[3][17] ), .B(key[536]), .Z(n4335) );
  XNOR U5857 ( .A(n4334), .B(n4335), .Z(n4336) );
  XNOR U5858 ( .A(n5812), .B(n4336), .Z(\w1[4][24] ) );
  XNOR U5859 ( .A(\w3[4][35] ), .B(\w3[4][59] ), .Z(n6291) );
  XNOR U5860 ( .A(\w3[4][67] ), .B(\w3[4][91] ), .Z(n6410) );
  XOR U5861 ( .A(key[533]), .B(n5805), .Z(n4337) );
  XNOR U5862 ( .A(\w3[3][13] ), .B(n5837), .Z(n4338) );
  XNOR U5863 ( .A(n4337), .B(n4338), .Z(\w1[4][21] ) );
  XOR U5864 ( .A(n6321), .B(\w3[4][42] ), .Z(n4339) );
  XNOR U5865 ( .A(n6320), .B(key[690]), .Z(n4340) );
  XNOR U5866 ( .A(n4339), .B(n4340), .Z(\w1[5][50] ) );
  XOR U5867 ( .A(n6460), .B(n6479), .Z(n4341) );
  XNOR U5868 ( .A(\w3[4][74] ), .B(key[713]), .Z(n4342) );
  XNOR U5869 ( .A(n4341), .B(n4342), .Z(n4343) );
  XNOR U5870 ( .A(\w3[4][65] ), .B(n4343), .Z(\w1[5][73] ) );
  XOR U5871 ( .A(\w3[4][96] ), .B(n6171), .Z(n4344) );
  XNOR U5872 ( .A(key[744]), .B(\w3[4][105] ), .Z(n4345) );
  XNOR U5873 ( .A(n4344), .B(n4345), .Z(n4346) );
  XOR U5874 ( .A(n4346), .B(n6502), .Z(\w1[5][104] ) );
  XOR U5875 ( .A(\w3[4][33] ), .B(\w3[4][41] ), .Z(n4347) );
  XNOR U5876 ( .A(\w3[4][32] ), .B(key[680]), .Z(n4348) );
  XNOR U5877 ( .A(n4347), .B(n4348), .Z(n4349) );
  XNOR U5878 ( .A(n6375), .B(n4349), .Z(\w1[5][40] ) );
  XNOR U5879 ( .A(\w3[5][67] ), .B(\w3[5][91] ), .Z(n6831) );
  XOR U5880 ( .A(\w3[4][25] ), .B(n6231), .Z(n4350) );
  XNOR U5881 ( .A(\w3[4][17] ), .B(key[664]), .Z(n4351) );
  XNOR U5882 ( .A(n4350), .B(n4351), .Z(n4352) );
  XNOR U5883 ( .A(n6232), .B(n4352), .Z(\w1[5][24] ) );
  XOR U5884 ( .A(n6861), .B(\w3[5][74] ), .Z(n4353) );
  XNOR U5885 ( .A(n6860), .B(key[850]), .Z(n4354) );
  XNOR U5886 ( .A(n4353), .B(n4354), .Z(\w1[6][82] ) );
  XOR U5887 ( .A(key[661]), .B(n6225), .Z(n4355) );
  XNOR U5888 ( .A(\w3[4][13] ), .B(n6257), .Z(n4356) );
  XNOR U5889 ( .A(n4355), .B(n4356), .Z(\w1[5][21] ) );
  XOR U5890 ( .A(\w3[5][96] ), .B(n6590), .Z(n4357) );
  XNOR U5891 ( .A(key[872]), .B(\w3[5][105] ), .Z(n4358) );
  XNOR U5892 ( .A(n4357), .B(n4358), .Z(n4359) );
  XOR U5893 ( .A(n4359), .B(n6920), .Z(\w1[6][104] ) );
  XOR U5894 ( .A(\w3[5][33] ), .B(\w3[5][41] ), .Z(n4360) );
  XNOR U5895 ( .A(\w3[5][32] ), .B(key[808]), .Z(n4361) );
  XNOR U5896 ( .A(n4360), .B(n4361), .Z(n4362) );
  XNOR U5897 ( .A(n6797), .B(n4362), .Z(\w1[6][40] ) );
  XOR U5898 ( .A(key[819]), .B(n6744), .Z(n4363) );
  XNOR U5899 ( .A(\w3[5][43] ), .B(n6775), .Z(n4364) );
  XNOR U5900 ( .A(n4363), .B(n4364), .Z(\w1[6][51] ) );
  XOR U5901 ( .A(\w3[5][65] ), .B(\w3[5][73] ), .Z(n4365) );
  XNOR U5902 ( .A(\w3[5][64] ), .B(key[840]), .Z(n4366) );
  XNOR U5903 ( .A(n4365), .B(n4366), .Z(n4367) );
  XNOR U5904 ( .A(n6916), .B(n4367), .Z(\w1[6][72] ) );
  XOR U5905 ( .A(\w3[5][25] ), .B(n6653), .Z(n4368) );
  XNOR U5906 ( .A(\w3[5][17] ), .B(key[792]), .Z(n4369) );
  XNOR U5907 ( .A(n4368), .B(n4369), .Z(n4370) );
  XNOR U5908 ( .A(n6654), .B(n4370), .Z(\w1[6][24] ) );
  XOR U5909 ( .A(key[979]), .B(n7276), .Z(n4371) );
  XNOR U5910 ( .A(\w3[6][75] ), .B(n7312), .Z(n4372) );
  XNOR U5911 ( .A(n4371), .B(n4372), .Z(\w1[7][83] ) );
  XOR U5912 ( .A(key[789]), .B(n6647), .Z(n4373) );
  XNOR U5913 ( .A(\w3[5][13] ), .B(n6679), .Z(n4374) );
  XNOR U5914 ( .A(n4373), .B(n4374), .Z(\w1[6][21] ) );
  XOR U5915 ( .A(\w3[6][96] ), .B(n7334), .Z(n4375) );
  XNOR U5916 ( .A(key[1000]), .B(\w3[6][105] ), .Z(n4376) );
  XNOR U5917 ( .A(n4375), .B(n4376), .Z(n4377) );
  XNOR U5918 ( .A(\w3[6][97] ), .B(n4377), .Z(\w1[7][104] ) );
  XOR U5919 ( .A(key[947]), .B(n7158), .Z(n4378) );
  XNOR U5920 ( .A(\w3[6][43] ), .B(n7189), .Z(n4379) );
  XNOR U5921 ( .A(n4378), .B(n4379), .Z(\w1[7][51] ) );
  XOR U5922 ( .A(\w3[6][33] ), .B(\w3[6][41] ), .Z(n4380) );
  XNOR U5923 ( .A(\w3[6][32] ), .B(key[936]), .Z(n4381) );
  XNOR U5924 ( .A(n4380), .B(n4381), .Z(n4382) );
  XNOR U5925 ( .A(n7211), .B(n4382), .Z(\w1[7][40] ) );
  XOR U5926 ( .A(\w3[6][65] ), .B(\w3[6][73] ), .Z(n4383) );
  XNOR U5927 ( .A(\w3[6][64] ), .B(key[968]), .Z(n4384) );
  XNOR U5928 ( .A(n4383), .B(n4384), .Z(n4385) );
  XNOR U5929 ( .A(n7330), .B(n4385), .Z(\w1[7][72] ) );
  XOR U5930 ( .A(\w3[6][25] ), .B(n7067), .Z(n4386) );
  XNOR U5931 ( .A(\w3[6][17] ), .B(key[920]), .Z(n4387) );
  XNOR U5932 ( .A(n4386), .B(n4387), .Z(n4388) );
  XNOR U5933 ( .A(n7068), .B(n4388), .Z(\w1[7][24] ) );
  XOR U5934 ( .A(key[1075]), .B(n7583), .Z(n4389) );
  XNOR U5935 ( .A(\w3[7][43] ), .B(n7614), .Z(n4390) );
  XNOR U5936 ( .A(n4389), .B(n4390), .Z(\w1[8][51] ) );
  XOR U5937 ( .A(key[917]), .B(n7061), .Z(n4391) );
  XNOR U5938 ( .A(\w3[6][13] ), .B(n7093), .Z(n4392) );
  XNOR U5939 ( .A(n4391), .B(n4392), .Z(\w1[7][21] ) );
  XOR U5940 ( .A(key[1107]), .B(n7701), .Z(n4393) );
  XNOR U5941 ( .A(\w3[7][75] ), .B(n7737), .Z(n4394) );
  XNOR U5942 ( .A(n4393), .B(n4394), .Z(\w1[8][83] ) );
  XOR U5943 ( .A(\w3[7][96] ), .B(n7425), .Z(n4395) );
  XNOR U5944 ( .A(key[1128]), .B(\w3[7][105] ), .Z(n4396) );
  XNOR U5945 ( .A(n4395), .B(n4396), .Z(n4397) );
  XOR U5946 ( .A(n4397), .B(n7759), .Z(\w1[8][104] ) );
  XOR U5947 ( .A(\w3[7][65] ), .B(\w3[7][73] ), .Z(n4398) );
  XNOR U5948 ( .A(\w3[7][64] ), .B(key[1096]), .Z(n4399) );
  XNOR U5949 ( .A(n4398), .B(n4399), .Z(n4400) );
  XNOR U5950 ( .A(n7755), .B(n4400), .Z(\w1[8][72] ) );
  XOR U5951 ( .A(\w3[7][25] ), .B(n7479), .Z(n4401) );
  XNOR U5952 ( .A(\w3[7][17] ), .B(key[1048]), .Z(n4402) );
  XNOR U5953 ( .A(n4401), .B(n4402), .Z(n4403) );
  XNOR U5954 ( .A(n7480), .B(n4403), .Z(\w1[8][24] ) );
  XNOR U5955 ( .A(\w3[8][80] ), .B(\w3[8][85] ), .Z(n8166) );
  XOR U5956 ( .A(key[1267]), .B(n7827), .Z(n4404) );
  XNOR U5957 ( .A(\w3[8][107] ), .B(n7856), .Z(n4405) );
  XNOR U5958 ( .A(n4404), .B(n4405), .Z(\w1[9][115] ) );
  XOR U5959 ( .A(key[1203]), .B(n8004), .Z(n4406) );
  XNOR U5960 ( .A(\w3[8][43] ), .B(n8033), .Z(n4407) );
  XNOR U5961 ( .A(n4406), .B(n4407), .Z(\w1[9][51] ) );
  XOR U5962 ( .A(key[1045]), .B(n7473), .Z(n4408) );
  XNOR U5963 ( .A(\w3[7][13] ), .B(n7510), .Z(n4409) );
  XNOR U5964 ( .A(n4408), .B(n4409), .Z(\w1[8][21] ) );
  XOR U5965 ( .A(key[1235]), .B(n8126), .Z(n4410) );
  XNOR U5966 ( .A(\w3[8][75] ), .B(n8161), .Z(n4411) );
  XNOR U5967 ( .A(n4410), .B(n4411), .Z(\w1[9][83] ) );
  XOR U5968 ( .A(n7852), .B(n8195), .Z(n4412) );
  XNOR U5969 ( .A(n7851), .B(key[1274]), .Z(n4413) );
  XNOR U5970 ( .A(n4412), .B(n4413), .Z(n4414) );
  XNOR U5971 ( .A(n4414), .B(\w3[8][98] ), .Z(\w1[9][122] ) );
  XOR U5972 ( .A(\w3[8][25] ), .B(n7905), .Z(n4415) );
  XNOR U5973 ( .A(\w3[8][17] ), .B(key[1176]), .Z(n4416) );
  XNOR U5974 ( .A(n4415), .B(n4416), .Z(n4417) );
  XNOR U5975 ( .A(n7906), .B(n4417), .Z(\w1[9][24] ) );
  XOR U5976 ( .A(n8148), .B(\w3[8][90] ), .Z(n4418) );
  XNOR U5977 ( .A(\w3[8][82] ), .B(key[1241]), .Z(n4419) );
  XNOR U5978 ( .A(n4418), .B(n4419), .Z(n4420) );
  XOR U5979 ( .A(n8149), .B(n4420), .Z(\w1[9][89] ) );
  XOR U5980 ( .A(n8026), .B(\w3[8][41] ), .Z(n4421) );
  XNOR U5981 ( .A(\w3[8][32] ), .B(key[1192]), .Z(n4422) );
  XNOR U5982 ( .A(n4421), .B(n4422), .Z(n4423) );
  XOR U5983 ( .A(n8055), .B(n4423), .Z(\w1[9][40] ) );
  XOR U5984 ( .A(key[1173]), .B(n7899), .Z(n4424) );
  XNOR U5985 ( .A(\w3[8][13] ), .B(n7936), .Z(n4425) );
  XNOR U5986 ( .A(n4424), .B(n4425), .Z(\w1[9][21] ) );
  XOR U5987 ( .A(key[1152]), .B(\w3[9][0] ), .Z(out[0]) );
  XOR U5988 ( .A(key[1252]), .B(\w3[9][100] ), .Z(out[100]) );
  XOR U5989 ( .A(key[1253]), .B(\w3[9][101] ), .Z(out[101]) );
  XOR U5990 ( .A(key[1254]), .B(\w3[9][102] ), .Z(out[102]) );
  XOR U5991 ( .A(key[1255]), .B(\w3[9][103] ), .Z(out[103]) );
  XOR U5992 ( .A(key[1256]), .B(\w3[9][104] ), .Z(out[104]) );
  XOR U5993 ( .A(key[1257]), .B(\w3[9][105] ), .Z(out[105]) );
  XOR U5994 ( .A(key[1258]), .B(\w3[9][106] ), .Z(out[106]) );
  XOR U5995 ( .A(key[1259]), .B(\w3[9][107] ), .Z(out[107]) );
  XOR U5996 ( .A(key[1260]), .B(\w3[9][108] ), .Z(out[108]) );
  XOR U5997 ( .A(key[1261]), .B(\w3[9][109] ), .Z(out[109]) );
  XOR U5998 ( .A(key[1162]), .B(\w3[9][10] ), .Z(out[10]) );
  XOR U5999 ( .A(key[1262]), .B(\w3[9][110] ), .Z(out[110]) );
  XOR U6000 ( .A(key[1263]), .B(\w3[9][111] ), .Z(out[111]) );
  XOR U6001 ( .A(key[1264]), .B(\w3[9][112] ), .Z(out[112]) );
  XOR U6002 ( .A(key[1265]), .B(\w3[9][113] ), .Z(out[113]) );
  XOR U6003 ( .A(key[1266]), .B(\w3[9][114] ), .Z(out[114]) );
  XOR U6004 ( .A(key[1267]), .B(\w3[9][115] ), .Z(out[115]) );
  XOR U6005 ( .A(key[1268]), .B(\w3[9][116] ), .Z(out[116]) );
  XOR U6006 ( .A(key[1269]), .B(\w3[9][117] ), .Z(out[117]) );
  XOR U6007 ( .A(key[1270]), .B(\w3[9][118] ), .Z(out[118]) );
  XOR U6008 ( .A(key[1271]), .B(\w3[9][119] ), .Z(out[119]) );
  XOR U6009 ( .A(key[1163]), .B(\w3[9][11] ), .Z(out[11]) );
  XOR U6010 ( .A(key[1272]), .B(\w3[9][120] ), .Z(out[120]) );
  XOR U6011 ( .A(key[1273]), .B(\w3[9][121] ), .Z(out[121]) );
  XOR U6012 ( .A(key[1274]), .B(\w3[9][122] ), .Z(out[122]) );
  XOR U6013 ( .A(key[1275]), .B(\w3[9][123] ), .Z(out[123]) );
  XOR U6014 ( .A(key[1276]), .B(\w3[9][124] ), .Z(out[124]) );
  XOR U6015 ( .A(key[1277]), .B(\w3[9][125] ), .Z(out[125]) );
  XOR U6016 ( .A(key[1278]), .B(\w3[9][126] ), .Z(out[126]) );
  XOR U6017 ( .A(key[1279]), .B(\w3[9][127] ), .Z(out[127]) );
  XOR U6018 ( .A(key[1164]), .B(\w3[9][12] ), .Z(out[12]) );
  XOR U6019 ( .A(key[1165]), .B(\w3[9][13] ), .Z(out[13]) );
  XOR U6020 ( .A(key[1166]), .B(\w3[9][14] ), .Z(out[14]) );
  XOR U6021 ( .A(key[1167]), .B(\w3[9][15] ), .Z(out[15]) );
  XOR U6022 ( .A(key[1168]), .B(\w3[9][16] ), .Z(out[16]) );
  XOR U6023 ( .A(key[1169]), .B(\w3[9][17] ), .Z(out[17]) );
  XOR U6024 ( .A(key[1170]), .B(\w3[9][18] ), .Z(out[18]) );
  XOR U6025 ( .A(key[1171]), .B(\w3[9][19] ), .Z(out[19]) );
  XOR U6026 ( .A(key[1153]), .B(\w3[9][1] ), .Z(out[1]) );
  XOR U6027 ( .A(key[1172]), .B(\w3[9][20] ), .Z(out[20]) );
  XOR U6028 ( .A(key[1173]), .B(\w3[9][21] ), .Z(out[21]) );
  XOR U6029 ( .A(key[1174]), .B(\w3[9][22] ), .Z(out[22]) );
  XOR U6030 ( .A(key[1175]), .B(\w3[9][23] ), .Z(out[23]) );
  XOR U6031 ( .A(key[1176]), .B(\w3[9][24] ), .Z(out[24]) );
  XOR U6032 ( .A(key[1177]), .B(\w3[9][25] ), .Z(out[25]) );
  XOR U6033 ( .A(key[1178]), .B(\w3[9][26] ), .Z(out[26]) );
  XOR U6034 ( .A(key[1179]), .B(\w3[9][27] ), .Z(out[27]) );
  XOR U6035 ( .A(key[1180]), .B(\w3[9][28] ), .Z(out[28]) );
  XOR U6036 ( .A(key[1181]), .B(\w3[9][29] ), .Z(out[29]) );
  XOR U6037 ( .A(key[1154]), .B(\w3[9][2] ), .Z(out[2]) );
  XOR U6038 ( .A(key[1182]), .B(\w3[9][30] ), .Z(out[30]) );
  XOR U6039 ( .A(key[1183]), .B(\w3[9][31] ), .Z(out[31]) );
  XOR U6040 ( .A(key[1184]), .B(\w3[9][32] ), .Z(out[32]) );
  XOR U6041 ( .A(key[1185]), .B(\w3[9][33] ), .Z(out[33]) );
  XOR U6042 ( .A(key[1186]), .B(\w3[9][34] ), .Z(out[34]) );
  XOR U6043 ( .A(key[1187]), .B(\w3[9][35] ), .Z(out[35]) );
  XOR U6044 ( .A(key[1188]), .B(\w3[9][36] ), .Z(out[36]) );
  XOR U6045 ( .A(key[1189]), .B(\w3[9][37] ), .Z(out[37]) );
  XOR U6046 ( .A(key[1190]), .B(\w3[9][38] ), .Z(out[38]) );
  XOR U6047 ( .A(key[1191]), .B(\w3[9][39] ), .Z(out[39]) );
  XOR U6048 ( .A(key[1155]), .B(\w3[9][3] ), .Z(out[3]) );
  XOR U6049 ( .A(key[1192]), .B(\w3[9][40] ), .Z(out[40]) );
  XOR U6050 ( .A(key[1193]), .B(\w3[9][41] ), .Z(out[41]) );
  XOR U6051 ( .A(key[1194]), .B(\w3[9][42] ), .Z(out[42]) );
  XOR U6052 ( .A(key[1195]), .B(\w3[9][43] ), .Z(out[43]) );
  XOR U6053 ( .A(key[1196]), .B(\w3[9][44] ), .Z(out[44]) );
  XOR U6054 ( .A(key[1197]), .B(\w3[9][45] ), .Z(out[45]) );
  XOR U6055 ( .A(key[1198]), .B(\w3[9][46] ), .Z(out[46]) );
  XOR U6056 ( .A(key[1199]), .B(\w3[9][47] ), .Z(out[47]) );
  XOR U6057 ( .A(key[1200]), .B(\w3[9][48] ), .Z(out[48]) );
  XOR U6058 ( .A(key[1201]), .B(\w3[9][49] ), .Z(out[49]) );
  XOR U6059 ( .A(key[1156]), .B(\w3[9][4] ), .Z(out[4]) );
  XOR U6060 ( .A(key[1202]), .B(\w3[9][50] ), .Z(out[50]) );
  XOR U6061 ( .A(key[1203]), .B(\w3[9][51] ), .Z(out[51]) );
  XOR U6062 ( .A(key[1204]), .B(\w3[9][52] ), .Z(out[52]) );
  XOR U6063 ( .A(key[1205]), .B(\w3[9][53] ), .Z(out[53]) );
  XOR U6064 ( .A(key[1206]), .B(\w3[9][54] ), .Z(out[54]) );
  XOR U6065 ( .A(key[1207]), .B(\w3[9][55] ), .Z(out[55]) );
  XOR U6066 ( .A(key[1208]), .B(\w3[9][56] ), .Z(out[56]) );
  XOR U6067 ( .A(key[1209]), .B(\w3[9][57] ), .Z(out[57]) );
  XOR U6068 ( .A(key[1210]), .B(\w3[9][58] ), .Z(out[58]) );
  XOR U6069 ( .A(key[1211]), .B(\w3[9][59] ), .Z(out[59]) );
  XOR U6070 ( .A(key[1157]), .B(\w3[9][5] ), .Z(out[5]) );
  XOR U6071 ( .A(key[1212]), .B(\w3[9][60] ), .Z(out[60]) );
  XOR U6072 ( .A(key[1213]), .B(\w3[9][61] ), .Z(out[61]) );
  XOR U6073 ( .A(key[1214]), .B(\w3[9][62] ), .Z(out[62]) );
  XOR U6074 ( .A(key[1215]), .B(\w3[9][63] ), .Z(out[63]) );
  XOR U6075 ( .A(key[1216]), .B(\w3[9][64] ), .Z(out[64]) );
  XOR U6076 ( .A(key[1217]), .B(\w3[9][65] ), .Z(out[65]) );
  XOR U6077 ( .A(key[1218]), .B(\w3[9][66] ), .Z(out[66]) );
  XOR U6078 ( .A(key[1219]), .B(\w3[9][67] ), .Z(out[67]) );
  XOR U6079 ( .A(key[1220]), .B(\w3[9][68] ), .Z(out[68]) );
  XOR U6080 ( .A(key[1221]), .B(\w3[9][69] ), .Z(out[69]) );
  XOR U6081 ( .A(key[1158]), .B(\w3[9][6] ), .Z(out[6]) );
  XOR U6082 ( .A(key[1222]), .B(\w3[9][70] ), .Z(out[70]) );
  XOR U6083 ( .A(key[1223]), .B(\w3[9][71] ), .Z(out[71]) );
  XOR U6084 ( .A(key[1224]), .B(\w3[9][72] ), .Z(out[72]) );
  XOR U6085 ( .A(key[1225]), .B(\w3[9][73] ), .Z(out[73]) );
  XOR U6086 ( .A(key[1226]), .B(\w3[9][74] ), .Z(out[74]) );
  XOR U6087 ( .A(key[1227]), .B(\w3[9][75] ), .Z(out[75]) );
  XOR U6088 ( .A(key[1228]), .B(\w3[9][76] ), .Z(out[76]) );
  XOR U6089 ( .A(key[1229]), .B(\w3[9][77] ), .Z(out[77]) );
  XOR U6090 ( .A(key[1230]), .B(\w3[9][78] ), .Z(out[78]) );
  XOR U6091 ( .A(key[1231]), .B(\w3[9][79] ), .Z(out[79]) );
  XOR U6092 ( .A(key[1159]), .B(\w3[9][7] ), .Z(out[7]) );
  XOR U6093 ( .A(key[1232]), .B(\w3[9][80] ), .Z(out[80]) );
  XOR U6094 ( .A(key[1233]), .B(\w3[9][81] ), .Z(out[81]) );
  XOR U6095 ( .A(key[1234]), .B(\w3[9][82] ), .Z(out[82]) );
  XOR U6096 ( .A(key[1235]), .B(\w3[9][83] ), .Z(out[83]) );
  XOR U6097 ( .A(key[1236]), .B(\w3[9][84] ), .Z(out[84]) );
  XOR U6098 ( .A(key[1237]), .B(\w3[9][85] ), .Z(out[85]) );
  XOR U6099 ( .A(key[1238]), .B(\w3[9][86] ), .Z(out[86]) );
  XOR U6100 ( .A(key[1239]), .B(\w3[9][87] ), .Z(out[87]) );
  XOR U6101 ( .A(key[1240]), .B(\w3[9][88] ), .Z(out[88]) );
  XOR U6102 ( .A(key[1241]), .B(\w3[9][89] ), .Z(out[89]) );
  XOR U6103 ( .A(key[1160]), .B(\w3[9][8] ), .Z(out[8]) );
  XOR U6104 ( .A(key[1242]), .B(\w3[9][90] ), .Z(out[90]) );
  XOR U6105 ( .A(key[1243]), .B(\w3[9][91] ), .Z(out[91]) );
  XOR U6106 ( .A(key[1244]), .B(\w3[9][92] ), .Z(out[92]) );
  XOR U6107 ( .A(key[1245]), .B(\w3[9][93] ), .Z(out[93]) );
  XOR U6108 ( .A(key[1246]), .B(\w3[9][94] ), .Z(out[94]) );
  XOR U6109 ( .A(key[1247]), .B(\w3[9][95] ), .Z(out[95]) );
  XOR U6110 ( .A(key[1248]), .B(\w3[9][96] ), .Z(out[96]) );
  XOR U6111 ( .A(key[1249]), .B(\w3[9][97] ), .Z(out[97]) );
  XOR U6112 ( .A(key[1250]), .B(\w3[9][98] ), .Z(out[98]) );
  XOR U6113 ( .A(key[1251]), .B(\w3[9][99] ), .Z(out[99]) );
  XOR U6114 ( .A(key[1161]), .B(\w3[9][9] ), .Z(out[9]) );
  XOR U6115 ( .A(key[0]), .B(msg[0]), .Z(\w1[0][0] ) );
  XOR U6116 ( .A(key[100]), .B(msg[100]), .Z(\w1[0][100] ) );
  XOR U6117 ( .A(key[101]), .B(msg[101]), .Z(\w1[0][101] ) );
  XOR U6118 ( .A(key[102]), .B(msg[102]), .Z(\w1[0][102] ) );
  XOR U6119 ( .A(key[103]), .B(msg[103]), .Z(\w1[0][103] ) );
  XOR U6120 ( .A(key[104]), .B(msg[104]), .Z(\w1[0][104] ) );
  XOR U6121 ( .A(key[105]), .B(msg[105]), .Z(\w1[0][105] ) );
  XOR U6122 ( .A(key[106]), .B(msg[106]), .Z(\w1[0][106] ) );
  XOR U6123 ( .A(key[107]), .B(msg[107]), .Z(\w1[0][107] ) );
  XOR U6124 ( .A(key[108]), .B(msg[108]), .Z(\w1[0][108] ) );
  XOR U6125 ( .A(key[109]), .B(msg[109]), .Z(\w1[0][109] ) );
  XOR U6126 ( .A(key[10]), .B(msg[10]), .Z(\w1[0][10] ) );
  XOR U6127 ( .A(key[110]), .B(msg[110]), .Z(\w1[0][110] ) );
  XOR U6128 ( .A(key[111]), .B(msg[111]), .Z(\w1[0][111] ) );
  XOR U6129 ( .A(key[112]), .B(msg[112]), .Z(\w1[0][112] ) );
  XOR U6130 ( .A(key[113]), .B(msg[113]), .Z(\w1[0][113] ) );
  XOR U6131 ( .A(key[114]), .B(msg[114]), .Z(\w1[0][114] ) );
  XOR U6132 ( .A(key[115]), .B(msg[115]), .Z(\w1[0][115] ) );
  XOR U6133 ( .A(key[116]), .B(msg[116]), .Z(\w1[0][116] ) );
  XOR U6134 ( .A(key[117]), .B(msg[117]), .Z(\w1[0][117] ) );
  XOR U6135 ( .A(key[118]), .B(msg[118]), .Z(\w1[0][118] ) );
  XOR U6136 ( .A(key[119]), .B(msg[119]), .Z(\w1[0][119] ) );
  XOR U6137 ( .A(key[11]), .B(msg[11]), .Z(\w1[0][11] ) );
  XOR U6138 ( .A(key[120]), .B(msg[120]), .Z(\w1[0][120] ) );
  XOR U6139 ( .A(key[121]), .B(msg[121]), .Z(\w1[0][121] ) );
  XOR U6140 ( .A(key[122]), .B(msg[122]), .Z(\w1[0][122] ) );
  XOR U6141 ( .A(key[123]), .B(msg[123]), .Z(\w1[0][123] ) );
  XOR U6142 ( .A(key[124]), .B(msg[124]), .Z(\w1[0][124] ) );
  XOR U6143 ( .A(key[125]), .B(msg[125]), .Z(\w1[0][125] ) );
  XOR U6144 ( .A(key[126]), .B(msg[126]), .Z(\w1[0][126] ) );
  XOR U6145 ( .A(key[127]), .B(msg[127]), .Z(\w1[0][127] ) );
  XOR U6146 ( .A(key[12]), .B(msg[12]), .Z(\w1[0][12] ) );
  XOR U6147 ( .A(key[13]), .B(msg[13]), .Z(\w1[0][13] ) );
  XOR U6148 ( .A(key[14]), .B(msg[14]), .Z(\w1[0][14] ) );
  XOR U6149 ( .A(key[15]), .B(msg[15]), .Z(\w1[0][15] ) );
  XOR U6150 ( .A(key[16]), .B(msg[16]), .Z(\w1[0][16] ) );
  XOR U6151 ( .A(key[17]), .B(msg[17]), .Z(\w1[0][17] ) );
  XOR U6152 ( .A(key[18]), .B(msg[18]), .Z(\w1[0][18] ) );
  XOR U6153 ( .A(key[19]), .B(msg[19]), .Z(\w1[0][19] ) );
  XOR U6154 ( .A(key[1]), .B(msg[1]), .Z(\w1[0][1] ) );
  XOR U6155 ( .A(key[20]), .B(msg[20]), .Z(\w1[0][20] ) );
  XOR U6156 ( .A(key[21]), .B(msg[21]), .Z(\w1[0][21] ) );
  XOR U6157 ( .A(key[22]), .B(msg[22]), .Z(\w1[0][22] ) );
  XOR U6158 ( .A(key[23]), .B(msg[23]), .Z(\w1[0][23] ) );
  XOR U6159 ( .A(key[24]), .B(msg[24]), .Z(\w1[0][24] ) );
  XOR U6160 ( .A(key[25]), .B(msg[25]), .Z(\w1[0][25] ) );
  XOR U6161 ( .A(key[26]), .B(msg[26]), .Z(\w1[0][26] ) );
  XOR U6162 ( .A(key[27]), .B(msg[27]), .Z(\w1[0][27] ) );
  XOR U6163 ( .A(key[28]), .B(msg[28]), .Z(\w1[0][28] ) );
  XOR U6164 ( .A(key[29]), .B(msg[29]), .Z(\w1[0][29] ) );
  XOR U6165 ( .A(key[2]), .B(msg[2]), .Z(\w1[0][2] ) );
  XOR U6166 ( .A(key[30]), .B(msg[30]), .Z(\w1[0][30] ) );
  XOR U6167 ( .A(key[31]), .B(msg[31]), .Z(\w1[0][31] ) );
  XOR U6168 ( .A(key[32]), .B(msg[32]), .Z(\w1[0][32] ) );
  XOR U6169 ( .A(key[33]), .B(msg[33]), .Z(\w1[0][33] ) );
  XOR U6170 ( .A(key[34]), .B(msg[34]), .Z(\w1[0][34] ) );
  XOR U6171 ( .A(key[35]), .B(msg[35]), .Z(\w1[0][35] ) );
  XOR U6172 ( .A(key[36]), .B(msg[36]), .Z(\w1[0][36] ) );
  XOR U6173 ( .A(key[37]), .B(msg[37]), .Z(\w1[0][37] ) );
  XOR U6174 ( .A(key[38]), .B(msg[38]), .Z(\w1[0][38] ) );
  XOR U6175 ( .A(key[39]), .B(msg[39]), .Z(\w1[0][39] ) );
  XOR U6176 ( .A(key[3]), .B(msg[3]), .Z(\w1[0][3] ) );
  XOR U6177 ( .A(key[40]), .B(msg[40]), .Z(\w1[0][40] ) );
  XOR U6178 ( .A(key[41]), .B(msg[41]), .Z(\w1[0][41] ) );
  XOR U6179 ( .A(key[42]), .B(msg[42]), .Z(\w1[0][42] ) );
  XOR U6180 ( .A(key[43]), .B(msg[43]), .Z(\w1[0][43] ) );
  XOR U6181 ( .A(key[44]), .B(msg[44]), .Z(\w1[0][44] ) );
  XOR U6182 ( .A(key[45]), .B(msg[45]), .Z(\w1[0][45] ) );
  XOR U6183 ( .A(key[46]), .B(msg[46]), .Z(\w1[0][46] ) );
  XOR U6184 ( .A(key[47]), .B(msg[47]), .Z(\w1[0][47] ) );
  XOR U6185 ( .A(key[48]), .B(msg[48]), .Z(\w1[0][48] ) );
  XOR U6186 ( .A(key[49]), .B(msg[49]), .Z(\w1[0][49] ) );
  XOR U6187 ( .A(key[4]), .B(msg[4]), .Z(\w1[0][4] ) );
  XOR U6188 ( .A(key[50]), .B(msg[50]), .Z(\w1[0][50] ) );
  XOR U6189 ( .A(key[51]), .B(msg[51]), .Z(\w1[0][51] ) );
  XOR U6190 ( .A(key[52]), .B(msg[52]), .Z(\w1[0][52] ) );
  XOR U6191 ( .A(key[53]), .B(msg[53]), .Z(\w1[0][53] ) );
  XOR U6192 ( .A(key[54]), .B(msg[54]), .Z(\w1[0][54] ) );
  XOR U6193 ( .A(key[55]), .B(msg[55]), .Z(\w1[0][55] ) );
  XOR U6194 ( .A(key[56]), .B(msg[56]), .Z(\w1[0][56] ) );
  XOR U6195 ( .A(key[57]), .B(msg[57]), .Z(\w1[0][57] ) );
  XOR U6196 ( .A(key[58]), .B(msg[58]), .Z(\w1[0][58] ) );
  XOR U6197 ( .A(key[59]), .B(msg[59]), .Z(\w1[0][59] ) );
  XOR U6198 ( .A(key[5]), .B(msg[5]), .Z(\w1[0][5] ) );
  XOR U6199 ( .A(key[60]), .B(msg[60]), .Z(\w1[0][60] ) );
  XOR U6200 ( .A(key[61]), .B(msg[61]), .Z(\w1[0][61] ) );
  XOR U6201 ( .A(key[62]), .B(msg[62]), .Z(\w1[0][62] ) );
  XOR U6202 ( .A(key[63]), .B(msg[63]), .Z(\w1[0][63] ) );
  XOR U6203 ( .A(key[64]), .B(msg[64]), .Z(\w1[0][64] ) );
  XOR U6204 ( .A(key[65]), .B(msg[65]), .Z(\w1[0][65] ) );
  XOR U6205 ( .A(key[66]), .B(msg[66]), .Z(\w1[0][66] ) );
  XOR U6206 ( .A(key[67]), .B(msg[67]), .Z(\w1[0][67] ) );
  XOR U6207 ( .A(key[68]), .B(msg[68]), .Z(\w1[0][68] ) );
  XOR U6208 ( .A(key[69]), .B(msg[69]), .Z(\w1[0][69] ) );
  XOR U6209 ( .A(key[6]), .B(msg[6]), .Z(\w1[0][6] ) );
  XOR U6210 ( .A(key[70]), .B(msg[70]), .Z(\w1[0][70] ) );
  XOR U6211 ( .A(key[71]), .B(msg[71]), .Z(\w1[0][71] ) );
  XOR U6212 ( .A(key[72]), .B(msg[72]), .Z(\w1[0][72] ) );
  XOR U6213 ( .A(key[73]), .B(msg[73]), .Z(\w1[0][73] ) );
  XOR U6214 ( .A(key[74]), .B(msg[74]), .Z(\w1[0][74] ) );
  XOR U6215 ( .A(key[75]), .B(msg[75]), .Z(\w1[0][75] ) );
  XOR U6216 ( .A(key[76]), .B(msg[76]), .Z(\w1[0][76] ) );
  XOR U6217 ( .A(key[77]), .B(msg[77]), .Z(\w1[0][77] ) );
  XOR U6218 ( .A(key[78]), .B(msg[78]), .Z(\w1[0][78] ) );
  XOR U6219 ( .A(key[79]), .B(msg[79]), .Z(\w1[0][79] ) );
  XOR U6220 ( .A(key[7]), .B(msg[7]), .Z(\w1[0][7] ) );
  XOR U6221 ( .A(key[80]), .B(msg[80]), .Z(\w1[0][80] ) );
  XOR U6222 ( .A(key[81]), .B(msg[81]), .Z(\w1[0][81] ) );
  XOR U6223 ( .A(key[82]), .B(msg[82]), .Z(\w1[0][82] ) );
  XOR U6224 ( .A(key[83]), .B(msg[83]), .Z(\w1[0][83] ) );
  XOR U6225 ( .A(key[84]), .B(msg[84]), .Z(\w1[0][84] ) );
  XOR U6226 ( .A(key[85]), .B(msg[85]), .Z(\w1[0][85] ) );
  XOR U6227 ( .A(key[86]), .B(msg[86]), .Z(\w1[0][86] ) );
  XOR U6228 ( .A(key[87]), .B(msg[87]), .Z(\w1[0][87] ) );
  XOR U6229 ( .A(key[88]), .B(msg[88]), .Z(\w1[0][88] ) );
  XOR U6230 ( .A(key[89]), .B(msg[89]), .Z(\w1[0][89] ) );
  XOR U6231 ( .A(key[8]), .B(msg[8]), .Z(\w1[0][8] ) );
  XOR U6232 ( .A(key[90]), .B(msg[90]), .Z(\w1[0][90] ) );
  XOR U6233 ( .A(key[91]), .B(msg[91]), .Z(\w1[0][91] ) );
  XOR U6234 ( .A(key[92]), .B(msg[92]), .Z(\w1[0][92] ) );
  XOR U6235 ( .A(key[93]), .B(msg[93]), .Z(\w1[0][93] ) );
  XOR U6236 ( .A(key[94]), .B(msg[94]), .Z(\w1[0][94] ) );
  XOR U6237 ( .A(key[95]), .B(msg[95]), .Z(\w1[0][95] ) );
  XOR U6238 ( .A(key[96]), .B(msg[96]), .Z(\w1[0][96] ) );
  XOR U6239 ( .A(key[97]), .B(msg[97]), .Z(\w1[0][97] ) );
  XOR U6240 ( .A(key[98]), .B(msg[98]), .Z(\w1[0][98] ) );
  XOR U6241 ( .A(key[99]), .B(msg[99]), .Z(\w1[0][99] ) );
  XOR U6242 ( .A(key[9]), .B(msg[9]), .Z(\w1[0][9] ) );
  XNOR U6243 ( .A(\w3[0][25] ), .B(\w3[0][1] ), .Z(n4844) );
  IV U6244 ( .A(\w3[0][16] ), .Z(n4555) );
  XOR U6245 ( .A(\w3[0][24] ), .B(n4555), .Z(n4796) );
  XNOR U6246 ( .A(\w3[0][8] ), .B(key[128]), .Z(n4426) );
  XNOR U6247 ( .A(n4796), .B(n4426), .Z(n4427) );
  XOR U6248 ( .A(n4844), .B(n4427), .Z(\w1[1][0] ) );
  XOR U6249 ( .A(\w3[0][96] ), .B(\w3[0][101] ), .Z(n4450) );
  XOR U6250 ( .A(\w3[0][116] ), .B(\w3[0][125] ), .Z(n4429) );
  IV U6251 ( .A(\w3[0][120] ), .Z(n4502) );
  XOR U6252 ( .A(n4502), .B(\w3[0][108] ), .Z(n4428) );
  XOR U6253 ( .A(n4429), .B(n4428), .Z(n4508) );
  XOR U6254 ( .A(n4508), .B(key[228]), .Z(n4430) );
  XOR U6255 ( .A(n4450), .B(n4430), .Z(n4431) );
  XNOR U6256 ( .A(\w3[0][124] ), .B(n4431), .Z(\w1[1][100] ) );
  XNOR U6257 ( .A(\w3[0][102] ), .B(\w3[0][126] ), .Z(n4459) );
  XNOR U6258 ( .A(n4459), .B(key[229]), .Z(n4433) );
  XNOR U6259 ( .A(\w3[0][109] ), .B(\w3[0][117] ), .Z(n4511) );
  XOR U6260 ( .A(\w3[0][125] ), .B(n4511), .Z(n4432) );
  XNOR U6261 ( .A(n4433), .B(n4432), .Z(\w1[1][101] ) );
  XOR U6262 ( .A(\w3[0][96] ), .B(\w3[0][103] ), .Z(n4460) );
  XOR U6263 ( .A(n4460), .B(key[230]), .Z(n4435) );
  XOR U6264 ( .A(n4502), .B(\w3[0][127] ), .Z(n4436) );
  XOR U6265 ( .A(\w3[0][110] ), .B(\w3[0][118] ), .Z(n4478) );
  XOR U6266 ( .A(n4436), .B(n4478), .Z(n4516) );
  XOR U6267 ( .A(\w3[0][126] ), .B(n4516), .Z(n4434) );
  XNOR U6268 ( .A(n4435), .B(n4434), .Z(\w1[1][102] ) );
  XNOR U6269 ( .A(\w3[0][111] ), .B(\w3[0][119] ), .Z(n4519) );
  XNOR U6270 ( .A(n4519), .B(key[231]), .Z(n4438) );
  XOR U6271 ( .A(\w3[0][96] ), .B(n4436), .Z(n4437) );
  XNOR U6272 ( .A(n4438), .B(n4437), .Z(\w1[1][103] ) );
  IV U6273 ( .A(\w3[0][97] ), .Z(n4498) );
  IV U6274 ( .A(\w3[0][112] ), .Z(n4494) );
  XOR U6275 ( .A(\w3[0][120] ), .B(n4494), .Z(n4825) );
  XOR U6276 ( .A(\w3[0][106] ), .B(\w3[0][113] ), .Z(n4440) );
  XNOR U6277 ( .A(\w3[0][97] ), .B(\w3[0][121] ), .Z(n4824) );
  XOR U6278 ( .A(n4824), .B(key[233]), .Z(n4439) );
  XNOR U6279 ( .A(n4440), .B(n4439), .Z(n4441) );
  XOR U6280 ( .A(\w3[0][98] ), .B(n4441), .Z(\w1[1][105] ) );
  XOR U6281 ( .A(\w3[0][107] ), .B(\w3[0][114] ), .Z(n4443) );
  XOR U6282 ( .A(\w3[0][98] ), .B(\w3[0][122] ), .Z(n4829) );
  XNOR U6283 ( .A(n4829), .B(key[234]), .Z(n4442) );
  XNOR U6284 ( .A(n4443), .B(n4442), .Z(n4444) );
  XOR U6285 ( .A(\w3[0][99] ), .B(n4444), .Z(\w1[1][106] ) );
  IV U6286 ( .A(\w3[0][123] ), .Z(n4837) );
  XOR U6287 ( .A(\w3[0][99] ), .B(n4837), .Z(n4833) );
  XOR U6288 ( .A(\w3[0][108] ), .B(n4833), .Z(n4445) );
  XOR U6289 ( .A(\w3[0][104] ), .B(n4445), .Z(n4471) );
  XNOR U6290 ( .A(n4471), .B(key[235]), .Z(n4447) );
  IV U6291 ( .A(\w3[0][100] ), .Z(n4507) );
  XOR U6292 ( .A(\w3[0][96] ), .B(n4507), .Z(n4838) );
  XOR U6293 ( .A(\w3[0][115] ), .B(n4838), .Z(n4446) );
  XNOR U6294 ( .A(n4447), .B(n4446), .Z(\w1[1][107] ) );
  XOR U6295 ( .A(\w3[0][100] ), .B(\w3[0][104] ), .Z(n4449) );
  XNOR U6296 ( .A(\w3[0][124] ), .B(\w3[0][109] ), .Z(n4448) );
  XOR U6297 ( .A(n4449), .B(n4448), .Z(n4474) );
  XNOR U6298 ( .A(n4474), .B(key[236]), .Z(n4452) );
  XNOR U6299 ( .A(\w3[0][116] ), .B(n4450), .Z(n4451) );
  XNOR U6300 ( .A(n4452), .B(n4451), .Z(\w1[1][108] ) );
  XNOR U6301 ( .A(\w3[0][125] ), .B(\w3[0][101] ), .Z(n4477) );
  XNOR U6302 ( .A(n4477), .B(key[237]), .Z(n4454) );
  XNOR U6303 ( .A(\w3[0][102] ), .B(\w3[0][110] ), .Z(n4453) );
  XNOR U6304 ( .A(n4454), .B(n4453), .Z(n4455) );
  XOR U6305 ( .A(\w3[0][117] ), .B(n4455), .Z(\w1[1][109] ) );
  XOR U6306 ( .A(\w3[0][11] ), .B(\w3[0][3] ), .Z(n4457) );
  XNOR U6307 ( .A(\w3[0][2] ), .B(\w3[0][26] ), .Z(n4542) );
  XOR U6308 ( .A(n4542), .B(key[138]), .Z(n4456) );
  XNOR U6309 ( .A(n4457), .B(n4456), .Z(n4458) );
  XOR U6310 ( .A(\w3[0][18] ), .B(n4458), .Z(\w1[1][10] ) );
  XOR U6311 ( .A(\w3[0][111] ), .B(\w3[0][104] ), .Z(n4485) );
  XOR U6312 ( .A(n4459), .B(n4485), .Z(n4481) );
  XNOR U6313 ( .A(n4481), .B(key[238]), .Z(n4462) );
  XNOR U6314 ( .A(\w3[0][118] ), .B(n4460), .Z(n4461) );
  XNOR U6315 ( .A(n4462), .B(n4461), .Z(\w1[1][110] ) );
  XOR U6316 ( .A(\w3[0][127] ), .B(\w3[0][103] ), .Z(n4484) );
  XOR U6317 ( .A(n4484), .B(key[239]), .Z(n4464) );
  XNOR U6318 ( .A(\w3[0][96] ), .B(\w3[0][104] ), .Z(n4490) );
  XOR U6319 ( .A(\w3[0][119] ), .B(n4490), .Z(n4463) );
  XNOR U6320 ( .A(n4464), .B(n4463), .Z(\w1[1][111] ) );
  XNOR U6321 ( .A(\w3[0][105] ), .B(\w3[0][113] ), .Z(n4828) );
  XNOR U6322 ( .A(n4828), .B(key[240]), .Z(n4466) );
  XNOR U6323 ( .A(n4502), .B(n4490), .Z(n4465) );
  XNOR U6324 ( .A(n4466), .B(n4465), .Z(\w1[1][112] ) );
  XNOR U6325 ( .A(\w3[0][106] ), .B(\w3[0][114] ), .Z(n4832) );
  XNOR U6326 ( .A(n4832), .B(key[241]), .Z(n4468) );
  XOR U6327 ( .A(\w3[0][105] ), .B(n4824), .Z(n4467) );
  XNOR U6328 ( .A(n4468), .B(n4467), .Z(\w1[1][113] ) );
  XNOR U6329 ( .A(\w3[0][107] ), .B(\w3[0][115] ), .Z(n4504) );
  XNOR U6330 ( .A(n4504), .B(key[242]), .Z(n4470) );
  XNOR U6331 ( .A(\w3[0][106] ), .B(n4829), .Z(n4469) );
  XNOR U6332 ( .A(n4470), .B(n4469), .Z(\w1[1][114] ) );
  XOR U6333 ( .A(\w3[0][116] ), .B(n4494), .Z(n4505) );
  XNOR U6334 ( .A(n4505), .B(key[243]), .Z(n4473) );
  XOR U6335 ( .A(\w3[0][107] ), .B(n4471), .Z(n4472) );
  XNOR U6336 ( .A(n4473), .B(n4472), .Z(\w1[1][115] ) );
  XOR U6337 ( .A(\w3[0][117] ), .B(n4494), .Z(n4506) );
  XNOR U6338 ( .A(n4506), .B(key[244]), .Z(n4476) );
  XOR U6339 ( .A(\w3[0][108] ), .B(n4474), .Z(n4475) );
  XNOR U6340 ( .A(n4476), .B(n4475), .Z(\w1[1][116] ) );
  XNOR U6341 ( .A(n4477), .B(key[245]), .Z(n4480) );
  XNOR U6342 ( .A(\w3[0][109] ), .B(n4478), .Z(n4479) );
  XNOR U6343 ( .A(n4480), .B(n4479), .Z(\w1[1][117] ) );
  XOR U6344 ( .A(\w3[0][119] ), .B(n4494), .Z(n4515) );
  XNOR U6345 ( .A(n4515), .B(key[246]), .Z(n4483) );
  XOR U6346 ( .A(\w3[0][110] ), .B(n4481), .Z(n4482) );
  XNOR U6347 ( .A(n4483), .B(n4482), .Z(\w1[1][118] ) );
  XOR U6348 ( .A(n4484), .B(key[247]), .Z(n4487) );
  XNOR U6349 ( .A(\w3[0][112] ), .B(n4485), .Z(n4486) );
  XNOR U6350 ( .A(n4487), .B(n4486), .Z(\w1[1][119] ) );
  XNOR U6351 ( .A(\w3[0][3] ), .B(\w3[0][27] ), .Z(n4576) );
  XNOR U6352 ( .A(n4539), .B(key[139]), .Z(n4489) );
  XNOR U6353 ( .A(\w3[0][0] ), .B(\w3[0][4] ), .Z(n4607) );
  XOR U6354 ( .A(\w3[0][19] ), .B(n4607), .Z(n4488) );
  XNOR U6355 ( .A(n4489), .B(n4488), .Z(\w1[1][11] ) );
  XNOR U6356 ( .A(n4490), .B(key[248]), .Z(n4492) );
  XNOR U6357 ( .A(\w3[0][121] ), .B(\w3[0][113] ), .Z(n4491) );
  XNOR U6358 ( .A(n4492), .B(n4491), .Z(n4493) );
  XNOR U6359 ( .A(n4494), .B(n4493), .Z(\w1[1][120] ) );
  XNOR U6360 ( .A(n4828), .B(key[249]), .Z(n4496) );
  XNOR U6361 ( .A(\w3[0][122] ), .B(\w3[0][114] ), .Z(n4495) );
  XNOR U6362 ( .A(n4496), .B(n4495), .Z(n4497) );
  XNOR U6363 ( .A(n4498), .B(n4497), .Z(\w1[1][121] ) );
  XNOR U6364 ( .A(n4832), .B(key[250]), .Z(n4500) );
  XNOR U6365 ( .A(\w3[0][115] ), .B(\w3[0][123] ), .Z(n4499) );
  XNOR U6366 ( .A(n4500), .B(n4499), .Z(n4501) );
  XOR U6367 ( .A(\w3[0][98] ), .B(n4501), .Z(\w1[1][122] ) );
  XOR U6368 ( .A(\w3[0][124] ), .B(n4502), .Z(n4503) );
  XOR U6369 ( .A(n4504), .B(n4503), .Z(n4836) );
  XNOR U6370 ( .A(n4506), .B(key[252]), .Z(n4510) );
  XNOR U6371 ( .A(n4508), .B(n4507), .Z(n4509) );
  XNOR U6372 ( .A(n4510), .B(n4509), .Z(\w1[1][124] ) );
  XOR U6373 ( .A(\w3[0][118] ), .B(key[253]), .Z(n4513) );
  XOR U6374 ( .A(n4511), .B(\w3[0][126] ), .Z(n4512) );
  XNOR U6375 ( .A(n4513), .B(n4512), .Z(n4514) );
  XOR U6376 ( .A(\w3[0][101] ), .B(n4514), .Z(\w1[1][125] ) );
  XNOR U6377 ( .A(n4515), .B(key[254]), .Z(n4518) );
  XOR U6378 ( .A(\w3[0][102] ), .B(n4516), .Z(n4517) );
  XNOR U6379 ( .A(n4518), .B(n4517), .Z(\w1[1][126] ) );
  XNOR U6380 ( .A(n4825), .B(key[255]), .Z(n4521) );
  XOR U6381 ( .A(\w3[0][103] ), .B(n4519), .Z(n4520) );
  XNOR U6382 ( .A(n4521), .B(n4520), .Z(\w1[1][127] ) );
  XOR U6383 ( .A(\w3[0][13] ), .B(\w3[0][28] ), .Z(n4523) );
  XNOR U6384 ( .A(\w3[0][8] ), .B(\w3[0][4] ), .Z(n4522) );
  XOR U6385 ( .A(n4523), .B(n4522), .Z(n4545) );
  XNOR U6386 ( .A(n4545), .B(key[140]), .Z(n4525) );
  XNOR U6387 ( .A(\w3[0][0] ), .B(\w3[0][5] ), .Z(n4641) );
  XOR U6388 ( .A(\w3[0][20] ), .B(n4641), .Z(n4524) );
  XNOR U6389 ( .A(n4525), .B(n4524), .Z(\w1[1][12] ) );
  IV U6390 ( .A(\w3[0][21] ), .Z(n4570) );
  XNOR U6391 ( .A(\w3[0][14] ), .B(n4570), .Z(n4527) );
  XNOR U6392 ( .A(\w3[0][5] ), .B(\w3[0][29] ), .Z(n4548) );
  XOR U6393 ( .A(n4548), .B(key[141]), .Z(n4526) );
  XNOR U6394 ( .A(n4527), .B(n4526), .Z(n4528) );
  XOR U6395 ( .A(\w3[0][6] ), .B(n4528), .Z(\w1[1][13] ) );
  IV U6396 ( .A(\w3[0][30] ), .Z(n4721) );
  XOR U6397 ( .A(\w3[0][6] ), .B(n4721), .Z(n4686) );
  XOR U6398 ( .A(\w3[0][8] ), .B(\w3[0][15] ), .Z(n4551) );
  XNOR U6399 ( .A(n4686), .B(n4551), .Z(n4549) );
  XOR U6400 ( .A(n4549), .B(key[142]), .Z(n4530) );
  XNOR U6401 ( .A(\w3[0][0] ), .B(\w3[0][7] ), .Z(n4722) );
  XOR U6402 ( .A(\w3[0][22] ), .B(n4722), .Z(n4529) );
  XNOR U6403 ( .A(n4530), .B(n4529), .Z(\w1[1][14] ) );
  XNOR U6404 ( .A(\w3[0][7] ), .B(\w3[0][31] ), .Z(n4550) );
  XNOR U6405 ( .A(n4550), .B(key[143]), .Z(n4532) );
  XOR U6406 ( .A(\w3[0][8] ), .B(\w3[0][0] ), .Z(n4554) );
  XNOR U6407 ( .A(\w3[0][23] ), .B(n4554), .Z(n4531) );
  XNOR U6408 ( .A(n4532), .B(n4531), .Z(\w1[1][15] ) );
  XNOR U6409 ( .A(\w3[0][17] ), .B(\w3[0][9] ), .Z(n4556) );
  XNOR U6410 ( .A(n4556), .B(key[144]), .Z(n4534) );
  XNOR U6411 ( .A(\w3[0][24] ), .B(n4554), .Z(n4533) );
  XNOR U6412 ( .A(n4534), .B(n4533), .Z(\w1[1][16] ) );
  XNOR U6413 ( .A(\w3[0][18] ), .B(\w3[0][10] ), .Z(n4575) );
  XNOR U6414 ( .A(n4575), .B(key[145]), .Z(n4536) );
  IV U6415 ( .A(\w3[0][9] ), .Z(n4793) );
  XNOR U6416 ( .A(n4844), .B(n4793), .Z(n4535) );
  XNOR U6417 ( .A(n4536), .B(n4535), .Z(\w1[1][17] ) );
  XNOR U6418 ( .A(\w3[0][11] ), .B(\w3[0][19] ), .Z(n4561) );
  XNOR U6419 ( .A(n4561), .B(key[146]), .Z(n4538) );
  XOR U6420 ( .A(n4542), .B(\w3[0][10] ), .Z(n4537) );
  XNOR U6421 ( .A(n4538), .B(n4537), .Z(\w1[1][18] ) );
  XOR U6422 ( .A(n4555), .B(\w3[0][20] ), .Z(n4562) );
  XNOR U6423 ( .A(n4562), .B(key[147]), .Z(n4541) );
  XOR U6424 ( .A(\w3[0][11] ), .B(n4539), .Z(n4540) );
  XNOR U6425 ( .A(n4541), .B(n4540), .Z(\w1[1][19] ) );
  XNOR U6426 ( .A(n4556), .B(key[129]), .Z(n4544) );
  XOR U6427 ( .A(\w3[0][25] ), .B(n4542), .Z(n4543) );
  XNOR U6428 ( .A(n4544), .B(n4543), .Z(\w1[1][1] ) );
  XOR U6429 ( .A(\w3[0][16] ), .B(n4570), .Z(n4567) );
  XNOR U6430 ( .A(n4567), .B(key[148]), .Z(n4547) );
  XOR U6431 ( .A(\w3[0][12] ), .B(n4545), .Z(n4546) );
  XNOR U6432 ( .A(n4547), .B(n4546), .Z(\w1[1][20] ) );
  IV U6433 ( .A(\w3[0][22] ), .Z(n4571) );
  XOR U6434 ( .A(\w3[0][14] ), .B(n4571), .Z(n4580) );
  XOR U6435 ( .A(n4555), .B(\w3[0][23] ), .Z(n4581) );
  XNOR U6436 ( .A(n4550), .B(key[151]), .Z(n4553) );
  XNOR U6437 ( .A(\w3[0][16] ), .B(n4551), .Z(n4552) );
  XNOR U6438 ( .A(n4553), .B(n4552), .Z(\w1[1][23] ) );
  XNOR U6439 ( .A(n4575), .B(key[154]), .Z(n4558) );
  XNOR U6440 ( .A(\w3[0][2] ), .B(\w3[0][19] ), .Z(n4557) );
  XNOR U6441 ( .A(n4558), .B(n4557), .Z(n4559) );
  XOR U6442 ( .A(\w3[0][27] ), .B(n4559), .Z(\w1[1][26] ) );
  IV U6443 ( .A(\w3[0][24] ), .Z(n4579) );
  XOR U6444 ( .A(n4579), .B(\w3[0][28] ), .Z(n4560) );
  XOR U6445 ( .A(n4561), .B(n4560), .Z(n4606) );
  XOR U6446 ( .A(n4606), .B(key[155]), .Z(n4564) );
  XOR U6447 ( .A(\w3[0][3] ), .B(n4562), .Z(n4563) );
  XNOR U6448 ( .A(n4564), .B(n4563), .Z(\w1[1][27] ) );
  XOR U6449 ( .A(\w3[0][20] ), .B(\w3[0][29] ), .Z(n4566) );
  XOR U6450 ( .A(n4579), .B(\w3[0][12] ), .Z(n4565) );
  XOR U6451 ( .A(n4566), .B(n4565), .Z(n4640) );
  XNOR U6452 ( .A(n4640), .B(key[156]), .Z(n4569) );
  XOR U6453 ( .A(\w3[0][4] ), .B(n4567), .Z(n4568) );
  XNOR U6454 ( .A(n4569), .B(n4568), .Z(\w1[1][28] ) );
  XOR U6455 ( .A(\w3[0][13] ), .B(n4570), .Z(n4685) );
  XNOR U6456 ( .A(n4685), .B(key[157]), .Z(n4573) );
  XNOR U6457 ( .A(n4571), .B(n4721), .Z(n4572) );
  XNOR U6458 ( .A(n4573), .B(n4572), .Z(n4574) );
  XOR U6459 ( .A(\w3[0][5] ), .B(n4574), .Z(\w1[1][29] ) );
  XNOR U6460 ( .A(n4575), .B(key[130]), .Z(n4578) );
  XOR U6461 ( .A(\w3[0][26] ), .B(n4576), .Z(n4577) );
  XNOR U6462 ( .A(n4578), .B(n4577), .Z(\w1[1][2] ) );
  XOR U6463 ( .A(n4579), .B(\w3[0][31] ), .Z(n4757) );
  XNOR U6464 ( .A(n4580), .B(n4757), .Z(n4720) );
  XNOR U6465 ( .A(\w3[0][15] ), .B(\w3[0][23] ), .Z(n4756) );
  XNOR U6466 ( .A(n4756), .B(key[159]), .Z(n4583) );
  XOR U6467 ( .A(n4796), .B(\w3[0][7] ), .Z(n4582) );
  XNOR U6468 ( .A(n4583), .B(n4582), .Z(\w1[1][31] ) );
  XOR U6469 ( .A(\w3[0][33] ), .B(\w3[0][57] ), .Z(n4585) );
  XNOR U6470 ( .A(\w3[0][40] ), .B(key[160]), .Z(n4584) );
  XNOR U6471 ( .A(n4585), .B(n4584), .Z(n4586) );
  IV U6472 ( .A(\w3[0][56] ), .Z(n4600) );
  XOR U6473 ( .A(\w3[0][48] ), .B(n4600), .Z(n4702) );
  XNOR U6474 ( .A(n4586), .B(n4702), .Z(\w1[1][32] ) );
  XNOR U6475 ( .A(\w3[0][34] ), .B(\w3[0][58] ), .Z(n4645) );
  XOR U6476 ( .A(\w3[0][57] ), .B(\w3[0][49] ), .Z(n4665) );
  XNOR U6477 ( .A(n4665), .B(key[161]), .Z(n4587) );
  XNOR U6478 ( .A(n4645), .B(n4587), .Z(n4588) );
  XNOR U6479 ( .A(\w3[0][41] ), .B(n4588), .Z(\w1[1][33] ) );
  XNOR U6480 ( .A(n4615), .B(key[162]), .Z(n4590) );
  XNOR U6481 ( .A(\w3[0][50] ), .B(\w3[0][42] ), .Z(n4675) );
  XOR U6482 ( .A(\w3[0][58] ), .B(n4675), .Z(n4589) );
  XNOR U6483 ( .A(n4590), .B(n4589), .Z(\w1[1][34] ) );
  XOR U6484 ( .A(\w3[0][36] ), .B(\w3[0][32] ), .Z(n4617) );
  XOR U6485 ( .A(n4617), .B(key[163]), .Z(n4593) );
  IV U6486 ( .A(\w3[0][51] ), .Z(n4674) );
  XOR U6487 ( .A(\w3[0][43] ), .B(n4674), .Z(n4644) );
  XNOR U6488 ( .A(n4600), .B(n4644), .Z(n4591) );
  XNOR U6489 ( .A(\w3[0][60] ), .B(n4591), .Z(n4681) );
  XNOR U6490 ( .A(\w3[0][59] ), .B(n4681), .Z(n4592) );
  XNOR U6491 ( .A(n4593), .B(n4592), .Z(\w1[1][35] ) );
  XOR U6492 ( .A(\w3[0][32] ), .B(\w3[0][37] ), .Z(n4623) );
  XOR U6493 ( .A(\w3[0][52] ), .B(\w3[0][61] ), .Z(n4595) );
  XOR U6494 ( .A(n4600), .B(\w3[0][44] ), .Z(n4594) );
  XOR U6495 ( .A(n4595), .B(n4594), .Z(n4690) );
  XOR U6496 ( .A(n4690), .B(key[164]), .Z(n4596) );
  XOR U6497 ( .A(n4623), .B(n4596), .Z(n4597) );
  XNOR U6498 ( .A(\w3[0][60] ), .B(n4597), .Z(\w1[1][36] ) );
  XNOR U6499 ( .A(\w3[0][38] ), .B(\w3[0][62] ), .Z(n4629) );
  XNOR U6500 ( .A(n4629), .B(key[165]), .Z(n4599) );
  IV U6501 ( .A(\w3[0][45] ), .Z(n4654) );
  XOR U6502 ( .A(\w3[0][53] ), .B(n4654), .Z(n4693) );
  XOR U6503 ( .A(\w3[0][61] ), .B(n4693), .Z(n4598) );
  XNOR U6504 ( .A(n4599), .B(n4598), .Z(\w1[1][37] ) );
  XOR U6505 ( .A(\w3[0][32] ), .B(\w3[0][39] ), .Z(n4630) );
  XOR U6506 ( .A(n4630), .B(key[166]), .Z(n4602) );
  XOR U6507 ( .A(n4600), .B(\w3[0][63] ), .Z(n4603) );
  XOR U6508 ( .A(\w3[0][46] ), .B(\w3[0][54] ), .Z(n4653) );
  XOR U6509 ( .A(n4603), .B(n4653), .Z(n4698) );
  XOR U6510 ( .A(\w3[0][62] ), .B(n4698), .Z(n4601) );
  XNOR U6511 ( .A(n4602), .B(n4601), .Z(\w1[1][38] ) );
  XNOR U6512 ( .A(\w3[0][55] ), .B(\w3[0][47] ), .Z(n4701) );
  XNOR U6513 ( .A(n4701), .B(key[167]), .Z(n4605) );
  XOR U6514 ( .A(\w3[0][32] ), .B(n4603), .Z(n4604) );
  XNOR U6515 ( .A(n4605), .B(n4604), .Z(\w1[1][39] ) );
  XOR U6516 ( .A(n4606), .B(key[131]), .Z(n4609) );
  XOR U6517 ( .A(n4607), .B(\w3[0][27] ), .Z(n4608) );
  XNOR U6518 ( .A(n4609), .B(n4608), .Z(\w1[1][3] ) );
  XNOR U6519 ( .A(\w3[0][33] ), .B(\w3[0][41] ), .Z(n4669) );
  XNOR U6520 ( .A(n4669), .B(key[168]), .Z(n4611) );
  XOR U6521 ( .A(n4702), .B(\w3[0][32] ), .Z(n4610) );
  XNOR U6522 ( .A(n4611), .B(n4610), .Z(\w1[1][40] ) );
  IV U6523 ( .A(\w3[0][34] ), .Z(n4679) );
  XOR U6524 ( .A(\w3[0][43] ), .B(key[170]), .Z(n4613) );
  IV U6525 ( .A(\w3[0][35] ), .Z(n4682) );
  XOR U6526 ( .A(\w3[0][50] ), .B(n4682), .Z(n4612) );
  XNOR U6527 ( .A(n4613), .B(n4612), .Z(n4614) );
  XNOR U6528 ( .A(n4614), .B(n4645), .Z(\w1[1][42] ) );
  IV U6529 ( .A(\w3[0][40] ), .Z(n4620) );
  XNOR U6530 ( .A(n4620), .B(n4615), .Z(n4616) );
  XOR U6531 ( .A(\w3[0][44] ), .B(n4616), .Z(n4648) );
  XNOR U6532 ( .A(n4648), .B(key[171]), .Z(n4619) );
  XNOR U6533 ( .A(\w3[0][51] ), .B(n4617), .Z(n4618) );
  XNOR U6534 ( .A(n4619), .B(n4618), .Z(\w1[1][43] ) );
  XOR U6535 ( .A(\w3[0][36] ), .B(\w3[0][45] ), .Z(n4622) );
  XOR U6536 ( .A(n4620), .B(\w3[0][60] ), .Z(n4621) );
  XOR U6537 ( .A(n4622), .B(n4621), .Z(n4649) );
  XNOR U6538 ( .A(n4649), .B(key[172]), .Z(n4625) );
  XNOR U6539 ( .A(\w3[0][52] ), .B(n4623), .Z(n4624) );
  XNOR U6540 ( .A(n4625), .B(n4624), .Z(\w1[1][44] ) );
  XNOR U6541 ( .A(\w3[0][61] ), .B(\w3[0][37] ), .Z(n4652) );
  XNOR U6542 ( .A(n4652), .B(key[173]), .Z(n4627) );
  XNOR U6543 ( .A(\w3[0][38] ), .B(\w3[0][46] ), .Z(n4626) );
  XNOR U6544 ( .A(n4627), .B(n4626), .Z(n4628) );
  XOR U6545 ( .A(\w3[0][53] ), .B(n4628), .Z(\w1[1][45] ) );
  XOR U6546 ( .A(\w3[0][40] ), .B(\w3[0][47] ), .Z(n4661) );
  XOR U6547 ( .A(n4629), .B(n4661), .Z(n4657) );
  XNOR U6548 ( .A(n4657), .B(key[174]), .Z(n4632) );
  XNOR U6549 ( .A(\w3[0][54] ), .B(n4630), .Z(n4631) );
  XNOR U6550 ( .A(n4632), .B(n4631), .Z(\w1[1][46] ) );
  XOR U6551 ( .A(\w3[0][63] ), .B(\w3[0][39] ), .Z(n4660) );
  XOR U6552 ( .A(n4660), .B(key[175]), .Z(n4634) );
  XNOR U6553 ( .A(\w3[0][40] ), .B(\w3[0][32] ), .Z(n4664) );
  XOR U6554 ( .A(\w3[0][55] ), .B(n4664), .Z(n4633) );
  XNOR U6555 ( .A(n4634), .B(n4633), .Z(\w1[1][47] ) );
  XNOR U6556 ( .A(n4664), .B(key[176]), .Z(n4636) );
  IV U6557 ( .A(\w3[0][49] ), .Z(n4670) );
  XOR U6558 ( .A(\w3[0][56] ), .B(n4670), .Z(n4635) );
  XNOR U6559 ( .A(n4636), .B(n4635), .Z(n4637) );
  XOR U6560 ( .A(\w3[0][41] ), .B(n4637), .Z(\w1[1][48] ) );
  XNOR U6561 ( .A(n4669), .B(key[177]), .Z(n4639) );
  XOR U6562 ( .A(\w3[0][57] ), .B(n4675), .Z(n4638) );
  XNOR U6563 ( .A(n4639), .B(n4638), .Z(\w1[1][49] ) );
  XNOR U6564 ( .A(n4640), .B(key[132]), .Z(n4643) );
  XOR U6565 ( .A(n4641), .B(\w3[0][28] ), .Z(n4642) );
  XNOR U6566 ( .A(n4643), .B(n4642), .Z(\w1[1][4] ) );
  XNOR U6567 ( .A(n4644), .B(key[178]), .Z(n4647) );
  XOR U6568 ( .A(n4645), .B(\w3[0][42] ), .Z(n4646) );
  XNOR U6569 ( .A(n4647), .B(n4646), .Z(\w1[1][50] ) );
  IV U6570 ( .A(\w3[0][48] ), .Z(n4666) );
  XOR U6571 ( .A(n4666), .B(\w3[0][52] ), .Z(n4680) );
  XNOR U6572 ( .A(n4689), .B(key[180]), .Z(n4651) );
  XOR U6573 ( .A(\w3[0][44] ), .B(n4649), .Z(n4650) );
  XNOR U6574 ( .A(n4651), .B(n4650), .Z(\w1[1][52] ) );
  XNOR U6575 ( .A(n4652), .B(key[181]), .Z(n4656) );
  XOR U6576 ( .A(n4654), .B(n4653), .Z(n4655) );
  XNOR U6577 ( .A(n4656), .B(n4655), .Z(\w1[1][53] ) );
  XOR U6578 ( .A(n4666), .B(\w3[0][55] ), .Z(n4697) );
  XNOR U6579 ( .A(n4697), .B(key[182]), .Z(n4659) );
  XOR U6580 ( .A(\w3[0][46] ), .B(n4657), .Z(n4658) );
  XNOR U6581 ( .A(n4659), .B(n4658), .Z(\w1[1][54] ) );
  XOR U6582 ( .A(n4660), .B(key[183]), .Z(n4663) );
  XNOR U6583 ( .A(\w3[0][48] ), .B(n4661), .Z(n4662) );
  XNOR U6584 ( .A(n4663), .B(n4662), .Z(\w1[1][55] ) );
  XNOR U6585 ( .A(n4664), .B(key[184]), .Z(n4668) );
  XOR U6586 ( .A(n4666), .B(n4665), .Z(n4667) );
  XNOR U6587 ( .A(n4668), .B(n4667), .Z(\w1[1][56] ) );
  XNOR U6588 ( .A(n4669), .B(key[185]), .Z(n4672) );
  XOR U6589 ( .A(n4670), .B(\w3[0][50] ), .Z(n4671) );
  XNOR U6590 ( .A(n4672), .B(n4671), .Z(n4673) );
  XOR U6591 ( .A(\w3[0][58] ), .B(n4673), .Z(\w1[1][57] ) );
  XNOR U6592 ( .A(n4674), .B(key[186]), .Z(n4677) );
  XOR U6593 ( .A(n4675), .B(\w3[0][59] ), .Z(n4676) );
  XNOR U6594 ( .A(n4677), .B(n4676), .Z(n4678) );
  XNOR U6595 ( .A(n4679), .B(n4678), .Z(\w1[1][58] ) );
  XNOR U6596 ( .A(n4680), .B(key[187]), .Z(n4684) );
  XOR U6597 ( .A(n4682), .B(n4681), .Z(n4683) );
  XNOR U6598 ( .A(n4684), .B(n4683), .Z(\w1[1][59] ) );
  XNOR U6599 ( .A(n4685), .B(key[133]), .Z(n4688) );
  XOR U6600 ( .A(\w3[0][29] ), .B(n4686), .Z(n4687) );
  XNOR U6601 ( .A(n4688), .B(n4687), .Z(\w1[1][5] ) );
  XNOR U6602 ( .A(n4689), .B(key[188]), .Z(n4692) );
  XOR U6603 ( .A(\w3[0][36] ), .B(n4690), .Z(n4691) );
  XNOR U6604 ( .A(n4692), .B(n4691), .Z(\w1[1][60] ) );
  XOR U6605 ( .A(\w3[0][54] ), .B(key[189]), .Z(n4695) );
  XOR U6606 ( .A(n4693), .B(\w3[0][62] ), .Z(n4694) );
  XNOR U6607 ( .A(n4695), .B(n4694), .Z(n4696) );
  XOR U6608 ( .A(\w3[0][37] ), .B(n4696), .Z(\w1[1][61] ) );
  XNOR U6609 ( .A(n4697), .B(key[190]), .Z(n4700) );
  XOR U6610 ( .A(\w3[0][38] ), .B(n4698), .Z(n4699) );
  XNOR U6611 ( .A(n4700), .B(n4699), .Z(\w1[1][62] ) );
  XNOR U6612 ( .A(n4701), .B(key[191]), .Z(n4704) );
  XOR U6613 ( .A(n4702), .B(\w3[0][39] ), .Z(n4703) );
  XNOR U6614 ( .A(n4704), .B(n4703), .Z(\w1[1][63] ) );
  XOR U6615 ( .A(\w3[0][65] ), .B(\w3[0][89] ), .Z(n4762) );
  XOR U6616 ( .A(n4762), .B(key[192]), .Z(n4706) );
  XNOR U6617 ( .A(\w3[0][80] ), .B(\w3[0][88] ), .Z(n4821) );
  XOR U6618 ( .A(n4821), .B(\w3[0][72] ), .Z(n4705) );
  XNOR U6619 ( .A(n4706), .B(n4705), .Z(\w1[1][64] ) );
  XNOR U6620 ( .A(\w3[0][66] ), .B(\w3[0][90] ), .Z(n4766) );
  XOR U6621 ( .A(\w3[0][89] ), .B(\w3[0][81] ), .Z(n4784) );
  XNOR U6622 ( .A(n4784), .B(key[193]), .Z(n4707) );
  XNOR U6623 ( .A(n4766), .B(n4707), .Z(n4708) );
  XNOR U6624 ( .A(\w3[0][73] ), .B(n4708), .Z(\w1[1][65] ) );
  XNOR U6625 ( .A(n4736), .B(key[194]), .Z(n4710) );
  XNOR U6626 ( .A(\w3[0][82] ), .B(\w3[0][74] ), .Z(n4799) );
  XOR U6627 ( .A(\w3[0][90] ), .B(n4799), .Z(n4709) );
  XNOR U6628 ( .A(n4710), .B(n4709), .Z(\w1[1][66] ) );
  XOR U6629 ( .A(\w3[0][68] ), .B(\w3[0][64] ), .Z(n4738) );
  XOR U6630 ( .A(n4738), .B(key[195]), .Z(n4713) );
  IV U6631 ( .A(\w3[0][83] ), .Z(n4798) );
  XOR U6632 ( .A(\w3[0][75] ), .B(n4798), .Z(n4765) );
  XOR U6633 ( .A(\w3[0][88] ), .B(n4765), .Z(n4711) );
  XNOR U6634 ( .A(\w3[0][92] ), .B(n4711), .Z(n4804) );
  XNOR U6635 ( .A(\w3[0][91] ), .B(n4804), .Z(n4712) );
  XNOR U6636 ( .A(n4713), .B(n4712), .Z(\w1[1][67] ) );
  XOR U6637 ( .A(\w3[0][64] ), .B(\w3[0][69] ), .Z(n4744) );
  XOR U6638 ( .A(\w3[0][84] ), .B(\w3[0][93] ), .Z(n4715) );
  XNOR U6639 ( .A(\w3[0][88] ), .B(\w3[0][76] ), .Z(n4714) );
  XOR U6640 ( .A(n4715), .B(n4714), .Z(n4809) );
  XOR U6641 ( .A(n4809), .B(key[196]), .Z(n4716) );
  XOR U6642 ( .A(n4744), .B(n4716), .Z(n4717) );
  XNOR U6643 ( .A(\w3[0][92] ), .B(n4717), .Z(\w1[1][68] ) );
  XNOR U6644 ( .A(\w3[0][70] ), .B(\w3[0][94] ), .Z(n4750) );
  XNOR U6645 ( .A(n4750), .B(key[197]), .Z(n4719) );
  IV U6646 ( .A(\w3[0][77] ), .Z(n4773) );
  XOR U6647 ( .A(\w3[0][85] ), .B(n4773), .Z(n4812) );
  XOR U6648 ( .A(\w3[0][93] ), .B(n4812), .Z(n4718) );
  XNOR U6649 ( .A(n4719), .B(n4718), .Z(\w1[1][69] ) );
  XNOR U6650 ( .A(n4720), .B(key[134]), .Z(n4724) );
  XNOR U6651 ( .A(n4722), .B(n4721), .Z(n4723) );
  XNOR U6652 ( .A(n4724), .B(n4723), .Z(\w1[1][6] ) );
  XOR U6653 ( .A(\w3[0][64] ), .B(\w3[0][71] ), .Z(n4751) );
  XOR U6654 ( .A(n4751), .B(key[198]), .Z(n4726) );
  XNOR U6655 ( .A(\w3[0][88] ), .B(\w3[0][95] ), .Z(n4727) );
  XOR U6656 ( .A(\w3[0][78] ), .B(\w3[0][86] ), .Z(n4772) );
  XOR U6657 ( .A(n4727), .B(n4772), .Z(n4817) );
  XOR U6658 ( .A(\w3[0][94] ), .B(n4817), .Z(n4725) );
  XNOR U6659 ( .A(n4726), .B(n4725), .Z(\w1[1][70] ) );
  XNOR U6660 ( .A(\w3[0][79] ), .B(\w3[0][87] ), .Z(n4820) );
  XNOR U6661 ( .A(n4820), .B(key[199]), .Z(n4729) );
  XOR U6662 ( .A(\w3[0][64] ), .B(n4727), .Z(n4728) );
  XNOR U6663 ( .A(n4729), .B(n4728), .Z(\w1[1][71] ) );
  IV U6664 ( .A(\w3[0][65] ), .Z(n4789) );
  XOR U6665 ( .A(\w3[0][74] ), .B(key[201]), .Z(n4731) );
  XNOR U6666 ( .A(n4784), .B(\w3[0][66] ), .Z(n4730) );
  XNOR U6667 ( .A(n4731), .B(n4730), .Z(n4732) );
  XNOR U6668 ( .A(n4789), .B(n4732), .Z(\w1[1][73] ) );
  XOR U6669 ( .A(\w3[0][75] ), .B(key[202]), .Z(n4734) );
  IV U6670 ( .A(\w3[0][67] ), .Z(n4805) );
  XOR U6671 ( .A(\w3[0][82] ), .B(n4805), .Z(n4733) );
  XNOR U6672 ( .A(n4734), .B(n4733), .Z(n4735) );
  XNOR U6673 ( .A(n4735), .B(n4766), .Z(\w1[1][74] ) );
  IV U6674 ( .A(\w3[0][72] ), .Z(n4741) );
  XNOR U6675 ( .A(n4741), .B(n4736), .Z(n4737) );
  XOR U6676 ( .A(\w3[0][76] ), .B(n4737), .Z(n4767) );
  XNOR U6677 ( .A(n4767), .B(key[203]), .Z(n4740) );
  XNOR U6678 ( .A(\w3[0][83] ), .B(n4738), .Z(n4739) );
  XNOR U6679 ( .A(n4740), .B(n4739), .Z(\w1[1][75] ) );
  XOR U6680 ( .A(\w3[0][68] ), .B(\w3[0][77] ), .Z(n4743) );
  XOR U6681 ( .A(n4741), .B(\w3[0][92] ), .Z(n4742) );
  XOR U6682 ( .A(n4743), .B(n4742), .Z(n4768) );
  XNOR U6683 ( .A(n4768), .B(key[204]), .Z(n4746) );
  XNOR U6684 ( .A(\w3[0][84] ), .B(n4744), .Z(n4745) );
  XNOR U6685 ( .A(n4746), .B(n4745), .Z(\w1[1][76] ) );
  XNOR U6686 ( .A(\w3[0][93] ), .B(\w3[0][69] ), .Z(n4771) );
  XNOR U6687 ( .A(n4771), .B(key[205]), .Z(n4748) );
  XNOR U6688 ( .A(\w3[0][70] ), .B(\w3[0][78] ), .Z(n4747) );
  XNOR U6689 ( .A(n4748), .B(n4747), .Z(n4749) );
  XOR U6690 ( .A(\w3[0][85] ), .B(n4749), .Z(\w1[1][77] ) );
  XOR U6691 ( .A(\w3[0][72] ), .B(\w3[0][79] ), .Z(n4780) );
  XOR U6692 ( .A(n4750), .B(n4780), .Z(n4776) );
  XNOR U6693 ( .A(n4776), .B(key[206]), .Z(n4753) );
  XNOR U6694 ( .A(\w3[0][86] ), .B(n4751), .Z(n4752) );
  XNOR U6695 ( .A(n4753), .B(n4752), .Z(\w1[1][78] ) );
  XOR U6696 ( .A(\w3[0][95] ), .B(\w3[0][71] ), .Z(n4779) );
  XOR U6697 ( .A(n4779), .B(key[207]), .Z(n4755) );
  XNOR U6698 ( .A(\w3[0][72] ), .B(\w3[0][64] ), .Z(n4783) );
  XOR U6699 ( .A(\w3[0][87] ), .B(n4783), .Z(n4754) );
  XNOR U6700 ( .A(n4755), .B(n4754), .Z(\w1[1][79] ) );
  XNOR U6701 ( .A(n4756), .B(key[135]), .Z(n4759) );
  XOR U6702 ( .A(\w3[0][0] ), .B(n4757), .Z(n4758) );
  XNOR U6703 ( .A(n4759), .B(n4758), .Z(\w1[1][7] ) );
  XNOR U6704 ( .A(\w3[0][73] ), .B(\w3[0][81] ), .Z(n4788) );
  XNOR U6705 ( .A(n4788), .B(key[208]), .Z(n4761) );
  XOR U6706 ( .A(\w3[0][88] ), .B(n4783), .Z(n4760) );
  XNOR U6707 ( .A(n4761), .B(n4760), .Z(\w1[1][80] ) );
  XNOR U6708 ( .A(n4799), .B(key[209]), .Z(n4764) );
  XNOR U6709 ( .A(n4762), .B(\w3[0][73] ), .Z(n4763) );
  XNOR U6710 ( .A(n4764), .B(n4763), .Z(\w1[1][81] ) );
  IV U6711 ( .A(\w3[0][80] ), .Z(n4785) );
  XOR U6712 ( .A(n4785), .B(\w3[0][84] ), .Z(n4803) );
  XNOR U6713 ( .A(n4808), .B(key[212]), .Z(n4770) );
  XOR U6714 ( .A(\w3[0][76] ), .B(n4768), .Z(n4769) );
  XNOR U6715 ( .A(n4770), .B(n4769), .Z(\w1[1][84] ) );
  XNOR U6716 ( .A(n4771), .B(key[213]), .Z(n4775) );
  XOR U6717 ( .A(n4773), .B(n4772), .Z(n4774) );
  XNOR U6718 ( .A(n4775), .B(n4774), .Z(\w1[1][85] ) );
  XOR U6719 ( .A(n4785), .B(\w3[0][87] ), .Z(n4816) );
  XNOR U6720 ( .A(n4816), .B(key[214]), .Z(n4778) );
  XOR U6721 ( .A(\w3[0][78] ), .B(n4776), .Z(n4777) );
  XNOR U6722 ( .A(n4778), .B(n4777), .Z(\w1[1][86] ) );
  XOR U6723 ( .A(n4779), .B(key[215]), .Z(n4782) );
  XNOR U6724 ( .A(\w3[0][80] ), .B(n4780), .Z(n4781) );
  XNOR U6725 ( .A(n4782), .B(n4781), .Z(\w1[1][87] ) );
  XNOR U6726 ( .A(n4783), .B(key[216]), .Z(n4787) );
  XOR U6727 ( .A(n4785), .B(n4784), .Z(n4786) );
  XNOR U6728 ( .A(n4787), .B(n4786), .Z(\w1[1][88] ) );
  XNOR U6729 ( .A(n4788), .B(key[217]), .Z(n4791) );
  XOR U6730 ( .A(n4789), .B(\w3[0][82] ), .Z(n4790) );
  XNOR U6731 ( .A(n4791), .B(n4790), .Z(n4792) );
  XOR U6732 ( .A(\w3[0][90] ), .B(n4792), .Z(\w1[1][89] ) );
  XNOR U6733 ( .A(n4793), .B(key[136]), .Z(n4795) );
  XNOR U6734 ( .A(\w3[0][1] ), .B(\w3[0][0] ), .Z(n4794) );
  XNOR U6735 ( .A(n4795), .B(n4794), .Z(n4797) );
  XNOR U6736 ( .A(n4797), .B(n4796), .Z(\w1[1][8] ) );
  XNOR U6737 ( .A(n4798), .B(key[218]), .Z(n4801) );
  XOR U6738 ( .A(n4799), .B(\w3[0][91] ), .Z(n4800) );
  XNOR U6739 ( .A(n4801), .B(n4800), .Z(n4802) );
  XOR U6740 ( .A(\w3[0][66] ), .B(n4802), .Z(\w1[1][90] ) );
  XNOR U6741 ( .A(n4803), .B(key[219]), .Z(n4807) );
  XOR U6742 ( .A(n4805), .B(n4804), .Z(n4806) );
  XNOR U6743 ( .A(n4807), .B(n4806), .Z(\w1[1][91] ) );
  XNOR U6744 ( .A(n4808), .B(key[220]), .Z(n4811) );
  XOR U6745 ( .A(\w3[0][68] ), .B(n4809), .Z(n4810) );
  XNOR U6746 ( .A(n4811), .B(n4810), .Z(\w1[1][92] ) );
  XOR U6747 ( .A(\w3[0][86] ), .B(key[221]), .Z(n4814) );
  XOR U6748 ( .A(n4812), .B(\w3[0][94] ), .Z(n4813) );
  XNOR U6749 ( .A(n4814), .B(n4813), .Z(n4815) );
  XOR U6750 ( .A(\w3[0][69] ), .B(n4815), .Z(\w1[1][93] ) );
  XNOR U6751 ( .A(n4816), .B(key[222]), .Z(n4819) );
  XOR U6752 ( .A(\w3[0][70] ), .B(n4817), .Z(n4818) );
  XNOR U6753 ( .A(n4819), .B(n4818), .Z(\w1[1][94] ) );
  XNOR U6754 ( .A(n4820), .B(key[223]), .Z(n4823) );
  XOR U6755 ( .A(n4821), .B(\w3[0][71] ), .Z(n4822) );
  XNOR U6756 ( .A(n4823), .B(n4822), .Z(\w1[1][95] ) );
  XOR U6757 ( .A(\w3[0][104] ), .B(key[224]), .Z(n4827) );
  XNOR U6758 ( .A(n4825), .B(n4824), .Z(n4826) );
  XNOR U6759 ( .A(n4827), .B(n4826), .Z(\w1[1][96] ) );
  XNOR U6760 ( .A(n4828), .B(key[225]), .Z(n4831) );
  XNOR U6761 ( .A(\w3[0][121] ), .B(n4829), .Z(n4830) );
  XNOR U6762 ( .A(n4831), .B(n4830), .Z(\w1[1][97] ) );
  XNOR U6763 ( .A(n4832), .B(key[226]), .Z(n4835) );
  XOR U6764 ( .A(\w3[0][122] ), .B(n4833), .Z(n4834) );
  XNOR U6765 ( .A(n4835), .B(n4834), .Z(\w1[1][98] ) );
  XOR U6766 ( .A(n4836), .B(key[227]), .Z(n4840) );
  XNOR U6767 ( .A(n4838), .B(n4837), .Z(n4839) );
  XNOR U6768 ( .A(n4840), .B(n4839), .Z(\w1[1][99] ) );
  XOR U6769 ( .A(\w3[0][10] ), .B(key[137]), .Z(n4842) );
  XNOR U6770 ( .A(\w3[0][2] ), .B(\w3[0][17] ), .Z(n4841) );
  XNOR U6771 ( .A(n4842), .B(n4841), .Z(n4843) );
  XNOR U6772 ( .A(n4844), .B(n4843), .Z(\w1[1][9] ) );
  XNOR U6773 ( .A(\w3[1][25] ), .B(\w3[1][1] ), .Z(n5264) );
  IV U6774 ( .A(\w3[1][16] ), .Z(n4976) );
  XOR U6775 ( .A(\w3[1][24] ), .B(n4976), .Z(n5216) );
  XNOR U6776 ( .A(\w3[1][8] ), .B(key[256]), .Z(n4845) );
  XNOR U6777 ( .A(n5216), .B(n4845), .Z(n4846) );
  XOR U6778 ( .A(n5264), .B(n4846), .Z(\w1[2][0] ) );
  XOR U6779 ( .A(\w3[1][96] ), .B(\w3[1][101] ), .Z(n4869) );
  XOR U6780 ( .A(\w3[1][116] ), .B(\w3[1][125] ), .Z(n4848) );
  IV U6781 ( .A(\w3[1][120] ), .Z(n4920) );
  XOR U6782 ( .A(n4920), .B(\w3[1][108] ), .Z(n4847) );
  XOR U6783 ( .A(n4848), .B(n4847), .Z(n4929) );
  XOR U6784 ( .A(n4929), .B(key[356]), .Z(n4849) );
  XOR U6785 ( .A(n4869), .B(n4849), .Z(n4850) );
  XNOR U6786 ( .A(\w3[1][124] ), .B(n4850), .Z(\w1[2][100] ) );
  XNOR U6787 ( .A(\w3[1][102] ), .B(\w3[1][126] ), .Z(n4878) );
  XNOR U6788 ( .A(n4878), .B(key[357]), .Z(n4852) );
  XNOR U6789 ( .A(\w3[1][109] ), .B(\w3[1][117] ), .Z(n4932) );
  XOR U6790 ( .A(\w3[1][125] ), .B(n4932), .Z(n4851) );
  XNOR U6791 ( .A(n4852), .B(n4851), .Z(\w1[2][101] ) );
  XOR U6792 ( .A(\w3[1][96] ), .B(\w3[1][103] ), .Z(n4879) );
  XOR U6793 ( .A(n4879), .B(key[358]), .Z(n4854) );
  XOR U6794 ( .A(n4920), .B(\w3[1][127] ), .Z(n4855) );
  XOR U6795 ( .A(\w3[1][110] ), .B(\w3[1][118] ), .Z(n4895) );
  XOR U6796 ( .A(n4855), .B(n4895), .Z(n4937) );
  XOR U6797 ( .A(\w3[1][126] ), .B(n4937), .Z(n4853) );
  XNOR U6798 ( .A(n4854), .B(n4853), .Z(\w1[2][102] ) );
  XNOR U6799 ( .A(\w3[1][111] ), .B(\w3[1][119] ), .Z(n4940) );
  XNOR U6800 ( .A(n4940), .B(key[359]), .Z(n4857) );
  XOR U6801 ( .A(\w3[1][96] ), .B(n4855), .Z(n4856) );
  XNOR U6802 ( .A(n4857), .B(n4856), .Z(\w1[2][103] ) );
  IV U6803 ( .A(\w3[1][97] ), .Z(n4915) );
  IV U6804 ( .A(\w3[1][112] ), .Z(n4911) );
  XOR U6805 ( .A(\w3[1][120] ), .B(n4911), .Z(n5245) );
  XOR U6806 ( .A(\w3[1][106] ), .B(\w3[1][98] ), .Z(n4859) );
  XNOR U6807 ( .A(\w3[1][97] ), .B(\w3[1][121] ), .Z(n5244) );
  XOR U6808 ( .A(n5244), .B(key[361]), .Z(n4858) );
  XNOR U6809 ( .A(n4859), .B(n4858), .Z(n4860) );
  XOR U6810 ( .A(\w3[1][113] ), .B(n4860), .Z(\w1[2][105] ) );
  IV U6811 ( .A(\w3[1][99] ), .Z(n4924) );
  XNOR U6812 ( .A(\w3[1][107] ), .B(n4924), .Z(n4862) );
  XOR U6813 ( .A(\w3[1][98] ), .B(\w3[1][122] ), .Z(n5249) );
  XNOR U6814 ( .A(n5249), .B(key[362]), .Z(n4861) );
  XNOR U6815 ( .A(n4862), .B(n4861), .Z(n4863) );
  XOR U6816 ( .A(\w3[1][114] ), .B(n4863), .Z(\w1[2][106] ) );
  IV U6817 ( .A(\w3[1][123] ), .Z(n5257) );
  XOR U6818 ( .A(\w3[1][99] ), .B(n5257), .Z(n5253) );
  XOR U6819 ( .A(\w3[1][108] ), .B(n5253), .Z(n4864) );
  XOR U6820 ( .A(\w3[1][104] ), .B(n4864), .Z(n4890) );
  XNOR U6821 ( .A(n4890), .B(key[363]), .Z(n4866) );
  IV U6822 ( .A(\w3[1][100] ), .Z(n4928) );
  XOR U6823 ( .A(\w3[1][96] ), .B(n4928), .Z(n5258) );
  XOR U6824 ( .A(\w3[1][115] ), .B(n5258), .Z(n4865) );
  XNOR U6825 ( .A(n4866), .B(n4865), .Z(\w1[2][107] ) );
  XOR U6826 ( .A(\w3[1][100] ), .B(\w3[1][104] ), .Z(n4868) );
  XNOR U6827 ( .A(\w3[1][124] ), .B(\w3[1][109] ), .Z(n4867) );
  XOR U6828 ( .A(n4868), .B(n4867), .Z(n4891) );
  XNOR U6829 ( .A(n4891), .B(key[364]), .Z(n4871) );
  XNOR U6830 ( .A(\w3[1][116] ), .B(n4869), .Z(n4870) );
  XNOR U6831 ( .A(n4871), .B(n4870), .Z(\w1[2][108] ) );
  XNOR U6832 ( .A(\w3[1][125] ), .B(\w3[1][101] ), .Z(n4894) );
  XNOR U6833 ( .A(n4894), .B(key[365]), .Z(n4873) );
  XNOR U6834 ( .A(\w3[1][102] ), .B(\w3[1][110] ), .Z(n4872) );
  XNOR U6835 ( .A(n4873), .B(n4872), .Z(n4874) );
  XOR U6836 ( .A(\w3[1][117] ), .B(n4874), .Z(\w1[2][109] ) );
  XOR U6837 ( .A(\w3[1][11] ), .B(\w3[1][3] ), .Z(n4876) );
  XNOR U6838 ( .A(\w3[1][2] ), .B(\w3[1][26] ), .Z(n4963) );
  XOR U6839 ( .A(n4963), .B(key[266]), .Z(n4875) );
  XNOR U6840 ( .A(n4876), .B(n4875), .Z(n4877) );
  XOR U6841 ( .A(\w3[1][18] ), .B(n4877), .Z(\w1[2][10] ) );
  XOR U6842 ( .A(\w3[1][111] ), .B(\w3[1][104] ), .Z(n4902) );
  XOR U6843 ( .A(n4878), .B(n4902), .Z(n4898) );
  XNOR U6844 ( .A(n4898), .B(key[366]), .Z(n4881) );
  XNOR U6845 ( .A(\w3[1][118] ), .B(n4879), .Z(n4880) );
  XNOR U6846 ( .A(n4881), .B(n4880), .Z(\w1[2][110] ) );
  XOR U6847 ( .A(\w3[1][127] ), .B(\w3[1][103] ), .Z(n4901) );
  XOR U6848 ( .A(n4901), .B(key[367]), .Z(n4883) );
  XNOR U6849 ( .A(\w3[1][96] ), .B(\w3[1][104] ), .Z(n4907) );
  XOR U6850 ( .A(\w3[1][119] ), .B(n4907), .Z(n4882) );
  XNOR U6851 ( .A(n4883), .B(n4882), .Z(\w1[2][111] ) );
  XNOR U6852 ( .A(\w3[1][105] ), .B(\w3[1][113] ), .Z(n5248) );
  XNOR U6853 ( .A(n5248), .B(key[368]), .Z(n4885) );
  XNOR U6854 ( .A(n4920), .B(n4907), .Z(n4884) );
  XNOR U6855 ( .A(n4885), .B(n4884), .Z(\w1[2][112] ) );
  XNOR U6856 ( .A(\w3[1][106] ), .B(\w3[1][114] ), .Z(n5252) );
  XNOR U6857 ( .A(n5252), .B(key[369]), .Z(n4887) );
  XOR U6858 ( .A(\w3[1][105] ), .B(n5244), .Z(n4886) );
  XNOR U6859 ( .A(n4887), .B(n4886), .Z(\w1[2][113] ) );
  IV U6860 ( .A(\w3[1][115] ), .Z(n4916) );
  XOR U6861 ( .A(\w3[1][107] ), .B(n4916), .Z(n4922) );
  XNOR U6862 ( .A(n4922), .B(key[370]), .Z(n4889) );
  XNOR U6863 ( .A(\w3[1][106] ), .B(n5249), .Z(n4888) );
  XNOR U6864 ( .A(n4889), .B(n4888), .Z(\w1[2][114] ) );
  XOR U6865 ( .A(\w3[1][116] ), .B(n4911), .Z(n4923) );
  XOR U6866 ( .A(\w3[1][117] ), .B(n4911), .Z(n4927) );
  XNOR U6867 ( .A(n4927), .B(key[372]), .Z(n4893) );
  XOR U6868 ( .A(\w3[1][108] ), .B(n4891), .Z(n4892) );
  XNOR U6869 ( .A(n4893), .B(n4892), .Z(\w1[2][116] ) );
  XNOR U6870 ( .A(n4894), .B(key[373]), .Z(n4897) );
  XNOR U6871 ( .A(\w3[1][109] ), .B(n4895), .Z(n4896) );
  XNOR U6872 ( .A(n4897), .B(n4896), .Z(\w1[2][117] ) );
  XOR U6873 ( .A(\w3[1][119] ), .B(n4911), .Z(n4936) );
  XNOR U6874 ( .A(n4936), .B(key[374]), .Z(n4900) );
  XOR U6875 ( .A(\w3[1][110] ), .B(n4898), .Z(n4899) );
  XNOR U6876 ( .A(n4900), .B(n4899), .Z(\w1[2][118] ) );
  XOR U6877 ( .A(n4901), .B(key[375]), .Z(n4904) );
  XNOR U6878 ( .A(\w3[1][112] ), .B(n4902), .Z(n4903) );
  XNOR U6879 ( .A(n4904), .B(n4903), .Z(\w1[2][119] ) );
  XNOR U6880 ( .A(\w3[1][3] ), .B(\w3[1][27] ), .Z(n4997) );
  XNOR U6881 ( .A(n4960), .B(key[267]), .Z(n4906) );
  XNOR U6882 ( .A(\w3[1][0] ), .B(\w3[1][4] ), .Z(n5029) );
  XOR U6883 ( .A(\w3[1][19] ), .B(n5029), .Z(n4905) );
  XNOR U6884 ( .A(n4906), .B(n4905), .Z(\w1[2][11] ) );
  XNOR U6885 ( .A(n4907), .B(key[376]), .Z(n4909) );
  XNOR U6886 ( .A(\w3[1][113] ), .B(\w3[1][121] ), .Z(n4908) );
  XNOR U6887 ( .A(n4909), .B(n4908), .Z(n4910) );
  XNOR U6888 ( .A(n4911), .B(n4910), .Z(\w1[2][120] ) );
  XNOR U6889 ( .A(n5248), .B(key[377]), .Z(n4913) );
  XNOR U6890 ( .A(\w3[1][114] ), .B(\w3[1][122] ), .Z(n4912) );
  XNOR U6891 ( .A(n4913), .B(n4912), .Z(n4914) );
  XNOR U6892 ( .A(n4915), .B(n4914), .Z(\w1[2][121] ) );
  XNOR U6893 ( .A(n5252), .B(key[378]), .Z(n4918) );
  XNOR U6894 ( .A(n4916), .B(n5257), .Z(n4917) );
  XNOR U6895 ( .A(n4918), .B(n4917), .Z(n4919) );
  XOR U6896 ( .A(\w3[1][98] ), .B(n4919), .Z(\w1[2][122] ) );
  XOR U6897 ( .A(\w3[1][124] ), .B(n4920), .Z(n4921) );
  XOR U6898 ( .A(n4922), .B(n4921), .Z(n5256) );
  XOR U6899 ( .A(n5256), .B(key[379]), .Z(n4926) );
  XNOR U6900 ( .A(n4924), .B(n4923), .Z(n4925) );
  XNOR U6901 ( .A(n4926), .B(n4925), .Z(\w1[2][123] ) );
  XNOR U6902 ( .A(n4927), .B(key[380]), .Z(n4931) );
  XNOR U6903 ( .A(n4929), .B(n4928), .Z(n4930) );
  XNOR U6904 ( .A(n4931), .B(n4930), .Z(\w1[2][124] ) );
  XOR U6905 ( .A(\w3[1][118] ), .B(key[381]), .Z(n4934) );
  XOR U6906 ( .A(n4932), .B(\w3[1][126] ), .Z(n4933) );
  XNOR U6907 ( .A(n4934), .B(n4933), .Z(n4935) );
  XOR U6908 ( .A(\w3[1][101] ), .B(n4935), .Z(\w1[2][125] ) );
  XNOR U6909 ( .A(n4936), .B(key[382]), .Z(n4939) );
  XOR U6910 ( .A(\w3[1][102] ), .B(n4937), .Z(n4938) );
  XNOR U6911 ( .A(n4939), .B(n4938), .Z(\w1[2][126] ) );
  XNOR U6912 ( .A(n5245), .B(key[383]), .Z(n4942) );
  XOR U6913 ( .A(\w3[1][103] ), .B(n4940), .Z(n4941) );
  XNOR U6914 ( .A(n4942), .B(n4941), .Z(\w1[2][127] ) );
  XOR U6915 ( .A(\w3[1][13] ), .B(\w3[1][28] ), .Z(n4944) );
  XNOR U6916 ( .A(\w3[1][8] ), .B(\w3[1][4] ), .Z(n4943) );
  XOR U6917 ( .A(n4944), .B(n4943), .Z(n4966) );
  XNOR U6918 ( .A(n4966), .B(key[268]), .Z(n4946) );
  XNOR U6919 ( .A(\w3[1][0] ), .B(\w3[1][5] ), .Z(n5064) );
  XOR U6920 ( .A(\w3[1][20] ), .B(n5064), .Z(n4945) );
  XNOR U6921 ( .A(n4946), .B(n4945), .Z(\w1[2][12] ) );
  IV U6922 ( .A(\w3[1][6] ), .Z(n5003) );
  XNOR U6923 ( .A(\w3[1][14] ), .B(n5003), .Z(n4948) );
  XNOR U6924 ( .A(\w3[1][5] ), .B(\w3[1][29] ), .Z(n4969) );
  XOR U6925 ( .A(n4969), .B(key[269]), .Z(n4947) );
  XNOR U6926 ( .A(n4948), .B(n4947), .Z(n4949) );
  XOR U6927 ( .A(\w3[1][21] ), .B(n4949), .Z(\w1[2][13] ) );
  IV U6928 ( .A(\w3[1][30] ), .Z(n5141) );
  XOR U6929 ( .A(\w3[1][6] ), .B(n5141), .Z(n5106) );
  XOR U6930 ( .A(\w3[1][8] ), .B(\w3[1][15] ), .Z(n4972) );
  XNOR U6931 ( .A(n5106), .B(n4972), .Z(n4970) );
  XOR U6932 ( .A(n4970), .B(key[270]), .Z(n4951) );
  XNOR U6933 ( .A(\w3[1][0] ), .B(\w3[1][7] ), .Z(n5142) );
  XOR U6934 ( .A(\w3[1][22] ), .B(n5142), .Z(n4950) );
  XNOR U6935 ( .A(n4951), .B(n4950), .Z(\w1[2][14] ) );
  XNOR U6936 ( .A(\w3[1][7] ), .B(\w3[1][31] ), .Z(n4971) );
  XNOR U6937 ( .A(n4971), .B(key[271]), .Z(n4953) );
  XOR U6938 ( .A(\w3[1][8] ), .B(\w3[1][0] ), .Z(n4975) );
  XNOR U6939 ( .A(\w3[1][23] ), .B(n4975), .Z(n4952) );
  XNOR U6940 ( .A(n4953), .B(n4952), .Z(\w1[2][15] ) );
  XNOR U6941 ( .A(\w3[1][17] ), .B(\w3[1][9] ), .Z(n4977) );
  XNOR U6942 ( .A(n4977), .B(key[272]), .Z(n4955) );
  XNOR U6943 ( .A(\w3[1][24] ), .B(n4975), .Z(n4954) );
  XNOR U6944 ( .A(n4955), .B(n4954), .Z(\w1[2][16] ) );
  XNOR U6945 ( .A(\w3[1][18] ), .B(\w3[1][10] ), .Z(n4996) );
  XNOR U6946 ( .A(n4996), .B(key[273]), .Z(n4957) );
  IV U6947 ( .A(\w3[1][9] ), .Z(n5213) );
  XNOR U6948 ( .A(n5264), .B(n5213), .Z(n4956) );
  XNOR U6949 ( .A(n4957), .B(n4956), .Z(\w1[2][17] ) );
  XNOR U6950 ( .A(\w3[1][11] ), .B(\w3[1][19] ), .Z(n4982) );
  XNOR U6951 ( .A(n4982), .B(key[274]), .Z(n4959) );
  XOR U6952 ( .A(n4963), .B(\w3[1][10] ), .Z(n4958) );
  XNOR U6953 ( .A(n4959), .B(n4958), .Z(\w1[2][18] ) );
  XOR U6954 ( .A(n4976), .B(\w3[1][20] ), .Z(n4983) );
  XNOR U6955 ( .A(n4983), .B(key[275]), .Z(n4962) );
  XOR U6956 ( .A(\w3[1][11] ), .B(n4960), .Z(n4961) );
  XNOR U6957 ( .A(n4962), .B(n4961), .Z(\w1[2][19] ) );
  XNOR U6958 ( .A(n4977), .B(key[257]), .Z(n4965) );
  XOR U6959 ( .A(\w3[1][25] ), .B(n4963), .Z(n4964) );
  XNOR U6960 ( .A(n4965), .B(n4964), .Z(\w1[2][1] ) );
  IV U6961 ( .A(\w3[1][21] ), .Z(n4991) );
  XOR U6962 ( .A(\w3[1][16] ), .B(n4991), .Z(n4988) );
  XNOR U6963 ( .A(n4988), .B(key[276]), .Z(n4968) );
  XOR U6964 ( .A(\w3[1][12] ), .B(n4966), .Z(n4967) );
  XNOR U6965 ( .A(n4968), .B(n4967), .Z(\w1[2][20] ) );
  IV U6966 ( .A(\w3[1][22] ), .Z(n4992) );
  XOR U6967 ( .A(\w3[1][14] ), .B(n4992), .Z(n5001) );
  XOR U6968 ( .A(n4976), .B(\w3[1][23] ), .Z(n5002) );
  XNOR U6969 ( .A(n4971), .B(key[279]), .Z(n4974) );
  XNOR U6970 ( .A(\w3[1][16] ), .B(n4972), .Z(n4973) );
  XNOR U6971 ( .A(n4974), .B(n4973), .Z(\w1[2][23] ) );
  XNOR U6972 ( .A(n4996), .B(key[282]), .Z(n4979) );
  XNOR U6973 ( .A(\w3[1][2] ), .B(\w3[1][19] ), .Z(n4978) );
  XNOR U6974 ( .A(n4979), .B(n4978), .Z(n4980) );
  XOR U6975 ( .A(\w3[1][27] ), .B(n4980), .Z(\w1[2][26] ) );
  IV U6976 ( .A(\w3[1][24] ), .Z(n5000) );
  XOR U6977 ( .A(n5000), .B(\w3[1][28] ), .Z(n4981) );
  XOR U6978 ( .A(n4982), .B(n4981), .Z(n5028) );
  XOR U6979 ( .A(n5028), .B(key[283]), .Z(n4985) );
  XOR U6980 ( .A(\w3[1][3] ), .B(n4983), .Z(n4984) );
  XNOR U6981 ( .A(n4985), .B(n4984), .Z(\w1[2][27] ) );
  XOR U6982 ( .A(\w3[1][20] ), .B(\w3[1][29] ), .Z(n4987) );
  XOR U6983 ( .A(n5000), .B(\w3[1][12] ), .Z(n4986) );
  XOR U6984 ( .A(n4987), .B(n4986), .Z(n5063) );
  XNOR U6985 ( .A(n5063), .B(key[284]), .Z(n4990) );
  XOR U6986 ( .A(\w3[1][4] ), .B(n4988), .Z(n4989) );
  XNOR U6987 ( .A(n4990), .B(n4989), .Z(\w1[2][28] ) );
  XOR U6988 ( .A(\w3[1][13] ), .B(n4991), .Z(n5105) );
  XNOR U6989 ( .A(n5105), .B(key[285]), .Z(n4994) );
  XNOR U6990 ( .A(n4992), .B(n5141), .Z(n4993) );
  XNOR U6991 ( .A(n4994), .B(n4993), .Z(n4995) );
  XOR U6992 ( .A(\w3[1][5] ), .B(n4995), .Z(\w1[2][29] ) );
  XNOR U6993 ( .A(n4996), .B(key[258]), .Z(n4999) );
  XOR U6994 ( .A(\w3[1][26] ), .B(n4997), .Z(n4998) );
  XNOR U6995 ( .A(n4999), .B(n4998), .Z(\w1[2][2] ) );
  XOR U6996 ( .A(n5000), .B(\w3[1][31] ), .Z(n5177) );
  XNOR U6997 ( .A(n5001), .B(n5177), .Z(n5140) );
  XNOR U6998 ( .A(n5140), .B(key[286]), .Z(n5005) );
  XNOR U6999 ( .A(n5003), .B(n5002), .Z(n5004) );
  XNOR U7000 ( .A(n5005), .B(n5004), .Z(\w1[2][30] ) );
  XNOR U7001 ( .A(\w3[1][15] ), .B(\w3[1][23] ), .Z(n5176) );
  XNOR U7002 ( .A(n5176), .B(key[287]), .Z(n5007) );
  XOR U7003 ( .A(n5216), .B(\w3[1][7] ), .Z(n5006) );
  XNOR U7004 ( .A(n5007), .B(n5006), .Z(\w1[2][31] ) );
  XOR U7005 ( .A(\w3[1][33] ), .B(\w3[1][57] ), .Z(n5060) );
  XOR U7006 ( .A(n5060), .B(key[288]), .Z(n5009) );
  XNOR U7007 ( .A(\w3[1][48] ), .B(\w3[1][56] ), .Z(n5122) );
  XOR U7008 ( .A(n5122), .B(\w3[1][40] ), .Z(n5008) );
  XNOR U7009 ( .A(n5009), .B(n5008), .Z(\w1[2][32] ) );
  XNOR U7010 ( .A(\w3[1][34] ), .B(\w3[1][58] ), .Z(n5068) );
  XOR U7011 ( .A(\w3[1][57] ), .B(\w3[1][49] ), .Z(n5086) );
  XNOR U7012 ( .A(n5086), .B(key[289]), .Z(n5010) );
  XNOR U7013 ( .A(n5068), .B(n5010), .Z(n5011) );
  XNOR U7014 ( .A(\w3[1][41] ), .B(n5011), .Z(\w1[2][33] ) );
  XNOR U7015 ( .A(n5038), .B(key[290]), .Z(n5013) );
  XNOR U7016 ( .A(\w3[1][50] ), .B(\w3[1][42] ), .Z(n5096) );
  XOR U7017 ( .A(\w3[1][58] ), .B(n5096), .Z(n5012) );
  XNOR U7018 ( .A(n5013), .B(n5012), .Z(\w1[2][34] ) );
  XOR U7019 ( .A(\w3[1][36] ), .B(\w3[1][32] ), .Z(n5040) );
  XOR U7020 ( .A(n5040), .B(key[291]), .Z(n5016) );
  IV U7021 ( .A(\w3[1][51] ), .Z(n5095) );
  XOR U7022 ( .A(\w3[1][43] ), .B(n5095), .Z(n5067) );
  XOR U7023 ( .A(\w3[1][56] ), .B(n5067), .Z(n5014) );
  XNOR U7024 ( .A(\w3[1][60] ), .B(n5014), .Z(n5101) );
  XNOR U7025 ( .A(\w3[1][59] ), .B(n5101), .Z(n5015) );
  XNOR U7026 ( .A(n5016), .B(n5015), .Z(\w1[2][35] ) );
  XOR U7027 ( .A(\w3[1][32] ), .B(\w3[1][37] ), .Z(n5046) );
  XOR U7028 ( .A(\w3[1][52] ), .B(\w3[1][61] ), .Z(n5018) );
  XNOR U7029 ( .A(\w3[1][56] ), .B(\w3[1][44] ), .Z(n5017) );
  XOR U7030 ( .A(n5018), .B(n5017), .Z(n5110) );
  XOR U7031 ( .A(n5110), .B(key[292]), .Z(n5019) );
  XOR U7032 ( .A(n5046), .B(n5019), .Z(n5020) );
  XNOR U7033 ( .A(\w3[1][60] ), .B(n5020), .Z(\w1[2][36] ) );
  XNOR U7034 ( .A(\w3[1][38] ), .B(\w3[1][62] ), .Z(n5052) );
  XNOR U7035 ( .A(n5052), .B(key[293]), .Z(n5022) );
  IV U7036 ( .A(\w3[1][45] ), .Z(n5075) );
  XOR U7037 ( .A(\w3[1][53] ), .B(n5075), .Z(n5113) );
  XOR U7038 ( .A(\w3[1][61] ), .B(n5113), .Z(n5021) );
  XNOR U7039 ( .A(n5022), .B(n5021), .Z(\w1[2][37] ) );
  XOR U7040 ( .A(\w3[1][32] ), .B(\w3[1][39] ), .Z(n5053) );
  XOR U7041 ( .A(n5053), .B(key[294]), .Z(n5024) );
  XNOR U7042 ( .A(\w3[1][46] ), .B(\w3[1][54] ), .Z(n5074) );
  XOR U7043 ( .A(\w3[1][56] ), .B(\w3[1][63] ), .Z(n5025) );
  XOR U7044 ( .A(n5074), .B(n5025), .Z(n5118) );
  XOR U7045 ( .A(\w3[1][62] ), .B(n5118), .Z(n5023) );
  XNOR U7046 ( .A(n5024), .B(n5023), .Z(\w1[2][38] ) );
  XNOR U7047 ( .A(\w3[1][55] ), .B(\w3[1][47] ), .Z(n5121) );
  XNOR U7048 ( .A(n5121), .B(key[295]), .Z(n5027) );
  XNOR U7049 ( .A(\w3[1][32] ), .B(n5025), .Z(n5026) );
  XNOR U7050 ( .A(n5027), .B(n5026), .Z(\w1[2][39] ) );
  XOR U7051 ( .A(n5028), .B(key[259]), .Z(n5031) );
  XOR U7052 ( .A(n5029), .B(\w3[1][27] ), .Z(n5030) );
  XNOR U7053 ( .A(n5031), .B(n5030), .Z(\w1[2][3] ) );
  IV U7054 ( .A(\w3[1][33] ), .Z(n5091) );
  XOR U7055 ( .A(\w3[1][42] ), .B(key[297]), .Z(n5033) );
  XNOR U7056 ( .A(n5086), .B(\w3[1][34] ), .Z(n5032) );
  XNOR U7057 ( .A(n5033), .B(n5032), .Z(n5034) );
  XNOR U7058 ( .A(n5091), .B(n5034), .Z(\w1[2][41] ) );
  XOR U7059 ( .A(\w3[1][43] ), .B(key[298]), .Z(n5036) );
  IV U7060 ( .A(\w3[1][35] ), .Z(n5102) );
  XOR U7061 ( .A(\w3[1][50] ), .B(n5102), .Z(n5035) );
  XNOR U7062 ( .A(n5036), .B(n5035), .Z(n5037) );
  XNOR U7063 ( .A(n5037), .B(n5068), .Z(\w1[2][42] ) );
  IV U7064 ( .A(\w3[1][40] ), .Z(n5043) );
  XNOR U7065 ( .A(n5043), .B(n5038), .Z(n5039) );
  XOR U7066 ( .A(\w3[1][44] ), .B(n5039), .Z(n5069) );
  XNOR U7067 ( .A(n5069), .B(key[299]), .Z(n5042) );
  XNOR U7068 ( .A(\w3[1][51] ), .B(n5040), .Z(n5041) );
  XNOR U7069 ( .A(n5042), .B(n5041), .Z(\w1[2][43] ) );
  XOR U7070 ( .A(\w3[1][36] ), .B(\w3[1][45] ), .Z(n5045) );
  XOR U7071 ( .A(n5043), .B(\w3[1][60] ), .Z(n5044) );
  XOR U7072 ( .A(n5045), .B(n5044), .Z(n5070) );
  XNOR U7073 ( .A(n5070), .B(key[300]), .Z(n5048) );
  XNOR U7074 ( .A(\w3[1][52] ), .B(n5046), .Z(n5047) );
  XNOR U7075 ( .A(n5048), .B(n5047), .Z(\w1[2][44] ) );
  XNOR U7076 ( .A(\w3[1][61] ), .B(\w3[1][37] ), .Z(n5073) );
  XNOR U7077 ( .A(n5073), .B(key[301]), .Z(n5050) );
  XNOR U7078 ( .A(\w3[1][38] ), .B(\w3[1][46] ), .Z(n5049) );
  XNOR U7079 ( .A(n5050), .B(n5049), .Z(n5051) );
  XOR U7080 ( .A(\w3[1][53] ), .B(n5051), .Z(\w1[2][45] ) );
  XOR U7081 ( .A(\w3[1][40] ), .B(\w3[1][47] ), .Z(n5082) );
  XOR U7082 ( .A(n5052), .B(n5082), .Z(n5078) );
  XNOR U7083 ( .A(n5078), .B(key[302]), .Z(n5055) );
  XNOR U7084 ( .A(\w3[1][54] ), .B(n5053), .Z(n5054) );
  XNOR U7085 ( .A(n5055), .B(n5054), .Z(\w1[2][46] ) );
  XOR U7086 ( .A(\w3[1][63] ), .B(\w3[1][39] ), .Z(n5081) );
  XOR U7087 ( .A(n5081), .B(key[303]), .Z(n5057) );
  XNOR U7088 ( .A(\w3[1][40] ), .B(\w3[1][32] ), .Z(n5085) );
  XOR U7089 ( .A(\w3[1][55] ), .B(n5085), .Z(n5056) );
  XNOR U7090 ( .A(n5057), .B(n5056), .Z(\w1[2][47] ) );
  XNOR U7091 ( .A(\w3[1][41] ), .B(\w3[1][49] ), .Z(n5090) );
  XNOR U7092 ( .A(n5090), .B(key[304]), .Z(n5059) );
  XOR U7093 ( .A(\w3[1][56] ), .B(n5085), .Z(n5058) );
  XNOR U7094 ( .A(n5059), .B(n5058), .Z(\w1[2][48] ) );
  XNOR U7095 ( .A(n5096), .B(key[305]), .Z(n5062) );
  XNOR U7096 ( .A(n5060), .B(\w3[1][41] ), .Z(n5061) );
  XNOR U7097 ( .A(n5062), .B(n5061), .Z(\w1[2][49] ) );
  XNOR U7098 ( .A(n5063), .B(key[260]), .Z(n5066) );
  XOR U7099 ( .A(n5064), .B(\w3[1][28] ), .Z(n5065) );
  XNOR U7100 ( .A(n5066), .B(n5065), .Z(\w1[2][4] ) );
  IV U7101 ( .A(\w3[1][48] ), .Z(n5087) );
  XOR U7102 ( .A(n5087), .B(\w3[1][52] ), .Z(n5100) );
  XNOR U7103 ( .A(n5109), .B(key[308]), .Z(n5072) );
  XOR U7104 ( .A(\w3[1][44] ), .B(n5070), .Z(n5071) );
  XNOR U7105 ( .A(n5072), .B(n5071), .Z(\w1[2][52] ) );
  XNOR U7106 ( .A(n5073), .B(key[309]), .Z(n5077) );
  XNOR U7107 ( .A(n5075), .B(n5074), .Z(n5076) );
  XNOR U7108 ( .A(n5077), .B(n5076), .Z(\w1[2][53] ) );
  XOR U7109 ( .A(n5087), .B(\w3[1][55] ), .Z(n5117) );
  XNOR U7110 ( .A(n5117), .B(key[310]), .Z(n5080) );
  XOR U7111 ( .A(\w3[1][46] ), .B(n5078), .Z(n5079) );
  XNOR U7112 ( .A(n5080), .B(n5079), .Z(\w1[2][54] ) );
  XOR U7113 ( .A(n5081), .B(key[311]), .Z(n5084) );
  XNOR U7114 ( .A(\w3[1][48] ), .B(n5082), .Z(n5083) );
  XNOR U7115 ( .A(n5084), .B(n5083), .Z(\w1[2][55] ) );
  XNOR U7116 ( .A(n5085), .B(key[312]), .Z(n5089) );
  XOR U7117 ( .A(n5087), .B(n5086), .Z(n5088) );
  XNOR U7118 ( .A(n5089), .B(n5088), .Z(\w1[2][56] ) );
  XNOR U7119 ( .A(n5090), .B(key[313]), .Z(n5093) );
  XOR U7120 ( .A(n5091), .B(\w3[1][50] ), .Z(n5092) );
  XNOR U7121 ( .A(n5093), .B(n5092), .Z(n5094) );
  XOR U7122 ( .A(\w3[1][58] ), .B(n5094), .Z(\w1[2][57] ) );
  XNOR U7123 ( .A(n5095), .B(key[314]), .Z(n5098) );
  XOR U7124 ( .A(n5096), .B(\w3[1][59] ), .Z(n5097) );
  XNOR U7125 ( .A(n5098), .B(n5097), .Z(n5099) );
  XOR U7126 ( .A(\w3[1][34] ), .B(n5099), .Z(\w1[2][58] ) );
  XNOR U7127 ( .A(n5100), .B(key[315]), .Z(n5104) );
  XOR U7128 ( .A(n5102), .B(n5101), .Z(n5103) );
  XNOR U7129 ( .A(n5104), .B(n5103), .Z(\w1[2][59] ) );
  XNOR U7130 ( .A(n5105), .B(key[261]), .Z(n5108) );
  XOR U7131 ( .A(\w3[1][29] ), .B(n5106), .Z(n5107) );
  XNOR U7132 ( .A(n5108), .B(n5107), .Z(\w1[2][5] ) );
  XNOR U7133 ( .A(n5109), .B(key[316]), .Z(n5112) );
  XOR U7134 ( .A(\w3[1][36] ), .B(n5110), .Z(n5111) );
  XNOR U7135 ( .A(n5112), .B(n5111), .Z(\w1[2][60] ) );
  XOR U7136 ( .A(\w3[1][54] ), .B(key[317]), .Z(n5115) );
  XOR U7137 ( .A(n5113), .B(\w3[1][62] ), .Z(n5114) );
  XNOR U7138 ( .A(n5115), .B(n5114), .Z(n5116) );
  XOR U7139 ( .A(\w3[1][37] ), .B(n5116), .Z(\w1[2][61] ) );
  XNOR U7140 ( .A(n5117), .B(key[318]), .Z(n5120) );
  XOR U7141 ( .A(\w3[1][38] ), .B(n5118), .Z(n5119) );
  XNOR U7142 ( .A(n5120), .B(n5119), .Z(\w1[2][62] ) );
  XNOR U7143 ( .A(n5121), .B(key[319]), .Z(n5124) );
  XOR U7144 ( .A(n5122), .B(\w3[1][39] ), .Z(n5123) );
  XNOR U7145 ( .A(n5124), .B(n5123), .Z(\w1[2][63] ) );
  XOR U7146 ( .A(\w3[1][65] ), .B(\w3[1][89] ), .Z(n5182) );
  XOR U7147 ( .A(n5182), .B(key[320]), .Z(n5126) );
  XNOR U7148 ( .A(\w3[1][80] ), .B(\w3[1][88] ), .Z(n5241) );
  XOR U7149 ( .A(n5241), .B(\w3[1][72] ), .Z(n5125) );
  XNOR U7150 ( .A(n5126), .B(n5125), .Z(\w1[2][64] ) );
  XNOR U7151 ( .A(\w3[1][66] ), .B(\w3[1][90] ), .Z(n5186) );
  XOR U7152 ( .A(\w3[1][89] ), .B(\w3[1][81] ), .Z(n5204) );
  XNOR U7153 ( .A(n5204), .B(key[321]), .Z(n5127) );
  XNOR U7154 ( .A(n5186), .B(n5127), .Z(n5128) );
  XNOR U7155 ( .A(\w3[1][73] ), .B(n5128), .Z(\w1[2][65] ) );
  XNOR U7156 ( .A(n5156), .B(key[322]), .Z(n5130) );
  XNOR U7157 ( .A(\w3[1][82] ), .B(\w3[1][74] ), .Z(n5219) );
  XOR U7158 ( .A(\w3[1][90] ), .B(n5219), .Z(n5129) );
  XNOR U7159 ( .A(n5130), .B(n5129), .Z(\w1[2][66] ) );
  XOR U7160 ( .A(\w3[1][68] ), .B(\w3[1][64] ), .Z(n5158) );
  XOR U7161 ( .A(n5158), .B(key[323]), .Z(n5133) );
  IV U7162 ( .A(\w3[1][83] ), .Z(n5218) );
  XOR U7163 ( .A(\w3[1][75] ), .B(n5218), .Z(n5185) );
  XOR U7164 ( .A(\w3[1][88] ), .B(n5185), .Z(n5131) );
  XNOR U7165 ( .A(\w3[1][92] ), .B(n5131), .Z(n5224) );
  XNOR U7166 ( .A(\w3[1][91] ), .B(n5224), .Z(n5132) );
  XNOR U7167 ( .A(n5133), .B(n5132), .Z(\w1[2][67] ) );
  XOR U7168 ( .A(\w3[1][64] ), .B(\w3[1][69] ), .Z(n5164) );
  XOR U7169 ( .A(\w3[1][84] ), .B(\w3[1][93] ), .Z(n5135) );
  XNOR U7170 ( .A(\w3[1][88] ), .B(\w3[1][76] ), .Z(n5134) );
  XOR U7171 ( .A(n5135), .B(n5134), .Z(n5229) );
  XOR U7172 ( .A(n5229), .B(key[324]), .Z(n5136) );
  XOR U7173 ( .A(n5164), .B(n5136), .Z(n5137) );
  XNOR U7174 ( .A(\w3[1][92] ), .B(n5137), .Z(\w1[2][68] ) );
  XNOR U7175 ( .A(\w3[1][70] ), .B(\w3[1][94] ), .Z(n5170) );
  XNOR U7176 ( .A(n5170), .B(key[325]), .Z(n5139) );
  IV U7177 ( .A(\w3[1][77] ), .Z(n5193) );
  XOR U7178 ( .A(\w3[1][85] ), .B(n5193), .Z(n5232) );
  XOR U7179 ( .A(\w3[1][93] ), .B(n5232), .Z(n5138) );
  XNOR U7180 ( .A(n5139), .B(n5138), .Z(\w1[2][69] ) );
  XNOR U7181 ( .A(n5140), .B(key[262]), .Z(n5144) );
  XNOR U7182 ( .A(n5142), .B(n5141), .Z(n5143) );
  XNOR U7183 ( .A(n5144), .B(n5143), .Z(\w1[2][6] ) );
  XOR U7184 ( .A(\w3[1][64] ), .B(\w3[1][71] ), .Z(n5171) );
  XOR U7185 ( .A(n5171), .B(key[326]), .Z(n5146) );
  XNOR U7186 ( .A(\w3[1][88] ), .B(\w3[1][95] ), .Z(n5147) );
  XOR U7187 ( .A(\w3[1][78] ), .B(\w3[1][86] ), .Z(n5192) );
  XOR U7188 ( .A(n5147), .B(n5192), .Z(n5237) );
  XOR U7189 ( .A(\w3[1][94] ), .B(n5237), .Z(n5145) );
  XNOR U7190 ( .A(n5146), .B(n5145), .Z(\w1[2][70] ) );
  XNOR U7191 ( .A(\w3[1][79] ), .B(\w3[1][87] ), .Z(n5240) );
  XNOR U7192 ( .A(n5240), .B(key[327]), .Z(n5149) );
  XOR U7193 ( .A(\w3[1][64] ), .B(n5147), .Z(n5148) );
  XNOR U7194 ( .A(n5149), .B(n5148), .Z(\w1[2][71] ) );
  IV U7195 ( .A(\w3[1][65] ), .Z(n5209) );
  XOR U7196 ( .A(\w3[1][74] ), .B(key[329]), .Z(n5151) );
  XNOR U7197 ( .A(n5204), .B(\w3[1][66] ), .Z(n5150) );
  XNOR U7198 ( .A(n5151), .B(n5150), .Z(n5152) );
  XNOR U7199 ( .A(n5209), .B(n5152), .Z(\w1[2][73] ) );
  XOR U7200 ( .A(\w3[1][75] ), .B(key[330]), .Z(n5154) );
  IV U7201 ( .A(\w3[1][67] ), .Z(n5225) );
  XOR U7202 ( .A(\w3[1][82] ), .B(n5225), .Z(n5153) );
  XNOR U7203 ( .A(n5154), .B(n5153), .Z(n5155) );
  XNOR U7204 ( .A(n5155), .B(n5186), .Z(\w1[2][74] ) );
  IV U7205 ( .A(\w3[1][72] ), .Z(n5161) );
  XNOR U7206 ( .A(n5161), .B(n5156), .Z(n5157) );
  XOR U7207 ( .A(\w3[1][76] ), .B(n5157), .Z(n5187) );
  XNOR U7208 ( .A(n5187), .B(key[331]), .Z(n5160) );
  XNOR U7209 ( .A(\w3[1][83] ), .B(n5158), .Z(n5159) );
  XNOR U7210 ( .A(n5160), .B(n5159), .Z(\w1[2][75] ) );
  XOR U7211 ( .A(\w3[1][68] ), .B(\w3[1][77] ), .Z(n5163) );
  XOR U7212 ( .A(n5161), .B(\w3[1][92] ), .Z(n5162) );
  XOR U7213 ( .A(n5163), .B(n5162), .Z(n5188) );
  XNOR U7214 ( .A(n5188), .B(key[332]), .Z(n5166) );
  XNOR U7215 ( .A(\w3[1][84] ), .B(n5164), .Z(n5165) );
  XNOR U7216 ( .A(n5166), .B(n5165), .Z(\w1[2][76] ) );
  XNOR U7217 ( .A(\w3[1][93] ), .B(\w3[1][69] ), .Z(n5191) );
  XNOR U7218 ( .A(n5191), .B(key[333]), .Z(n5168) );
  XNOR U7219 ( .A(\w3[1][70] ), .B(\w3[1][78] ), .Z(n5167) );
  XNOR U7220 ( .A(n5168), .B(n5167), .Z(n5169) );
  XOR U7221 ( .A(\w3[1][85] ), .B(n5169), .Z(\w1[2][77] ) );
  XOR U7222 ( .A(\w3[1][72] ), .B(\w3[1][79] ), .Z(n5200) );
  XOR U7223 ( .A(n5170), .B(n5200), .Z(n5196) );
  XNOR U7224 ( .A(n5196), .B(key[334]), .Z(n5173) );
  XNOR U7225 ( .A(\w3[1][86] ), .B(n5171), .Z(n5172) );
  XNOR U7226 ( .A(n5173), .B(n5172), .Z(\w1[2][78] ) );
  XOR U7227 ( .A(\w3[1][95] ), .B(\w3[1][71] ), .Z(n5199) );
  XOR U7228 ( .A(n5199), .B(key[335]), .Z(n5175) );
  XNOR U7229 ( .A(\w3[1][72] ), .B(\w3[1][64] ), .Z(n5203) );
  XOR U7230 ( .A(\w3[1][87] ), .B(n5203), .Z(n5174) );
  XNOR U7231 ( .A(n5175), .B(n5174), .Z(\w1[2][79] ) );
  XNOR U7232 ( .A(n5176), .B(key[263]), .Z(n5179) );
  XOR U7233 ( .A(\w3[1][0] ), .B(n5177), .Z(n5178) );
  XNOR U7234 ( .A(n5179), .B(n5178), .Z(\w1[2][7] ) );
  XNOR U7235 ( .A(\w3[1][73] ), .B(\w3[1][81] ), .Z(n5208) );
  XNOR U7236 ( .A(n5208), .B(key[336]), .Z(n5181) );
  XOR U7237 ( .A(\w3[1][88] ), .B(n5203), .Z(n5180) );
  XNOR U7238 ( .A(n5181), .B(n5180), .Z(\w1[2][80] ) );
  XNOR U7239 ( .A(n5219), .B(key[337]), .Z(n5184) );
  XNOR U7240 ( .A(n5182), .B(\w3[1][73] ), .Z(n5183) );
  XNOR U7241 ( .A(n5184), .B(n5183), .Z(\w1[2][81] ) );
  IV U7242 ( .A(\w3[1][80] ), .Z(n5205) );
  XOR U7243 ( .A(n5205), .B(\w3[1][84] ), .Z(n5223) );
  XNOR U7244 ( .A(n5228), .B(key[340]), .Z(n5190) );
  XOR U7245 ( .A(\w3[1][76] ), .B(n5188), .Z(n5189) );
  XNOR U7246 ( .A(n5190), .B(n5189), .Z(\w1[2][84] ) );
  XNOR U7247 ( .A(n5191), .B(key[341]), .Z(n5195) );
  XOR U7248 ( .A(n5193), .B(n5192), .Z(n5194) );
  XNOR U7249 ( .A(n5195), .B(n5194), .Z(\w1[2][85] ) );
  XOR U7250 ( .A(n5205), .B(\w3[1][87] ), .Z(n5236) );
  XNOR U7251 ( .A(n5236), .B(key[342]), .Z(n5198) );
  XOR U7252 ( .A(\w3[1][78] ), .B(n5196), .Z(n5197) );
  XNOR U7253 ( .A(n5198), .B(n5197), .Z(\w1[2][86] ) );
  XOR U7254 ( .A(n5199), .B(key[343]), .Z(n5202) );
  XNOR U7255 ( .A(\w3[1][80] ), .B(n5200), .Z(n5201) );
  XNOR U7256 ( .A(n5202), .B(n5201), .Z(\w1[2][87] ) );
  XNOR U7257 ( .A(n5203), .B(key[344]), .Z(n5207) );
  XOR U7258 ( .A(n5205), .B(n5204), .Z(n5206) );
  XNOR U7259 ( .A(n5207), .B(n5206), .Z(\w1[2][88] ) );
  XNOR U7260 ( .A(n5208), .B(key[345]), .Z(n5211) );
  XOR U7261 ( .A(n5209), .B(\w3[1][82] ), .Z(n5210) );
  XNOR U7262 ( .A(n5211), .B(n5210), .Z(n5212) );
  XOR U7263 ( .A(\w3[1][90] ), .B(n5212), .Z(\w1[2][89] ) );
  XNOR U7264 ( .A(n5213), .B(key[264]), .Z(n5215) );
  XNOR U7265 ( .A(\w3[1][1] ), .B(\w3[1][0] ), .Z(n5214) );
  XNOR U7266 ( .A(n5215), .B(n5214), .Z(n5217) );
  XNOR U7267 ( .A(n5217), .B(n5216), .Z(\w1[2][8] ) );
  XNOR U7268 ( .A(n5218), .B(key[346]), .Z(n5221) );
  XOR U7269 ( .A(n5219), .B(\w3[1][91] ), .Z(n5220) );
  XNOR U7270 ( .A(n5221), .B(n5220), .Z(n5222) );
  XOR U7271 ( .A(\w3[1][66] ), .B(n5222), .Z(\w1[2][90] ) );
  XNOR U7272 ( .A(n5223), .B(key[347]), .Z(n5227) );
  XOR U7273 ( .A(n5225), .B(n5224), .Z(n5226) );
  XNOR U7274 ( .A(n5227), .B(n5226), .Z(\w1[2][91] ) );
  XNOR U7275 ( .A(n5228), .B(key[348]), .Z(n5231) );
  XOR U7276 ( .A(\w3[1][68] ), .B(n5229), .Z(n5230) );
  XNOR U7277 ( .A(n5231), .B(n5230), .Z(\w1[2][92] ) );
  XOR U7278 ( .A(\w3[1][86] ), .B(key[349]), .Z(n5234) );
  XOR U7279 ( .A(n5232), .B(\w3[1][94] ), .Z(n5233) );
  XNOR U7280 ( .A(n5234), .B(n5233), .Z(n5235) );
  XOR U7281 ( .A(\w3[1][69] ), .B(n5235), .Z(\w1[2][93] ) );
  XNOR U7282 ( .A(n5236), .B(key[350]), .Z(n5239) );
  XOR U7283 ( .A(\w3[1][70] ), .B(n5237), .Z(n5238) );
  XNOR U7284 ( .A(n5239), .B(n5238), .Z(\w1[2][94] ) );
  XNOR U7285 ( .A(n5240), .B(key[351]), .Z(n5243) );
  XOR U7286 ( .A(n5241), .B(\w3[1][71] ), .Z(n5242) );
  XNOR U7287 ( .A(n5243), .B(n5242), .Z(\w1[2][95] ) );
  XOR U7288 ( .A(\w3[1][104] ), .B(key[352]), .Z(n5247) );
  XNOR U7289 ( .A(n5245), .B(n5244), .Z(n5246) );
  XNOR U7290 ( .A(n5247), .B(n5246), .Z(\w1[2][96] ) );
  XNOR U7291 ( .A(n5248), .B(key[353]), .Z(n5251) );
  XNOR U7292 ( .A(\w3[1][121] ), .B(n5249), .Z(n5250) );
  XNOR U7293 ( .A(n5251), .B(n5250), .Z(\w1[2][97] ) );
  XNOR U7294 ( .A(n5252), .B(key[354]), .Z(n5255) );
  XOR U7295 ( .A(\w3[1][122] ), .B(n5253), .Z(n5254) );
  XNOR U7296 ( .A(n5255), .B(n5254), .Z(\w1[2][98] ) );
  XOR U7297 ( .A(n5256), .B(key[355]), .Z(n5260) );
  XNOR U7298 ( .A(n5258), .B(n5257), .Z(n5259) );
  XNOR U7299 ( .A(n5260), .B(n5259), .Z(\w1[2][99] ) );
  XOR U7300 ( .A(\w3[1][10] ), .B(key[265]), .Z(n5262) );
  XNOR U7301 ( .A(\w3[1][2] ), .B(\w3[1][17] ), .Z(n5261) );
  XNOR U7302 ( .A(n5262), .B(n5261), .Z(n5263) );
  XNOR U7303 ( .A(n5264), .B(n5263), .Z(\w1[2][9] ) );
  XNOR U7304 ( .A(\w3[2][25] ), .B(\w3[2][1] ), .Z(n5686) );
  IV U7305 ( .A(\w3[2][16] ), .Z(n5394) );
  XOR U7306 ( .A(\w3[2][24] ), .B(n5394), .Z(n5639) );
  XNOR U7307 ( .A(\w3[2][8] ), .B(key[384]), .Z(n5265) );
  XNOR U7308 ( .A(n5639), .B(n5265), .Z(n5266) );
  XOR U7309 ( .A(n5686), .B(n5266), .Z(\w1[3][0] ) );
  XOR U7310 ( .A(\w3[2][96] ), .B(\w3[2][101] ), .Z(n5288) );
  XOR U7311 ( .A(\w3[2][116] ), .B(\w3[2][125] ), .Z(n5268) );
  IV U7312 ( .A(\w3[2][120] ), .Z(n5341) );
  XOR U7313 ( .A(n5341), .B(\w3[2][108] ), .Z(n5267) );
  XOR U7314 ( .A(n5268), .B(n5267), .Z(n5349) );
  XOR U7315 ( .A(n5349), .B(key[484]), .Z(n5269) );
  XOR U7316 ( .A(n5288), .B(n5269), .Z(n5270) );
  XNOR U7317 ( .A(\w3[2][124] ), .B(n5270), .Z(\w1[3][100] ) );
  XNOR U7318 ( .A(\w3[2][102] ), .B(\w3[2][126] ), .Z(n5297) );
  XNOR U7319 ( .A(n5297), .B(key[485]), .Z(n5272) );
  XNOR U7320 ( .A(\w3[2][109] ), .B(\w3[2][117] ), .Z(n5352) );
  XOR U7321 ( .A(\w3[2][125] ), .B(n5352), .Z(n5271) );
  XNOR U7322 ( .A(n5272), .B(n5271), .Z(\w1[3][101] ) );
  XOR U7323 ( .A(\w3[2][96] ), .B(\w3[2][103] ), .Z(n5298) );
  XOR U7324 ( .A(n5298), .B(key[486]), .Z(n5274) );
  XOR U7325 ( .A(n5341), .B(\w3[2][127] ), .Z(n5275) );
  XOR U7326 ( .A(\w3[2][110] ), .B(\w3[2][118] ), .Z(n5316) );
  XOR U7327 ( .A(n5275), .B(n5316), .Z(n5357) );
  XOR U7328 ( .A(\w3[2][126] ), .B(n5357), .Z(n5273) );
  XNOR U7329 ( .A(n5274), .B(n5273), .Z(\w1[3][102] ) );
  XNOR U7330 ( .A(\w3[2][111] ), .B(\w3[2][119] ), .Z(n5360) );
  XNOR U7331 ( .A(n5360), .B(key[487]), .Z(n5277) );
  XOR U7332 ( .A(\w3[2][96] ), .B(n5275), .Z(n5276) );
  XNOR U7333 ( .A(n5277), .B(n5276), .Z(\w1[3][103] ) );
  IV U7334 ( .A(\w3[2][97] ), .Z(n5336) );
  IV U7335 ( .A(\w3[2][112] ), .Z(n5332) );
  XOR U7336 ( .A(\w3[2][120] ), .B(n5332), .Z(n5668) );
  XOR U7337 ( .A(\w3[2][106] ), .B(\w3[2][98] ), .Z(n5339) );
  XNOR U7338 ( .A(\w3[2][97] ), .B(\w3[2][121] ), .Z(n5667) );
  XOR U7339 ( .A(n5667), .B(key[489]), .Z(n5278) );
  XOR U7340 ( .A(n5339), .B(n5278), .Z(n5279) );
  XNOR U7341 ( .A(\w3[2][113] ), .B(n5279), .Z(\w1[3][105] ) );
  XOR U7342 ( .A(\w3[2][107] ), .B(\w3[2][99] ), .Z(n5281) );
  XNOR U7343 ( .A(\w3[2][98] ), .B(\w3[2][122] ), .Z(n5672) );
  XOR U7344 ( .A(n5672), .B(key[490]), .Z(n5280) );
  XNOR U7345 ( .A(n5281), .B(n5280), .Z(n5282) );
  XOR U7346 ( .A(\w3[2][114] ), .B(n5282), .Z(\w1[3][106] ) );
  XNOR U7347 ( .A(\w3[2][99] ), .B(\w3[2][123] ), .Z(n5676) );
  XOR U7348 ( .A(\w3[2][108] ), .B(n5676), .Z(n5283) );
  XOR U7349 ( .A(\w3[2][104] ), .B(n5283), .Z(n5309) );
  XNOR U7350 ( .A(n5309), .B(key[491]), .Z(n5285) );
  IV U7351 ( .A(\w3[2][100] ), .Z(n5348) );
  XOR U7352 ( .A(\w3[2][96] ), .B(n5348), .Z(n5680) );
  XOR U7353 ( .A(\w3[2][115] ), .B(n5680), .Z(n5284) );
  XNOR U7354 ( .A(n5285), .B(n5284), .Z(\w1[3][107] ) );
  XOR U7355 ( .A(\w3[2][100] ), .B(\w3[2][104] ), .Z(n5287) );
  XNOR U7356 ( .A(\w3[2][124] ), .B(\w3[2][109] ), .Z(n5286) );
  XOR U7357 ( .A(n5287), .B(n5286), .Z(n5312) );
  XNOR U7358 ( .A(n5312), .B(key[492]), .Z(n5290) );
  XNOR U7359 ( .A(\w3[2][116] ), .B(n5288), .Z(n5289) );
  XNOR U7360 ( .A(n5290), .B(n5289), .Z(\w1[3][108] ) );
  XNOR U7361 ( .A(\w3[2][125] ), .B(\w3[2][101] ), .Z(n5315) );
  XNOR U7362 ( .A(n5315), .B(key[493]), .Z(n5292) );
  XNOR U7363 ( .A(\w3[2][102] ), .B(\w3[2][110] ), .Z(n5291) );
  XNOR U7364 ( .A(n5292), .B(n5291), .Z(n5293) );
  XOR U7365 ( .A(\w3[2][117] ), .B(n5293), .Z(\w1[3][109] ) );
  IV U7366 ( .A(\w3[2][18] ), .Z(n5399) );
  XNOR U7367 ( .A(\w3[2][11] ), .B(n5399), .Z(n5295) );
  XNOR U7368 ( .A(\w3[2][2] ), .B(\w3[2][26] ), .Z(n5381) );
  XOR U7369 ( .A(n5381), .B(key[394]), .Z(n5294) );
  XNOR U7370 ( .A(n5295), .B(n5294), .Z(n5296) );
  XOR U7371 ( .A(\w3[2][3] ), .B(n5296), .Z(\w1[3][10] ) );
  XOR U7372 ( .A(\w3[2][111] ), .B(\w3[2][104] ), .Z(n5323) );
  XOR U7373 ( .A(n5297), .B(n5323), .Z(n5319) );
  XNOR U7374 ( .A(n5319), .B(key[494]), .Z(n5300) );
  XNOR U7375 ( .A(\w3[2][118] ), .B(n5298), .Z(n5299) );
  XNOR U7376 ( .A(n5300), .B(n5299), .Z(\w1[3][110] ) );
  XOR U7377 ( .A(\w3[2][127] ), .B(\w3[2][103] ), .Z(n5322) );
  XOR U7378 ( .A(n5322), .B(key[495]), .Z(n5302) );
  XNOR U7379 ( .A(\w3[2][96] ), .B(\w3[2][104] ), .Z(n5328) );
  XOR U7380 ( .A(\w3[2][119] ), .B(n5328), .Z(n5301) );
  XNOR U7381 ( .A(n5302), .B(n5301), .Z(\w1[3][111] ) );
  XNOR U7382 ( .A(\w3[2][105] ), .B(\w3[2][113] ), .Z(n5671) );
  XNOR U7383 ( .A(n5671), .B(key[496]), .Z(n5304) );
  XNOR U7384 ( .A(n5341), .B(n5328), .Z(n5303) );
  XNOR U7385 ( .A(n5304), .B(n5303), .Z(\w1[3][112] ) );
  XNOR U7386 ( .A(\w3[2][106] ), .B(\w3[2][114] ), .Z(n5675) );
  XNOR U7387 ( .A(n5675), .B(key[497]), .Z(n5306) );
  XOR U7388 ( .A(\w3[2][105] ), .B(n5667), .Z(n5305) );
  XNOR U7389 ( .A(n5306), .B(n5305), .Z(\w1[3][113] ) );
  XNOR U7390 ( .A(\w3[2][107] ), .B(\w3[2][115] ), .Z(n5343) );
  XNOR U7391 ( .A(n5343), .B(key[498]), .Z(n5308) );
  XNOR U7392 ( .A(n5339), .B(\w3[2][122] ), .Z(n5307) );
  XNOR U7393 ( .A(n5308), .B(n5307), .Z(\w1[3][114] ) );
  XOR U7394 ( .A(\w3[2][116] ), .B(n5332), .Z(n5344) );
  XNOR U7395 ( .A(n5344), .B(key[499]), .Z(n5311) );
  XOR U7396 ( .A(\w3[2][107] ), .B(n5309), .Z(n5310) );
  XNOR U7397 ( .A(n5311), .B(n5310), .Z(\w1[3][115] ) );
  XOR U7398 ( .A(\w3[2][117] ), .B(n5332), .Z(n5347) );
  XNOR U7399 ( .A(n5347), .B(key[500]), .Z(n5314) );
  XOR U7400 ( .A(\w3[2][108] ), .B(n5312), .Z(n5313) );
  XNOR U7401 ( .A(n5314), .B(n5313), .Z(\w1[3][116] ) );
  XNOR U7402 ( .A(n5315), .B(key[501]), .Z(n5318) );
  XNOR U7403 ( .A(\w3[2][109] ), .B(n5316), .Z(n5317) );
  XNOR U7404 ( .A(n5318), .B(n5317), .Z(\w1[3][117] ) );
  XOR U7405 ( .A(\w3[2][119] ), .B(n5332), .Z(n5356) );
  XNOR U7406 ( .A(n5356), .B(key[502]), .Z(n5321) );
  XOR U7407 ( .A(\w3[2][110] ), .B(n5319), .Z(n5320) );
  XNOR U7408 ( .A(n5321), .B(n5320), .Z(\w1[3][118] ) );
  XOR U7409 ( .A(n5322), .B(key[503]), .Z(n5325) );
  XNOR U7410 ( .A(\w3[2][112] ), .B(n5323), .Z(n5324) );
  XNOR U7411 ( .A(n5325), .B(n5324), .Z(\w1[3][119] ) );
  XNOR U7412 ( .A(\w3[2][3] ), .B(\w3[2][27] ), .Z(n5420) );
  XNOR U7413 ( .A(n5380), .B(key[395]), .Z(n5327) );
  XNOR U7414 ( .A(\w3[2][0] ), .B(\w3[2][4] ), .Z(n5452) );
  XOR U7415 ( .A(\w3[2][19] ), .B(n5452), .Z(n5326) );
  XNOR U7416 ( .A(n5327), .B(n5326), .Z(\w1[3][11] ) );
  XNOR U7417 ( .A(n5328), .B(key[504]), .Z(n5330) );
  XNOR U7418 ( .A(\w3[2][113] ), .B(\w3[2][121] ), .Z(n5329) );
  XNOR U7419 ( .A(n5330), .B(n5329), .Z(n5331) );
  XNOR U7420 ( .A(n5332), .B(n5331), .Z(\w1[3][120] ) );
  XNOR U7421 ( .A(n5671), .B(key[505]), .Z(n5334) );
  XNOR U7422 ( .A(\w3[2][114] ), .B(\w3[2][122] ), .Z(n5333) );
  XNOR U7423 ( .A(n5334), .B(n5333), .Z(n5335) );
  XNOR U7424 ( .A(n5336), .B(n5335), .Z(\w1[3][121] ) );
  XOR U7425 ( .A(\w3[2][123] ), .B(key[506]), .Z(n5338) );
  XNOR U7426 ( .A(\w3[2][114] ), .B(\w3[2][115] ), .Z(n5337) );
  XNOR U7427 ( .A(n5338), .B(n5337), .Z(n5340) );
  XOR U7428 ( .A(n5340), .B(n5339), .Z(\w1[3][122] ) );
  XOR U7429 ( .A(\w3[2][124] ), .B(n5341), .Z(n5342) );
  XOR U7430 ( .A(n5343), .B(n5342), .Z(n5679) );
  XOR U7431 ( .A(n5679), .B(key[507]), .Z(n5346) );
  XOR U7432 ( .A(\w3[2][99] ), .B(n5344), .Z(n5345) );
  XNOR U7433 ( .A(n5346), .B(n5345), .Z(\w1[3][123] ) );
  XNOR U7434 ( .A(n5347), .B(key[508]), .Z(n5351) );
  XNOR U7435 ( .A(n5349), .B(n5348), .Z(n5350) );
  XNOR U7436 ( .A(n5351), .B(n5350), .Z(\w1[3][124] ) );
  XOR U7437 ( .A(\w3[2][118] ), .B(key[509]), .Z(n5354) );
  XOR U7438 ( .A(n5352), .B(\w3[2][126] ), .Z(n5353) );
  XNOR U7439 ( .A(n5354), .B(n5353), .Z(n5355) );
  XOR U7440 ( .A(\w3[2][101] ), .B(n5355), .Z(\w1[3][125] ) );
  XNOR U7441 ( .A(n5356), .B(key[510]), .Z(n5359) );
  XOR U7442 ( .A(\w3[2][102] ), .B(n5357), .Z(n5358) );
  XNOR U7443 ( .A(n5359), .B(n5358), .Z(\w1[3][126] ) );
  XNOR U7444 ( .A(n5668), .B(key[511]), .Z(n5362) );
  XOR U7445 ( .A(\w3[2][103] ), .B(n5360), .Z(n5361) );
  XNOR U7446 ( .A(n5362), .B(n5361), .Z(\w1[3][127] ) );
  XOR U7447 ( .A(\w3[2][13] ), .B(\w3[2][28] ), .Z(n5364) );
  XNOR U7448 ( .A(\w3[2][8] ), .B(\w3[2][4] ), .Z(n5363) );
  XOR U7449 ( .A(n5364), .B(n5363), .Z(n5384) );
  XNOR U7450 ( .A(n5384), .B(key[396]), .Z(n5366) );
  XNOR U7451 ( .A(\w3[2][0] ), .B(\w3[2][5] ), .Z(n5487) );
  XOR U7452 ( .A(\w3[2][20] ), .B(n5487), .Z(n5365) );
  XNOR U7453 ( .A(n5366), .B(n5365), .Z(\w1[3][12] ) );
  IV U7454 ( .A(\w3[2][6] ), .Z(n5426) );
  XNOR U7455 ( .A(\w3[2][14] ), .B(n5426), .Z(n5368) );
  XNOR U7456 ( .A(\w3[2][5] ), .B(\w3[2][29] ), .Z(n5387) );
  XOR U7457 ( .A(n5387), .B(key[397]), .Z(n5367) );
  XNOR U7458 ( .A(n5368), .B(n5367), .Z(n5369) );
  XOR U7459 ( .A(\w3[2][21] ), .B(n5369), .Z(\w1[3][13] ) );
  IV U7460 ( .A(\w3[2][30] ), .Z(n5564) );
  XOR U7461 ( .A(\w3[2][6] ), .B(n5564), .Z(n5529) );
  XOR U7462 ( .A(\w3[2][8] ), .B(\w3[2][15] ), .Z(n5390) );
  XNOR U7463 ( .A(n5529), .B(n5390), .Z(n5388) );
  XOR U7464 ( .A(n5388), .B(key[398]), .Z(n5371) );
  XNOR U7465 ( .A(\w3[2][0] ), .B(\w3[2][7] ), .Z(n5565) );
  XOR U7466 ( .A(\w3[2][22] ), .B(n5565), .Z(n5370) );
  XNOR U7467 ( .A(n5371), .B(n5370), .Z(\w1[3][14] ) );
  XNOR U7468 ( .A(\w3[2][7] ), .B(\w3[2][31] ), .Z(n5389) );
  XNOR U7469 ( .A(n5389), .B(key[399]), .Z(n5373) );
  XOR U7470 ( .A(\w3[2][8] ), .B(\w3[2][0] ), .Z(n5393) );
  XNOR U7471 ( .A(\w3[2][23] ), .B(n5393), .Z(n5372) );
  XNOR U7472 ( .A(n5373), .B(n5372), .Z(\w1[3][15] ) );
  XNOR U7473 ( .A(\w3[2][17] ), .B(\w3[2][9] ), .Z(n5395) );
  XNOR U7474 ( .A(n5395), .B(key[400]), .Z(n5375) );
  XNOR U7475 ( .A(\w3[2][24] ), .B(n5393), .Z(n5374) );
  XNOR U7476 ( .A(n5375), .B(n5374), .Z(\w1[3][16] ) );
  XNOR U7477 ( .A(\w3[2][18] ), .B(\w3[2][10] ), .Z(n5419) );
  XNOR U7478 ( .A(n5419), .B(key[401]), .Z(n5377) );
  IV U7479 ( .A(\w3[2][9] ), .Z(n5636) );
  XNOR U7480 ( .A(n5686), .B(n5636), .Z(n5376) );
  XNOR U7481 ( .A(n5377), .B(n5376), .Z(\w1[3][17] ) );
  IV U7482 ( .A(\w3[2][19] ), .Z(n5400) );
  XOR U7483 ( .A(\w3[2][11] ), .B(n5400), .Z(n5405) );
  XNOR U7484 ( .A(n5405), .B(key[402]), .Z(n5379) );
  XOR U7485 ( .A(n5381), .B(\w3[2][10] ), .Z(n5378) );
  XNOR U7486 ( .A(n5379), .B(n5378), .Z(\w1[3][18] ) );
  XOR U7487 ( .A(n5394), .B(\w3[2][20] ), .Z(n5406) );
  XNOR U7488 ( .A(n5395), .B(key[385]), .Z(n5383) );
  XOR U7489 ( .A(\w3[2][25] ), .B(n5381), .Z(n5382) );
  XNOR U7490 ( .A(n5383), .B(n5382), .Z(\w1[3][1] ) );
  IV U7491 ( .A(\w3[2][21] ), .Z(n5414) );
  XOR U7492 ( .A(\w3[2][16] ), .B(n5414), .Z(n5411) );
  XNOR U7493 ( .A(n5411), .B(key[404]), .Z(n5386) );
  XOR U7494 ( .A(\w3[2][12] ), .B(n5384), .Z(n5385) );
  XNOR U7495 ( .A(n5386), .B(n5385), .Z(\w1[3][20] ) );
  IV U7496 ( .A(\w3[2][22] ), .Z(n5415) );
  XOR U7497 ( .A(\w3[2][14] ), .B(n5415), .Z(n5424) );
  XOR U7498 ( .A(n5394), .B(\w3[2][23] ), .Z(n5425) );
  XNOR U7499 ( .A(n5389), .B(key[407]), .Z(n5392) );
  XNOR U7500 ( .A(\w3[2][16] ), .B(n5390), .Z(n5391) );
  XNOR U7501 ( .A(n5392), .B(n5391), .Z(\w1[3][23] ) );
  XNOR U7502 ( .A(n5395), .B(key[409]), .Z(n5397) );
  XNOR U7503 ( .A(\w3[2][1] ), .B(\w3[2][26] ), .Z(n5396) );
  XNOR U7504 ( .A(n5397), .B(n5396), .Z(n5398) );
  XNOR U7505 ( .A(n5399), .B(n5398), .Z(\w1[3][25] ) );
  XNOR U7506 ( .A(n5419), .B(key[410]), .Z(n5402) );
  XOR U7507 ( .A(\w3[2][2] ), .B(n5400), .Z(n5401) );
  XNOR U7508 ( .A(n5402), .B(n5401), .Z(n5403) );
  XOR U7509 ( .A(\w3[2][27] ), .B(n5403), .Z(\w1[3][26] ) );
  IV U7510 ( .A(\w3[2][24] ), .Z(n5423) );
  XOR U7511 ( .A(n5423), .B(\w3[2][28] ), .Z(n5404) );
  XOR U7512 ( .A(n5405), .B(n5404), .Z(n5451) );
  XOR U7513 ( .A(n5451), .B(key[411]), .Z(n5408) );
  XOR U7514 ( .A(\w3[2][3] ), .B(n5406), .Z(n5407) );
  XNOR U7515 ( .A(n5408), .B(n5407), .Z(\w1[3][27] ) );
  XOR U7516 ( .A(\w3[2][20] ), .B(\w3[2][29] ), .Z(n5410) );
  XOR U7517 ( .A(n5423), .B(\w3[2][12] ), .Z(n5409) );
  XOR U7518 ( .A(n5410), .B(n5409), .Z(n5486) );
  XNOR U7519 ( .A(n5486), .B(key[412]), .Z(n5413) );
  XOR U7520 ( .A(\w3[2][4] ), .B(n5411), .Z(n5412) );
  XNOR U7521 ( .A(n5413), .B(n5412), .Z(\w1[3][28] ) );
  XOR U7522 ( .A(\w3[2][13] ), .B(n5414), .Z(n5528) );
  XNOR U7523 ( .A(n5528), .B(key[413]), .Z(n5417) );
  XNOR U7524 ( .A(n5415), .B(n5564), .Z(n5416) );
  XNOR U7525 ( .A(n5417), .B(n5416), .Z(n5418) );
  XOR U7526 ( .A(\w3[2][5] ), .B(n5418), .Z(\w1[3][29] ) );
  XNOR U7527 ( .A(n5419), .B(key[386]), .Z(n5422) );
  XOR U7528 ( .A(\w3[2][26] ), .B(n5420), .Z(n5421) );
  XNOR U7529 ( .A(n5422), .B(n5421), .Z(\w1[3][2] ) );
  XOR U7530 ( .A(n5423), .B(\w3[2][31] ), .Z(n5600) );
  XNOR U7531 ( .A(n5424), .B(n5600), .Z(n5563) );
  XNOR U7532 ( .A(n5563), .B(key[414]), .Z(n5428) );
  XNOR U7533 ( .A(n5426), .B(n5425), .Z(n5427) );
  XNOR U7534 ( .A(n5428), .B(n5427), .Z(\w1[3][30] ) );
  XNOR U7535 ( .A(\w3[2][15] ), .B(\w3[2][23] ), .Z(n5599) );
  XNOR U7536 ( .A(n5599), .B(key[415]), .Z(n5430) );
  XOR U7537 ( .A(n5639), .B(\w3[2][7] ), .Z(n5429) );
  XNOR U7538 ( .A(n5430), .B(n5429), .Z(\w1[3][31] ) );
  XOR U7539 ( .A(\w3[2][33] ), .B(\w3[2][57] ), .Z(n5483) );
  XOR U7540 ( .A(n5483), .B(key[416]), .Z(n5432) );
  XNOR U7541 ( .A(\w3[2][48] ), .B(\w3[2][56] ), .Z(n5545) );
  XOR U7542 ( .A(n5545), .B(\w3[2][40] ), .Z(n5431) );
  XNOR U7543 ( .A(n5432), .B(n5431), .Z(\w1[3][32] ) );
  XNOR U7544 ( .A(\w3[2][34] ), .B(\w3[2][58] ), .Z(n5491) );
  XOR U7545 ( .A(\w3[2][57] ), .B(\w3[2][49] ), .Z(n5509) );
  XNOR U7546 ( .A(n5509), .B(key[417]), .Z(n5433) );
  XNOR U7547 ( .A(n5491), .B(n5433), .Z(n5434) );
  XNOR U7548 ( .A(\w3[2][41] ), .B(n5434), .Z(\w1[3][33] ) );
  XNOR U7549 ( .A(n5461), .B(key[418]), .Z(n5436) );
  XNOR U7550 ( .A(\w3[2][50] ), .B(\w3[2][42] ), .Z(n5519) );
  XOR U7551 ( .A(\w3[2][58] ), .B(n5519), .Z(n5435) );
  XNOR U7552 ( .A(n5436), .B(n5435), .Z(\w1[3][34] ) );
  XOR U7553 ( .A(\w3[2][36] ), .B(\w3[2][32] ), .Z(n5463) );
  XOR U7554 ( .A(n5463), .B(key[419]), .Z(n5439) );
  IV U7555 ( .A(\w3[2][51] ), .Z(n5518) );
  XOR U7556 ( .A(\w3[2][43] ), .B(n5518), .Z(n5490) );
  XOR U7557 ( .A(\w3[2][56] ), .B(n5490), .Z(n5437) );
  XNOR U7558 ( .A(\w3[2][60] ), .B(n5437), .Z(n5524) );
  XNOR U7559 ( .A(\w3[2][59] ), .B(n5524), .Z(n5438) );
  XNOR U7560 ( .A(n5439), .B(n5438), .Z(\w1[3][35] ) );
  XOR U7561 ( .A(\w3[2][32] ), .B(\w3[2][37] ), .Z(n5469) );
  XOR U7562 ( .A(\w3[2][52] ), .B(\w3[2][61] ), .Z(n5441) );
  XNOR U7563 ( .A(\w3[2][56] ), .B(\w3[2][44] ), .Z(n5440) );
  XOR U7564 ( .A(n5441), .B(n5440), .Z(n5533) );
  XOR U7565 ( .A(n5533), .B(key[420]), .Z(n5442) );
  XOR U7566 ( .A(n5469), .B(n5442), .Z(n5443) );
  XNOR U7567 ( .A(\w3[2][60] ), .B(n5443), .Z(\w1[3][36] ) );
  XNOR U7568 ( .A(\w3[2][38] ), .B(\w3[2][62] ), .Z(n5475) );
  XNOR U7569 ( .A(n5475), .B(key[421]), .Z(n5445) );
  IV U7570 ( .A(\w3[2][45] ), .Z(n5498) );
  XOR U7571 ( .A(\w3[2][53] ), .B(n5498), .Z(n5536) );
  XOR U7572 ( .A(\w3[2][61] ), .B(n5536), .Z(n5444) );
  XNOR U7573 ( .A(n5445), .B(n5444), .Z(\w1[3][37] ) );
  XOR U7574 ( .A(\w3[2][32] ), .B(\w3[2][39] ), .Z(n5476) );
  XOR U7575 ( .A(n5476), .B(key[422]), .Z(n5447) );
  XNOR U7576 ( .A(\w3[2][46] ), .B(\w3[2][54] ), .Z(n5497) );
  XOR U7577 ( .A(\w3[2][56] ), .B(\w3[2][63] ), .Z(n5448) );
  XOR U7578 ( .A(n5497), .B(n5448), .Z(n5541) );
  XOR U7579 ( .A(\w3[2][62] ), .B(n5541), .Z(n5446) );
  XNOR U7580 ( .A(n5447), .B(n5446), .Z(\w1[3][38] ) );
  XNOR U7581 ( .A(\w3[2][55] ), .B(\w3[2][47] ), .Z(n5544) );
  XNOR U7582 ( .A(n5544), .B(key[423]), .Z(n5450) );
  XNOR U7583 ( .A(\w3[2][32] ), .B(n5448), .Z(n5449) );
  XNOR U7584 ( .A(n5450), .B(n5449), .Z(\w1[3][39] ) );
  XOR U7585 ( .A(n5451), .B(key[387]), .Z(n5454) );
  XOR U7586 ( .A(n5452), .B(\w3[2][27] ), .Z(n5453) );
  XNOR U7587 ( .A(n5454), .B(n5453), .Z(\w1[3][3] ) );
  IV U7588 ( .A(\w3[2][33] ), .Z(n5514) );
  XOR U7589 ( .A(\w3[2][42] ), .B(key[425]), .Z(n5456) );
  XNOR U7590 ( .A(n5509), .B(\w3[2][34] ), .Z(n5455) );
  XNOR U7591 ( .A(n5456), .B(n5455), .Z(n5457) );
  XNOR U7592 ( .A(n5514), .B(n5457), .Z(\w1[3][41] ) );
  XOR U7593 ( .A(\w3[2][43] ), .B(key[426]), .Z(n5459) );
  IV U7594 ( .A(\w3[2][35] ), .Z(n5525) );
  XOR U7595 ( .A(\w3[2][50] ), .B(n5525), .Z(n5458) );
  XNOR U7596 ( .A(n5459), .B(n5458), .Z(n5460) );
  XNOR U7597 ( .A(n5460), .B(n5491), .Z(\w1[3][42] ) );
  IV U7598 ( .A(\w3[2][40] ), .Z(n5466) );
  XNOR U7599 ( .A(n5466), .B(n5461), .Z(n5462) );
  XOR U7600 ( .A(\w3[2][44] ), .B(n5462), .Z(n5492) );
  XNOR U7601 ( .A(n5492), .B(key[427]), .Z(n5465) );
  XNOR U7602 ( .A(\w3[2][51] ), .B(n5463), .Z(n5464) );
  XNOR U7603 ( .A(n5465), .B(n5464), .Z(\w1[3][43] ) );
  XOR U7604 ( .A(\w3[2][36] ), .B(\w3[2][45] ), .Z(n5468) );
  XOR U7605 ( .A(n5466), .B(\w3[2][60] ), .Z(n5467) );
  XOR U7606 ( .A(n5468), .B(n5467), .Z(n5493) );
  XNOR U7607 ( .A(n5493), .B(key[428]), .Z(n5471) );
  XNOR U7608 ( .A(\w3[2][52] ), .B(n5469), .Z(n5470) );
  XNOR U7609 ( .A(n5471), .B(n5470), .Z(\w1[3][44] ) );
  XNOR U7610 ( .A(\w3[2][61] ), .B(\w3[2][37] ), .Z(n5496) );
  XNOR U7611 ( .A(n5496), .B(key[429]), .Z(n5473) );
  XNOR U7612 ( .A(\w3[2][38] ), .B(\w3[2][46] ), .Z(n5472) );
  XNOR U7613 ( .A(n5473), .B(n5472), .Z(n5474) );
  XOR U7614 ( .A(\w3[2][53] ), .B(n5474), .Z(\w1[3][45] ) );
  XOR U7615 ( .A(\w3[2][40] ), .B(\w3[2][47] ), .Z(n5505) );
  XOR U7616 ( .A(n5475), .B(n5505), .Z(n5501) );
  XNOR U7617 ( .A(n5501), .B(key[430]), .Z(n5478) );
  XNOR U7618 ( .A(\w3[2][54] ), .B(n5476), .Z(n5477) );
  XNOR U7619 ( .A(n5478), .B(n5477), .Z(\w1[3][46] ) );
  XOR U7620 ( .A(\w3[2][63] ), .B(\w3[2][39] ), .Z(n5504) );
  XOR U7621 ( .A(n5504), .B(key[431]), .Z(n5480) );
  XNOR U7622 ( .A(\w3[2][40] ), .B(\w3[2][32] ), .Z(n5508) );
  XOR U7623 ( .A(\w3[2][55] ), .B(n5508), .Z(n5479) );
  XNOR U7624 ( .A(n5480), .B(n5479), .Z(\w1[3][47] ) );
  XNOR U7625 ( .A(\w3[2][41] ), .B(\w3[2][49] ), .Z(n5513) );
  XNOR U7626 ( .A(n5513), .B(key[432]), .Z(n5482) );
  XOR U7627 ( .A(\w3[2][56] ), .B(n5508), .Z(n5481) );
  XNOR U7628 ( .A(n5482), .B(n5481), .Z(\w1[3][48] ) );
  XNOR U7629 ( .A(n5519), .B(key[433]), .Z(n5485) );
  XNOR U7630 ( .A(n5483), .B(\w3[2][41] ), .Z(n5484) );
  XNOR U7631 ( .A(n5485), .B(n5484), .Z(\w1[3][49] ) );
  XNOR U7632 ( .A(n5486), .B(key[388]), .Z(n5489) );
  XOR U7633 ( .A(n5487), .B(\w3[2][28] ), .Z(n5488) );
  XNOR U7634 ( .A(n5489), .B(n5488), .Z(\w1[3][4] ) );
  IV U7635 ( .A(\w3[2][48] ), .Z(n5510) );
  XOR U7636 ( .A(n5510), .B(\w3[2][52] ), .Z(n5523) );
  XNOR U7637 ( .A(n5532), .B(key[436]), .Z(n5495) );
  XOR U7638 ( .A(\w3[2][44] ), .B(n5493), .Z(n5494) );
  XNOR U7639 ( .A(n5495), .B(n5494), .Z(\w1[3][52] ) );
  XNOR U7640 ( .A(n5496), .B(key[437]), .Z(n5500) );
  XNOR U7641 ( .A(n5498), .B(n5497), .Z(n5499) );
  XNOR U7642 ( .A(n5500), .B(n5499), .Z(\w1[3][53] ) );
  XOR U7643 ( .A(n5510), .B(\w3[2][55] ), .Z(n5540) );
  XNOR U7644 ( .A(n5540), .B(key[438]), .Z(n5503) );
  XOR U7645 ( .A(\w3[2][46] ), .B(n5501), .Z(n5502) );
  XNOR U7646 ( .A(n5503), .B(n5502), .Z(\w1[3][54] ) );
  XOR U7647 ( .A(n5504), .B(key[439]), .Z(n5507) );
  XNOR U7648 ( .A(\w3[2][48] ), .B(n5505), .Z(n5506) );
  XNOR U7649 ( .A(n5507), .B(n5506), .Z(\w1[3][55] ) );
  XNOR U7650 ( .A(n5508), .B(key[440]), .Z(n5512) );
  XOR U7651 ( .A(n5510), .B(n5509), .Z(n5511) );
  XNOR U7652 ( .A(n5512), .B(n5511), .Z(\w1[3][56] ) );
  XNOR U7653 ( .A(n5513), .B(key[441]), .Z(n5516) );
  XOR U7654 ( .A(n5514), .B(\w3[2][50] ), .Z(n5515) );
  XNOR U7655 ( .A(n5516), .B(n5515), .Z(n5517) );
  XOR U7656 ( .A(\w3[2][58] ), .B(n5517), .Z(\w1[3][57] ) );
  XNOR U7657 ( .A(n5518), .B(key[442]), .Z(n5521) );
  XOR U7658 ( .A(n5519), .B(\w3[2][59] ), .Z(n5520) );
  XNOR U7659 ( .A(n5521), .B(n5520), .Z(n5522) );
  XOR U7660 ( .A(\w3[2][34] ), .B(n5522), .Z(\w1[3][58] ) );
  XNOR U7661 ( .A(n5523), .B(key[443]), .Z(n5527) );
  XOR U7662 ( .A(n5525), .B(n5524), .Z(n5526) );
  XNOR U7663 ( .A(n5527), .B(n5526), .Z(\w1[3][59] ) );
  XNOR U7664 ( .A(n5528), .B(key[389]), .Z(n5531) );
  XOR U7665 ( .A(\w3[2][29] ), .B(n5529), .Z(n5530) );
  XNOR U7666 ( .A(n5531), .B(n5530), .Z(\w1[3][5] ) );
  XNOR U7667 ( .A(n5532), .B(key[444]), .Z(n5535) );
  XOR U7668 ( .A(\w3[2][36] ), .B(n5533), .Z(n5534) );
  XNOR U7669 ( .A(n5535), .B(n5534), .Z(\w1[3][60] ) );
  XOR U7670 ( .A(\w3[2][54] ), .B(key[445]), .Z(n5538) );
  XOR U7671 ( .A(n5536), .B(\w3[2][62] ), .Z(n5537) );
  XNOR U7672 ( .A(n5538), .B(n5537), .Z(n5539) );
  XOR U7673 ( .A(\w3[2][37] ), .B(n5539), .Z(\w1[3][61] ) );
  XNOR U7674 ( .A(n5540), .B(key[446]), .Z(n5543) );
  XOR U7675 ( .A(\w3[2][38] ), .B(n5541), .Z(n5542) );
  XNOR U7676 ( .A(n5543), .B(n5542), .Z(\w1[3][62] ) );
  XNOR U7677 ( .A(n5544), .B(key[447]), .Z(n5547) );
  XOR U7678 ( .A(n5545), .B(\w3[2][39] ), .Z(n5546) );
  XNOR U7679 ( .A(n5547), .B(n5546), .Z(\w1[3][63] ) );
  XOR U7680 ( .A(\w3[2][65] ), .B(\w3[2][89] ), .Z(n5605) );
  XOR U7681 ( .A(n5605), .B(key[448]), .Z(n5549) );
  XNOR U7682 ( .A(\w3[2][80] ), .B(\w3[2][88] ), .Z(n5664) );
  XOR U7683 ( .A(n5664), .B(\w3[2][72] ), .Z(n5548) );
  XNOR U7684 ( .A(n5549), .B(n5548), .Z(\w1[3][64] ) );
  XNOR U7685 ( .A(\w3[2][66] ), .B(\w3[2][90] ), .Z(n5609) );
  XOR U7686 ( .A(\w3[2][89] ), .B(\w3[2][81] ), .Z(n5627) );
  XNOR U7687 ( .A(n5627), .B(key[449]), .Z(n5550) );
  XNOR U7688 ( .A(n5609), .B(n5550), .Z(n5551) );
  XNOR U7689 ( .A(\w3[2][73] ), .B(n5551), .Z(\w1[3][65] ) );
  XNOR U7690 ( .A(n5579), .B(key[450]), .Z(n5553) );
  XNOR U7691 ( .A(\w3[2][82] ), .B(\w3[2][74] ), .Z(n5642) );
  XOR U7692 ( .A(\w3[2][90] ), .B(n5642), .Z(n5552) );
  XNOR U7693 ( .A(n5553), .B(n5552), .Z(\w1[3][66] ) );
  XOR U7694 ( .A(\w3[2][68] ), .B(\w3[2][64] ), .Z(n5581) );
  XOR U7695 ( .A(n5581), .B(key[451]), .Z(n5556) );
  IV U7696 ( .A(\w3[2][83] ), .Z(n5641) );
  XOR U7697 ( .A(\w3[2][75] ), .B(n5641), .Z(n5608) );
  XOR U7698 ( .A(\w3[2][88] ), .B(n5608), .Z(n5554) );
  XNOR U7699 ( .A(\w3[2][92] ), .B(n5554), .Z(n5647) );
  XNOR U7700 ( .A(\w3[2][91] ), .B(n5647), .Z(n5555) );
  XNOR U7701 ( .A(n5556), .B(n5555), .Z(\w1[3][67] ) );
  XOR U7702 ( .A(\w3[2][64] ), .B(\w3[2][69] ), .Z(n5587) );
  XOR U7703 ( .A(\w3[2][84] ), .B(\w3[2][93] ), .Z(n5558) );
  XNOR U7704 ( .A(\w3[2][88] ), .B(\w3[2][76] ), .Z(n5557) );
  XOR U7705 ( .A(n5558), .B(n5557), .Z(n5652) );
  XOR U7706 ( .A(n5652), .B(key[452]), .Z(n5559) );
  XOR U7707 ( .A(n5587), .B(n5559), .Z(n5560) );
  XNOR U7708 ( .A(\w3[2][92] ), .B(n5560), .Z(\w1[3][68] ) );
  XNOR U7709 ( .A(\w3[2][70] ), .B(\w3[2][94] ), .Z(n5593) );
  XNOR U7710 ( .A(n5593), .B(key[453]), .Z(n5562) );
  IV U7711 ( .A(\w3[2][77] ), .Z(n5616) );
  XOR U7712 ( .A(\w3[2][85] ), .B(n5616), .Z(n5655) );
  XOR U7713 ( .A(\w3[2][93] ), .B(n5655), .Z(n5561) );
  XNOR U7714 ( .A(n5562), .B(n5561), .Z(\w1[3][69] ) );
  XNOR U7715 ( .A(n5563), .B(key[390]), .Z(n5567) );
  XNOR U7716 ( .A(n5565), .B(n5564), .Z(n5566) );
  XNOR U7717 ( .A(n5567), .B(n5566), .Z(\w1[3][6] ) );
  XOR U7718 ( .A(\w3[2][64] ), .B(\w3[2][71] ), .Z(n5594) );
  XOR U7719 ( .A(n5594), .B(key[454]), .Z(n5569) );
  XNOR U7720 ( .A(\w3[2][88] ), .B(\w3[2][95] ), .Z(n5570) );
  XOR U7721 ( .A(\w3[2][78] ), .B(\w3[2][86] ), .Z(n5615) );
  XOR U7722 ( .A(n5570), .B(n5615), .Z(n5660) );
  XOR U7723 ( .A(\w3[2][94] ), .B(n5660), .Z(n5568) );
  XNOR U7724 ( .A(n5569), .B(n5568), .Z(\w1[3][70] ) );
  XNOR U7725 ( .A(\w3[2][79] ), .B(\w3[2][87] ), .Z(n5663) );
  XNOR U7726 ( .A(n5663), .B(key[455]), .Z(n5572) );
  XOR U7727 ( .A(\w3[2][64] ), .B(n5570), .Z(n5571) );
  XNOR U7728 ( .A(n5572), .B(n5571), .Z(\w1[3][71] ) );
  IV U7729 ( .A(\w3[2][65] ), .Z(n5632) );
  XOR U7730 ( .A(\w3[2][74] ), .B(key[457]), .Z(n5574) );
  XNOR U7731 ( .A(n5627), .B(\w3[2][66] ), .Z(n5573) );
  XNOR U7732 ( .A(n5574), .B(n5573), .Z(n5575) );
  XNOR U7733 ( .A(n5632), .B(n5575), .Z(\w1[3][73] ) );
  XOR U7734 ( .A(\w3[2][75] ), .B(key[458]), .Z(n5577) );
  IV U7735 ( .A(\w3[2][67] ), .Z(n5648) );
  XOR U7736 ( .A(\w3[2][82] ), .B(n5648), .Z(n5576) );
  XNOR U7737 ( .A(n5577), .B(n5576), .Z(n5578) );
  XNOR U7738 ( .A(n5578), .B(n5609), .Z(\w1[3][74] ) );
  IV U7739 ( .A(\w3[2][72] ), .Z(n5584) );
  XNOR U7740 ( .A(n5584), .B(n5579), .Z(n5580) );
  XOR U7741 ( .A(\w3[2][76] ), .B(n5580), .Z(n5610) );
  XNOR U7742 ( .A(n5610), .B(key[459]), .Z(n5583) );
  XNOR U7743 ( .A(\w3[2][83] ), .B(n5581), .Z(n5582) );
  XNOR U7744 ( .A(n5583), .B(n5582), .Z(\w1[3][75] ) );
  XOR U7745 ( .A(\w3[2][68] ), .B(\w3[2][77] ), .Z(n5586) );
  XOR U7746 ( .A(n5584), .B(\w3[2][92] ), .Z(n5585) );
  XOR U7747 ( .A(n5586), .B(n5585), .Z(n5611) );
  XNOR U7748 ( .A(n5611), .B(key[460]), .Z(n5589) );
  XNOR U7749 ( .A(\w3[2][84] ), .B(n5587), .Z(n5588) );
  XNOR U7750 ( .A(n5589), .B(n5588), .Z(\w1[3][76] ) );
  XNOR U7751 ( .A(\w3[2][93] ), .B(\w3[2][69] ), .Z(n5614) );
  XNOR U7752 ( .A(n5614), .B(key[461]), .Z(n5591) );
  XNOR U7753 ( .A(\w3[2][70] ), .B(\w3[2][78] ), .Z(n5590) );
  XNOR U7754 ( .A(n5591), .B(n5590), .Z(n5592) );
  XOR U7755 ( .A(\w3[2][85] ), .B(n5592), .Z(\w1[3][77] ) );
  XOR U7756 ( .A(\w3[2][72] ), .B(\w3[2][79] ), .Z(n5623) );
  XOR U7757 ( .A(n5593), .B(n5623), .Z(n5619) );
  XNOR U7758 ( .A(n5619), .B(key[462]), .Z(n5596) );
  XNOR U7759 ( .A(\w3[2][86] ), .B(n5594), .Z(n5595) );
  XNOR U7760 ( .A(n5596), .B(n5595), .Z(\w1[3][78] ) );
  XOR U7761 ( .A(\w3[2][95] ), .B(\w3[2][71] ), .Z(n5622) );
  XOR U7762 ( .A(n5622), .B(key[463]), .Z(n5598) );
  XNOR U7763 ( .A(\w3[2][72] ), .B(\w3[2][64] ), .Z(n5626) );
  XOR U7764 ( .A(\w3[2][87] ), .B(n5626), .Z(n5597) );
  XNOR U7765 ( .A(n5598), .B(n5597), .Z(\w1[3][79] ) );
  XNOR U7766 ( .A(n5599), .B(key[391]), .Z(n5602) );
  XOR U7767 ( .A(\w3[2][0] ), .B(n5600), .Z(n5601) );
  XNOR U7768 ( .A(n5602), .B(n5601), .Z(\w1[3][7] ) );
  XNOR U7769 ( .A(\w3[2][73] ), .B(\w3[2][81] ), .Z(n5631) );
  XNOR U7770 ( .A(n5631), .B(key[464]), .Z(n5604) );
  XOR U7771 ( .A(\w3[2][88] ), .B(n5626), .Z(n5603) );
  XNOR U7772 ( .A(n5604), .B(n5603), .Z(\w1[3][80] ) );
  XNOR U7773 ( .A(n5642), .B(key[465]), .Z(n5607) );
  XNOR U7774 ( .A(n5605), .B(\w3[2][73] ), .Z(n5606) );
  XNOR U7775 ( .A(n5607), .B(n5606), .Z(\w1[3][81] ) );
  IV U7776 ( .A(\w3[2][80] ), .Z(n5628) );
  XOR U7777 ( .A(n5628), .B(\w3[2][84] ), .Z(n5646) );
  XNOR U7778 ( .A(n5651), .B(key[468]), .Z(n5613) );
  XOR U7779 ( .A(\w3[2][76] ), .B(n5611), .Z(n5612) );
  XNOR U7780 ( .A(n5613), .B(n5612), .Z(\w1[3][84] ) );
  XNOR U7781 ( .A(n5614), .B(key[469]), .Z(n5618) );
  XOR U7782 ( .A(n5616), .B(n5615), .Z(n5617) );
  XNOR U7783 ( .A(n5618), .B(n5617), .Z(\w1[3][85] ) );
  XOR U7784 ( .A(n5628), .B(\w3[2][87] ), .Z(n5659) );
  XNOR U7785 ( .A(n5659), .B(key[470]), .Z(n5621) );
  XOR U7786 ( .A(\w3[2][78] ), .B(n5619), .Z(n5620) );
  XNOR U7787 ( .A(n5621), .B(n5620), .Z(\w1[3][86] ) );
  XOR U7788 ( .A(n5622), .B(key[471]), .Z(n5625) );
  XNOR U7789 ( .A(\w3[2][80] ), .B(n5623), .Z(n5624) );
  XNOR U7790 ( .A(n5625), .B(n5624), .Z(\w1[3][87] ) );
  XNOR U7791 ( .A(n5626), .B(key[472]), .Z(n5630) );
  XOR U7792 ( .A(n5628), .B(n5627), .Z(n5629) );
  XNOR U7793 ( .A(n5630), .B(n5629), .Z(\w1[3][88] ) );
  XNOR U7794 ( .A(n5631), .B(key[473]), .Z(n5634) );
  XOR U7795 ( .A(n5632), .B(\w3[2][82] ), .Z(n5633) );
  XNOR U7796 ( .A(n5634), .B(n5633), .Z(n5635) );
  XOR U7797 ( .A(\w3[2][90] ), .B(n5635), .Z(\w1[3][89] ) );
  XNOR U7798 ( .A(n5636), .B(key[392]), .Z(n5638) );
  XNOR U7799 ( .A(\w3[2][1] ), .B(\w3[2][0] ), .Z(n5637) );
  XNOR U7800 ( .A(n5638), .B(n5637), .Z(n5640) );
  XNOR U7801 ( .A(n5640), .B(n5639), .Z(\w1[3][8] ) );
  XNOR U7802 ( .A(n5641), .B(key[474]), .Z(n5644) );
  XOR U7803 ( .A(n5642), .B(\w3[2][91] ), .Z(n5643) );
  XNOR U7804 ( .A(n5644), .B(n5643), .Z(n5645) );
  XOR U7805 ( .A(\w3[2][66] ), .B(n5645), .Z(\w1[3][90] ) );
  XNOR U7806 ( .A(n5646), .B(key[475]), .Z(n5650) );
  XOR U7807 ( .A(n5648), .B(n5647), .Z(n5649) );
  XNOR U7808 ( .A(n5650), .B(n5649), .Z(\w1[3][91] ) );
  XNOR U7809 ( .A(n5651), .B(key[476]), .Z(n5654) );
  XOR U7810 ( .A(\w3[2][68] ), .B(n5652), .Z(n5653) );
  XNOR U7811 ( .A(n5654), .B(n5653), .Z(\w1[3][92] ) );
  XOR U7812 ( .A(\w3[2][86] ), .B(key[477]), .Z(n5657) );
  XOR U7813 ( .A(n5655), .B(\w3[2][94] ), .Z(n5656) );
  XNOR U7814 ( .A(n5657), .B(n5656), .Z(n5658) );
  XOR U7815 ( .A(\w3[2][69] ), .B(n5658), .Z(\w1[3][93] ) );
  XNOR U7816 ( .A(n5659), .B(key[478]), .Z(n5662) );
  XOR U7817 ( .A(\w3[2][70] ), .B(n5660), .Z(n5661) );
  XNOR U7818 ( .A(n5662), .B(n5661), .Z(\w1[3][94] ) );
  XNOR U7819 ( .A(n5663), .B(key[479]), .Z(n5666) );
  XOR U7820 ( .A(n5664), .B(\w3[2][71] ), .Z(n5665) );
  XNOR U7821 ( .A(n5666), .B(n5665), .Z(\w1[3][95] ) );
  XOR U7822 ( .A(\w3[2][104] ), .B(key[480]), .Z(n5670) );
  XNOR U7823 ( .A(n5668), .B(n5667), .Z(n5669) );
  XNOR U7824 ( .A(n5670), .B(n5669), .Z(\w1[3][96] ) );
  XNOR U7825 ( .A(n5671), .B(key[481]), .Z(n5674) );
  XOR U7826 ( .A(\w3[2][121] ), .B(n5672), .Z(n5673) );
  XNOR U7827 ( .A(n5674), .B(n5673), .Z(\w1[3][97] ) );
  XNOR U7828 ( .A(n5675), .B(key[482]), .Z(n5678) );
  XOR U7829 ( .A(\w3[2][122] ), .B(n5676), .Z(n5677) );
  XNOR U7830 ( .A(n5678), .B(n5677), .Z(\w1[3][98] ) );
  XOR U7831 ( .A(n5679), .B(key[483]), .Z(n5682) );
  XOR U7832 ( .A(n5680), .B(\w3[2][123] ), .Z(n5681) );
  XNOR U7833 ( .A(n5682), .B(n5681), .Z(\w1[3][99] ) );
  XOR U7834 ( .A(\w3[2][10] ), .B(key[393]), .Z(n5684) );
  XNOR U7835 ( .A(\w3[2][2] ), .B(\w3[2][17] ), .Z(n5683) );
  XNOR U7836 ( .A(n5684), .B(n5683), .Z(n5685) );
  XNOR U7837 ( .A(n5686), .B(n5685), .Z(\w1[3][9] ) );
  XNOR U7838 ( .A(\w3[3][25] ), .B(\w3[3][1] ), .Z(n6100) );
  IV U7839 ( .A(\w3[3][16] ), .Z(n5812) );
  XOR U7840 ( .A(\w3[3][24] ), .B(n5812), .Z(n6052) );
  XNOR U7841 ( .A(\w3[3][8] ), .B(key[512]), .Z(n5687) );
  XNOR U7842 ( .A(n6052), .B(n5687), .Z(n5688) );
  XOR U7843 ( .A(n6100), .B(n5688), .Z(\w1[4][0] ) );
  XOR U7844 ( .A(\w3[3][96] ), .B(\w3[3][101] ), .Z(n5711) );
  XOR U7845 ( .A(\w3[3][116] ), .B(\w3[3][125] ), .Z(n5690) );
  IV U7846 ( .A(\w3[3][120] ), .Z(n5759) );
  XOR U7847 ( .A(n5759), .B(\w3[3][108] ), .Z(n5689) );
  XOR U7848 ( .A(n5690), .B(n5689), .Z(n5765) );
  XOR U7849 ( .A(n5765), .B(key[612]), .Z(n5691) );
  XOR U7850 ( .A(n5711), .B(n5691), .Z(n5692) );
  XNOR U7851 ( .A(\w3[3][124] ), .B(n5692), .Z(\w1[4][100] ) );
  XNOR U7852 ( .A(\w3[3][102] ), .B(\w3[3][126] ), .Z(n5720) );
  XNOR U7853 ( .A(n5720), .B(key[613]), .Z(n5694) );
  XNOR U7854 ( .A(\w3[3][109] ), .B(\w3[3][117] ), .Z(n5768) );
  XOR U7855 ( .A(\w3[3][125] ), .B(n5768), .Z(n5693) );
  XNOR U7856 ( .A(n5694), .B(n5693), .Z(\w1[4][101] ) );
  XOR U7857 ( .A(\w3[3][96] ), .B(\w3[3][103] ), .Z(n5721) );
  XOR U7858 ( .A(n5721), .B(key[614]), .Z(n5696) );
  XNOR U7859 ( .A(\w3[3][110] ), .B(\w3[3][118] ), .Z(n5737) );
  XNOR U7860 ( .A(n5759), .B(\w3[3][127] ), .Z(n5697) );
  XOR U7861 ( .A(n5737), .B(n5697), .Z(n5773) );
  XOR U7862 ( .A(\w3[3][126] ), .B(n5773), .Z(n5695) );
  XNOR U7863 ( .A(n5696), .B(n5695), .Z(\w1[4][102] ) );
  XNOR U7864 ( .A(\w3[3][111] ), .B(\w3[3][119] ), .Z(n5776) );
  XNOR U7865 ( .A(n5776), .B(key[615]), .Z(n5699) );
  XNOR U7866 ( .A(\w3[3][96] ), .B(n5697), .Z(n5698) );
  XNOR U7867 ( .A(n5699), .B(n5698), .Z(\w1[4][103] ) );
  XNOR U7868 ( .A(\w3[3][120] ), .B(\w3[3][112] ), .Z(n6081) );
  XOR U7869 ( .A(\w3[3][106] ), .B(\w3[3][98] ), .Z(n5701) );
  XOR U7870 ( .A(\w3[3][97] ), .B(\w3[3][121] ), .Z(n6080) );
  XNOR U7871 ( .A(n6080), .B(key[617]), .Z(n5700) );
  XNOR U7872 ( .A(n5701), .B(n5700), .Z(n5702) );
  XOR U7873 ( .A(\w3[3][113] ), .B(n5702), .Z(\w1[4][105] ) );
  XOR U7874 ( .A(\w3[3][107] ), .B(\w3[3][114] ), .Z(n5704) );
  XOR U7875 ( .A(\w3[3][98] ), .B(\w3[3][122] ), .Z(n6085) );
  XNOR U7876 ( .A(n6085), .B(key[618]), .Z(n5703) );
  XNOR U7877 ( .A(n5704), .B(n5703), .Z(n5705) );
  XOR U7878 ( .A(\w3[3][99] ), .B(n5705), .Z(\w1[4][106] ) );
  IV U7879 ( .A(\w3[3][123] ), .Z(n6093) );
  XOR U7880 ( .A(\w3[3][99] ), .B(n6093), .Z(n6089) );
  XOR U7881 ( .A(\w3[3][108] ), .B(n6089), .Z(n5706) );
  XOR U7882 ( .A(\w3[3][104] ), .B(n5706), .Z(n5730) );
  XNOR U7883 ( .A(n5730), .B(key[619]), .Z(n5708) );
  IV U7884 ( .A(\w3[3][100] ), .Z(n5764) );
  XOR U7885 ( .A(\w3[3][96] ), .B(n5764), .Z(n6094) );
  XOR U7886 ( .A(\w3[3][115] ), .B(n6094), .Z(n5707) );
  XNOR U7887 ( .A(n5708), .B(n5707), .Z(\w1[4][107] ) );
  XOR U7888 ( .A(\w3[3][100] ), .B(\w3[3][104] ), .Z(n5710) );
  XNOR U7889 ( .A(\w3[3][124] ), .B(\w3[3][109] ), .Z(n5709) );
  XOR U7890 ( .A(n5710), .B(n5709), .Z(n5733) );
  XNOR U7891 ( .A(n5733), .B(key[620]), .Z(n5713) );
  XNOR U7892 ( .A(\w3[3][116] ), .B(n5711), .Z(n5712) );
  XNOR U7893 ( .A(n5713), .B(n5712), .Z(\w1[4][108] ) );
  XNOR U7894 ( .A(\w3[3][125] ), .B(\w3[3][101] ), .Z(n5736) );
  XNOR U7895 ( .A(n5736), .B(key[621]), .Z(n5715) );
  XNOR U7896 ( .A(\w3[3][102] ), .B(\w3[3][110] ), .Z(n5714) );
  XNOR U7897 ( .A(n5715), .B(n5714), .Z(n5716) );
  XOR U7898 ( .A(\w3[3][117] ), .B(n5716), .Z(\w1[4][109] ) );
  XOR U7899 ( .A(\w3[3][11] ), .B(\w3[3][3] ), .Z(n5718) );
  XNOR U7900 ( .A(\w3[3][2] ), .B(\w3[3][26] ), .Z(n5799) );
  XOR U7901 ( .A(n5799), .B(key[522]), .Z(n5717) );
  XNOR U7902 ( .A(n5718), .B(n5717), .Z(n5719) );
  XOR U7903 ( .A(\w3[3][18] ), .B(n5719), .Z(\w1[4][10] ) );
  XOR U7904 ( .A(\w3[3][111] ), .B(\w3[3][104] ), .Z(n5744) );
  XOR U7905 ( .A(n5720), .B(n5744), .Z(n5740) );
  XNOR U7906 ( .A(n5740), .B(key[622]), .Z(n5723) );
  XNOR U7907 ( .A(\w3[3][118] ), .B(n5721), .Z(n5722) );
  XNOR U7908 ( .A(n5723), .B(n5722), .Z(\w1[4][110] ) );
  XOR U7909 ( .A(\w3[3][127] ), .B(\w3[3][103] ), .Z(n5743) );
  XOR U7910 ( .A(n5743), .B(key[623]), .Z(n5725) );
  XNOR U7911 ( .A(\w3[3][96] ), .B(\w3[3][104] ), .Z(n5749) );
  XOR U7912 ( .A(\w3[3][119] ), .B(n5749), .Z(n5724) );
  XNOR U7913 ( .A(n5725), .B(n5724), .Z(\w1[4][111] ) );
  XNOR U7914 ( .A(\w3[3][105] ), .B(\w3[3][113] ), .Z(n6084) );
  XNOR U7915 ( .A(n6084), .B(key[624]), .Z(n5727) );
  XNOR U7916 ( .A(n5759), .B(n5749), .Z(n5726) );
  XNOR U7917 ( .A(n5727), .B(n5726), .Z(\w1[4][112] ) );
  XNOR U7918 ( .A(\w3[3][106] ), .B(\w3[3][114] ), .Z(n6088) );
  XNOR U7919 ( .A(\w3[3][107] ), .B(\w3[3][115] ), .Z(n5761) );
  XNOR U7920 ( .A(n5761), .B(key[626]), .Z(n5729) );
  XNOR U7921 ( .A(\w3[3][106] ), .B(n6085), .Z(n5728) );
  XNOR U7922 ( .A(n5729), .B(n5728), .Z(\w1[4][114] ) );
  XNOR U7923 ( .A(\w3[3][116] ), .B(\w3[3][112] ), .Z(n5762) );
  XNOR U7924 ( .A(n5762), .B(key[627]), .Z(n5732) );
  XOR U7925 ( .A(\w3[3][107] ), .B(n5730), .Z(n5731) );
  XNOR U7926 ( .A(n5732), .B(n5731), .Z(\w1[4][115] ) );
  XNOR U7927 ( .A(\w3[3][117] ), .B(\w3[3][112] ), .Z(n5763) );
  XNOR U7928 ( .A(n5763), .B(key[628]), .Z(n5735) );
  XOR U7929 ( .A(\w3[3][108] ), .B(n5733), .Z(n5734) );
  XNOR U7930 ( .A(n5735), .B(n5734), .Z(\w1[4][116] ) );
  XNOR U7931 ( .A(n5736), .B(key[629]), .Z(n5739) );
  XOR U7932 ( .A(\w3[3][109] ), .B(n5737), .Z(n5738) );
  XNOR U7933 ( .A(n5739), .B(n5738), .Z(\w1[4][117] ) );
  XNOR U7934 ( .A(\w3[3][119] ), .B(\w3[3][112] ), .Z(n5772) );
  XNOR U7935 ( .A(n5772), .B(key[630]), .Z(n5742) );
  XOR U7936 ( .A(\w3[3][110] ), .B(n5740), .Z(n5741) );
  XNOR U7937 ( .A(n5742), .B(n5741), .Z(\w1[4][118] ) );
  XOR U7938 ( .A(n5743), .B(key[631]), .Z(n5746) );
  XNOR U7939 ( .A(\w3[3][112] ), .B(n5744), .Z(n5745) );
  XNOR U7940 ( .A(n5746), .B(n5745), .Z(\w1[4][119] ) );
  XNOR U7941 ( .A(\w3[3][3] ), .B(\w3[3][27] ), .Z(n5833) );
  XNOR U7942 ( .A(n5796), .B(key[523]), .Z(n5748) );
  XNOR U7943 ( .A(\w3[3][0] ), .B(\w3[3][4] ), .Z(n5862) );
  XOR U7944 ( .A(\w3[3][19] ), .B(n5862), .Z(n5747) );
  XNOR U7945 ( .A(n5748), .B(n5747), .Z(\w1[4][11] ) );
  XNOR U7946 ( .A(n5749), .B(key[632]), .Z(n5751) );
  XNOR U7947 ( .A(\w3[3][113] ), .B(\w3[3][121] ), .Z(n5750) );
  XNOR U7948 ( .A(n5751), .B(n5750), .Z(n5752) );
  XOR U7949 ( .A(\w3[3][112] ), .B(n5752), .Z(\w1[4][120] ) );
  XNOR U7950 ( .A(n6084), .B(key[633]), .Z(n5754) );
  XNOR U7951 ( .A(\w3[3][122] ), .B(\w3[3][114] ), .Z(n5753) );
  XNOR U7952 ( .A(n5754), .B(n5753), .Z(n5755) );
  XOR U7953 ( .A(\w3[3][97] ), .B(n5755), .Z(\w1[4][121] ) );
  XNOR U7954 ( .A(n6088), .B(key[634]), .Z(n5757) );
  XNOR U7955 ( .A(\w3[3][115] ), .B(\w3[3][123] ), .Z(n5756) );
  XNOR U7956 ( .A(n5757), .B(n5756), .Z(n5758) );
  XOR U7957 ( .A(\w3[3][98] ), .B(n5758), .Z(\w1[4][122] ) );
  XOR U7958 ( .A(\w3[3][124] ), .B(n5759), .Z(n5760) );
  XOR U7959 ( .A(n5761), .B(n5760), .Z(n6092) );
  XNOR U7960 ( .A(n5763), .B(key[636]), .Z(n5767) );
  XNOR U7961 ( .A(n5765), .B(n5764), .Z(n5766) );
  XNOR U7962 ( .A(n5767), .B(n5766), .Z(\w1[4][124] ) );
  XOR U7963 ( .A(\w3[3][118] ), .B(key[637]), .Z(n5770) );
  XOR U7964 ( .A(n5768), .B(\w3[3][126] ), .Z(n5769) );
  XNOR U7965 ( .A(n5770), .B(n5769), .Z(n5771) );
  XOR U7966 ( .A(\w3[3][101] ), .B(n5771), .Z(\w1[4][125] ) );
  XNOR U7967 ( .A(n5772), .B(key[638]), .Z(n5775) );
  XOR U7968 ( .A(\w3[3][102] ), .B(n5773), .Z(n5774) );
  XNOR U7969 ( .A(n5775), .B(n5774), .Z(\w1[4][126] ) );
  XNOR U7970 ( .A(n6081), .B(key[639]), .Z(n5778) );
  XOR U7971 ( .A(\w3[3][103] ), .B(n5776), .Z(n5777) );
  XNOR U7972 ( .A(n5778), .B(n5777), .Z(\w1[4][127] ) );
  XOR U7973 ( .A(\w3[3][13] ), .B(\w3[3][28] ), .Z(n5780) );
  XNOR U7974 ( .A(\w3[3][8] ), .B(\w3[3][4] ), .Z(n5779) );
  XOR U7975 ( .A(n5780), .B(n5779), .Z(n5802) );
  XNOR U7976 ( .A(n5802), .B(key[524]), .Z(n5782) );
  XNOR U7977 ( .A(\w3[3][0] ), .B(\w3[3][5] ), .Z(n5897) );
  XOR U7978 ( .A(\w3[3][20] ), .B(n5897), .Z(n5781) );
  XNOR U7979 ( .A(n5782), .B(n5781), .Z(\w1[4][12] ) );
  IV U7980 ( .A(\w3[3][21] ), .Z(n5827) );
  XNOR U7981 ( .A(\w3[3][14] ), .B(n5827), .Z(n5784) );
  XNOR U7982 ( .A(\w3[3][5] ), .B(\w3[3][29] ), .Z(n5805) );
  XOR U7983 ( .A(n5805), .B(key[525]), .Z(n5783) );
  XNOR U7984 ( .A(n5784), .B(n5783), .Z(n5785) );
  XOR U7985 ( .A(\w3[3][6] ), .B(n5785), .Z(\w1[4][13] ) );
  IV U7986 ( .A(\w3[3][30] ), .Z(n5977) );
  XOR U7987 ( .A(\w3[3][6] ), .B(n5977), .Z(n5942) );
  XOR U7988 ( .A(\w3[3][8] ), .B(\w3[3][15] ), .Z(n5808) );
  XNOR U7989 ( .A(n5942), .B(n5808), .Z(n5806) );
  XOR U7990 ( .A(n5806), .B(key[526]), .Z(n5787) );
  XNOR U7991 ( .A(\w3[3][0] ), .B(\w3[3][7] ), .Z(n5978) );
  XOR U7992 ( .A(\w3[3][22] ), .B(n5978), .Z(n5786) );
  XNOR U7993 ( .A(n5787), .B(n5786), .Z(\w1[4][14] ) );
  XNOR U7994 ( .A(\w3[3][7] ), .B(\w3[3][31] ), .Z(n5807) );
  XNOR U7995 ( .A(n5807), .B(key[527]), .Z(n5789) );
  XOR U7996 ( .A(\w3[3][8] ), .B(\w3[3][0] ), .Z(n5811) );
  XNOR U7997 ( .A(\w3[3][23] ), .B(n5811), .Z(n5788) );
  XNOR U7998 ( .A(n5789), .B(n5788), .Z(\w1[4][15] ) );
  XNOR U7999 ( .A(\w3[3][17] ), .B(\w3[3][9] ), .Z(n5813) );
  XNOR U8000 ( .A(n5813), .B(key[528]), .Z(n5791) );
  XNOR U8001 ( .A(\w3[3][24] ), .B(n5811), .Z(n5790) );
  XNOR U8002 ( .A(n5791), .B(n5790), .Z(\w1[4][16] ) );
  XNOR U8003 ( .A(\w3[3][18] ), .B(\w3[3][10] ), .Z(n5832) );
  XNOR U8004 ( .A(n5832), .B(key[529]), .Z(n5793) );
  IV U8005 ( .A(\w3[3][9] ), .Z(n6049) );
  XNOR U8006 ( .A(n6100), .B(n6049), .Z(n5792) );
  XNOR U8007 ( .A(n5793), .B(n5792), .Z(\w1[4][17] ) );
  XNOR U8008 ( .A(\w3[3][11] ), .B(\w3[3][19] ), .Z(n5818) );
  XNOR U8009 ( .A(n5818), .B(key[530]), .Z(n5795) );
  XOR U8010 ( .A(n5799), .B(\w3[3][10] ), .Z(n5794) );
  XNOR U8011 ( .A(n5795), .B(n5794), .Z(\w1[4][18] ) );
  XOR U8012 ( .A(n5812), .B(\w3[3][20] ), .Z(n5819) );
  XNOR U8013 ( .A(n5819), .B(key[531]), .Z(n5798) );
  XOR U8014 ( .A(\w3[3][11] ), .B(n5796), .Z(n5797) );
  XNOR U8015 ( .A(n5798), .B(n5797), .Z(\w1[4][19] ) );
  XNOR U8016 ( .A(n5813), .B(key[513]), .Z(n5801) );
  XOR U8017 ( .A(\w3[3][25] ), .B(n5799), .Z(n5800) );
  XNOR U8018 ( .A(n5801), .B(n5800), .Z(\w1[4][1] ) );
  XOR U8019 ( .A(\w3[3][16] ), .B(n5827), .Z(n5824) );
  XNOR U8020 ( .A(n5824), .B(key[532]), .Z(n5804) );
  XOR U8021 ( .A(\w3[3][12] ), .B(n5802), .Z(n5803) );
  XNOR U8022 ( .A(n5804), .B(n5803), .Z(\w1[4][20] ) );
  IV U8023 ( .A(\w3[3][22] ), .Z(n5828) );
  XOR U8024 ( .A(\w3[3][14] ), .B(n5828), .Z(n5837) );
  XOR U8025 ( .A(n5812), .B(\w3[3][23] ), .Z(n5838) );
  XNOR U8026 ( .A(n5807), .B(key[535]), .Z(n5810) );
  XNOR U8027 ( .A(\w3[3][16] ), .B(n5808), .Z(n5809) );
  XNOR U8028 ( .A(n5810), .B(n5809), .Z(\w1[4][23] ) );
  XNOR U8029 ( .A(n5832), .B(key[538]), .Z(n5815) );
  XNOR U8030 ( .A(\w3[3][2] ), .B(\w3[3][19] ), .Z(n5814) );
  XNOR U8031 ( .A(n5815), .B(n5814), .Z(n5816) );
  XOR U8032 ( .A(\w3[3][27] ), .B(n5816), .Z(\w1[4][26] ) );
  IV U8033 ( .A(\w3[3][24] ), .Z(n5836) );
  XOR U8034 ( .A(n5836), .B(\w3[3][28] ), .Z(n5817) );
  XOR U8035 ( .A(n5818), .B(n5817), .Z(n5861) );
  XOR U8036 ( .A(n5861), .B(key[539]), .Z(n5821) );
  XOR U8037 ( .A(\w3[3][3] ), .B(n5819), .Z(n5820) );
  XNOR U8038 ( .A(n5821), .B(n5820), .Z(\w1[4][27] ) );
  XOR U8039 ( .A(\w3[3][20] ), .B(\w3[3][29] ), .Z(n5823) );
  XOR U8040 ( .A(n5836), .B(\w3[3][12] ), .Z(n5822) );
  XOR U8041 ( .A(n5823), .B(n5822), .Z(n5896) );
  XNOR U8042 ( .A(n5896), .B(key[540]), .Z(n5826) );
  XOR U8043 ( .A(\w3[3][4] ), .B(n5824), .Z(n5825) );
  XNOR U8044 ( .A(n5826), .B(n5825), .Z(\w1[4][28] ) );
  XOR U8045 ( .A(\w3[3][13] ), .B(n5827), .Z(n5941) );
  XNOR U8046 ( .A(n5941), .B(key[541]), .Z(n5830) );
  XNOR U8047 ( .A(n5828), .B(n5977), .Z(n5829) );
  XNOR U8048 ( .A(n5830), .B(n5829), .Z(n5831) );
  XOR U8049 ( .A(\w3[3][5] ), .B(n5831), .Z(\w1[4][29] ) );
  XNOR U8050 ( .A(n5832), .B(key[514]), .Z(n5835) );
  XOR U8051 ( .A(\w3[3][26] ), .B(n5833), .Z(n5834) );
  XNOR U8052 ( .A(n5835), .B(n5834), .Z(\w1[4][2] ) );
  XOR U8053 ( .A(n5836), .B(\w3[3][31] ), .Z(n6013) );
  XNOR U8054 ( .A(n5837), .B(n6013), .Z(n5976) );
  XNOR U8055 ( .A(\w3[3][15] ), .B(\w3[3][23] ), .Z(n6012) );
  XNOR U8056 ( .A(n6012), .B(key[543]), .Z(n5840) );
  XOR U8057 ( .A(n6052), .B(\w3[3][7] ), .Z(n5839) );
  XNOR U8058 ( .A(n5840), .B(n5839), .Z(\w1[4][31] ) );
  XOR U8059 ( .A(\w3[3][33] ), .B(\w3[3][57] ), .Z(n5893) );
  XOR U8060 ( .A(n5893), .B(key[544]), .Z(n5842) );
  XNOR U8061 ( .A(\w3[3][48] ), .B(\w3[3][56] ), .Z(n5958) );
  XOR U8062 ( .A(n5958), .B(\w3[3][40] ), .Z(n5841) );
  XNOR U8063 ( .A(n5842), .B(n5841), .Z(\w1[4][32] ) );
  XNOR U8064 ( .A(\w3[3][34] ), .B(\w3[3][58] ), .Z(n5901) );
  XOR U8065 ( .A(\w3[3][57] ), .B(\w3[3][49] ), .Z(n5921) );
  XNOR U8066 ( .A(n5921), .B(key[545]), .Z(n5843) );
  XNOR U8067 ( .A(n5901), .B(n5843), .Z(n5844) );
  XNOR U8068 ( .A(\w3[3][41] ), .B(n5844), .Z(\w1[4][33] ) );
  XNOR U8069 ( .A(n5870), .B(key[546]), .Z(n5846) );
  XNOR U8070 ( .A(\w3[3][50] ), .B(\w3[3][42] ), .Z(n5931) );
  XOR U8071 ( .A(\w3[3][58] ), .B(n5931), .Z(n5845) );
  XNOR U8072 ( .A(n5846), .B(n5845), .Z(\w1[4][34] ) );
  XOR U8073 ( .A(\w3[3][36] ), .B(\w3[3][32] ), .Z(n5872) );
  XOR U8074 ( .A(n5872), .B(key[547]), .Z(n5849) );
  IV U8075 ( .A(\w3[3][51] ), .Z(n5930) );
  XOR U8076 ( .A(\w3[3][43] ), .B(n5930), .Z(n5900) );
  XOR U8077 ( .A(\w3[3][56] ), .B(n5900), .Z(n5847) );
  XNOR U8078 ( .A(\w3[3][60] ), .B(n5847), .Z(n5937) );
  XNOR U8079 ( .A(\w3[3][59] ), .B(n5937), .Z(n5848) );
  XNOR U8080 ( .A(n5849), .B(n5848), .Z(\w1[4][35] ) );
  XOR U8081 ( .A(\w3[3][32] ), .B(\w3[3][37] ), .Z(n5878) );
  XOR U8082 ( .A(\w3[3][52] ), .B(\w3[3][61] ), .Z(n5851) );
  XNOR U8083 ( .A(\w3[3][56] ), .B(\w3[3][44] ), .Z(n5850) );
  XOR U8084 ( .A(n5851), .B(n5850), .Z(n5946) );
  XOR U8085 ( .A(n5946), .B(key[548]), .Z(n5852) );
  XOR U8086 ( .A(n5878), .B(n5852), .Z(n5853) );
  XNOR U8087 ( .A(\w3[3][60] ), .B(n5853), .Z(\w1[4][36] ) );
  XNOR U8088 ( .A(\w3[3][38] ), .B(\w3[3][62] ), .Z(n5884) );
  XNOR U8089 ( .A(n5884), .B(key[549]), .Z(n5855) );
  IV U8090 ( .A(\w3[3][45] ), .Z(n5910) );
  XOR U8091 ( .A(\w3[3][53] ), .B(n5910), .Z(n5949) );
  XOR U8092 ( .A(\w3[3][61] ), .B(n5949), .Z(n5854) );
  XNOR U8093 ( .A(n5855), .B(n5854), .Z(\w1[4][37] ) );
  XOR U8094 ( .A(\w3[3][32] ), .B(\w3[3][39] ), .Z(n5885) );
  XOR U8095 ( .A(n5885), .B(key[550]), .Z(n5857) );
  XNOR U8096 ( .A(\w3[3][56] ), .B(\w3[3][63] ), .Z(n5858) );
  XOR U8097 ( .A(\w3[3][46] ), .B(\w3[3][54] ), .Z(n5909) );
  XOR U8098 ( .A(n5858), .B(n5909), .Z(n5954) );
  XOR U8099 ( .A(\w3[3][62] ), .B(n5954), .Z(n5856) );
  XNOR U8100 ( .A(n5857), .B(n5856), .Z(\w1[4][38] ) );
  XNOR U8101 ( .A(\w3[3][55] ), .B(\w3[3][47] ), .Z(n5957) );
  XNOR U8102 ( .A(n5957), .B(key[551]), .Z(n5860) );
  XOR U8103 ( .A(\w3[3][32] ), .B(n5858), .Z(n5859) );
  XNOR U8104 ( .A(n5860), .B(n5859), .Z(\w1[4][39] ) );
  XOR U8105 ( .A(n5861), .B(key[515]), .Z(n5864) );
  XOR U8106 ( .A(n5862), .B(\w3[3][27] ), .Z(n5863) );
  XNOR U8107 ( .A(n5864), .B(n5863), .Z(\w1[4][3] ) );
  XNOR U8108 ( .A(\w3[3][33] ), .B(\w3[3][41] ), .Z(n5925) );
  XNOR U8109 ( .A(n5925), .B(key[552]), .Z(n5866) );
  XOR U8110 ( .A(n5958), .B(\w3[3][32] ), .Z(n5865) );
  XNOR U8111 ( .A(n5866), .B(n5865), .Z(\w1[4][40] ) );
  IV U8112 ( .A(\w3[3][34] ), .Z(n5935) );
  XOR U8113 ( .A(\w3[3][43] ), .B(key[554]), .Z(n5868) );
  IV U8114 ( .A(\w3[3][35] ), .Z(n5938) );
  XOR U8115 ( .A(\w3[3][50] ), .B(n5938), .Z(n5867) );
  XNOR U8116 ( .A(n5868), .B(n5867), .Z(n5869) );
  XNOR U8117 ( .A(n5869), .B(n5901), .Z(\w1[4][42] ) );
  IV U8118 ( .A(\w3[3][40] ), .Z(n5875) );
  XNOR U8119 ( .A(n5875), .B(n5870), .Z(n5871) );
  XOR U8120 ( .A(\w3[3][44] ), .B(n5871), .Z(n5904) );
  XNOR U8121 ( .A(n5904), .B(key[555]), .Z(n5874) );
  XNOR U8122 ( .A(\w3[3][51] ), .B(n5872), .Z(n5873) );
  XNOR U8123 ( .A(n5874), .B(n5873), .Z(\w1[4][43] ) );
  XOR U8124 ( .A(\w3[3][36] ), .B(\w3[3][45] ), .Z(n5877) );
  XOR U8125 ( .A(n5875), .B(\w3[3][60] ), .Z(n5876) );
  XOR U8126 ( .A(n5877), .B(n5876), .Z(n5905) );
  XNOR U8127 ( .A(n5905), .B(key[556]), .Z(n5880) );
  XNOR U8128 ( .A(\w3[3][52] ), .B(n5878), .Z(n5879) );
  XNOR U8129 ( .A(n5880), .B(n5879), .Z(\w1[4][44] ) );
  XNOR U8130 ( .A(\w3[3][61] ), .B(\w3[3][37] ), .Z(n5908) );
  XNOR U8131 ( .A(n5908), .B(key[557]), .Z(n5882) );
  XNOR U8132 ( .A(\w3[3][38] ), .B(\w3[3][46] ), .Z(n5881) );
  XNOR U8133 ( .A(n5882), .B(n5881), .Z(n5883) );
  XOR U8134 ( .A(\w3[3][53] ), .B(n5883), .Z(\w1[4][45] ) );
  XOR U8135 ( .A(\w3[3][40] ), .B(\w3[3][47] ), .Z(n5917) );
  XOR U8136 ( .A(n5884), .B(n5917), .Z(n5913) );
  XNOR U8137 ( .A(n5913), .B(key[558]), .Z(n5887) );
  XNOR U8138 ( .A(\w3[3][54] ), .B(n5885), .Z(n5886) );
  XNOR U8139 ( .A(n5887), .B(n5886), .Z(\w1[4][46] ) );
  XOR U8140 ( .A(\w3[3][63] ), .B(\w3[3][39] ), .Z(n5916) );
  XOR U8141 ( .A(n5916), .B(key[559]), .Z(n5889) );
  XNOR U8142 ( .A(\w3[3][40] ), .B(\w3[3][32] ), .Z(n5920) );
  XOR U8143 ( .A(\w3[3][55] ), .B(n5920), .Z(n5888) );
  XNOR U8144 ( .A(n5889), .B(n5888), .Z(\w1[4][47] ) );
  XNOR U8145 ( .A(n5920), .B(key[560]), .Z(n5891) );
  IV U8146 ( .A(\w3[3][49] ), .Z(n5926) );
  XOR U8147 ( .A(\w3[3][56] ), .B(n5926), .Z(n5890) );
  XNOR U8148 ( .A(n5891), .B(n5890), .Z(n5892) );
  XOR U8149 ( .A(\w3[3][41] ), .B(n5892), .Z(\w1[4][48] ) );
  XNOR U8150 ( .A(n5931), .B(key[561]), .Z(n5895) );
  XNOR U8151 ( .A(n5893), .B(\w3[3][41] ), .Z(n5894) );
  XNOR U8152 ( .A(n5895), .B(n5894), .Z(\w1[4][49] ) );
  XNOR U8153 ( .A(n5896), .B(key[516]), .Z(n5899) );
  XOR U8154 ( .A(n5897), .B(\w3[3][28] ), .Z(n5898) );
  XNOR U8155 ( .A(n5899), .B(n5898), .Z(\w1[4][4] ) );
  XNOR U8156 ( .A(n5900), .B(key[562]), .Z(n5903) );
  XOR U8157 ( .A(n5901), .B(\w3[3][42] ), .Z(n5902) );
  XNOR U8158 ( .A(n5903), .B(n5902), .Z(\w1[4][50] ) );
  IV U8159 ( .A(\w3[3][48] ), .Z(n5922) );
  XOR U8160 ( .A(n5922), .B(\w3[3][52] ), .Z(n5936) );
  XNOR U8161 ( .A(n5945), .B(key[564]), .Z(n5907) );
  XOR U8162 ( .A(\w3[3][44] ), .B(n5905), .Z(n5906) );
  XNOR U8163 ( .A(n5907), .B(n5906), .Z(\w1[4][52] ) );
  XNOR U8164 ( .A(n5908), .B(key[565]), .Z(n5912) );
  XOR U8165 ( .A(n5910), .B(n5909), .Z(n5911) );
  XNOR U8166 ( .A(n5912), .B(n5911), .Z(\w1[4][53] ) );
  XOR U8167 ( .A(n5922), .B(\w3[3][55] ), .Z(n5953) );
  XNOR U8168 ( .A(n5953), .B(key[566]), .Z(n5915) );
  XOR U8169 ( .A(\w3[3][46] ), .B(n5913), .Z(n5914) );
  XNOR U8170 ( .A(n5915), .B(n5914), .Z(\w1[4][54] ) );
  XOR U8171 ( .A(n5916), .B(key[567]), .Z(n5919) );
  XNOR U8172 ( .A(\w3[3][48] ), .B(n5917), .Z(n5918) );
  XNOR U8173 ( .A(n5919), .B(n5918), .Z(\w1[4][55] ) );
  XNOR U8174 ( .A(n5920), .B(key[568]), .Z(n5924) );
  XOR U8175 ( .A(n5922), .B(n5921), .Z(n5923) );
  XNOR U8176 ( .A(n5924), .B(n5923), .Z(\w1[4][56] ) );
  XNOR U8177 ( .A(n5925), .B(key[569]), .Z(n5928) );
  XOR U8178 ( .A(n5926), .B(\w3[3][50] ), .Z(n5927) );
  XNOR U8179 ( .A(n5928), .B(n5927), .Z(n5929) );
  XOR U8180 ( .A(\w3[3][58] ), .B(n5929), .Z(\w1[4][57] ) );
  XNOR U8181 ( .A(n5930), .B(key[570]), .Z(n5933) );
  XOR U8182 ( .A(n5931), .B(\w3[3][59] ), .Z(n5932) );
  XNOR U8183 ( .A(n5933), .B(n5932), .Z(n5934) );
  XNOR U8184 ( .A(n5935), .B(n5934), .Z(\w1[4][58] ) );
  XNOR U8185 ( .A(n5936), .B(key[571]), .Z(n5940) );
  XOR U8186 ( .A(n5938), .B(n5937), .Z(n5939) );
  XNOR U8187 ( .A(n5940), .B(n5939), .Z(\w1[4][59] ) );
  XNOR U8188 ( .A(n5941), .B(key[517]), .Z(n5944) );
  XOR U8189 ( .A(\w3[3][29] ), .B(n5942), .Z(n5943) );
  XNOR U8190 ( .A(n5944), .B(n5943), .Z(\w1[4][5] ) );
  XNOR U8191 ( .A(n5945), .B(key[572]), .Z(n5948) );
  XOR U8192 ( .A(\w3[3][36] ), .B(n5946), .Z(n5947) );
  XNOR U8193 ( .A(n5948), .B(n5947), .Z(\w1[4][60] ) );
  XOR U8194 ( .A(\w3[3][54] ), .B(key[573]), .Z(n5951) );
  XOR U8195 ( .A(n5949), .B(\w3[3][62] ), .Z(n5950) );
  XNOR U8196 ( .A(n5951), .B(n5950), .Z(n5952) );
  XOR U8197 ( .A(\w3[3][37] ), .B(n5952), .Z(\w1[4][61] ) );
  XNOR U8198 ( .A(n5953), .B(key[574]), .Z(n5956) );
  XOR U8199 ( .A(\w3[3][38] ), .B(n5954), .Z(n5955) );
  XNOR U8200 ( .A(n5956), .B(n5955), .Z(\w1[4][62] ) );
  XNOR U8201 ( .A(n5957), .B(key[575]), .Z(n5960) );
  XOR U8202 ( .A(n5958), .B(\w3[3][39] ), .Z(n5959) );
  XNOR U8203 ( .A(n5960), .B(n5959), .Z(\w1[4][63] ) );
  XOR U8204 ( .A(\w3[3][65] ), .B(\w3[3][89] ), .Z(n6018) );
  XOR U8205 ( .A(n6018), .B(key[576]), .Z(n5962) );
  XNOR U8206 ( .A(\w3[3][80] ), .B(\w3[3][88] ), .Z(n6077) );
  XOR U8207 ( .A(n6077), .B(\w3[3][72] ), .Z(n5961) );
  XNOR U8208 ( .A(n5962), .B(n5961), .Z(\w1[4][64] ) );
  XNOR U8209 ( .A(\w3[3][66] ), .B(\w3[3][90] ), .Z(n6022) );
  XOR U8210 ( .A(\w3[3][89] ), .B(\w3[3][81] ), .Z(n6040) );
  XNOR U8211 ( .A(n6040), .B(key[577]), .Z(n5963) );
  XNOR U8212 ( .A(n6022), .B(n5963), .Z(n5964) );
  XNOR U8213 ( .A(\w3[3][73] ), .B(n5964), .Z(\w1[4][65] ) );
  XNOR U8214 ( .A(n5992), .B(key[578]), .Z(n5966) );
  XNOR U8215 ( .A(\w3[3][82] ), .B(\w3[3][74] ), .Z(n6055) );
  XOR U8216 ( .A(\w3[3][90] ), .B(n6055), .Z(n5965) );
  XNOR U8217 ( .A(n5966), .B(n5965), .Z(\w1[4][66] ) );
  XOR U8218 ( .A(\w3[3][68] ), .B(\w3[3][64] ), .Z(n5994) );
  XOR U8219 ( .A(n5994), .B(key[579]), .Z(n5969) );
  IV U8220 ( .A(\w3[3][83] ), .Z(n6054) );
  XOR U8221 ( .A(\w3[3][75] ), .B(n6054), .Z(n6021) );
  XOR U8222 ( .A(\w3[3][88] ), .B(n6021), .Z(n5967) );
  XNOR U8223 ( .A(\w3[3][92] ), .B(n5967), .Z(n6060) );
  XNOR U8224 ( .A(\w3[3][91] ), .B(n6060), .Z(n5968) );
  XNOR U8225 ( .A(n5969), .B(n5968), .Z(\w1[4][67] ) );
  XOR U8226 ( .A(\w3[3][64] ), .B(\w3[3][69] ), .Z(n6000) );
  XOR U8227 ( .A(\w3[3][84] ), .B(\w3[3][93] ), .Z(n5971) );
  XNOR U8228 ( .A(\w3[3][88] ), .B(\w3[3][76] ), .Z(n5970) );
  XOR U8229 ( .A(n5971), .B(n5970), .Z(n6065) );
  XOR U8230 ( .A(n6065), .B(key[580]), .Z(n5972) );
  XOR U8231 ( .A(n6000), .B(n5972), .Z(n5973) );
  XNOR U8232 ( .A(\w3[3][92] ), .B(n5973), .Z(\w1[4][68] ) );
  XNOR U8233 ( .A(\w3[3][70] ), .B(\w3[3][94] ), .Z(n6006) );
  XNOR U8234 ( .A(n6006), .B(key[581]), .Z(n5975) );
  IV U8235 ( .A(\w3[3][77] ), .Z(n6029) );
  XOR U8236 ( .A(\w3[3][85] ), .B(n6029), .Z(n6068) );
  XOR U8237 ( .A(\w3[3][93] ), .B(n6068), .Z(n5974) );
  XNOR U8238 ( .A(n5975), .B(n5974), .Z(\w1[4][69] ) );
  XNOR U8239 ( .A(n5976), .B(key[518]), .Z(n5980) );
  XNOR U8240 ( .A(n5978), .B(n5977), .Z(n5979) );
  XNOR U8241 ( .A(n5980), .B(n5979), .Z(\w1[4][6] ) );
  XOR U8242 ( .A(\w3[3][64] ), .B(\w3[3][71] ), .Z(n6007) );
  XOR U8243 ( .A(n6007), .B(key[582]), .Z(n5982) );
  XNOR U8244 ( .A(\w3[3][78] ), .B(\w3[3][86] ), .Z(n6028) );
  XOR U8245 ( .A(\w3[3][88] ), .B(\w3[3][95] ), .Z(n5983) );
  XOR U8246 ( .A(n6028), .B(n5983), .Z(n6073) );
  XOR U8247 ( .A(\w3[3][94] ), .B(n6073), .Z(n5981) );
  XNOR U8248 ( .A(n5982), .B(n5981), .Z(\w1[4][70] ) );
  XNOR U8249 ( .A(\w3[3][79] ), .B(\w3[3][87] ), .Z(n6076) );
  XNOR U8250 ( .A(n6076), .B(key[583]), .Z(n5985) );
  XNOR U8251 ( .A(\w3[3][64] ), .B(n5983), .Z(n5984) );
  XNOR U8252 ( .A(n5985), .B(n5984), .Z(\w1[4][71] ) );
  IV U8253 ( .A(\w3[3][65] ), .Z(n6045) );
  XOR U8254 ( .A(\w3[3][74] ), .B(key[585]), .Z(n5987) );
  XNOR U8255 ( .A(n6040), .B(\w3[3][66] ), .Z(n5986) );
  XNOR U8256 ( .A(n5987), .B(n5986), .Z(n5988) );
  XNOR U8257 ( .A(n6045), .B(n5988), .Z(\w1[4][73] ) );
  XOR U8258 ( .A(\w3[3][75] ), .B(key[586]), .Z(n5990) );
  IV U8259 ( .A(\w3[3][67] ), .Z(n6061) );
  XOR U8260 ( .A(\w3[3][82] ), .B(n6061), .Z(n5989) );
  XNOR U8261 ( .A(n5990), .B(n5989), .Z(n5991) );
  XNOR U8262 ( .A(n5991), .B(n6022), .Z(\w1[4][74] ) );
  IV U8263 ( .A(\w3[3][72] ), .Z(n5997) );
  XNOR U8264 ( .A(n5997), .B(n5992), .Z(n5993) );
  XOR U8265 ( .A(\w3[3][76] ), .B(n5993), .Z(n6023) );
  XNOR U8266 ( .A(n6023), .B(key[587]), .Z(n5996) );
  XNOR U8267 ( .A(\w3[3][83] ), .B(n5994), .Z(n5995) );
  XNOR U8268 ( .A(n5996), .B(n5995), .Z(\w1[4][75] ) );
  XOR U8269 ( .A(\w3[3][68] ), .B(\w3[3][77] ), .Z(n5999) );
  XOR U8270 ( .A(n5997), .B(\w3[3][92] ), .Z(n5998) );
  XOR U8271 ( .A(n5999), .B(n5998), .Z(n6024) );
  XNOR U8272 ( .A(n6024), .B(key[588]), .Z(n6002) );
  XNOR U8273 ( .A(\w3[3][84] ), .B(n6000), .Z(n6001) );
  XNOR U8274 ( .A(n6002), .B(n6001), .Z(\w1[4][76] ) );
  XNOR U8275 ( .A(\w3[3][93] ), .B(\w3[3][69] ), .Z(n6027) );
  XNOR U8276 ( .A(n6027), .B(key[589]), .Z(n6004) );
  XNOR U8277 ( .A(\w3[3][70] ), .B(\w3[3][78] ), .Z(n6003) );
  XNOR U8278 ( .A(n6004), .B(n6003), .Z(n6005) );
  XOR U8279 ( .A(\w3[3][85] ), .B(n6005), .Z(\w1[4][77] ) );
  XOR U8280 ( .A(\w3[3][72] ), .B(\w3[3][79] ), .Z(n6036) );
  XOR U8281 ( .A(n6006), .B(n6036), .Z(n6032) );
  XNOR U8282 ( .A(n6032), .B(key[590]), .Z(n6009) );
  XNOR U8283 ( .A(\w3[3][86] ), .B(n6007), .Z(n6008) );
  XNOR U8284 ( .A(n6009), .B(n6008), .Z(\w1[4][78] ) );
  XOR U8285 ( .A(\w3[3][95] ), .B(\w3[3][71] ), .Z(n6035) );
  XOR U8286 ( .A(n6035), .B(key[591]), .Z(n6011) );
  XNOR U8287 ( .A(\w3[3][72] ), .B(\w3[3][64] ), .Z(n6039) );
  XOR U8288 ( .A(\w3[3][87] ), .B(n6039), .Z(n6010) );
  XNOR U8289 ( .A(n6011), .B(n6010), .Z(\w1[4][79] ) );
  XNOR U8290 ( .A(n6012), .B(key[519]), .Z(n6015) );
  XOR U8291 ( .A(\w3[3][0] ), .B(n6013), .Z(n6014) );
  XNOR U8292 ( .A(n6015), .B(n6014), .Z(\w1[4][7] ) );
  XNOR U8293 ( .A(\w3[3][73] ), .B(\w3[3][81] ), .Z(n6044) );
  XNOR U8294 ( .A(n6044), .B(key[592]), .Z(n6017) );
  XOR U8295 ( .A(\w3[3][88] ), .B(n6039), .Z(n6016) );
  XNOR U8296 ( .A(n6017), .B(n6016), .Z(\w1[4][80] ) );
  XNOR U8297 ( .A(n6055), .B(key[593]), .Z(n6020) );
  XNOR U8298 ( .A(n6018), .B(\w3[3][73] ), .Z(n6019) );
  XNOR U8299 ( .A(n6020), .B(n6019), .Z(\w1[4][81] ) );
  IV U8300 ( .A(\w3[3][80] ), .Z(n6041) );
  XOR U8301 ( .A(n6041), .B(\w3[3][84] ), .Z(n6059) );
  XNOR U8302 ( .A(n6064), .B(key[596]), .Z(n6026) );
  XOR U8303 ( .A(\w3[3][76] ), .B(n6024), .Z(n6025) );
  XNOR U8304 ( .A(n6026), .B(n6025), .Z(\w1[4][84] ) );
  XNOR U8305 ( .A(n6027), .B(key[597]), .Z(n6031) );
  XNOR U8306 ( .A(n6029), .B(n6028), .Z(n6030) );
  XNOR U8307 ( .A(n6031), .B(n6030), .Z(\w1[4][85] ) );
  XOR U8308 ( .A(n6041), .B(\w3[3][87] ), .Z(n6072) );
  XNOR U8309 ( .A(n6072), .B(key[598]), .Z(n6034) );
  XOR U8310 ( .A(\w3[3][78] ), .B(n6032), .Z(n6033) );
  XNOR U8311 ( .A(n6034), .B(n6033), .Z(\w1[4][86] ) );
  XOR U8312 ( .A(n6035), .B(key[599]), .Z(n6038) );
  XNOR U8313 ( .A(\w3[3][80] ), .B(n6036), .Z(n6037) );
  XNOR U8314 ( .A(n6038), .B(n6037), .Z(\w1[4][87] ) );
  XNOR U8315 ( .A(n6039), .B(key[600]), .Z(n6043) );
  XOR U8316 ( .A(n6041), .B(n6040), .Z(n6042) );
  XNOR U8317 ( .A(n6043), .B(n6042), .Z(\w1[4][88] ) );
  XNOR U8318 ( .A(n6044), .B(key[601]), .Z(n6047) );
  XOR U8319 ( .A(n6045), .B(\w3[3][82] ), .Z(n6046) );
  XNOR U8320 ( .A(n6047), .B(n6046), .Z(n6048) );
  XOR U8321 ( .A(\w3[3][90] ), .B(n6048), .Z(\w1[4][89] ) );
  XNOR U8322 ( .A(n6049), .B(key[520]), .Z(n6051) );
  XNOR U8323 ( .A(\w3[3][1] ), .B(\w3[3][0] ), .Z(n6050) );
  XNOR U8324 ( .A(n6051), .B(n6050), .Z(n6053) );
  XNOR U8325 ( .A(n6053), .B(n6052), .Z(\w1[4][8] ) );
  XNOR U8326 ( .A(n6054), .B(key[602]), .Z(n6057) );
  XOR U8327 ( .A(n6055), .B(\w3[3][91] ), .Z(n6056) );
  XNOR U8328 ( .A(n6057), .B(n6056), .Z(n6058) );
  XOR U8329 ( .A(\w3[3][66] ), .B(n6058), .Z(\w1[4][90] ) );
  XNOR U8330 ( .A(n6059), .B(key[603]), .Z(n6063) );
  XOR U8331 ( .A(n6061), .B(n6060), .Z(n6062) );
  XNOR U8332 ( .A(n6063), .B(n6062), .Z(\w1[4][91] ) );
  XNOR U8333 ( .A(n6064), .B(key[604]), .Z(n6067) );
  XOR U8334 ( .A(\w3[3][68] ), .B(n6065), .Z(n6066) );
  XNOR U8335 ( .A(n6067), .B(n6066), .Z(\w1[4][92] ) );
  XOR U8336 ( .A(\w3[3][86] ), .B(key[605]), .Z(n6070) );
  XOR U8337 ( .A(n6068), .B(\w3[3][94] ), .Z(n6069) );
  XNOR U8338 ( .A(n6070), .B(n6069), .Z(n6071) );
  XOR U8339 ( .A(\w3[3][69] ), .B(n6071), .Z(\w1[4][93] ) );
  XNOR U8340 ( .A(n6072), .B(key[606]), .Z(n6075) );
  XOR U8341 ( .A(\w3[3][70] ), .B(n6073), .Z(n6074) );
  XNOR U8342 ( .A(n6075), .B(n6074), .Z(\w1[4][94] ) );
  XNOR U8343 ( .A(n6076), .B(key[607]), .Z(n6079) );
  XOR U8344 ( .A(n6077), .B(\w3[3][71] ), .Z(n6078) );
  XNOR U8345 ( .A(n6079), .B(n6078), .Z(\w1[4][95] ) );
  XOR U8346 ( .A(\w3[3][104] ), .B(key[608]), .Z(n6083) );
  XOR U8347 ( .A(n6081), .B(n6080), .Z(n6082) );
  XNOR U8348 ( .A(n6083), .B(n6082), .Z(\w1[4][96] ) );
  XNOR U8349 ( .A(n6084), .B(key[609]), .Z(n6087) );
  XNOR U8350 ( .A(\w3[3][121] ), .B(n6085), .Z(n6086) );
  XNOR U8351 ( .A(n6087), .B(n6086), .Z(\w1[4][97] ) );
  XNOR U8352 ( .A(n6088), .B(key[610]), .Z(n6091) );
  XOR U8353 ( .A(\w3[3][122] ), .B(n6089), .Z(n6090) );
  XNOR U8354 ( .A(n6091), .B(n6090), .Z(\w1[4][98] ) );
  XOR U8355 ( .A(n6092), .B(key[611]), .Z(n6096) );
  XNOR U8356 ( .A(n6094), .B(n6093), .Z(n6095) );
  XNOR U8357 ( .A(n6096), .B(n6095), .Z(\w1[4][99] ) );
  XOR U8358 ( .A(\w3[3][10] ), .B(key[521]), .Z(n6098) );
  XNOR U8359 ( .A(\w3[3][2] ), .B(\w3[3][17] ), .Z(n6097) );
  XNOR U8360 ( .A(n6098), .B(n6097), .Z(n6099) );
  XNOR U8361 ( .A(n6100), .B(n6099), .Z(\w1[4][9] ) );
  XNOR U8362 ( .A(\w3[4][25] ), .B(\w3[4][1] ), .Z(n6521) );
  IV U8363 ( .A(\w3[4][16] ), .Z(n6232) );
  XOR U8364 ( .A(\w3[4][24] ), .B(n6232), .Z(n6472) );
  XNOR U8365 ( .A(\w3[4][8] ), .B(key[640]), .Z(n6101) );
  XNOR U8366 ( .A(n6472), .B(n6101), .Z(n6102) );
  XOR U8367 ( .A(n6521), .B(n6102), .Z(\w1[5][0] ) );
  XOR U8368 ( .A(\w3[4][96] ), .B(\w3[4][101] ), .Z(n6125) );
  XOR U8369 ( .A(\w3[4][116] ), .B(\w3[4][125] ), .Z(n6104) );
  IV U8370 ( .A(\w3[4][120] ), .Z(n6176) );
  XOR U8371 ( .A(n6176), .B(\w3[4][108] ), .Z(n6103) );
  XOR U8372 ( .A(n6104), .B(n6103), .Z(n6185) );
  XOR U8373 ( .A(n6185), .B(key[740]), .Z(n6105) );
  XOR U8374 ( .A(n6125), .B(n6105), .Z(n6106) );
  XNOR U8375 ( .A(\w3[4][124] ), .B(n6106), .Z(\w1[5][100] ) );
  XNOR U8376 ( .A(\w3[4][102] ), .B(\w3[4][126] ), .Z(n6134) );
  XNOR U8377 ( .A(n6134), .B(key[741]), .Z(n6108) );
  XNOR U8378 ( .A(\w3[4][109] ), .B(\w3[4][117] ), .Z(n6188) );
  XOR U8379 ( .A(\w3[4][125] ), .B(n6188), .Z(n6107) );
  XNOR U8380 ( .A(n6108), .B(n6107), .Z(\w1[5][101] ) );
  XOR U8381 ( .A(\w3[4][96] ), .B(\w3[4][103] ), .Z(n6135) );
  XOR U8382 ( .A(n6135), .B(key[742]), .Z(n6110) );
  XNOR U8383 ( .A(\w3[4][110] ), .B(\w3[4][118] ), .Z(n6151) );
  XNOR U8384 ( .A(n6176), .B(\w3[4][127] ), .Z(n6111) );
  XOR U8385 ( .A(n6151), .B(n6111), .Z(n6193) );
  XOR U8386 ( .A(\w3[4][126] ), .B(n6193), .Z(n6109) );
  XNOR U8387 ( .A(n6110), .B(n6109), .Z(\w1[5][102] ) );
  XNOR U8388 ( .A(\w3[4][111] ), .B(\w3[4][119] ), .Z(n6196) );
  XNOR U8389 ( .A(n6196), .B(key[743]), .Z(n6113) );
  XNOR U8390 ( .A(\w3[4][96] ), .B(n6111), .Z(n6112) );
  XNOR U8391 ( .A(n6113), .B(n6112), .Z(\w1[5][103] ) );
  IV U8392 ( .A(\w3[4][97] ), .Z(n6171) );
  IV U8393 ( .A(\w3[4][112] ), .Z(n6167) );
  XOR U8394 ( .A(\w3[4][120] ), .B(n6167), .Z(n6502) );
  XOR U8395 ( .A(\w3[4][106] ), .B(\w3[4][98] ), .Z(n6115) );
  XNOR U8396 ( .A(\w3[4][97] ), .B(\w3[4][121] ), .Z(n6501) );
  XOR U8397 ( .A(n6501), .B(key[745]), .Z(n6114) );
  XNOR U8398 ( .A(n6115), .B(n6114), .Z(n6116) );
  XOR U8399 ( .A(\w3[4][113] ), .B(n6116), .Z(\w1[5][105] ) );
  IV U8400 ( .A(\w3[4][99] ), .Z(n6180) );
  XNOR U8401 ( .A(\w3[4][107] ), .B(n6180), .Z(n6118) );
  XOR U8402 ( .A(\w3[4][98] ), .B(\w3[4][122] ), .Z(n6506) );
  XNOR U8403 ( .A(n6506), .B(key[746]), .Z(n6117) );
  XNOR U8404 ( .A(n6118), .B(n6117), .Z(n6119) );
  XOR U8405 ( .A(\w3[4][114] ), .B(n6119), .Z(\w1[5][106] ) );
  IV U8406 ( .A(\w3[4][123] ), .Z(n6514) );
  XOR U8407 ( .A(\w3[4][99] ), .B(n6514), .Z(n6510) );
  XOR U8408 ( .A(\w3[4][108] ), .B(n6510), .Z(n6120) );
  XOR U8409 ( .A(\w3[4][104] ), .B(n6120), .Z(n6146) );
  XNOR U8410 ( .A(n6146), .B(key[747]), .Z(n6122) );
  IV U8411 ( .A(\w3[4][100] ), .Z(n6184) );
  XOR U8412 ( .A(\w3[4][96] ), .B(n6184), .Z(n6515) );
  XOR U8413 ( .A(\w3[4][115] ), .B(n6515), .Z(n6121) );
  XNOR U8414 ( .A(n6122), .B(n6121), .Z(\w1[5][107] ) );
  XOR U8415 ( .A(\w3[4][100] ), .B(\w3[4][104] ), .Z(n6124) );
  XNOR U8416 ( .A(\w3[4][124] ), .B(\w3[4][109] ), .Z(n6123) );
  XOR U8417 ( .A(n6124), .B(n6123), .Z(n6147) );
  XNOR U8418 ( .A(n6147), .B(key[748]), .Z(n6127) );
  XNOR U8419 ( .A(\w3[4][116] ), .B(n6125), .Z(n6126) );
  XNOR U8420 ( .A(n6127), .B(n6126), .Z(\w1[5][108] ) );
  XNOR U8421 ( .A(\w3[4][125] ), .B(\w3[4][101] ), .Z(n6150) );
  XNOR U8422 ( .A(n6150), .B(key[749]), .Z(n6129) );
  XNOR U8423 ( .A(\w3[4][102] ), .B(\w3[4][110] ), .Z(n6128) );
  XNOR U8424 ( .A(n6129), .B(n6128), .Z(n6130) );
  XOR U8425 ( .A(\w3[4][117] ), .B(n6130), .Z(\w1[5][109] ) );
  XOR U8426 ( .A(\w3[4][11] ), .B(\w3[4][3] ), .Z(n6132) );
  XNOR U8427 ( .A(\w3[4][2] ), .B(\w3[4][26] ), .Z(n6219) );
  XOR U8428 ( .A(n6219), .B(key[650]), .Z(n6131) );
  XNOR U8429 ( .A(n6132), .B(n6131), .Z(n6133) );
  XOR U8430 ( .A(\w3[4][18] ), .B(n6133), .Z(\w1[5][10] ) );
  XOR U8431 ( .A(\w3[4][111] ), .B(\w3[4][104] ), .Z(n6158) );
  XOR U8432 ( .A(n6134), .B(n6158), .Z(n6154) );
  XNOR U8433 ( .A(n6154), .B(key[750]), .Z(n6137) );
  XNOR U8434 ( .A(\w3[4][118] ), .B(n6135), .Z(n6136) );
  XNOR U8435 ( .A(n6137), .B(n6136), .Z(\w1[5][110] ) );
  XOR U8436 ( .A(\w3[4][127] ), .B(\w3[4][103] ), .Z(n6157) );
  XOR U8437 ( .A(n6157), .B(key[751]), .Z(n6139) );
  XNOR U8438 ( .A(\w3[4][96] ), .B(\w3[4][104] ), .Z(n6163) );
  XOR U8439 ( .A(\w3[4][119] ), .B(n6163), .Z(n6138) );
  XNOR U8440 ( .A(n6139), .B(n6138), .Z(\w1[5][111] ) );
  XNOR U8441 ( .A(\w3[4][105] ), .B(\w3[4][113] ), .Z(n6505) );
  XNOR U8442 ( .A(n6505), .B(key[752]), .Z(n6141) );
  XNOR U8443 ( .A(n6176), .B(n6163), .Z(n6140) );
  XNOR U8444 ( .A(n6141), .B(n6140), .Z(\w1[5][112] ) );
  XNOR U8445 ( .A(\w3[4][106] ), .B(\w3[4][114] ), .Z(n6509) );
  XNOR U8446 ( .A(n6509), .B(key[753]), .Z(n6143) );
  XOR U8447 ( .A(\w3[4][105] ), .B(n6501), .Z(n6142) );
  XNOR U8448 ( .A(n6143), .B(n6142), .Z(\w1[5][113] ) );
  IV U8449 ( .A(\w3[4][115] ), .Z(n6172) );
  XOR U8450 ( .A(\w3[4][107] ), .B(n6172), .Z(n6178) );
  XNOR U8451 ( .A(n6178), .B(key[754]), .Z(n6145) );
  XNOR U8452 ( .A(\w3[4][106] ), .B(n6506), .Z(n6144) );
  XNOR U8453 ( .A(n6145), .B(n6144), .Z(\w1[5][114] ) );
  XOR U8454 ( .A(\w3[4][116] ), .B(n6167), .Z(n6179) );
  XOR U8455 ( .A(\w3[4][117] ), .B(n6167), .Z(n6183) );
  XNOR U8456 ( .A(n6183), .B(key[756]), .Z(n6149) );
  XOR U8457 ( .A(\w3[4][108] ), .B(n6147), .Z(n6148) );
  XNOR U8458 ( .A(n6149), .B(n6148), .Z(\w1[5][116] ) );
  XNOR U8459 ( .A(n6150), .B(key[757]), .Z(n6153) );
  XOR U8460 ( .A(\w3[4][109] ), .B(n6151), .Z(n6152) );
  XNOR U8461 ( .A(n6153), .B(n6152), .Z(\w1[5][117] ) );
  XOR U8462 ( .A(\w3[4][119] ), .B(n6167), .Z(n6192) );
  XNOR U8463 ( .A(n6192), .B(key[758]), .Z(n6156) );
  XOR U8464 ( .A(\w3[4][110] ), .B(n6154), .Z(n6155) );
  XNOR U8465 ( .A(n6156), .B(n6155), .Z(\w1[5][118] ) );
  XOR U8466 ( .A(n6157), .B(key[759]), .Z(n6160) );
  XNOR U8467 ( .A(\w3[4][112] ), .B(n6158), .Z(n6159) );
  XNOR U8468 ( .A(n6160), .B(n6159), .Z(\w1[5][119] ) );
  XNOR U8469 ( .A(\w3[4][3] ), .B(\w3[4][27] ), .Z(n6253) );
  XNOR U8470 ( .A(n6216), .B(key[651]), .Z(n6162) );
  XNOR U8471 ( .A(\w3[4][0] ), .B(\w3[4][4] ), .Z(n6282) );
  XOR U8472 ( .A(\w3[4][19] ), .B(n6282), .Z(n6161) );
  XNOR U8473 ( .A(n6162), .B(n6161), .Z(\w1[5][11] ) );
  XNOR U8474 ( .A(n6163), .B(key[760]), .Z(n6165) );
  XNOR U8475 ( .A(\w3[4][113] ), .B(\w3[4][121] ), .Z(n6164) );
  XNOR U8476 ( .A(n6165), .B(n6164), .Z(n6166) );
  XNOR U8477 ( .A(n6167), .B(n6166), .Z(\w1[5][120] ) );
  XNOR U8478 ( .A(n6505), .B(key[761]), .Z(n6169) );
  XNOR U8479 ( .A(\w3[4][114] ), .B(\w3[4][122] ), .Z(n6168) );
  XNOR U8480 ( .A(n6169), .B(n6168), .Z(n6170) );
  XNOR U8481 ( .A(n6171), .B(n6170), .Z(\w1[5][121] ) );
  XNOR U8482 ( .A(n6509), .B(key[762]), .Z(n6174) );
  XNOR U8483 ( .A(n6172), .B(n6514), .Z(n6173) );
  XNOR U8484 ( .A(n6174), .B(n6173), .Z(n6175) );
  XOR U8485 ( .A(\w3[4][98] ), .B(n6175), .Z(\w1[5][122] ) );
  XOR U8486 ( .A(\w3[4][124] ), .B(n6176), .Z(n6177) );
  XOR U8487 ( .A(n6178), .B(n6177), .Z(n6513) );
  XOR U8488 ( .A(n6513), .B(key[763]), .Z(n6182) );
  XNOR U8489 ( .A(n6180), .B(n6179), .Z(n6181) );
  XNOR U8490 ( .A(n6182), .B(n6181), .Z(\w1[5][123] ) );
  XNOR U8491 ( .A(n6183), .B(key[764]), .Z(n6187) );
  XNOR U8492 ( .A(n6185), .B(n6184), .Z(n6186) );
  XNOR U8493 ( .A(n6187), .B(n6186), .Z(\w1[5][124] ) );
  XOR U8494 ( .A(\w3[4][118] ), .B(key[765]), .Z(n6190) );
  XOR U8495 ( .A(n6188), .B(\w3[4][126] ), .Z(n6189) );
  XNOR U8496 ( .A(n6190), .B(n6189), .Z(n6191) );
  XOR U8497 ( .A(\w3[4][101] ), .B(n6191), .Z(\w1[5][125] ) );
  XNOR U8498 ( .A(n6192), .B(key[766]), .Z(n6195) );
  XOR U8499 ( .A(\w3[4][102] ), .B(n6193), .Z(n6194) );
  XNOR U8500 ( .A(n6195), .B(n6194), .Z(\w1[5][126] ) );
  XNOR U8501 ( .A(n6502), .B(key[767]), .Z(n6198) );
  XOR U8502 ( .A(\w3[4][103] ), .B(n6196), .Z(n6197) );
  XNOR U8503 ( .A(n6198), .B(n6197), .Z(\w1[5][127] ) );
  XOR U8504 ( .A(\w3[4][13] ), .B(\w3[4][28] ), .Z(n6200) );
  XNOR U8505 ( .A(\w3[4][8] ), .B(\w3[4][4] ), .Z(n6199) );
  XOR U8506 ( .A(n6200), .B(n6199), .Z(n6222) );
  XNOR U8507 ( .A(n6222), .B(key[652]), .Z(n6202) );
  XNOR U8508 ( .A(\w3[4][0] ), .B(\w3[4][5] ), .Z(n6317) );
  XOR U8509 ( .A(\w3[4][20] ), .B(n6317), .Z(n6201) );
  XNOR U8510 ( .A(n6202), .B(n6201), .Z(\w1[5][12] ) );
  IV U8511 ( .A(\w3[4][21] ), .Z(n6247) );
  XNOR U8512 ( .A(\w3[4][14] ), .B(n6247), .Z(n6204) );
  XNOR U8513 ( .A(\w3[4][5] ), .B(\w3[4][29] ), .Z(n6225) );
  XOR U8514 ( .A(n6225), .B(key[653]), .Z(n6203) );
  XNOR U8515 ( .A(n6204), .B(n6203), .Z(n6205) );
  XOR U8516 ( .A(\w3[4][6] ), .B(n6205), .Z(\w1[5][13] ) );
  IV U8517 ( .A(\w3[4][30] ), .Z(n6395) );
  XOR U8518 ( .A(\w3[4][6] ), .B(n6395), .Z(n6359) );
  XOR U8519 ( .A(\w3[4][8] ), .B(\w3[4][15] ), .Z(n6228) );
  XNOR U8520 ( .A(n6359), .B(n6228), .Z(n6226) );
  XOR U8521 ( .A(n6226), .B(key[654]), .Z(n6207) );
  XNOR U8522 ( .A(\w3[4][0] ), .B(\w3[4][7] ), .Z(n6396) );
  XOR U8523 ( .A(\w3[4][22] ), .B(n6396), .Z(n6206) );
  XNOR U8524 ( .A(n6207), .B(n6206), .Z(\w1[5][14] ) );
  XNOR U8525 ( .A(\w3[4][7] ), .B(\w3[4][31] ), .Z(n6227) );
  XNOR U8526 ( .A(n6227), .B(key[655]), .Z(n6209) );
  XOR U8527 ( .A(\w3[4][8] ), .B(\w3[4][0] ), .Z(n6231) );
  XNOR U8528 ( .A(\w3[4][23] ), .B(n6231), .Z(n6208) );
  XNOR U8529 ( .A(n6209), .B(n6208), .Z(\w1[5][15] ) );
  XNOR U8530 ( .A(\w3[4][17] ), .B(\w3[4][9] ), .Z(n6233) );
  XNOR U8531 ( .A(n6233), .B(key[656]), .Z(n6211) );
  XNOR U8532 ( .A(\w3[4][24] ), .B(n6231), .Z(n6210) );
  XNOR U8533 ( .A(n6211), .B(n6210), .Z(\w1[5][16] ) );
  XNOR U8534 ( .A(\w3[4][18] ), .B(\w3[4][10] ), .Z(n6252) );
  XNOR U8535 ( .A(n6252), .B(key[657]), .Z(n6213) );
  IV U8536 ( .A(\w3[4][9] ), .Z(n6469) );
  XNOR U8537 ( .A(n6521), .B(n6469), .Z(n6212) );
  XNOR U8538 ( .A(n6213), .B(n6212), .Z(\w1[5][17] ) );
  XNOR U8539 ( .A(\w3[4][11] ), .B(\w3[4][19] ), .Z(n6238) );
  XNOR U8540 ( .A(n6238), .B(key[658]), .Z(n6215) );
  XOR U8541 ( .A(n6219), .B(\w3[4][10] ), .Z(n6214) );
  XNOR U8542 ( .A(n6215), .B(n6214), .Z(\w1[5][18] ) );
  XOR U8543 ( .A(n6232), .B(\w3[4][20] ), .Z(n6239) );
  XNOR U8544 ( .A(n6239), .B(key[659]), .Z(n6218) );
  XOR U8545 ( .A(\w3[4][11] ), .B(n6216), .Z(n6217) );
  XNOR U8546 ( .A(n6218), .B(n6217), .Z(\w1[5][19] ) );
  XNOR U8547 ( .A(n6233), .B(key[641]), .Z(n6221) );
  XOR U8548 ( .A(\w3[4][25] ), .B(n6219), .Z(n6220) );
  XNOR U8549 ( .A(n6221), .B(n6220), .Z(\w1[5][1] ) );
  XOR U8550 ( .A(\w3[4][16] ), .B(n6247), .Z(n6244) );
  XNOR U8551 ( .A(n6244), .B(key[660]), .Z(n6224) );
  XOR U8552 ( .A(\w3[4][12] ), .B(n6222), .Z(n6223) );
  XNOR U8553 ( .A(n6224), .B(n6223), .Z(\w1[5][20] ) );
  IV U8554 ( .A(\w3[4][22] ), .Z(n6248) );
  XOR U8555 ( .A(\w3[4][14] ), .B(n6248), .Z(n6257) );
  XOR U8556 ( .A(n6232), .B(\w3[4][23] ), .Z(n6258) );
  XNOR U8557 ( .A(n6227), .B(key[663]), .Z(n6230) );
  XNOR U8558 ( .A(\w3[4][16] ), .B(n6228), .Z(n6229) );
  XNOR U8559 ( .A(n6230), .B(n6229), .Z(\w1[5][23] ) );
  XNOR U8560 ( .A(n6252), .B(key[666]), .Z(n6235) );
  XNOR U8561 ( .A(\w3[4][2] ), .B(\w3[4][19] ), .Z(n6234) );
  XNOR U8562 ( .A(n6235), .B(n6234), .Z(n6236) );
  XOR U8563 ( .A(\w3[4][27] ), .B(n6236), .Z(\w1[5][26] ) );
  IV U8564 ( .A(\w3[4][24] ), .Z(n6256) );
  XOR U8565 ( .A(n6256), .B(\w3[4][28] ), .Z(n6237) );
  XOR U8566 ( .A(n6238), .B(n6237), .Z(n6281) );
  XOR U8567 ( .A(n6281), .B(key[667]), .Z(n6241) );
  XOR U8568 ( .A(\w3[4][3] ), .B(n6239), .Z(n6240) );
  XNOR U8569 ( .A(n6241), .B(n6240), .Z(\w1[5][27] ) );
  XOR U8570 ( .A(\w3[4][20] ), .B(\w3[4][29] ), .Z(n6243) );
  XOR U8571 ( .A(n6256), .B(\w3[4][12] ), .Z(n6242) );
  XOR U8572 ( .A(n6243), .B(n6242), .Z(n6316) );
  XNOR U8573 ( .A(n6316), .B(key[668]), .Z(n6246) );
  XOR U8574 ( .A(\w3[4][4] ), .B(n6244), .Z(n6245) );
  XNOR U8575 ( .A(n6246), .B(n6245), .Z(\w1[5][28] ) );
  XOR U8576 ( .A(\w3[4][13] ), .B(n6247), .Z(n6358) );
  XNOR U8577 ( .A(n6358), .B(key[669]), .Z(n6250) );
  XNOR U8578 ( .A(n6248), .B(n6395), .Z(n6249) );
  XNOR U8579 ( .A(n6250), .B(n6249), .Z(n6251) );
  XOR U8580 ( .A(\w3[4][5] ), .B(n6251), .Z(\w1[5][29] ) );
  XNOR U8581 ( .A(n6252), .B(key[642]), .Z(n6255) );
  XOR U8582 ( .A(\w3[4][26] ), .B(n6253), .Z(n6254) );
  XNOR U8583 ( .A(n6255), .B(n6254), .Z(\w1[5][2] ) );
  XOR U8584 ( .A(n6256), .B(\w3[4][31] ), .Z(n6431) );
  XNOR U8585 ( .A(n6257), .B(n6431), .Z(n6394) );
  XNOR U8586 ( .A(\w3[4][15] ), .B(\w3[4][23] ), .Z(n6430) );
  XNOR U8587 ( .A(n6430), .B(key[671]), .Z(n6260) );
  XOR U8588 ( .A(n6472), .B(\w3[4][7] ), .Z(n6259) );
  XNOR U8589 ( .A(n6260), .B(n6259), .Z(\w1[5][31] ) );
  XOR U8590 ( .A(\w3[4][33] ), .B(\w3[4][57] ), .Z(n6313) );
  XOR U8591 ( .A(n6313), .B(key[672]), .Z(n6262) );
  XNOR U8592 ( .A(\w3[4][48] ), .B(\w3[4][56] ), .Z(n6375) );
  XOR U8593 ( .A(n6375), .B(\w3[4][40] ), .Z(n6261) );
  XNOR U8594 ( .A(n6262), .B(n6261), .Z(\w1[5][32] ) );
  XNOR U8595 ( .A(\w3[4][34] ), .B(\w3[4][58] ), .Z(n6321) );
  XOR U8596 ( .A(\w3[4][57] ), .B(\w3[4][49] ), .Z(n6339) );
  XNOR U8597 ( .A(n6339), .B(key[673]), .Z(n6263) );
  XNOR U8598 ( .A(n6321), .B(n6263), .Z(n6264) );
  XNOR U8599 ( .A(\w3[4][41] ), .B(n6264), .Z(\w1[5][33] ) );
  XNOR U8600 ( .A(n6291), .B(key[674]), .Z(n6266) );
  XNOR U8601 ( .A(\w3[4][50] ), .B(\w3[4][42] ), .Z(n6349) );
  XOR U8602 ( .A(\w3[4][58] ), .B(n6349), .Z(n6265) );
  XNOR U8603 ( .A(n6266), .B(n6265), .Z(\w1[5][34] ) );
  XOR U8604 ( .A(\w3[4][36] ), .B(\w3[4][32] ), .Z(n6293) );
  XOR U8605 ( .A(n6293), .B(key[675]), .Z(n6269) );
  IV U8606 ( .A(\w3[4][51] ), .Z(n6348) );
  XOR U8607 ( .A(\w3[4][43] ), .B(n6348), .Z(n6320) );
  XOR U8608 ( .A(\w3[4][56] ), .B(n6320), .Z(n6267) );
  XNOR U8609 ( .A(\w3[4][60] ), .B(n6267), .Z(n6354) );
  XNOR U8610 ( .A(\w3[4][59] ), .B(n6354), .Z(n6268) );
  XNOR U8611 ( .A(n6269), .B(n6268), .Z(\w1[5][35] ) );
  XOR U8612 ( .A(\w3[4][32] ), .B(\w3[4][37] ), .Z(n6299) );
  XOR U8613 ( .A(\w3[4][52] ), .B(\w3[4][61] ), .Z(n6271) );
  XNOR U8614 ( .A(\w3[4][56] ), .B(\w3[4][44] ), .Z(n6270) );
  XOR U8615 ( .A(n6271), .B(n6270), .Z(n6363) );
  XOR U8616 ( .A(n6363), .B(key[676]), .Z(n6272) );
  XOR U8617 ( .A(n6299), .B(n6272), .Z(n6273) );
  XNOR U8618 ( .A(\w3[4][60] ), .B(n6273), .Z(\w1[5][36] ) );
  XNOR U8619 ( .A(\w3[4][38] ), .B(\w3[4][62] ), .Z(n6305) );
  XNOR U8620 ( .A(n6305), .B(key[677]), .Z(n6275) );
  IV U8621 ( .A(\w3[4][45] ), .Z(n6328) );
  XOR U8622 ( .A(\w3[4][53] ), .B(n6328), .Z(n6366) );
  XOR U8623 ( .A(\w3[4][61] ), .B(n6366), .Z(n6274) );
  XNOR U8624 ( .A(n6275), .B(n6274), .Z(\w1[5][37] ) );
  XOR U8625 ( .A(\w3[4][32] ), .B(\w3[4][39] ), .Z(n6306) );
  XOR U8626 ( .A(n6306), .B(key[678]), .Z(n6277) );
  XNOR U8627 ( .A(\w3[4][46] ), .B(\w3[4][54] ), .Z(n6327) );
  XOR U8628 ( .A(\w3[4][56] ), .B(\w3[4][63] ), .Z(n6278) );
  XOR U8629 ( .A(n6327), .B(n6278), .Z(n6371) );
  XOR U8630 ( .A(\w3[4][62] ), .B(n6371), .Z(n6276) );
  XNOR U8631 ( .A(n6277), .B(n6276), .Z(\w1[5][38] ) );
  XNOR U8632 ( .A(\w3[4][55] ), .B(\w3[4][47] ), .Z(n6374) );
  XNOR U8633 ( .A(n6374), .B(key[679]), .Z(n6280) );
  XNOR U8634 ( .A(\w3[4][32] ), .B(n6278), .Z(n6279) );
  XNOR U8635 ( .A(n6280), .B(n6279), .Z(\w1[5][39] ) );
  XOR U8636 ( .A(n6281), .B(key[643]), .Z(n6284) );
  XOR U8637 ( .A(n6282), .B(\w3[4][27] ), .Z(n6283) );
  XNOR U8638 ( .A(n6284), .B(n6283), .Z(\w1[5][3] ) );
  IV U8639 ( .A(\w3[4][33] ), .Z(n6344) );
  XOR U8640 ( .A(\w3[4][42] ), .B(key[681]), .Z(n6286) );
  XNOR U8641 ( .A(n6339), .B(\w3[4][34] ), .Z(n6285) );
  XNOR U8642 ( .A(n6286), .B(n6285), .Z(n6287) );
  XNOR U8643 ( .A(n6344), .B(n6287), .Z(\w1[5][41] ) );
  XOR U8644 ( .A(\w3[4][43] ), .B(key[682]), .Z(n6289) );
  IV U8645 ( .A(\w3[4][35] ), .Z(n6355) );
  XOR U8646 ( .A(\w3[4][50] ), .B(n6355), .Z(n6288) );
  XNOR U8647 ( .A(n6289), .B(n6288), .Z(n6290) );
  XNOR U8648 ( .A(n6290), .B(n6321), .Z(\w1[5][42] ) );
  IV U8649 ( .A(\w3[4][40] ), .Z(n6296) );
  XNOR U8650 ( .A(n6296), .B(n6291), .Z(n6292) );
  XOR U8651 ( .A(\w3[4][44] ), .B(n6292), .Z(n6322) );
  XNOR U8652 ( .A(n6322), .B(key[683]), .Z(n6295) );
  XNOR U8653 ( .A(\w3[4][51] ), .B(n6293), .Z(n6294) );
  XNOR U8654 ( .A(n6295), .B(n6294), .Z(\w1[5][43] ) );
  XOR U8655 ( .A(\w3[4][36] ), .B(\w3[4][45] ), .Z(n6298) );
  XOR U8656 ( .A(n6296), .B(\w3[4][60] ), .Z(n6297) );
  XOR U8657 ( .A(n6298), .B(n6297), .Z(n6323) );
  XNOR U8658 ( .A(n6323), .B(key[684]), .Z(n6301) );
  XNOR U8659 ( .A(\w3[4][52] ), .B(n6299), .Z(n6300) );
  XNOR U8660 ( .A(n6301), .B(n6300), .Z(\w1[5][44] ) );
  XNOR U8661 ( .A(\w3[4][61] ), .B(\w3[4][37] ), .Z(n6326) );
  XNOR U8662 ( .A(n6326), .B(key[685]), .Z(n6303) );
  XNOR U8663 ( .A(\w3[4][38] ), .B(\w3[4][46] ), .Z(n6302) );
  XNOR U8664 ( .A(n6303), .B(n6302), .Z(n6304) );
  XOR U8665 ( .A(\w3[4][53] ), .B(n6304), .Z(\w1[5][45] ) );
  XOR U8666 ( .A(\w3[4][40] ), .B(\w3[4][47] ), .Z(n6335) );
  XOR U8667 ( .A(n6305), .B(n6335), .Z(n6331) );
  XNOR U8668 ( .A(n6331), .B(key[686]), .Z(n6308) );
  XNOR U8669 ( .A(\w3[4][54] ), .B(n6306), .Z(n6307) );
  XNOR U8670 ( .A(n6308), .B(n6307), .Z(\w1[5][46] ) );
  XOR U8671 ( .A(\w3[4][63] ), .B(\w3[4][39] ), .Z(n6334) );
  XOR U8672 ( .A(n6334), .B(key[687]), .Z(n6310) );
  XNOR U8673 ( .A(\w3[4][40] ), .B(\w3[4][32] ), .Z(n6338) );
  XOR U8674 ( .A(\w3[4][55] ), .B(n6338), .Z(n6309) );
  XNOR U8675 ( .A(n6310), .B(n6309), .Z(\w1[5][47] ) );
  XNOR U8676 ( .A(\w3[4][41] ), .B(\w3[4][49] ), .Z(n6343) );
  XNOR U8677 ( .A(n6343), .B(key[688]), .Z(n6312) );
  XOR U8678 ( .A(\w3[4][56] ), .B(n6338), .Z(n6311) );
  XNOR U8679 ( .A(n6312), .B(n6311), .Z(\w1[5][48] ) );
  XNOR U8680 ( .A(n6349), .B(key[689]), .Z(n6315) );
  XNOR U8681 ( .A(n6313), .B(\w3[4][41] ), .Z(n6314) );
  XNOR U8682 ( .A(n6315), .B(n6314), .Z(\w1[5][49] ) );
  XNOR U8683 ( .A(n6316), .B(key[644]), .Z(n6319) );
  XOR U8684 ( .A(n6317), .B(\w3[4][28] ), .Z(n6318) );
  XNOR U8685 ( .A(n6319), .B(n6318), .Z(\w1[5][4] ) );
  IV U8686 ( .A(\w3[4][48] ), .Z(n6340) );
  XOR U8687 ( .A(n6340), .B(\w3[4][52] ), .Z(n6353) );
  XNOR U8688 ( .A(n6362), .B(key[692]), .Z(n6325) );
  XOR U8689 ( .A(\w3[4][44] ), .B(n6323), .Z(n6324) );
  XNOR U8690 ( .A(n6325), .B(n6324), .Z(\w1[5][52] ) );
  XNOR U8691 ( .A(n6326), .B(key[693]), .Z(n6330) );
  XNOR U8692 ( .A(n6328), .B(n6327), .Z(n6329) );
  XNOR U8693 ( .A(n6330), .B(n6329), .Z(\w1[5][53] ) );
  XOR U8694 ( .A(n6340), .B(\w3[4][55] ), .Z(n6370) );
  XNOR U8695 ( .A(n6370), .B(key[694]), .Z(n6333) );
  XOR U8696 ( .A(\w3[4][46] ), .B(n6331), .Z(n6332) );
  XNOR U8697 ( .A(n6333), .B(n6332), .Z(\w1[5][54] ) );
  XOR U8698 ( .A(n6334), .B(key[695]), .Z(n6337) );
  XNOR U8699 ( .A(\w3[4][48] ), .B(n6335), .Z(n6336) );
  XNOR U8700 ( .A(n6337), .B(n6336), .Z(\w1[5][55] ) );
  XNOR U8701 ( .A(n6338), .B(key[696]), .Z(n6342) );
  XOR U8702 ( .A(n6340), .B(n6339), .Z(n6341) );
  XNOR U8703 ( .A(n6342), .B(n6341), .Z(\w1[5][56] ) );
  XNOR U8704 ( .A(n6343), .B(key[697]), .Z(n6346) );
  XOR U8705 ( .A(n6344), .B(\w3[4][50] ), .Z(n6345) );
  XNOR U8706 ( .A(n6346), .B(n6345), .Z(n6347) );
  XOR U8707 ( .A(\w3[4][58] ), .B(n6347), .Z(\w1[5][57] ) );
  XNOR U8708 ( .A(n6348), .B(key[698]), .Z(n6351) );
  XOR U8709 ( .A(n6349), .B(\w3[4][59] ), .Z(n6350) );
  XNOR U8710 ( .A(n6351), .B(n6350), .Z(n6352) );
  XOR U8711 ( .A(\w3[4][34] ), .B(n6352), .Z(\w1[5][58] ) );
  XNOR U8712 ( .A(n6353), .B(key[699]), .Z(n6357) );
  XOR U8713 ( .A(n6355), .B(n6354), .Z(n6356) );
  XNOR U8714 ( .A(n6357), .B(n6356), .Z(\w1[5][59] ) );
  XNOR U8715 ( .A(n6358), .B(key[645]), .Z(n6361) );
  XOR U8716 ( .A(\w3[4][29] ), .B(n6359), .Z(n6360) );
  XNOR U8717 ( .A(n6361), .B(n6360), .Z(\w1[5][5] ) );
  XNOR U8718 ( .A(n6362), .B(key[700]), .Z(n6365) );
  XOR U8719 ( .A(\w3[4][36] ), .B(n6363), .Z(n6364) );
  XNOR U8720 ( .A(n6365), .B(n6364), .Z(\w1[5][60] ) );
  XOR U8721 ( .A(\w3[4][54] ), .B(key[701]), .Z(n6368) );
  XOR U8722 ( .A(n6366), .B(\w3[4][62] ), .Z(n6367) );
  XNOR U8723 ( .A(n6368), .B(n6367), .Z(n6369) );
  XOR U8724 ( .A(\w3[4][37] ), .B(n6369), .Z(\w1[5][61] ) );
  XNOR U8725 ( .A(n6370), .B(key[702]), .Z(n6373) );
  XOR U8726 ( .A(\w3[4][38] ), .B(n6371), .Z(n6372) );
  XNOR U8727 ( .A(n6373), .B(n6372), .Z(\w1[5][62] ) );
  XNOR U8728 ( .A(n6374), .B(key[703]), .Z(n6377) );
  XOR U8729 ( .A(n6375), .B(\w3[4][39] ), .Z(n6376) );
  XNOR U8730 ( .A(n6377), .B(n6376), .Z(\w1[5][63] ) );
  XOR U8731 ( .A(\w3[4][65] ), .B(\w3[4][89] ), .Z(n6379) );
  XNOR U8732 ( .A(\w3[4][72] ), .B(key[704]), .Z(n6378) );
  XNOR U8733 ( .A(n6379), .B(n6378), .Z(n6380) );
  IV U8734 ( .A(\w3[4][88] ), .Z(n6399) );
  XOR U8735 ( .A(\w3[4][80] ), .B(n6399), .Z(n6498) );
  XNOR U8736 ( .A(n6380), .B(n6498), .Z(\w1[5][64] ) );
  XNOR U8737 ( .A(\w3[4][66] ), .B(\w3[4][90] ), .Z(n6440) );
  XOR U8738 ( .A(\w3[4][89] ), .B(\w3[4][81] ), .Z(n6460) );
  XNOR U8739 ( .A(n6460), .B(key[705]), .Z(n6381) );
  XNOR U8740 ( .A(n6440), .B(n6381), .Z(n6382) );
  XNOR U8741 ( .A(\w3[4][73] ), .B(n6382), .Z(\w1[5][65] ) );
  XNOR U8742 ( .A(n6410), .B(key[706]), .Z(n6384) );
  XNOR U8743 ( .A(\w3[4][82] ), .B(\w3[4][74] ), .Z(n6475) );
  XOR U8744 ( .A(\w3[4][90] ), .B(n6475), .Z(n6383) );
  XNOR U8745 ( .A(n6384), .B(n6383), .Z(\w1[5][66] ) );
  XOR U8746 ( .A(\w3[4][68] ), .B(\w3[4][64] ), .Z(n6412) );
  XOR U8747 ( .A(n6412), .B(key[707]), .Z(n6387) );
  IV U8748 ( .A(\w3[4][83] ), .Z(n6474) );
  XOR U8749 ( .A(\w3[4][75] ), .B(n6474), .Z(n6439) );
  XNOR U8750 ( .A(n6399), .B(n6439), .Z(n6385) );
  XNOR U8751 ( .A(\w3[4][92] ), .B(n6385), .Z(n6481) );
  XNOR U8752 ( .A(\w3[4][91] ), .B(n6481), .Z(n6386) );
  XNOR U8753 ( .A(n6387), .B(n6386), .Z(\w1[5][67] ) );
  XOR U8754 ( .A(\w3[4][64] ), .B(\w3[4][69] ), .Z(n6418) );
  XOR U8755 ( .A(\w3[4][84] ), .B(\w3[4][93] ), .Z(n6389) );
  XOR U8756 ( .A(n6399), .B(\w3[4][76] ), .Z(n6388) );
  XOR U8757 ( .A(n6389), .B(n6388), .Z(n6486) );
  XOR U8758 ( .A(n6486), .B(key[708]), .Z(n6390) );
  XOR U8759 ( .A(n6418), .B(n6390), .Z(n6391) );
  XNOR U8760 ( .A(\w3[4][92] ), .B(n6391), .Z(\w1[5][68] ) );
  XNOR U8761 ( .A(\w3[4][70] ), .B(\w3[4][94] ), .Z(n6424) );
  XNOR U8762 ( .A(n6424), .B(key[709]), .Z(n6393) );
  IV U8763 ( .A(\w3[4][77] ), .Z(n6449) );
  XOR U8764 ( .A(\w3[4][85] ), .B(n6449), .Z(n6489) );
  XOR U8765 ( .A(\w3[4][93] ), .B(n6489), .Z(n6392) );
  XNOR U8766 ( .A(n6393), .B(n6392), .Z(\w1[5][69] ) );
  XNOR U8767 ( .A(n6394), .B(key[646]), .Z(n6398) );
  XNOR U8768 ( .A(n6396), .B(n6395), .Z(n6397) );
  XNOR U8769 ( .A(n6398), .B(n6397), .Z(\w1[5][6] ) );
  XOR U8770 ( .A(\w3[4][64] ), .B(\w3[4][71] ), .Z(n6425) );
  XOR U8771 ( .A(n6425), .B(key[710]), .Z(n6401) );
  XNOR U8772 ( .A(\w3[4][78] ), .B(\w3[4][86] ), .Z(n6448) );
  XNOR U8773 ( .A(n6399), .B(\w3[4][95] ), .Z(n6402) );
  XOR U8774 ( .A(n6448), .B(n6402), .Z(n6494) );
  XOR U8775 ( .A(\w3[4][94] ), .B(n6494), .Z(n6400) );
  XNOR U8776 ( .A(n6401), .B(n6400), .Z(\w1[5][70] ) );
  XNOR U8777 ( .A(\w3[4][79] ), .B(\w3[4][87] ), .Z(n6497) );
  XNOR U8778 ( .A(n6497), .B(key[711]), .Z(n6404) );
  XNOR U8779 ( .A(\w3[4][64] ), .B(n6402), .Z(n6403) );
  XNOR U8780 ( .A(n6404), .B(n6403), .Z(\w1[5][71] ) );
  XNOR U8781 ( .A(\w3[4][65] ), .B(\w3[4][73] ), .Z(n6464) );
  XNOR U8782 ( .A(n6464), .B(key[712]), .Z(n6406) );
  XOR U8783 ( .A(n6498), .B(\w3[4][64] ), .Z(n6405) );
  XNOR U8784 ( .A(n6406), .B(n6405), .Z(\w1[5][72] ) );
  IV U8785 ( .A(\w3[4][66] ), .Z(n6479) );
  XOR U8786 ( .A(\w3[4][75] ), .B(key[714]), .Z(n6408) );
  IV U8787 ( .A(\w3[4][67] ), .Z(n6482) );
  XOR U8788 ( .A(\w3[4][82] ), .B(n6482), .Z(n6407) );
  XNOR U8789 ( .A(n6408), .B(n6407), .Z(n6409) );
  XNOR U8790 ( .A(n6409), .B(n6440), .Z(\w1[5][74] ) );
  IV U8791 ( .A(\w3[4][72] ), .Z(n6415) );
  XNOR U8792 ( .A(n6415), .B(n6410), .Z(n6411) );
  XOR U8793 ( .A(\w3[4][76] ), .B(n6411), .Z(n6443) );
  XNOR U8794 ( .A(n6443), .B(key[715]), .Z(n6414) );
  XNOR U8795 ( .A(\w3[4][83] ), .B(n6412), .Z(n6413) );
  XNOR U8796 ( .A(n6414), .B(n6413), .Z(\w1[5][75] ) );
  XOR U8797 ( .A(\w3[4][68] ), .B(\w3[4][77] ), .Z(n6417) );
  XOR U8798 ( .A(n6415), .B(\w3[4][92] ), .Z(n6416) );
  XOR U8799 ( .A(n6417), .B(n6416), .Z(n6444) );
  XNOR U8800 ( .A(n6444), .B(key[716]), .Z(n6420) );
  XNOR U8801 ( .A(\w3[4][84] ), .B(n6418), .Z(n6419) );
  XNOR U8802 ( .A(n6420), .B(n6419), .Z(\w1[5][76] ) );
  XNOR U8803 ( .A(\w3[4][93] ), .B(\w3[4][69] ), .Z(n6447) );
  XNOR U8804 ( .A(n6447), .B(key[717]), .Z(n6422) );
  XNOR U8805 ( .A(\w3[4][70] ), .B(\w3[4][78] ), .Z(n6421) );
  XNOR U8806 ( .A(n6422), .B(n6421), .Z(n6423) );
  XOR U8807 ( .A(\w3[4][85] ), .B(n6423), .Z(\w1[5][77] ) );
  XOR U8808 ( .A(\w3[4][72] ), .B(\w3[4][79] ), .Z(n6456) );
  XOR U8809 ( .A(n6424), .B(n6456), .Z(n6452) );
  XNOR U8810 ( .A(n6452), .B(key[718]), .Z(n6427) );
  XNOR U8811 ( .A(\w3[4][86] ), .B(n6425), .Z(n6426) );
  XNOR U8812 ( .A(n6427), .B(n6426), .Z(\w1[5][78] ) );
  XOR U8813 ( .A(\w3[4][95] ), .B(\w3[4][71] ), .Z(n6455) );
  XOR U8814 ( .A(n6455), .B(key[719]), .Z(n6429) );
  XNOR U8815 ( .A(\w3[4][72] ), .B(\w3[4][64] ), .Z(n6459) );
  XOR U8816 ( .A(\w3[4][87] ), .B(n6459), .Z(n6428) );
  XNOR U8817 ( .A(n6429), .B(n6428), .Z(\w1[5][79] ) );
  XNOR U8818 ( .A(n6430), .B(key[647]), .Z(n6433) );
  XOR U8819 ( .A(\w3[4][0] ), .B(n6431), .Z(n6432) );
  XNOR U8820 ( .A(n6433), .B(n6432), .Z(\w1[5][7] ) );
  XNOR U8821 ( .A(n6459), .B(key[720]), .Z(n6435) );
  IV U8822 ( .A(\w3[4][81] ), .Z(n6465) );
  XOR U8823 ( .A(\w3[4][88] ), .B(n6465), .Z(n6434) );
  XNOR U8824 ( .A(n6435), .B(n6434), .Z(n6436) );
  XOR U8825 ( .A(\w3[4][73] ), .B(n6436), .Z(\w1[5][80] ) );
  XNOR U8826 ( .A(n6464), .B(key[721]), .Z(n6438) );
  XOR U8827 ( .A(\w3[4][89] ), .B(n6475), .Z(n6437) );
  XNOR U8828 ( .A(n6438), .B(n6437), .Z(\w1[5][81] ) );
  XNOR U8829 ( .A(n6439), .B(key[722]), .Z(n6442) );
  XOR U8830 ( .A(n6440), .B(\w3[4][74] ), .Z(n6441) );
  XNOR U8831 ( .A(n6442), .B(n6441), .Z(\w1[5][82] ) );
  IV U8832 ( .A(\w3[4][80] ), .Z(n6461) );
  XOR U8833 ( .A(n6461), .B(\w3[4][84] ), .Z(n6480) );
  XNOR U8834 ( .A(n6485), .B(key[724]), .Z(n6446) );
  XOR U8835 ( .A(\w3[4][76] ), .B(n6444), .Z(n6445) );
  XNOR U8836 ( .A(n6446), .B(n6445), .Z(\w1[5][84] ) );
  XNOR U8837 ( .A(n6447), .B(key[725]), .Z(n6451) );
  XNOR U8838 ( .A(n6449), .B(n6448), .Z(n6450) );
  XNOR U8839 ( .A(n6451), .B(n6450), .Z(\w1[5][85] ) );
  XOR U8840 ( .A(n6461), .B(\w3[4][87] ), .Z(n6493) );
  XNOR U8841 ( .A(n6493), .B(key[726]), .Z(n6454) );
  XOR U8842 ( .A(\w3[4][78] ), .B(n6452), .Z(n6453) );
  XNOR U8843 ( .A(n6454), .B(n6453), .Z(\w1[5][86] ) );
  XOR U8844 ( .A(n6455), .B(key[727]), .Z(n6458) );
  XNOR U8845 ( .A(\w3[4][80] ), .B(n6456), .Z(n6457) );
  XNOR U8846 ( .A(n6458), .B(n6457), .Z(\w1[5][87] ) );
  XNOR U8847 ( .A(n6459), .B(key[728]), .Z(n6463) );
  XOR U8848 ( .A(n6461), .B(n6460), .Z(n6462) );
  XNOR U8849 ( .A(n6463), .B(n6462), .Z(\w1[5][88] ) );
  XNOR U8850 ( .A(n6464), .B(key[729]), .Z(n6467) );
  XOR U8851 ( .A(n6465), .B(\w3[4][82] ), .Z(n6466) );
  XNOR U8852 ( .A(n6467), .B(n6466), .Z(n6468) );
  XOR U8853 ( .A(\w3[4][90] ), .B(n6468), .Z(\w1[5][89] ) );
  XNOR U8854 ( .A(n6469), .B(key[648]), .Z(n6471) );
  XNOR U8855 ( .A(\w3[4][1] ), .B(\w3[4][0] ), .Z(n6470) );
  XNOR U8856 ( .A(n6471), .B(n6470), .Z(n6473) );
  XNOR U8857 ( .A(n6473), .B(n6472), .Z(\w1[5][8] ) );
  XNOR U8858 ( .A(n6474), .B(key[730]), .Z(n6477) );
  XOR U8859 ( .A(n6475), .B(\w3[4][91] ), .Z(n6476) );
  XNOR U8860 ( .A(n6477), .B(n6476), .Z(n6478) );
  XNOR U8861 ( .A(n6479), .B(n6478), .Z(\w1[5][90] ) );
  XNOR U8862 ( .A(n6480), .B(key[731]), .Z(n6484) );
  XOR U8863 ( .A(n6482), .B(n6481), .Z(n6483) );
  XNOR U8864 ( .A(n6484), .B(n6483), .Z(\w1[5][91] ) );
  XNOR U8865 ( .A(n6485), .B(key[732]), .Z(n6488) );
  XOR U8866 ( .A(\w3[4][68] ), .B(n6486), .Z(n6487) );
  XNOR U8867 ( .A(n6488), .B(n6487), .Z(\w1[5][92] ) );
  XOR U8868 ( .A(\w3[4][86] ), .B(key[733]), .Z(n6491) );
  XOR U8869 ( .A(n6489), .B(\w3[4][94] ), .Z(n6490) );
  XNOR U8870 ( .A(n6491), .B(n6490), .Z(n6492) );
  XOR U8871 ( .A(\w3[4][69] ), .B(n6492), .Z(\w1[5][93] ) );
  XNOR U8872 ( .A(n6493), .B(key[734]), .Z(n6496) );
  XOR U8873 ( .A(\w3[4][70] ), .B(n6494), .Z(n6495) );
  XNOR U8874 ( .A(n6496), .B(n6495), .Z(\w1[5][94] ) );
  XNOR U8875 ( .A(n6497), .B(key[735]), .Z(n6500) );
  XOR U8876 ( .A(n6498), .B(\w3[4][71] ), .Z(n6499) );
  XNOR U8877 ( .A(n6500), .B(n6499), .Z(\w1[5][95] ) );
  XOR U8878 ( .A(\w3[4][104] ), .B(key[736]), .Z(n6504) );
  XNOR U8879 ( .A(n6502), .B(n6501), .Z(n6503) );
  XNOR U8880 ( .A(n6504), .B(n6503), .Z(\w1[5][96] ) );
  XNOR U8881 ( .A(n6505), .B(key[737]), .Z(n6508) );
  XNOR U8882 ( .A(\w3[4][121] ), .B(n6506), .Z(n6507) );
  XNOR U8883 ( .A(n6508), .B(n6507), .Z(\w1[5][97] ) );
  XNOR U8884 ( .A(n6509), .B(key[738]), .Z(n6512) );
  XOR U8885 ( .A(\w3[4][122] ), .B(n6510), .Z(n6511) );
  XNOR U8886 ( .A(n6512), .B(n6511), .Z(\w1[5][98] ) );
  XOR U8887 ( .A(n6513), .B(key[739]), .Z(n6517) );
  XNOR U8888 ( .A(n6515), .B(n6514), .Z(n6516) );
  XNOR U8889 ( .A(n6517), .B(n6516), .Z(\w1[5][99] ) );
  XOR U8890 ( .A(\w3[4][10] ), .B(key[649]), .Z(n6519) );
  XNOR U8891 ( .A(\w3[4][2] ), .B(\w3[4][17] ), .Z(n6518) );
  XNOR U8892 ( .A(n6519), .B(n6518), .Z(n6520) );
  XNOR U8893 ( .A(n6521), .B(n6520), .Z(\w1[5][9] ) );
  XNOR U8894 ( .A(\w3[5][25] ), .B(\w3[5][1] ), .Z(n6940) );
  IV U8895 ( .A(\w3[5][16] ), .Z(n6654) );
  XOR U8896 ( .A(\w3[5][24] ), .B(n6654), .Z(n6891) );
  XNOR U8897 ( .A(\w3[5][8] ), .B(key[768]), .Z(n6522) );
  XNOR U8898 ( .A(n6891), .B(n6522), .Z(n6523) );
  XOR U8899 ( .A(n6940), .B(n6523), .Z(\w1[6][0] ) );
  XOR U8900 ( .A(\w3[5][96] ), .B(\w3[5][101] ), .Z(n6546) );
  XOR U8901 ( .A(\w3[5][116] ), .B(\w3[5][125] ), .Z(n6525) );
  IV U8902 ( .A(\w3[5][120] ), .Z(n6598) );
  XOR U8903 ( .A(n6598), .B(\w3[5][108] ), .Z(n6524) );
  XOR U8904 ( .A(n6525), .B(n6524), .Z(n6607) );
  XOR U8905 ( .A(n6607), .B(key[868]), .Z(n6526) );
  XOR U8906 ( .A(n6546), .B(n6526), .Z(n6527) );
  XNOR U8907 ( .A(\w3[5][124] ), .B(n6527), .Z(\w1[6][100] ) );
  XNOR U8908 ( .A(\w3[5][102] ), .B(\w3[5][126] ), .Z(n6555) );
  XNOR U8909 ( .A(n6555), .B(key[869]), .Z(n6529) );
  XNOR U8910 ( .A(\w3[5][109] ), .B(\w3[5][117] ), .Z(n6610) );
  XOR U8911 ( .A(\w3[5][125] ), .B(n6610), .Z(n6528) );
  XNOR U8912 ( .A(n6529), .B(n6528), .Z(\w1[6][101] ) );
  XOR U8913 ( .A(\w3[5][96] ), .B(\w3[5][103] ), .Z(n6556) );
  XOR U8914 ( .A(n6556), .B(key[870]), .Z(n6531) );
  XOR U8915 ( .A(n6598), .B(\w3[5][127] ), .Z(n6532) );
  XOR U8916 ( .A(\w3[5][110] ), .B(\w3[5][118] ), .Z(n6572) );
  XOR U8917 ( .A(n6532), .B(n6572), .Z(n6615) );
  XOR U8918 ( .A(\w3[5][126] ), .B(n6615), .Z(n6530) );
  XNOR U8919 ( .A(n6531), .B(n6530), .Z(\w1[6][102] ) );
  XNOR U8920 ( .A(\w3[5][111] ), .B(\w3[5][119] ), .Z(n6618) );
  XNOR U8921 ( .A(n6618), .B(key[871]), .Z(n6534) );
  XOR U8922 ( .A(\w3[5][96] ), .B(n6532), .Z(n6533) );
  XNOR U8923 ( .A(n6534), .B(n6533), .Z(\w1[6][103] ) );
  IV U8924 ( .A(\w3[5][97] ), .Z(n6590) );
  IV U8925 ( .A(\w3[5][112] ), .Z(n6588) );
  XOR U8926 ( .A(\w3[5][120] ), .B(n6588), .Z(n6920) );
  XOR U8927 ( .A(\w3[5][106] ), .B(\w3[5][113] ), .Z(n6536) );
  XNOR U8928 ( .A(\w3[5][97] ), .B(\w3[5][121] ), .Z(n6919) );
  XOR U8929 ( .A(n6919), .B(key[873]), .Z(n6535) );
  XNOR U8930 ( .A(n6536), .B(n6535), .Z(n6537) );
  XOR U8931 ( .A(\w3[5][98] ), .B(n6537), .Z(\w1[6][105] ) );
  IV U8932 ( .A(\w3[5][98] ), .Z(n6597) );
  IV U8933 ( .A(\w3[5][99] ), .Z(n6602) );
  XNOR U8934 ( .A(\w3[5][107] ), .B(n6602), .Z(n6539) );
  IV U8935 ( .A(\w3[5][122] ), .Z(n6929) );
  XOR U8936 ( .A(n6929), .B(\w3[5][114] ), .Z(n6589) );
  XOR U8937 ( .A(n6589), .B(key[874]), .Z(n6538) );
  XNOR U8938 ( .A(n6539), .B(n6538), .Z(n6540) );
  XNOR U8939 ( .A(n6597), .B(n6540), .Z(\w1[6][106] ) );
  IV U8940 ( .A(\w3[5][123] ), .Z(n6933) );
  XOR U8941 ( .A(\w3[5][99] ), .B(n6933), .Z(n6928) );
  XOR U8942 ( .A(\w3[5][108] ), .B(n6928), .Z(n6541) );
  XOR U8943 ( .A(\w3[5][104] ), .B(n6541), .Z(n6567) );
  XNOR U8944 ( .A(n6567), .B(key[875]), .Z(n6543) );
  IV U8945 ( .A(\w3[5][100] ), .Z(n6606) );
  XOR U8946 ( .A(\w3[5][96] ), .B(n6606), .Z(n6934) );
  XOR U8947 ( .A(\w3[5][115] ), .B(n6934), .Z(n6542) );
  XNOR U8948 ( .A(n6543), .B(n6542), .Z(\w1[6][107] ) );
  XOR U8949 ( .A(\w3[5][100] ), .B(\w3[5][104] ), .Z(n6545) );
  XNOR U8950 ( .A(\w3[5][124] ), .B(\w3[5][109] ), .Z(n6544) );
  XOR U8951 ( .A(n6545), .B(n6544), .Z(n6568) );
  XNOR U8952 ( .A(n6568), .B(key[876]), .Z(n6548) );
  XNOR U8953 ( .A(\w3[5][116] ), .B(n6546), .Z(n6547) );
  XNOR U8954 ( .A(n6548), .B(n6547), .Z(\w1[6][108] ) );
  XNOR U8955 ( .A(\w3[5][125] ), .B(\w3[5][101] ), .Z(n6571) );
  XNOR U8956 ( .A(n6571), .B(key[877]), .Z(n6550) );
  XNOR U8957 ( .A(\w3[5][102] ), .B(\w3[5][110] ), .Z(n6549) );
  XNOR U8958 ( .A(n6550), .B(n6549), .Z(n6551) );
  XOR U8959 ( .A(\w3[5][117] ), .B(n6551), .Z(\w1[6][109] ) );
  XOR U8960 ( .A(\w3[5][11] ), .B(\w3[5][3] ), .Z(n6553) );
  XNOR U8961 ( .A(\w3[5][2] ), .B(\w3[5][26] ), .Z(n6641) );
  XOR U8962 ( .A(n6641), .B(key[778]), .Z(n6552) );
  XNOR U8963 ( .A(n6553), .B(n6552), .Z(n6554) );
  XOR U8964 ( .A(\w3[5][18] ), .B(n6554), .Z(\w1[6][10] ) );
  XOR U8965 ( .A(\w3[5][111] ), .B(\w3[5][104] ), .Z(n6579) );
  XOR U8966 ( .A(n6555), .B(n6579), .Z(n6575) );
  XNOR U8967 ( .A(n6575), .B(key[878]), .Z(n6558) );
  XNOR U8968 ( .A(\w3[5][118] ), .B(n6556), .Z(n6557) );
  XNOR U8969 ( .A(n6558), .B(n6557), .Z(\w1[6][110] ) );
  XOR U8970 ( .A(\w3[5][127] ), .B(\w3[5][103] ), .Z(n6578) );
  XOR U8971 ( .A(n6578), .B(key[879]), .Z(n6560) );
  XNOR U8972 ( .A(\w3[5][96] ), .B(\w3[5][104] ), .Z(n6584) );
  XOR U8973 ( .A(\w3[5][119] ), .B(n6584), .Z(n6559) );
  XNOR U8974 ( .A(n6560), .B(n6559), .Z(\w1[6][111] ) );
  XOR U8975 ( .A(\w3[5][105] ), .B(\w3[5][113] ), .Z(n6924) );
  XOR U8976 ( .A(n6924), .B(key[880]), .Z(n6562) );
  XNOR U8977 ( .A(n6598), .B(n6584), .Z(n6561) );
  XNOR U8978 ( .A(n6562), .B(n6561), .Z(\w1[6][112] ) );
  XNOR U8979 ( .A(\w3[5][106] ), .B(\w3[5][114] ), .Z(n6927) );
  XNOR U8980 ( .A(n6927), .B(key[881]), .Z(n6564) );
  XOR U8981 ( .A(\w3[5][105] ), .B(n6919), .Z(n6563) );
  XNOR U8982 ( .A(n6564), .B(n6563), .Z(\w1[6][113] ) );
  XOR U8983 ( .A(\w3[5][98] ), .B(n6929), .Z(n6923) );
  XNOR U8984 ( .A(n6923), .B(key[882]), .Z(n6566) );
  IV U8985 ( .A(\w3[5][115] ), .Z(n6593) );
  XOR U8986 ( .A(\w3[5][107] ), .B(n6593), .Z(n6600) );
  XOR U8987 ( .A(\w3[5][106] ), .B(n6600), .Z(n6565) );
  XNOR U8988 ( .A(n6566), .B(n6565), .Z(\w1[6][114] ) );
  XOR U8989 ( .A(\w3[5][116] ), .B(n6588), .Z(n6601) );
  XOR U8990 ( .A(\w3[5][117] ), .B(n6588), .Z(n6605) );
  XNOR U8991 ( .A(n6605), .B(key[884]), .Z(n6570) );
  XOR U8992 ( .A(\w3[5][108] ), .B(n6568), .Z(n6569) );
  XNOR U8993 ( .A(n6570), .B(n6569), .Z(\w1[6][116] ) );
  XNOR U8994 ( .A(n6571), .B(key[885]), .Z(n6574) );
  XNOR U8995 ( .A(\w3[5][109] ), .B(n6572), .Z(n6573) );
  XNOR U8996 ( .A(n6574), .B(n6573), .Z(\w1[6][117] ) );
  XOR U8997 ( .A(\w3[5][119] ), .B(n6588), .Z(n6614) );
  XNOR U8998 ( .A(n6614), .B(key[886]), .Z(n6577) );
  XOR U8999 ( .A(\w3[5][110] ), .B(n6575), .Z(n6576) );
  XNOR U9000 ( .A(n6577), .B(n6576), .Z(\w1[6][118] ) );
  XOR U9001 ( .A(n6578), .B(key[887]), .Z(n6581) );
  XNOR U9002 ( .A(\w3[5][112] ), .B(n6579), .Z(n6580) );
  XNOR U9003 ( .A(n6581), .B(n6580), .Z(\w1[6][119] ) );
  XNOR U9004 ( .A(\w3[5][3] ), .B(\w3[5][27] ), .Z(n6675) );
  XNOR U9005 ( .A(n6638), .B(key[779]), .Z(n6583) );
  XNOR U9006 ( .A(\w3[5][0] ), .B(\w3[5][4] ), .Z(n6704) );
  XOR U9007 ( .A(\w3[5][19] ), .B(n6704), .Z(n6582) );
  XNOR U9008 ( .A(n6583), .B(n6582), .Z(\w1[6][11] ) );
  XNOR U9009 ( .A(n6584), .B(key[888]), .Z(n6586) );
  XNOR U9010 ( .A(\w3[5][121] ), .B(\w3[5][113] ), .Z(n6585) );
  XNOR U9011 ( .A(n6586), .B(n6585), .Z(n6587) );
  XNOR U9012 ( .A(n6588), .B(n6587), .Z(\w1[6][120] ) );
  XOR U9013 ( .A(n6924), .B(key[889]), .Z(n6592) );
  XNOR U9014 ( .A(n6590), .B(n6589), .Z(n6591) );
  XNOR U9015 ( .A(n6592), .B(n6591), .Z(\w1[6][121] ) );
  XNOR U9016 ( .A(n6927), .B(key[890]), .Z(n6595) );
  XNOR U9017 ( .A(n6593), .B(n6933), .Z(n6594) );
  XNOR U9018 ( .A(n6595), .B(n6594), .Z(n6596) );
  XNOR U9019 ( .A(n6597), .B(n6596), .Z(\w1[6][122] ) );
  XOR U9020 ( .A(\w3[5][124] ), .B(n6598), .Z(n6599) );
  XOR U9021 ( .A(n6600), .B(n6599), .Z(n6932) );
  XOR U9022 ( .A(n6932), .B(key[891]), .Z(n6604) );
  XNOR U9023 ( .A(n6602), .B(n6601), .Z(n6603) );
  XNOR U9024 ( .A(n6604), .B(n6603), .Z(\w1[6][123] ) );
  XNOR U9025 ( .A(n6605), .B(key[892]), .Z(n6609) );
  XNOR U9026 ( .A(n6607), .B(n6606), .Z(n6608) );
  XNOR U9027 ( .A(n6609), .B(n6608), .Z(\w1[6][124] ) );
  XOR U9028 ( .A(\w3[5][118] ), .B(key[893]), .Z(n6612) );
  XOR U9029 ( .A(n6610), .B(\w3[5][126] ), .Z(n6611) );
  XNOR U9030 ( .A(n6612), .B(n6611), .Z(n6613) );
  XOR U9031 ( .A(\w3[5][101] ), .B(n6613), .Z(\w1[6][125] ) );
  XNOR U9032 ( .A(n6614), .B(key[894]), .Z(n6617) );
  XOR U9033 ( .A(\w3[5][102] ), .B(n6615), .Z(n6616) );
  XNOR U9034 ( .A(n6617), .B(n6616), .Z(\w1[6][126] ) );
  XNOR U9035 ( .A(n6920), .B(key[895]), .Z(n6620) );
  XOR U9036 ( .A(\w3[5][103] ), .B(n6618), .Z(n6619) );
  XNOR U9037 ( .A(n6620), .B(n6619), .Z(\w1[6][127] ) );
  XOR U9038 ( .A(\w3[5][13] ), .B(\w3[5][28] ), .Z(n6622) );
  XNOR U9039 ( .A(\w3[5][8] ), .B(\w3[5][4] ), .Z(n6621) );
  XOR U9040 ( .A(n6622), .B(n6621), .Z(n6644) );
  XNOR U9041 ( .A(n6644), .B(key[780]), .Z(n6624) );
  XNOR U9042 ( .A(\w3[5][0] ), .B(\w3[5][5] ), .Z(n6739) );
  XOR U9043 ( .A(\w3[5][20] ), .B(n6739), .Z(n6623) );
  XNOR U9044 ( .A(n6624), .B(n6623), .Z(\w1[6][12] ) );
  IV U9045 ( .A(\w3[5][21] ), .Z(n6669) );
  XNOR U9046 ( .A(\w3[5][14] ), .B(n6669), .Z(n6626) );
  XNOR U9047 ( .A(\w3[5][5] ), .B(\w3[5][29] ), .Z(n6647) );
  XOR U9048 ( .A(n6647), .B(key[781]), .Z(n6625) );
  XNOR U9049 ( .A(n6626), .B(n6625), .Z(n6627) );
  XOR U9050 ( .A(\w3[5][6] ), .B(n6627), .Z(\w1[6][13] ) );
  IV U9051 ( .A(\w3[5][30] ), .Z(n6816) );
  XOR U9052 ( .A(\w3[5][6] ), .B(n6816), .Z(n6781) );
  XOR U9053 ( .A(\w3[5][8] ), .B(\w3[5][15] ), .Z(n6650) );
  XNOR U9054 ( .A(n6781), .B(n6650), .Z(n6648) );
  XOR U9055 ( .A(n6648), .B(key[782]), .Z(n6629) );
  XNOR U9056 ( .A(\w3[5][0] ), .B(\w3[5][7] ), .Z(n6817) );
  XOR U9057 ( .A(\w3[5][22] ), .B(n6817), .Z(n6628) );
  XNOR U9058 ( .A(n6629), .B(n6628), .Z(\w1[6][14] ) );
  XNOR U9059 ( .A(\w3[5][7] ), .B(\w3[5][31] ), .Z(n6649) );
  XNOR U9060 ( .A(n6649), .B(key[783]), .Z(n6631) );
  XOR U9061 ( .A(\w3[5][8] ), .B(\w3[5][0] ), .Z(n6653) );
  XNOR U9062 ( .A(\w3[5][23] ), .B(n6653), .Z(n6630) );
  XNOR U9063 ( .A(n6631), .B(n6630), .Z(\w1[6][15] ) );
  XNOR U9064 ( .A(\w3[5][17] ), .B(\w3[5][9] ), .Z(n6655) );
  XNOR U9065 ( .A(n6655), .B(key[784]), .Z(n6633) );
  XNOR U9066 ( .A(\w3[5][24] ), .B(n6653), .Z(n6632) );
  XNOR U9067 ( .A(n6633), .B(n6632), .Z(\w1[6][16] ) );
  XNOR U9068 ( .A(\w3[5][18] ), .B(\w3[5][10] ), .Z(n6674) );
  XNOR U9069 ( .A(n6674), .B(key[785]), .Z(n6635) );
  IV U9070 ( .A(\w3[5][9] ), .Z(n6888) );
  XNOR U9071 ( .A(n6940), .B(n6888), .Z(n6634) );
  XNOR U9072 ( .A(n6635), .B(n6634), .Z(\w1[6][17] ) );
  XNOR U9073 ( .A(\w3[5][11] ), .B(\w3[5][19] ), .Z(n6660) );
  XNOR U9074 ( .A(n6660), .B(key[786]), .Z(n6637) );
  XOR U9075 ( .A(n6641), .B(\w3[5][10] ), .Z(n6636) );
  XNOR U9076 ( .A(n6637), .B(n6636), .Z(\w1[6][18] ) );
  XOR U9077 ( .A(n6654), .B(\w3[5][20] ), .Z(n6661) );
  XNOR U9078 ( .A(n6661), .B(key[787]), .Z(n6640) );
  XOR U9079 ( .A(\w3[5][11] ), .B(n6638), .Z(n6639) );
  XNOR U9080 ( .A(n6640), .B(n6639), .Z(\w1[6][19] ) );
  XNOR U9081 ( .A(n6655), .B(key[769]), .Z(n6643) );
  XOR U9082 ( .A(\w3[5][25] ), .B(n6641), .Z(n6642) );
  XNOR U9083 ( .A(n6643), .B(n6642), .Z(\w1[6][1] ) );
  XOR U9084 ( .A(\w3[5][16] ), .B(n6669), .Z(n6666) );
  XNOR U9085 ( .A(n6666), .B(key[788]), .Z(n6646) );
  XOR U9086 ( .A(\w3[5][12] ), .B(n6644), .Z(n6645) );
  XNOR U9087 ( .A(n6646), .B(n6645), .Z(\w1[6][20] ) );
  IV U9088 ( .A(\w3[5][22] ), .Z(n6670) );
  XOR U9089 ( .A(\w3[5][14] ), .B(n6670), .Z(n6679) );
  XOR U9090 ( .A(n6654), .B(\w3[5][23] ), .Z(n6680) );
  XNOR U9091 ( .A(n6649), .B(key[791]), .Z(n6652) );
  XNOR U9092 ( .A(\w3[5][16] ), .B(n6650), .Z(n6651) );
  XNOR U9093 ( .A(n6652), .B(n6651), .Z(\w1[6][23] ) );
  XNOR U9094 ( .A(n6674), .B(key[794]), .Z(n6657) );
  XNOR U9095 ( .A(\w3[5][2] ), .B(\w3[5][19] ), .Z(n6656) );
  XNOR U9096 ( .A(n6657), .B(n6656), .Z(n6658) );
  XOR U9097 ( .A(\w3[5][27] ), .B(n6658), .Z(\w1[6][26] ) );
  IV U9098 ( .A(\w3[5][24] ), .Z(n6678) );
  XOR U9099 ( .A(n6678), .B(\w3[5][28] ), .Z(n6659) );
  XOR U9100 ( .A(n6660), .B(n6659), .Z(n6703) );
  XOR U9101 ( .A(n6703), .B(key[795]), .Z(n6663) );
  XOR U9102 ( .A(\w3[5][3] ), .B(n6661), .Z(n6662) );
  XNOR U9103 ( .A(n6663), .B(n6662), .Z(\w1[6][27] ) );
  XOR U9104 ( .A(\w3[5][20] ), .B(\w3[5][29] ), .Z(n6665) );
  XOR U9105 ( .A(n6678), .B(\w3[5][12] ), .Z(n6664) );
  XOR U9106 ( .A(n6665), .B(n6664), .Z(n6738) );
  XNOR U9107 ( .A(n6738), .B(key[796]), .Z(n6668) );
  XOR U9108 ( .A(\w3[5][4] ), .B(n6666), .Z(n6667) );
  XNOR U9109 ( .A(n6668), .B(n6667), .Z(\w1[6][28] ) );
  XOR U9110 ( .A(\w3[5][13] ), .B(n6669), .Z(n6780) );
  XNOR U9111 ( .A(n6780), .B(key[797]), .Z(n6672) );
  XNOR U9112 ( .A(n6670), .B(n6816), .Z(n6671) );
  XNOR U9113 ( .A(n6672), .B(n6671), .Z(n6673) );
  XOR U9114 ( .A(\w3[5][5] ), .B(n6673), .Z(\w1[6][29] ) );
  XNOR U9115 ( .A(n6674), .B(key[770]), .Z(n6677) );
  XOR U9116 ( .A(\w3[5][26] ), .B(n6675), .Z(n6676) );
  XNOR U9117 ( .A(n6677), .B(n6676), .Z(\w1[6][2] ) );
  XOR U9118 ( .A(n6678), .B(\w3[5][31] ), .Z(n6852) );
  XNOR U9119 ( .A(n6679), .B(n6852), .Z(n6815) );
  XNOR U9120 ( .A(\w3[5][15] ), .B(\w3[5][23] ), .Z(n6851) );
  XNOR U9121 ( .A(n6851), .B(key[799]), .Z(n6682) );
  XOR U9122 ( .A(n6891), .B(\w3[5][7] ), .Z(n6681) );
  XNOR U9123 ( .A(n6682), .B(n6681), .Z(\w1[6][31] ) );
  XOR U9124 ( .A(\w3[5][33] ), .B(\w3[5][57] ), .Z(n6735) );
  XOR U9125 ( .A(n6735), .B(key[800]), .Z(n6684) );
  XNOR U9126 ( .A(\w3[5][48] ), .B(\w3[5][56] ), .Z(n6797) );
  XOR U9127 ( .A(n6797), .B(\w3[5][40] ), .Z(n6683) );
  XNOR U9128 ( .A(n6684), .B(n6683), .Z(\w1[6][32] ) );
  XNOR U9129 ( .A(\w3[5][34] ), .B(\w3[5][58] ), .Z(n6743) );
  XOR U9130 ( .A(\w3[5][57] ), .B(\w3[5][49] ), .Z(n6761) );
  XNOR U9131 ( .A(n6761), .B(key[801]), .Z(n6685) );
  XNOR U9132 ( .A(n6743), .B(n6685), .Z(n6686) );
  XNOR U9133 ( .A(\w3[5][41] ), .B(n6686), .Z(\w1[6][33] ) );
  XNOR U9134 ( .A(n6713), .B(key[802]), .Z(n6688) );
  XNOR U9135 ( .A(\w3[5][50] ), .B(\w3[5][42] ), .Z(n6771) );
  XOR U9136 ( .A(\w3[5][58] ), .B(n6771), .Z(n6687) );
  XNOR U9137 ( .A(n6688), .B(n6687), .Z(\w1[6][34] ) );
  XOR U9138 ( .A(\w3[5][36] ), .B(\w3[5][32] ), .Z(n6715) );
  XOR U9139 ( .A(n6715), .B(key[803]), .Z(n6691) );
  IV U9140 ( .A(\w3[5][51] ), .Z(n6770) );
  XOR U9141 ( .A(\w3[5][43] ), .B(n6770), .Z(n6742) );
  XOR U9142 ( .A(\w3[5][56] ), .B(n6742), .Z(n6689) );
  XNOR U9143 ( .A(\w3[5][60] ), .B(n6689), .Z(n6776) );
  XNOR U9144 ( .A(\w3[5][59] ), .B(n6776), .Z(n6690) );
  XNOR U9145 ( .A(n6691), .B(n6690), .Z(\w1[6][35] ) );
  XOR U9146 ( .A(\w3[5][32] ), .B(\w3[5][37] ), .Z(n6721) );
  XOR U9147 ( .A(\w3[5][52] ), .B(\w3[5][61] ), .Z(n6693) );
  XNOR U9148 ( .A(\w3[5][56] ), .B(\w3[5][44] ), .Z(n6692) );
  XOR U9149 ( .A(n6693), .B(n6692), .Z(n6785) );
  XOR U9150 ( .A(n6785), .B(key[804]), .Z(n6694) );
  XOR U9151 ( .A(n6721), .B(n6694), .Z(n6695) );
  XNOR U9152 ( .A(\w3[5][60] ), .B(n6695), .Z(\w1[6][36] ) );
  XNOR U9153 ( .A(\w3[5][38] ), .B(\w3[5][62] ), .Z(n6727) );
  XNOR U9154 ( .A(n6727), .B(key[805]), .Z(n6697) );
  IV U9155 ( .A(\w3[5][45] ), .Z(n6750) );
  XOR U9156 ( .A(\w3[5][53] ), .B(n6750), .Z(n6788) );
  XOR U9157 ( .A(\w3[5][61] ), .B(n6788), .Z(n6696) );
  XNOR U9158 ( .A(n6697), .B(n6696), .Z(\w1[6][37] ) );
  XOR U9159 ( .A(\w3[5][32] ), .B(\w3[5][39] ), .Z(n6728) );
  XOR U9160 ( .A(n6728), .B(key[806]), .Z(n6699) );
  XNOR U9161 ( .A(\w3[5][56] ), .B(\w3[5][63] ), .Z(n6700) );
  XOR U9162 ( .A(\w3[5][46] ), .B(\w3[5][54] ), .Z(n6749) );
  XOR U9163 ( .A(n6700), .B(n6749), .Z(n6793) );
  XOR U9164 ( .A(\w3[5][62] ), .B(n6793), .Z(n6698) );
  XNOR U9165 ( .A(n6699), .B(n6698), .Z(\w1[6][38] ) );
  XNOR U9166 ( .A(\w3[5][55] ), .B(\w3[5][47] ), .Z(n6796) );
  XNOR U9167 ( .A(n6796), .B(key[807]), .Z(n6702) );
  XOR U9168 ( .A(\w3[5][32] ), .B(n6700), .Z(n6701) );
  XNOR U9169 ( .A(n6702), .B(n6701), .Z(\w1[6][39] ) );
  XOR U9170 ( .A(n6703), .B(key[771]), .Z(n6706) );
  XOR U9171 ( .A(n6704), .B(\w3[5][27] ), .Z(n6705) );
  XNOR U9172 ( .A(n6706), .B(n6705), .Z(\w1[6][3] ) );
  IV U9173 ( .A(\w3[5][33] ), .Z(n6766) );
  XOR U9174 ( .A(\w3[5][42] ), .B(key[809]), .Z(n6708) );
  XNOR U9175 ( .A(n6761), .B(\w3[5][34] ), .Z(n6707) );
  XNOR U9176 ( .A(n6708), .B(n6707), .Z(n6709) );
  XNOR U9177 ( .A(n6766), .B(n6709), .Z(\w1[6][41] ) );
  XOR U9178 ( .A(\w3[5][43] ), .B(key[810]), .Z(n6711) );
  IV U9179 ( .A(\w3[5][35] ), .Z(n6777) );
  XOR U9180 ( .A(\w3[5][50] ), .B(n6777), .Z(n6710) );
  XNOR U9181 ( .A(n6711), .B(n6710), .Z(n6712) );
  XNOR U9182 ( .A(n6712), .B(n6743), .Z(\w1[6][42] ) );
  IV U9183 ( .A(\w3[5][40] ), .Z(n6718) );
  XNOR U9184 ( .A(n6718), .B(n6713), .Z(n6714) );
  XOR U9185 ( .A(\w3[5][44] ), .B(n6714), .Z(n6744) );
  XNOR U9186 ( .A(n6744), .B(key[811]), .Z(n6717) );
  XNOR U9187 ( .A(\w3[5][51] ), .B(n6715), .Z(n6716) );
  XNOR U9188 ( .A(n6717), .B(n6716), .Z(\w1[6][43] ) );
  XOR U9189 ( .A(\w3[5][36] ), .B(\w3[5][45] ), .Z(n6720) );
  XOR U9190 ( .A(n6718), .B(\w3[5][60] ), .Z(n6719) );
  XOR U9191 ( .A(n6720), .B(n6719), .Z(n6745) );
  XNOR U9192 ( .A(n6745), .B(key[812]), .Z(n6723) );
  XNOR U9193 ( .A(\w3[5][52] ), .B(n6721), .Z(n6722) );
  XNOR U9194 ( .A(n6723), .B(n6722), .Z(\w1[6][44] ) );
  XNOR U9195 ( .A(\w3[5][61] ), .B(\w3[5][37] ), .Z(n6748) );
  XNOR U9196 ( .A(n6748), .B(key[813]), .Z(n6725) );
  XNOR U9197 ( .A(\w3[5][38] ), .B(\w3[5][46] ), .Z(n6724) );
  XNOR U9198 ( .A(n6725), .B(n6724), .Z(n6726) );
  XOR U9199 ( .A(\w3[5][53] ), .B(n6726), .Z(\w1[6][45] ) );
  XOR U9200 ( .A(\w3[5][40] ), .B(\w3[5][47] ), .Z(n6757) );
  XOR U9201 ( .A(n6727), .B(n6757), .Z(n6753) );
  XNOR U9202 ( .A(n6753), .B(key[814]), .Z(n6730) );
  XNOR U9203 ( .A(\w3[5][54] ), .B(n6728), .Z(n6729) );
  XNOR U9204 ( .A(n6730), .B(n6729), .Z(\w1[6][46] ) );
  XOR U9205 ( .A(\w3[5][63] ), .B(\w3[5][39] ), .Z(n6756) );
  XOR U9206 ( .A(n6756), .B(key[815]), .Z(n6732) );
  XNOR U9207 ( .A(\w3[5][40] ), .B(\w3[5][32] ), .Z(n6760) );
  XOR U9208 ( .A(\w3[5][55] ), .B(n6760), .Z(n6731) );
  XNOR U9209 ( .A(n6732), .B(n6731), .Z(\w1[6][47] ) );
  XNOR U9210 ( .A(\w3[5][41] ), .B(\w3[5][49] ), .Z(n6765) );
  XNOR U9211 ( .A(n6765), .B(key[816]), .Z(n6734) );
  XOR U9212 ( .A(\w3[5][56] ), .B(n6760), .Z(n6733) );
  XNOR U9213 ( .A(n6734), .B(n6733), .Z(\w1[6][48] ) );
  XNOR U9214 ( .A(n6771), .B(key[817]), .Z(n6737) );
  XNOR U9215 ( .A(n6735), .B(\w3[5][41] ), .Z(n6736) );
  XNOR U9216 ( .A(n6737), .B(n6736), .Z(\w1[6][49] ) );
  XNOR U9217 ( .A(n6738), .B(key[772]), .Z(n6741) );
  XOR U9218 ( .A(n6739), .B(\w3[5][28] ), .Z(n6740) );
  XNOR U9219 ( .A(n6741), .B(n6740), .Z(\w1[6][4] ) );
  IV U9220 ( .A(\w3[5][48] ), .Z(n6762) );
  XOR U9221 ( .A(n6762), .B(\w3[5][52] ), .Z(n6775) );
  XNOR U9222 ( .A(n6784), .B(key[820]), .Z(n6747) );
  XOR U9223 ( .A(\w3[5][44] ), .B(n6745), .Z(n6746) );
  XNOR U9224 ( .A(n6747), .B(n6746), .Z(\w1[6][52] ) );
  XNOR U9225 ( .A(n6748), .B(key[821]), .Z(n6752) );
  XOR U9226 ( .A(n6750), .B(n6749), .Z(n6751) );
  XNOR U9227 ( .A(n6752), .B(n6751), .Z(\w1[6][53] ) );
  XOR U9228 ( .A(n6762), .B(\w3[5][55] ), .Z(n6792) );
  XNOR U9229 ( .A(n6792), .B(key[822]), .Z(n6755) );
  XOR U9230 ( .A(\w3[5][46] ), .B(n6753), .Z(n6754) );
  XNOR U9231 ( .A(n6755), .B(n6754), .Z(\w1[6][54] ) );
  XOR U9232 ( .A(n6756), .B(key[823]), .Z(n6759) );
  XNOR U9233 ( .A(\w3[5][48] ), .B(n6757), .Z(n6758) );
  XNOR U9234 ( .A(n6759), .B(n6758), .Z(\w1[6][55] ) );
  XNOR U9235 ( .A(n6760), .B(key[824]), .Z(n6764) );
  XOR U9236 ( .A(n6762), .B(n6761), .Z(n6763) );
  XNOR U9237 ( .A(n6764), .B(n6763), .Z(\w1[6][56] ) );
  XNOR U9238 ( .A(n6765), .B(key[825]), .Z(n6768) );
  XOR U9239 ( .A(n6766), .B(\w3[5][50] ), .Z(n6767) );
  XNOR U9240 ( .A(n6768), .B(n6767), .Z(n6769) );
  XOR U9241 ( .A(\w3[5][58] ), .B(n6769), .Z(\w1[6][57] ) );
  XNOR U9242 ( .A(n6770), .B(key[826]), .Z(n6773) );
  XOR U9243 ( .A(n6771), .B(\w3[5][59] ), .Z(n6772) );
  XNOR U9244 ( .A(n6773), .B(n6772), .Z(n6774) );
  XOR U9245 ( .A(\w3[5][34] ), .B(n6774), .Z(\w1[6][58] ) );
  XNOR U9246 ( .A(n6775), .B(key[827]), .Z(n6779) );
  XOR U9247 ( .A(n6777), .B(n6776), .Z(n6778) );
  XNOR U9248 ( .A(n6779), .B(n6778), .Z(\w1[6][59] ) );
  XNOR U9249 ( .A(n6780), .B(key[773]), .Z(n6783) );
  XOR U9250 ( .A(\w3[5][29] ), .B(n6781), .Z(n6782) );
  XNOR U9251 ( .A(n6783), .B(n6782), .Z(\w1[6][5] ) );
  XNOR U9252 ( .A(n6784), .B(key[828]), .Z(n6787) );
  XOR U9253 ( .A(\w3[5][36] ), .B(n6785), .Z(n6786) );
  XNOR U9254 ( .A(n6787), .B(n6786), .Z(\w1[6][60] ) );
  XOR U9255 ( .A(\w3[5][54] ), .B(key[829]), .Z(n6790) );
  XOR U9256 ( .A(n6788), .B(\w3[5][62] ), .Z(n6789) );
  XNOR U9257 ( .A(n6790), .B(n6789), .Z(n6791) );
  XOR U9258 ( .A(\w3[5][37] ), .B(n6791), .Z(\w1[6][61] ) );
  XNOR U9259 ( .A(n6792), .B(key[830]), .Z(n6795) );
  XOR U9260 ( .A(\w3[5][38] ), .B(n6793), .Z(n6794) );
  XNOR U9261 ( .A(n6795), .B(n6794), .Z(\w1[6][62] ) );
  XNOR U9262 ( .A(n6796), .B(key[831]), .Z(n6799) );
  XOR U9263 ( .A(n6797), .B(\w3[5][39] ), .Z(n6798) );
  XNOR U9264 ( .A(n6799), .B(n6798), .Z(\w1[6][63] ) );
  XOR U9265 ( .A(\w3[5][65] ), .B(\w3[5][89] ), .Z(n6857) );
  XOR U9266 ( .A(n6857), .B(key[832]), .Z(n6801) );
  XNOR U9267 ( .A(\w3[5][80] ), .B(\w3[5][88] ), .Z(n6916) );
  XOR U9268 ( .A(n6916), .B(\w3[5][72] ), .Z(n6800) );
  XNOR U9269 ( .A(n6801), .B(n6800), .Z(\w1[6][64] ) );
  XNOR U9270 ( .A(\w3[5][66] ), .B(\w3[5][90] ), .Z(n6861) );
  XOR U9271 ( .A(\w3[5][89] ), .B(\w3[5][81] ), .Z(n6879) );
  XNOR U9272 ( .A(n6879), .B(key[833]), .Z(n6802) );
  XNOR U9273 ( .A(n6861), .B(n6802), .Z(n6803) );
  XNOR U9274 ( .A(\w3[5][73] ), .B(n6803), .Z(\w1[6][65] ) );
  XNOR U9275 ( .A(n6831), .B(key[834]), .Z(n6805) );
  XNOR U9276 ( .A(\w3[5][82] ), .B(\w3[5][74] ), .Z(n6894) );
  XOR U9277 ( .A(\w3[5][90] ), .B(n6894), .Z(n6804) );
  XNOR U9278 ( .A(n6805), .B(n6804), .Z(\w1[6][66] ) );
  XOR U9279 ( .A(\w3[5][68] ), .B(\w3[5][64] ), .Z(n6833) );
  XOR U9280 ( .A(n6833), .B(key[835]), .Z(n6808) );
  IV U9281 ( .A(\w3[5][83] ), .Z(n6893) );
  XOR U9282 ( .A(\w3[5][75] ), .B(n6893), .Z(n6860) );
  XOR U9283 ( .A(\w3[5][88] ), .B(n6860), .Z(n6806) );
  XNOR U9284 ( .A(\w3[5][92] ), .B(n6806), .Z(n6899) );
  XNOR U9285 ( .A(\w3[5][91] ), .B(n6899), .Z(n6807) );
  XNOR U9286 ( .A(n6808), .B(n6807), .Z(\w1[6][67] ) );
  XOR U9287 ( .A(\w3[5][64] ), .B(\w3[5][69] ), .Z(n6839) );
  XOR U9288 ( .A(\w3[5][84] ), .B(\w3[5][93] ), .Z(n6810) );
  XNOR U9289 ( .A(\w3[5][88] ), .B(\w3[5][76] ), .Z(n6809) );
  XOR U9290 ( .A(n6810), .B(n6809), .Z(n6904) );
  XOR U9291 ( .A(n6904), .B(key[836]), .Z(n6811) );
  XOR U9292 ( .A(n6839), .B(n6811), .Z(n6812) );
  XNOR U9293 ( .A(\w3[5][92] ), .B(n6812), .Z(\w1[6][68] ) );
  XNOR U9294 ( .A(\w3[5][70] ), .B(\w3[5][94] ), .Z(n6845) );
  XNOR U9295 ( .A(n6845), .B(key[837]), .Z(n6814) );
  IV U9296 ( .A(\w3[5][77] ), .Z(n6868) );
  XOR U9297 ( .A(\w3[5][85] ), .B(n6868), .Z(n6907) );
  XOR U9298 ( .A(\w3[5][93] ), .B(n6907), .Z(n6813) );
  XNOR U9299 ( .A(n6814), .B(n6813), .Z(\w1[6][69] ) );
  XNOR U9300 ( .A(n6815), .B(key[774]), .Z(n6819) );
  XNOR U9301 ( .A(n6817), .B(n6816), .Z(n6818) );
  XNOR U9302 ( .A(n6819), .B(n6818), .Z(\w1[6][6] ) );
  XOR U9303 ( .A(\w3[5][64] ), .B(\w3[5][71] ), .Z(n6846) );
  XOR U9304 ( .A(n6846), .B(key[838]), .Z(n6821) );
  XNOR U9305 ( .A(\w3[5][88] ), .B(\w3[5][95] ), .Z(n6822) );
  XOR U9306 ( .A(\w3[5][78] ), .B(\w3[5][86] ), .Z(n6867) );
  XOR U9307 ( .A(n6822), .B(n6867), .Z(n6912) );
  XOR U9308 ( .A(\w3[5][94] ), .B(n6912), .Z(n6820) );
  XNOR U9309 ( .A(n6821), .B(n6820), .Z(\w1[6][70] ) );
  XNOR U9310 ( .A(\w3[5][79] ), .B(\w3[5][87] ), .Z(n6915) );
  XNOR U9311 ( .A(n6915), .B(key[839]), .Z(n6824) );
  XOR U9312 ( .A(\w3[5][64] ), .B(n6822), .Z(n6823) );
  XNOR U9313 ( .A(n6824), .B(n6823), .Z(\w1[6][71] ) );
  IV U9314 ( .A(\w3[5][65] ), .Z(n6884) );
  XOR U9315 ( .A(\w3[5][74] ), .B(key[841]), .Z(n6826) );
  XNOR U9316 ( .A(n6879), .B(\w3[5][66] ), .Z(n6825) );
  XNOR U9317 ( .A(n6826), .B(n6825), .Z(n6827) );
  XNOR U9318 ( .A(n6884), .B(n6827), .Z(\w1[6][73] ) );
  XOR U9319 ( .A(\w3[5][75] ), .B(key[842]), .Z(n6829) );
  IV U9320 ( .A(\w3[5][67] ), .Z(n6900) );
  XOR U9321 ( .A(\w3[5][82] ), .B(n6900), .Z(n6828) );
  XNOR U9322 ( .A(n6829), .B(n6828), .Z(n6830) );
  XNOR U9323 ( .A(n6830), .B(n6861), .Z(\w1[6][74] ) );
  IV U9324 ( .A(\w3[5][72] ), .Z(n6836) );
  XNOR U9325 ( .A(n6836), .B(n6831), .Z(n6832) );
  XOR U9326 ( .A(\w3[5][76] ), .B(n6832), .Z(n6862) );
  XNOR U9327 ( .A(n6862), .B(key[843]), .Z(n6835) );
  XNOR U9328 ( .A(\w3[5][83] ), .B(n6833), .Z(n6834) );
  XNOR U9329 ( .A(n6835), .B(n6834), .Z(\w1[6][75] ) );
  XOR U9330 ( .A(\w3[5][68] ), .B(\w3[5][77] ), .Z(n6838) );
  XOR U9331 ( .A(n6836), .B(\w3[5][92] ), .Z(n6837) );
  XOR U9332 ( .A(n6838), .B(n6837), .Z(n6863) );
  XNOR U9333 ( .A(n6863), .B(key[844]), .Z(n6841) );
  XNOR U9334 ( .A(\w3[5][84] ), .B(n6839), .Z(n6840) );
  XNOR U9335 ( .A(n6841), .B(n6840), .Z(\w1[6][76] ) );
  XNOR U9336 ( .A(\w3[5][93] ), .B(\w3[5][69] ), .Z(n6866) );
  XNOR U9337 ( .A(n6866), .B(key[845]), .Z(n6843) );
  XNOR U9338 ( .A(\w3[5][70] ), .B(\w3[5][78] ), .Z(n6842) );
  XNOR U9339 ( .A(n6843), .B(n6842), .Z(n6844) );
  XOR U9340 ( .A(\w3[5][85] ), .B(n6844), .Z(\w1[6][77] ) );
  XOR U9341 ( .A(\w3[5][72] ), .B(\w3[5][79] ), .Z(n6875) );
  XOR U9342 ( .A(n6845), .B(n6875), .Z(n6871) );
  XNOR U9343 ( .A(n6871), .B(key[846]), .Z(n6848) );
  XNOR U9344 ( .A(\w3[5][86] ), .B(n6846), .Z(n6847) );
  XNOR U9345 ( .A(n6848), .B(n6847), .Z(\w1[6][78] ) );
  XOR U9346 ( .A(\w3[5][95] ), .B(\w3[5][71] ), .Z(n6874) );
  XOR U9347 ( .A(n6874), .B(key[847]), .Z(n6850) );
  XNOR U9348 ( .A(\w3[5][72] ), .B(\w3[5][64] ), .Z(n6878) );
  XOR U9349 ( .A(\w3[5][87] ), .B(n6878), .Z(n6849) );
  XNOR U9350 ( .A(n6850), .B(n6849), .Z(\w1[6][79] ) );
  XNOR U9351 ( .A(n6851), .B(key[775]), .Z(n6854) );
  XOR U9352 ( .A(\w3[5][0] ), .B(n6852), .Z(n6853) );
  XNOR U9353 ( .A(n6854), .B(n6853), .Z(\w1[6][7] ) );
  XNOR U9354 ( .A(\w3[5][73] ), .B(\w3[5][81] ), .Z(n6883) );
  XNOR U9355 ( .A(n6883), .B(key[848]), .Z(n6856) );
  XOR U9356 ( .A(\w3[5][88] ), .B(n6878), .Z(n6855) );
  XNOR U9357 ( .A(n6856), .B(n6855), .Z(\w1[6][80] ) );
  XNOR U9358 ( .A(n6894), .B(key[849]), .Z(n6859) );
  XNOR U9359 ( .A(n6857), .B(\w3[5][73] ), .Z(n6858) );
  XNOR U9360 ( .A(n6859), .B(n6858), .Z(\w1[6][81] ) );
  IV U9361 ( .A(\w3[5][80] ), .Z(n6880) );
  XOR U9362 ( .A(n6880), .B(\w3[5][84] ), .Z(n6898) );
  XNOR U9363 ( .A(n6903), .B(key[852]), .Z(n6865) );
  XOR U9364 ( .A(\w3[5][76] ), .B(n6863), .Z(n6864) );
  XNOR U9365 ( .A(n6865), .B(n6864), .Z(\w1[6][84] ) );
  XNOR U9366 ( .A(n6866), .B(key[853]), .Z(n6870) );
  XOR U9367 ( .A(n6868), .B(n6867), .Z(n6869) );
  XNOR U9368 ( .A(n6870), .B(n6869), .Z(\w1[6][85] ) );
  XOR U9369 ( .A(n6880), .B(\w3[5][87] ), .Z(n6911) );
  XNOR U9370 ( .A(n6911), .B(key[854]), .Z(n6873) );
  XOR U9371 ( .A(\w3[5][78] ), .B(n6871), .Z(n6872) );
  XNOR U9372 ( .A(n6873), .B(n6872), .Z(\w1[6][86] ) );
  XOR U9373 ( .A(n6874), .B(key[855]), .Z(n6877) );
  XNOR U9374 ( .A(\w3[5][80] ), .B(n6875), .Z(n6876) );
  XNOR U9375 ( .A(n6877), .B(n6876), .Z(\w1[6][87] ) );
  XNOR U9376 ( .A(n6878), .B(key[856]), .Z(n6882) );
  XOR U9377 ( .A(n6880), .B(n6879), .Z(n6881) );
  XNOR U9378 ( .A(n6882), .B(n6881), .Z(\w1[6][88] ) );
  XNOR U9379 ( .A(n6883), .B(key[857]), .Z(n6886) );
  XOR U9380 ( .A(n6884), .B(\w3[5][82] ), .Z(n6885) );
  XNOR U9381 ( .A(n6886), .B(n6885), .Z(n6887) );
  XOR U9382 ( .A(\w3[5][90] ), .B(n6887), .Z(\w1[6][89] ) );
  XNOR U9383 ( .A(n6888), .B(key[776]), .Z(n6890) );
  XNOR U9384 ( .A(\w3[5][1] ), .B(\w3[5][0] ), .Z(n6889) );
  XNOR U9385 ( .A(n6890), .B(n6889), .Z(n6892) );
  XNOR U9386 ( .A(n6892), .B(n6891), .Z(\w1[6][8] ) );
  XNOR U9387 ( .A(n6893), .B(key[858]), .Z(n6896) );
  XOR U9388 ( .A(n6894), .B(\w3[5][91] ), .Z(n6895) );
  XNOR U9389 ( .A(n6896), .B(n6895), .Z(n6897) );
  XOR U9390 ( .A(\w3[5][66] ), .B(n6897), .Z(\w1[6][90] ) );
  XNOR U9391 ( .A(n6898), .B(key[859]), .Z(n6902) );
  XOR U9392 ( .A(n6900), .B(n6899), .Z(n6901) );
  XNOR U9393 ( .A(n6902), .B(n6901), .Z(\w1[6][91] ) );
  XNOR U9394 ( .A(n6903), .B(key[860]), .Z(n6906) );
  XOR U9395 ( .A(\w3[5][68] ), .B(n6904), .Z(n6905) );
  XNOR U9396 ( .A(n6906), .B(n6905), .Z(\w1[6][92] ) );
  XOR U9397 ( .A(\w3[5][86] ), .B(key[861]), .Z(n6909) );
  XOR U9398 ( .A(n6907), .B(\w3[5][94] ), .Z(n6908) );
  XNOR U9399 ( .A(n6909), .B(n6908), .Z(n6910) );
  XOR U9400 ( .A(\w3[5][69] ), .B(n6910), .Z(\w1[6][93] ) );
  XNOR U9401 ( .A(n6911), .B(key[862]), .Z(n6914) );
  XOR U9402 ( .A(\w3[5][70] ), .B(n6912), .Z(n6913) );
  XNOR U9403 ( .A(n6914), .B(n6913), .Z(\w1[6][94] ) );
  XNOR U9404 ( .A(n6915), .B(key[863]), .Z(n6918) );
  XOR U9405 ( .A(n6916), .B(\w3[5][71] ), .Z(n6917) );
  XNOR U9406 ( .A(n6918), .B(n6917), .Z(\w1[6][95] ) );
  XOR U9407 ( .A(\w3[5][104] ), .B(key[864]), .Z(n6922) );
  XNOR U9408 ( .A(n6920), .B(n6919), .Z(n6921) );
  XNOR U9409 ( .A(n6922), .B(n6921), .Z(\w1[6][96] ) );
  XNOR U9410 ( .A(n6923), .B(key[865]), .Z(n6926) );
  XNOR U9411 ( .A(\w3[5][121] ), .B(n6924), .Z(n6925) );
  XNOR U9412 ( .A(n6926), .B(n6925), .Z(\w1[6][97] ) );
  XNOR U9413 ( .A(n6927), .B(key[866]), .Z(n6931) );
  XNOR U9414 ( .A(n6929), .B(n6928), .Z(n6930) );
  XNOR U9415 ( .A(n6931), .B(n6930), .Z(\w1[6][98] ) );
  XOR U9416 ( .A(n6932), .B(key[867]), .Z(n6936) );
  XNOR U9417 ( .A(n6934), .B(n6933), .Z(n6935) );
  XNOR U9418 ( .A(n6936), .B(n6935), .Z(\w1[6][99] ) );
  XOR U9419 ( .A(\w3[5][10] ), .B(key[777]), .Z(n6938) );
  XNOR U9420 ( .A(\w3[5][2] ), .B(\w3[5][17] ), .Z(n6937) );
  XNOR U9421 ( .A(n6938), .B(n6937), .Z(n6939) );
  XNOR U9422 ( .A(n6940), .B(n6939), .Z(\w1[6][9] ) );
  XNOR U9423 ( .A(\w3[6][25] ), .B(\w3[6][1] ), .Z(n7352) );
  IV U9424 ( .A(\w3[6][16] ), .Z(n7068) );
  XOR U9425 ( .A(\w3[6][24] ), .B(n7068), .Z(n7305) );
  XNOR U9426 ( .A(\w3[6][8] ), .B(key[896]), .Z(n6941) );
  XNOR U9427 ( .A(n7305), .B(n6941), .Z(n6942) );
  XOR U9428 ( .A(n7352), .B(n6942), .Z(\w1[7][0] ) );
  XOR U9429 ( .A(\w3[6][96] ), .B(\w3[6][101] ), .Z(n6964) );
  XOR U9430 ( .A(\w3[6][116] ), .B(\w3[6][125] ), .Z(n6944) );
  IV U9431 ( .A(\w3[6][120] ), .Z(n7013) );
  XOR U9432 ( .A(n7013), .B(\w3[6][108] ), .Z(n6943) );
  XOR U9433 ( .A(n6944), .B(n6943), .Z(n7021) );
  XOR U9434 ( .A(n7021), .B(key[996]), .Z(n6945) );
  XOR U9435 ( .A(n6964), .B(n6945), .Z(n6946) );
  XNOR U9436 ( .A(\w3[6][124] ), .B(n6946), .Z(\w1[7][100] ) );
  XNOR U9437 ( .A(\w3[6][102] ), .B(\w3[6][126] ), .Z(n6973) );
  XNOR U9438 ( .A(n6973), .B(key[997]), .Z(n6948) );
  XNOR U9439 ( .A(\w3[6][109] ), .B(\w3[6][117] ), .Z(n7024) );
  XOR U9440 ( .A(\w3[6][125] ), .B(n7024), .Z(n6947) );
  XNOR U9441 ( .A(n6948), .B(n6947), .Z(\w1[7][101] ) );
  XOR U9442 ( .A(\w3[6][96] ), .B(\w3[6][103] ), .Z(n6974) );
  XOR U9443 ( .A(n6974), .B(key[998]), .Z(n6950) );
  XOR U9444 ( .A(n7013), .B(\w3[6][127] ), .Z(n6951) );
  XOR U9445 ( .A(\w3[6][110] ), .B(\w3[6][118] ), .Z(n6990) );
  XOR U9446 ( .A(n6951), .B(n6990), .Z(n7029) );
  XOR U9447 ( .A(\w3[6][126] ), .B(n7029), .Z(n6949) );
  XNOR U9448 ( .A(n6950), .B(n6949), .Z(\w1[7][102] ) );
  XNOR U9449 ( .A(\w3[6][111] ), .B(\w3[6][119] ), .Z(n7032) );
  XNOR U9450 ( .A(n7032), .B(key[999]), .Z(n6953) );
  XOR U9451 ( .A(\w3[6][96] ), .B(n6951), .Z(n6952) );
  XNOR U9452 ( .A(n6953), .B(n6952), .Z(\w1[7][103] ) );
  XNOR U9453 ( .A(\w3[6][120] ), .B(\w3[6][112] ), .Z(n7334) );
  XOR U9454 ( .A(\w3[6][106] ), .B(\w3[6][98] ), .Z(n7011) );
  XOR U9455 ( .A(\w3[6][97] ), .B(\w3[6][121] ), .Z(n7333) );
  XNOR U9456 ( .A(n7333), .B(key[1001]), .Z(n6954) );
  XOR U9457 ( .A(n7011), .B(n6954), .Z(n6955) );
  XNOR U9458 ( .A(\w3[6][113] ), .B(n6955), .Z(\w1[7][105] ) );
  XOR U9459 ( .A(\w3[6][107] ), .B(\w3[6][99] ), .Z(n6957) );
  XNOR U9460 ( .A(\w3[6][98] ), .B(\w3[6][122] ), .Z(n7338) );
  XOR U9461 ( .A(n7338), .B(key[1002]), .Z(n6956) );
  XNOR U9462 ( .A(n6957), .B(n6956), .Z(n6958) );
  XOR U9463 ( .A(\w3[6][114] ), .B(n6958), .Z(\w1[7][106] ) );
  XNOR U9464 ( .A(\w3[6][99] ), .B(\w3[6][123] ), .Z(n7342) );
  XOR U9465 ( .A(\w3[6][108] ), .B(n7342), .Z(n6959) );
  XOR U9466 ( .A(\w3[6][104] ), .B(n6959), .Z(n6983) );
  XNOR U9467 ( .A(n6983), .B(key[1003]), .Z(n6961) );
  IV U9468 ( .A(\w3[6][100] ), .Z(n7020) );
  XOR U9469 ( .A(\w3[6][96] ), .B(n7020), .Z(n7346) );
  XOR U9470 ( .A(\w3[6][115] ), .B(n7346), .Z(n6960) );
  XNOR U9471 ( .A(n6961), .B(n6960), .Z(\w1[7][107] ) );
  XOR U9472 ( .A(\w3[6][100] ), .B(\w3[6][104] ), .Z(n6963) );
  XNOR U9473 ( .A(\w3[6][124] ), .B(\w3[6][109] ), .Z(n6962) );
  XOR U9474 ( .A(n6963), .B(n6962), .Z(n6986) );
  XNOR U9475 ( .A(n6986), .B(key[1004]), .Z(n6966) );
  XNOR U9476 ( .A(\w3[6][116] ), .B(n6964), .Z(n6965) );
  XNOR U9477 ( .A(n6966), .B(n6965), .Z(\w1[7][108] ) );
  XNOR U9478 ( .A(\w3[6][125] ), .B(\w3[6][101] ), .Z(n6989) );
  XNOR U9479 ( .A(n6989), .B(key[1005]), .Z(n6968) );
  XNOR U9480 ( .A(\w3[6][102] ), .B(\w3[6][110] ), .Z(n6967) );
  XNOR U9481 ( .A(n6968), .B(n6967), .Z(n6969) );
  XOR U9482 ( .A(\w3[6][117] ), .B(n6969), .Z(\w1[7][109] ) );
  XOR U9483 ( .A(\w3[6][11] ), .B(\w3[6][3] ), .Z(n6971) );
  XNOR U9484 ( .A(\w3[6][2] ), .B(\w3[6][26] ), .Z(n7055) );
  XOR U9485 ( .A(n7055), .B(key[906]), .Z(n6970) );
  XNOR U9486 ( .A(n6971), .B(n6970), .Z(n6972) );
  XOR U9487 ( .A(\w3[6][18] ), .B(n6972), .Z(\w1[7][10] ) );
  XOR U9488 ( .A(\w3[6][111] ), .B(\w3[6][104] ), .Z(n6997) );
  XOR U9489 ( .A(n6973), .B(n6997), .Z(n6993) );
  XNOR U9490 ( .A(n6993), .B(key[1006]), .Z(n6976) );
  XNOR U9491 ( .A(\w3[6][118] ), .B(n6974), .Z(n6975) );
  XNOR U9492 ( .A(n6976), .B(n6975), .Z(\w1[7][110] ) );
  XOR U9493 ( .A(\w3[6][127] ), .B(\w3[6][103] ), .Z(n6996) );
  XOR U9494 ( .A(n6996), .B(key[1007]), .Z(n6978) );
  XNOR U9495 ( .A(\w3[6][96] ), .B(\w3[6][104] ), .Z(n7002) );
  XOR U9496 ( .A(\w3[6][119] ), .B(n7002), .Z(n6977) );
  XNOR U9497 ( .A(n6978), .B(n6977), .Z(\w1[7][111] ) );
  XNOR U9498 ( .A(\w3[6][105] ), .B(\w3[6][113] ), .Z(n7337) );
  XNOR U9499 ( .A(n7337), .B(key[1008]), .Z(n6980) );
  XNOR U9500 ( .A(n7013), .B(n7002), .Z(n6979) );
  XNOR U9501 ( .A(n6980), .B(n6979), .Z(\w1[7][112] ) );
  XNOR U9502 ( .A(\w3[6][106] ), .B(\w3[6][114] ), .Z(n7341) );
  XNOR U9503 ( .A(\w3[6][107] ), .B(\w3[6][115] ), .Z(n7015) );
  XNOR U9504 ( .A(n7015), .B(key[1010]), .Z(n6982) );
  XNOR U9505 ( .A(n7011), .B(\w3[6][122] ), .Z(n6981) );
  XNOR U9506 ( .A(n6982), .B(n6981), .Z(\w1[7][114] ) );
  XNOR U9507 ( .A(\w3[6][116] ), .B(\w3[6][112] ), .Z(n7016) );
  XNOR U9508 ( .A(n7016), .B(key[1011]), .Z(n6985) );
  XOR U9509 ( .A(\w3[6][107] ), .B(n6983), .Z(n6984) );
  XNOR U9510 ( .A(n6985), .B(n6984), .Z(\w1[7][115] ) );
  XNOR U9511 ( .A(\w3[6][117] ), .B(\w3[6][112] ), .Z(n7019) );
  XNOR U9512 ( .A(n7019), .B(key[1012]), .Z(n6988) );
  XOR U9513 ( .A(\w3[6][108] ), .B(n6986), .Z(n6987) );
  XNOR U9514 ( .A(n6988), .B(n6987), .Z(\w1[7][116] ) );
  XNOR U9515 ( .A(n6989), .B(key[1013]), .Z(n6992) );
  XNOR U9516 ( .A(\w3[6][109] ), .B(n6990), .Z(n6991) );
  XNOR U9517 ( .A(n6992), .B(n6991), .Z(\w1[7][117] ) );
  XNOR U9518 ( .A(\w3[6][119] ), .B(\w3[6][112] ), .Z(n7028) );
  XNOR U9519 ( .A(n7028), .B(key[1014]), .Z(n6995) );
  XOR U9520 ( .A(\w3[6][110] ), .B(n6993), .Z(n6994) );
  XNOR U9521 ( .A(n6995), .B(n6994), .Z(\w1[7][118] ) );
  XOR U9522 ( .A(n6996), .B(key[1015]), .Z(n6999) );
  XNOR U9523 ( .A(\w3[6][112] ), .B(n6997), .Z(n6998) );
  XNOR U9524 ( .A(n6999), .B(n6998), .Z(\w1[7][119] ) );
  XNOR U9525 ( .A(\w3[6][3] ), .B(\w3[6][27] ), .Z(n7089) );
  XNOR U9526 ( .A(n7052), .B(key[907]), .Z(n7001) );
  XNOR U9527 ( .A(\w3[6][0] ), .B(\w3[6][4] ), .Z(n7118) );
  XOR U9528 ( .A(\w3[6][19] ), .B(n7118), .Z(n7000) );
  XNOR U9529 ( .A(n7001), .B(n7000), .Z(\w1[7][11] ) );
  XNOR U9530 ( .A(n7002), .B(key[1016]), .Z(n7004) );
  XNOR U9531 ( .A(\w3[6][113] ), .B(\w3[6][121] ), .Z(n7003) );
  XNOR U9532 ( .A(n7004), .B(n7003), .Z(n7005) );
  XOR U9533 ( .A(\w3[6][112] ), .B(n7005), .Z(\w1[7][120] ) );
  XNOR U9534 ( .A(n7337), .B(key[1017]), .Z(n7007) );
  XNOR U9535 ( .A(\w3[6][114] ), .B(\w3[6][122] ), .Z(n7006) );
  XNOR U9536 ( .A(n7007), .B(n7006), .Z(n7008) );
  XOR U9537 ( .A(\w3[6][97] ), .B(n7008), .Z(\w1[7][121] ) );
  XOR U9538 ( .A(\w3[6][123] ), .B(key[1018]), .Z(n7010) );
  XNOR U9539 ( .A(\w3[6][114] ), .B(\w3[6][115] ), .Z(n7009) );
  XNOR U9540 ( .A(n7010), .B(n7009), .Z(n7012) );
  XOR U9541 ( .A(n7012), .B(n7011), .Z(\w1[7][122] ) );
  XOR U9542 ( .A(\w3[6][124] ), .B(n7013), .Z(n7014) );
  XOR U9543 ( .A(n7015), .B(n7014), .Z(n7345) );
  XOR U9544 ( .A(n7345), .B(key[1019]), .Z(n7018) );
  XOR U9545 ( .A(\w3[6][99] ), .B(n7016), .Z(n7017) );
  XNOR U9546 ( .A(n7018), .B(n7017), .Z(\w1[7][123] ) );
  XNOR U9547 ( .A(n7019), .B(key[1020]), .Z(n7023) );
  XNOR U9548 ( .A(n7021), .B(n7020), .Z(n7022) );
  XNOR U9549 ( .A(n7023), .B(n7022), .Z(\w1[7][124] ) );
  XOR U9550 ( .A(\w3[6][118] ), .B(key[1021]), .Z(n7026) );
  XOR U9551 ( .A(n7024), .B(\w3[6][126] ), .Z(n7025) );
  XNOR U9552 ( .A(n7026), .B(n7025), .Z(n7027) );
  XOR U9553 ( .A(\w3[6][101] ), .B(n7027), .Z(\w1[7][125] ) );
  XNOR U9554 ( .A(n7028), .B(key[1022]), .Z(n7031) );
  XOR U9555 ( .A(\w3[6][102] ), .B(n7029), .Z(n7030) );
  XNOR U9556 ( .A(n7031), .B(n7030), .Z(\w1[7][126] ) );
  XNOR U9557 ( .A(n7334), .B(key[1023]), .Z(n7034) );
  XOR U9558 ( .A(\w3[6][103] ), .B(n7032), .Z(n7033) );
  XNOR U9559 ( .A(n7034), .B(n7033), .Z(\w1[7][127] ) );
  XOR U9560 ( .A(\w3[6][13] ), .B(\w3[6][28] ), .Z(n7036) );
  XNOR U9561 ( .A(\w3[6][8] ), .B(\w3[6][4] ), .Z(n7035) );
  XOR U9562 ( .A(n7036), .B(n7035), .Z(n7058) );
  XNOR U9563 ( .A(n7058), .B(key[908]), .Z(n7038) );
  XNOR U9564 ( .A(\w3[6][0] ), .B(\w3[6][5] ), .Z(n7153) );
  XOR U9565 ( .A(\w3[6][20] ), .B(n7153), .Z(n7037) );
  XNOR U9566 ( .A(n7038), .B(n7037), .Z(\w1[7][12] ) );
  IV U9567 ( .A(\w3[6][21] ), .Z(n7083) );
  XNOR U9568 ( .A(\w3[6][14] ), .B(n7083), .Z(n7040) );
  XNOR U9569 ( .A(\w3[6][5] ), .B(\w3[6][29] ), .Z(n7061) );
  XOR U9570 ( .A(n7061), .B(key[909]), .Z(n7039) );
  XNOR U9571 ( .A(n7040), .B(n7039), .Z(n7041) );
  XOR U9572 ( .A(\w3[6][6] ), .B(n7041), .Z(\w1[7][13] ) );
  IV U9573 ( .A(\w3[6][30] ), .Z(n7230) );
  XOR U9574 ( .A(\w3[6][6] ), .B(n7230), .Z(n7195) );
  XOR U9575 ( .A(\w3[6][8] ), .B(\w3[6][15] ), .Z(n7064) );
  XNOR U9576 ( .A(n7195), .B(n7064), .Z(n7062) );
  XOR U9577 ( .A(n7062), .B(key[910]), .Z(n7043) );
  XNOR U9578 ( .A(\w3[6][0] ), .B(\w3[6][7] ), .Z(n7231) );
  XOR U9579 ( .A(\w3[6][22] ), .B(n7231), .Z(n7042) );
  XNOR U9580 ( .A(n7043), .B(n7042), .Z(\w1[7][14] ) );
  XNOR U9581 ( .A(\w3[6][7] ), .B(\w3[6][31] ), .Z(n7063) );
  XNOR U9582 ( .A(n7063), .B(key[911]), .Z(n7045) );
  XOR U9583 ( .A(\w3[6][8] ), .B(\w3[6][0] ), .Z(n7067) );
  XNOR U9584 ( .A(\w3[6][23] ), .B(n7067), .Z(n7044) );
  XNOR U9585 ( .A(n7045), .B(n7044), .Z(\w1[7][15] ) );
  XNOR U9586 ( .A(\w3[6][17] ), .B(\w3[6][9] ), .Z(n7069) );
  XNOR U9587 ( .A(n7069), .B(key[912]), .Z(n7047) );
  XNOR U9588 ( .A(\w3[6][24] ), .B(n7067), .Z(n7046) );
  XNOR U9589 ( .A(n7047), .B(n7046), .Z(\w1[7][16] ) );
  XNOR U9590 ( .A(\w3[6][18] ), .B(\w3[6][10] ), .Z(n7088) );
  XNOR U9591 ( .A(n7088), .B(key[913]), .Z(n7049) );
  IV U9592 ( .A(\w3[6][9] ), .Z(n7302) );
  XNOR U9593 ( .A(n7352), .B(n7302), .Z(n7048) );
  XNOR U9594 ( .A(n7049), .B(n7048), .Z(\w1[7][17] ) );
  XNOR U9595 ( .A(\w3[6][11] ), .B(\w3[6][19] ), .Z(n7074) );
  XNOR U9596 ( .A(n7074), .B(key[914]), .Z(n7051) );
  XOR U9597 ( .A(n7055), .B(\w3[6][10] ), .Z(n7050) );
  XNOR U9598 ( .A(n7051), .B(n7050), .Z(\w1[7][18] ) );
  XOR U9599 ( .A(n7068), .B(\w3[6][20] ), .Z(n7075) );
  XNOR U9600 ( .A(n7075), .B(key[915]), .Z(n7054) );
  XOR U9601 ( .A(\w3[6][11] ), .B(n7052), .Z(n7053) );
  XNOR U9602 ( .A(n7054), .B(n7053), .Z(\w1[7][19] ) );
  XNOR U9603 ( .A(n7069), .B(key[897]), .Z(n7057) );
  XOR U9604 ( .A(\w3[6][25] ), .B(n7055), .Z(n7056) );
  XNOR U9605 ( .A(n7057), .B(n7056), .Z(\w1[7][1] ) );
  XOR U9606 ( .A(\w3[6][16] ), .B(n7083), .Z(n7080) );
  XNOR U9607 ( .A(n7080), .B(key[916]), .Z(n7060) );
  XOR U9608 ( .A(\w3[6][12] ), .B(n7058), .Z(n7059) );
  XNOR U9609 ( .A(n7060), .B(n7059), .Z(\w1[7][20] ) );
  IV U9610 ( .A(\w3[6][22] ), .Z(n7084) );
  XOR U9611 ( .A(\w3[6][14] ), .B(n7084), .Z(n7093) );
  XOR U9612 ( .A(n7068), .B(\w3[6][23] ), .Z(n7094) );
  XNOR U9613 ( .A(n7063), .B(key[919]), .Z(n7066) );
  XNOR U9614 ( .A(\w3[6][16] ), .B(n7064), .Z(n7065) );
  XNOR U9615 ( .A(n7066), .B(n7065), .Z(\w1[7][23] ) );
  XNOR U9616 ( .A(n7088), .B(key[922]), .Z(n7071) );
  XNOR U9617 ( .A(\w3[6][2] ), .B(\w3[6][19] ), .Z(n7070) );
  XNOR U9618 ( .A(n7071), .B(n7070), .Z(n7072) );
  XOR U9619 ( .A(\w3[6][27] ), .B(n7072), .Z(\w1[7][26] ) );
  IV U9620 ( .A(\w3[6][24] ), .Z(n7092) );
  XOR U9621 ( .A(n7092), .B(\w3[6][28] ), .Z(n7073) );
  XOR U9622 ( .A(n7074), .B(n7073), .Z(n7117) );
  XOR U9623 ( .A(n7117), .B(key[923]), .Z(n7077) );
  XOR U9624 ( .A(\w3[6][3] ), .B(n7075), .Z(n7076) );
  XNOR U9625 ( .A(n7077), .B(n7076), .Z(\w1[7][27] ) );
  XOR U9626 ( .A(\w3[6][20] ), .B(\w3[6][29] ), .Z(n7079) );
  XOR U9627 ( .A(n7092), .B(\w3[6][12] ), .Z(n7078) );
  XOR U9628 ( .A(n7079), .B(n7078), .Z(n7152) );
  XNOR U9629 ( .A(n7152), .B(key[924]), .Z(n7082) );
  XOR U9630 ( .A(\w3[6][4] ), .B(n7080), .Z(n7081) );
  XNOR U9631 ( .A(n7082), .B(n7081), .Z(\w1[7][28] ) );
  XOR U9632 ( .A(\w3[6][13] ), .B(n7083), .Z(n7194) );
  XNOR U9633 ( .A(n7194), .B(key[925]), .Z(n7086) );
  XNOR U9634 ( .A(n7084), .B(n7230), .Z(n7085) );
  XNOR U9635 ( .A(n7086), .B(n7085), .Z(n7087) );
  XOR U9636 ( .A(\w3[6][5] ), .B(n7087), .Z(\w1[7][29] ) );
  XNOR U9637 ( .A(n7088), .B(key[898]), .Z(n7091) );
  XOR U9638 ( .A(\w3[6][26] ), .B(n7089), .Z(n7090) );
  XNOR U9639 ( .A(n7091), .B(n7090), .Z(\w1[7][2] ) );
  XOR U9640 ( .A(n7092), .B(\w3[6][31] ), .Z(n7266) );
  XNOR U9641 ( .A(n7093), .B(n7266), .Z(n7229) );
  XNOR U9642 ( .A(\w3[6][15] ), .B(\w3[6][23] ), .Z(n7265) );
  XNOR U9643 ( .A(n7265), .B(key[927]), .Z(n7096) );
  XOR U9644 ( .A(n7305), .B(\w3[6][7] ), .Z(n7095) );
  XNOR U9645 ( .A(n7096), .B(n7095), .Z(\w1[7][31] ) );
  XOR U9646 ( .A(\w3[6][33] ), .B(\w3[6][57] ), .Z(n7149) );
  XOR U9647 ( .A(n7149), .B(key[928]), .Z(n7098) );
  XNOR U9648 ( .A(\w3[6][48] ), .B(\w3[6][56] ), .Z(n7211) );
  XOR U9649 ( .A(n7211), .B(\w3[6][40] ), .Z(n7097) );
  XNOR U9650 ( .A(n7098), .B(n7097), .Z(\w1[7][32] ) );
  XNOR U9651 ( .A(\w3[6][34] ), .B(\w3[6][58] ), .Z(n7157) );
  XOR U9652 ( .A(\w3[6][57] ), .B(\w3[6][49] ), .Z(n7175) );
  XNOR U9653 ( .A(n7175), .B(key[929]), .Z(n7099) );
  XNOR U9654 ( .A(n7157), .B(n7099), .Z(n7100) );
  XNOR U9655 ( .A(\w3[6][41] ), .B(n7100), .Z(\w1[7][33] ) );
  XNOR U9656 ( .A(n7127), .B(key[930]), .Z(n7102) );
  XNOR U9657 ( .A(\w3[6][50] ), .B(\w3[6][42] ), .Z(n7185) );
  XOR U9658 ( .A(\w3[6][58] ), .B(n7185), .Z(n7101) );
  XNOR U9659 ( .A(n7102), .B(n7101), .Z(\w1[7][34] ) );
  XOR U9660 ( .A(\w3[6][36] ), .B(\w3[6][32] ), .Z(n7129) );
  XOR U9661 ( .A(n7129), .B(key[931]), .Z(n7105) );
  IV U9662 ( .A(\w3[6][51] ), .Z(n7184) );
  XOR U9663 ( .A(\w3[6][43] ), .B(n7184), .Z(n7156) );
  XOR U9664 ( .A(\w3[6][56] ), .B(n7156), .Z(n7103) );
  XNOR U9665 ( .A(\w3[6][60] ), .B(n7103), .Z(n7190) );
  XNOR U9666 ( .A(\w3[6][59] ), .B(n7190), .Z(n7104) );
  XNOR U9667 ( .A(n7105), .B(n7104), .Z(\w1[7][35] ) );
  XOR U9668 ( .A(\w3[6][32] ), .B(\w3[6][37] ), .Z(n7135) );
  XOR U9669 ( .A(\w3[6][52] ), .B(\w3[6][61] ), .Z(n7107) );
  XNOR U9670 ( .A(\w3[6][56] ), .B(\w3[6][44] ), .Z(n7106) );
  XOR U9671 ( .A(n7107), .B(n7106), .Z(n7199) );
  XOR U9672 ( .A(n7199), .B(key[932]), .Z(n7108) );
  XOR U9673 ( .A(n7135), .B(n7108), .Z(n7109) );
  XNOR U9674 ( .A(\w3[6][60] ), .B(n7109), .Z(\w1[7][36] ) );
  XNOR U9675 ( .A(\w3[6][38] ), .B(\w3[6][62] ), .Z(n7141) );
  XNOR U9676 ( .A(n7141), .B(key[933]), .Z(n7111) );
  IV U9677 ( .A(\w3[6][45] ), .Z(n7164) );
  XOR U9678 ( .A(\w3[6][53] ), .B(n7164), .Z(n7202) );
  XOR U9679 ( .A(\w3[6][61] ), .B(n7202), .Z(n7110) );
  XNOR U9680 ( .A(n7111), .B(n7110), .Z(\w1[7][37] ) );
  XOR U9681 ( .A(\w3[6][32] ), .B(\w3[6][39] ), .Z(n7142) );
  XOR U9682 ( .A(n7142), .B(key[934]), .Z(n7113) );
  XNOR U9683 ( .A(\w3[6][56] ), .B(\w3[6][63] ), .Z(n7114) );
  XOR U9684 ( .A(\w3[6][46] ), .B(\w3[6][54] ), .Z(n7163) );
  XOR U9685 ( .A(n7114), .B(n7163), .Z(n7207) );
  XOR U9686 ( .A(\w3[6][62] ), .B(n7207), .Z(n7112) );
  XNOR U9687 ( .A(n7113), .B(n7112), .Z(\w1[7][38] ) );
  XNOR U9688 ( .A(\w3[6][55] ), .B(\w3[6][47] ), .Z(n7210) );
  XNOR U9689 ( .A(n7210), .B(key[935]), .Z(n7116) );
  XOR U9690 ( .A(\w3[6][32] ), .B(n7114), .Z(n7115) );
  XNOR U9691 ( .A(n7116), .B(n7115), .Z(\w1[7][39] ) );
  XOR U9692 ( .A(n7117), .B(key[899]), .Z(n7120) );
  XOR U9693 ( .A(n7118), .B(\w3[6][27] ), .Z(n7119) );
  XNOR U9694 ( .A(n7120), .B(n7119), .Z(\w1[7][3] ) );
  IV U9695 ( .A(\w3[6][33] ), .Z(n7180) );
  XOR U9696 ( .A(\w3[6][42] ), .B(key[937]), .Z(n7122) );
  XNOR U9697 ( .A(n7175), .B(\w3[6][34] ), .Z(n7121) );
  XNOR U9698 ( .A(n7122), .B(n7121), .Z(n7123) );
  XNOR U9699 ( .A(n7180), .B(n7123), .Z(\w1[7][41] ) );
  XOR U9700 ( .A(\w3[6][43] ), .B(key[938]), .Z(n7125) );
  IV U9701 ( .A(\w3[6][35] ), .Z(n7191) );
  XOR U9702 ( .A(\w3[6][50] ), .B(n7191), .Z(n7124) );
  XNOR U9703 ( .A(n7125), .B(n7124), .Z(n7126) );
  XNOR U9704 ( .A(n7126), .B(n7157), .Z(\w1[7][42] ) );
  IV U9705 ( .A(\w3[6][40] ), .Z(n7132) );
  XNOR U9706 ( .A(n7132), .B(n7127), .Z(n7128) );
  XOR U9707 ( .A(\w3[6][44] ), .B(n7128), .Z(n7158) );
  XNOR U9708 ( .A(n7158), .B(key[939]), .Z(n7131) );
  XNOR U9709 ( .A(\w3[6][51] ), .B(n7129), .Z(n7130) );
  XNOR U9710 ( .A(n7131), .B(n7130), .Z(\w1[7][43] ) );
  XOR U9711 ( .A(\w3[6][36] ), .B(\w3[6][45] ), .Z(n7134) );
  XOR U9712 ( .A(n7132), .B(\w3[6][60] ), .Z(n7133) );
  XOR U9713 ( .A(n7134), .B(n7133), .Z(n7159) );
  XNOR U9714 ( .A(n7159), .B(key[940]), .Z(n7137) );
  XNOR U9715 ( .A(\w3[6][52] ), .B(n7135), .Z(n7136) );
  XNOR U9716 ( .A(n7137), .B(n7136), .Z(\w1[7][44] ) );
  XNOR U9717 ( .A(\w3[6][61] ), .B(\w3[6][37] ), .Z(n7162) );
  XNOR U9718 ( .A(n7162), .B(key[941]), .Z(n7139) );
  XNOR U9719 ( .A(\w3[6][38] ), .B(\w3[6][46] ), .Z(n7138) );
  XNOR U9720 ( .A(n7139), .B(n7138), .Z(n7140) );
  XOR U9721 ( .A(\w3[6][53] ), .B(n7140), .Z(\w1[7][45] ) );
  XOR U9722 ( .A(\w3[6][40] ), .B(\w3[6][47] ), .Z(n7171) );
  XOR U9723 ( .A(n7141), .B(n7171), .Z(n7167) );
  XNOR U9724 ( .A(n7167), .B(key[942]), .Z(n7144) );
  XNOR U9725 ( .A(\w3[6][54] ), .B(n7142), .Z(n7143) );
  XNOR U9726 ( .A(n7144), .B(n7143), .Z(\w1[7][46] ) );
  XOR U9727 ( .A(\w3[6][63] ), .B(\w3[6][39] ), .Z(n7170) );
  XOR U9728 ( .A(n7170), .B(key[943]), .Z(n7146) );
  XNOR U9729 ( .A(\w3[6][40] ), .B(\w3[6][32] ), .Z(n7174) );
  XOR U9730 ( .A(\w3[6][55] ), .B(n7174), .Z(n7145) );
  XNOR U9731 ( .A(n7146), .B(n7145), .Z(\w1[7][47] ) );
  XNOR U9732 ( .A(\w3[6][41] ), .B(\w3[6][49] ), .Z(n7179) );
  XNOR U9733 ( .A(n7179), .B(key[944]), .Z(n7148) );
  XOR U9734 ( .A(\w3[6][56] ), .B(n7174), .Z(n7147) );
  XNOR U9735 ( .A(n7148), .B(n7147), .Z(\w1[7][48] ) );
  XNOR U9736 ( .A(n7185), .B(key[945]), .Z(n7151) );
  XNOR U9737 ( .A(n7149), .B(\w3[6][41] ), .Z(n7150) );
  XNOR U9738 ( .A(n7151), .B(n7150), .Z(\w1[7][49] ) );
  XNOR U9739 ( .A(n7152), .B(key[900]), .Z(n7155) );
  XOR U9740 ( .A(n7153), .B(\w3[6][28] ), .Z(n7154) );
  XNOR U9741 ( .A(n7155), .B(n7154), .Z(\w1[7][4] ) );
  IV U9742 ( .A(\w3[6][48] ), .Z(n7176) );
  XOR U9743 ( .A(n7176), .B(\w3[6][52] ), .Z(n7189) );
  XNOR U9744 ( .A(n7198), .B(key[948]), .Z(n7161) );
  XOR U9745 ( .A(\w3[6][44] ), .B(n7159), .Z(n7160) );
  XNOR U9746 ( .A(n7161), .B(n7160), .Z(\w1[7][52] ) );
  XNOR U9747 ( .A(n7162), .B(key[949]), .Z(n7166) );
  XOR U9748 ( .A(n7164), .B(n7163), .Z(n7165) );
  XNOR U9749 ( .A(n7166), .B(n7165), .Z(\w1[7][53] ) );
  XOR U9750 ( .A(n7176), .B(\w3[6][55] ), .Z(n7206) );
  XNOR U9751 ( .A(n7206), .B(key[950]), .Z(n7169) );
  XOR U9752 ( .A(\w3[6][46] ), .B(n7167), .Z(n7168) );
  XNOR U9753 ( .A(n7169), .B(n7168), .Z(\w1[7][54] ) );
  XOR U9754 ( .A(n7170), .B(key[951]), .Z(n7173) );
  XNOR U9755 ( .A(\w3[6][48] ), .B(n7171), .Z(n7172) );
  XNOR U9756 ( .A(n7173), .B(n7172), .Z(\w1[7][55] ) );
  XNOR U9757 ( .A(n7174), .B(key[952]), .Z(n7178) );
  XOR U9758 ( .A(n7176), .B(n7175), .Z(n7177) );
  XNOR U9759 ( .A(n7178), .B(n7177), .Z(\w1[7][56] ) );
  XNOR U9760 ( .A(n7179), .B(key[953]), .Z(n7182) );
  XOR U9761 ( .A(n7180), .B(\w3[6][50] ), .Z(n7181) );
  XNOR U9762 ( .A(n7182), .B(n7181), .Z(n7183) );
  XOR U9763 ( .A(\w3[6][58] ), .B(n7183), .Z(\w1[7][57] ) );
  XNOR U9764 ( .A(n7184), .B(key[954]), .Z(n7187) );
  XOR U9765 ( .A(n7185), .B(\w3[6][59] ), .Z(n7186) );
  XNOR U9766 ( .A(n7187), .B(n7186), .Z(n7188) );
  XOR U9767 ( .A(\w3[6][34] ), .B(n7188), .Z(\w1[7][58] ) );
  XNOR U9768 ( .A(n7189), .B(key[955]), .Z(n7193) );
  XOR U9769 ( .A(n7191), .B(n7190), .Z(n7192) );
  XNOR U9770 ( .A(n7193), .B(n7192), .Z(\w1[7][59] ) );
  XNOR U9771 ( .A(n7194), .B(key[901]), .Z(n7197) );
  XOR U9772 ( .A(\w3[6][29] ), .B(n7195), .Z(n7196) );
  XNOR U9773 ( .A(n7197), .B(n7196), .Z(\w1[7][5] ) );
  XNOR U9774 ( .A(n7198), .B(key[956]), .Z(n7201) );
  XOR U9775 ( .A(\w3[6][36] ), .B(n7199), .Z(n7200) );
  XNOR U9776 ( .A(n7201), .B(n7200), .Z(\w1[7][60] ) );
  XOR U9777 ( .A(\w3[6][54] ), .B(key[957]), .Z(n7204) );
  XOR U9778 ( .A(n7202), .B(\w3[6][62] ), .Z(n7203) );
  XNOR U9779 ( .A(n7204), .B(n7203), .Z(n7205) );
  XOR U9780 ( .A(\w3[6][37] ), .B(n7205), .Z(\w1[7][61] ) );
  XNOR U9781 ( .A(n7206), .B(key[958]), .Z(n7209) );
  XOR U9782 ( .A(\w3[6][38] ), .B(n7207), .Z(n7208) );
  XNOR U9783 ( .A(n7209), .B(n7208), .Z(\w1[7][62] ) );
  XNOR U9784 ( .A(n7210), .B(key[959]), .Z(n7213) );
  XOR U9785 ( .A(n7211), .B(\w3[6][39] ), .Z(n7212) );
  XNOR U9786 ( .A(n7213), .B(n7212), .Z(\w1[7][63] ) );
  XOR U9787 ( .A(\w3[6][65] ), .B(\w3[6][89] ), .Z(n7271) );
  XOR U9788 ( .A(n7271), .B(key[960]), .Z(n7215) );
  XNOR U9789 ( .A(\w3[6][80] ), .B(\w3[6][88] ), .Z(n7330) );
  XOR U9790 ( .A(n7330), .B(\w3[6][72] ), .Z(n7214) );
  XNOR U9791 ( .A(n7215), .B(n7214), .Z(\w1[7][64] ) );
  XNOR U9792 ( .A(\w3[6][66] ), .B(\w3[6][90] ), .Z(n7275) );
  XOR U9793 ( .A(\w3[6][89] ), .B(\w3[6][81] ), .Z(n7293) );
  XNOR U9794 ( .A(n7293), .B(key[961]), .Z(n7216) );
  XNOR U9795 ( .A(n7275), .B(n7216), .Z(n7217) );
  XNOR U9796 ( .A(\w3[6][73] ), .B(n7217), .Z(\w1[7][65] ) );
  XNOR U9797 ( .A(n7245), .B(key[962]), .Z(n7219) );
  XNOR U9798 ( .A(\w3[6][82] ), .B(\w3[6][74] ), .Z(n7308) );
  XOR U9799 ( .A(\w3[6][90] ), .B(n7308), .Z(n7218) );
  XNOR U9800 ( .A(n7219), .B(n7218), .Z(\w1[7][66] ) );
  XOR U9801 ( .A(\w3[6][68] ), .B(\w3[6][64] ), .Z(n7247) );
  XOR U9802 ( .A(n7247), .B(key[963]), .Z(n7222) );
  IV U9803 ( .A(\w3[6][83] ), .Z(n7307) );
  XOR U9804 ( .A(\w3[6][75] ), .B(n7307), .Z(n7274) );
  XOR U9805 ( .A(\w3[6][88] ), .B(n7274), .Z(n7220) );
  XNOR U9806 ( .A(\w3[6][92] ), .B(n7220), .Z(n7313) );
  XNOR U9807 ( .A(\w3[6][91] ), .B(n7313), .Z(n7221) );
  XNOR U9808 ( .A(n7222), .B(n7221), .Z(\w1[7][67] ) );
  XOR U9809 ( .A(\w3[6][64] ), .B(\w3[6][69] ), .Z(n7253) );
  XOR U9810 ( .A(\w3[6][84] ), .B(\w3[6][93] ), .Z(n7224) );
  XNOR U9811 ( .A(\w3[6][88] ), .B(\w3[6][76] ), .Z(n7223) );
  XOR U9812 ( .A(n7224), .B(n7223), .Z(n7318) );
  XOR U9813 ( .A(n7318), .B(key[964]), .Z(n7225) );
  XOR U9814 ( .A(n7253), .B(n7225), .Z(n7226) );
  XNOR U9815 ( .A(\w3[6][92] ), .B(n7226), .Z(\w1[7][68] ) );
  XNOR U9816 ( .A(\w3[6][70] ), .B(\w3[6][94] ), .Z(n7259) );
  XNOR U9817 ( .A(n7259), .B(key[965]), .Z(n7228) );
  IV U9818 ( .A(\w3[6][77] ), .Z(n7282) );
  XOR U9819 ( .A(\w3[6][85] ), .B(n7282), .Z(n7321) );
  XOR U9820 ( .A(\w3[6][93] ), .B(n7321), .Z(n7227) );
  XNOR U9821 ( .A(n7228), .B(n7227), .Z(\w1[7][69] ) );
  XNOR U9822 ( .A(n7229), .B(key[902]), .Z(n7233) );
  XNOR U9823 ( .A(n7231), .B(n7230), .Z(n7232) );
  XNOR U9824 ( .A(n7233), .B(n7232), .Z(\w1[7][6] ) );
  XOR U9825 ( .A(\w3[6][64] ), .B(\w3[6][71] ), .Z(n7260) );
  XOR U9826 ( .A(n7260), .B(key[966]), .Z(n7235) );
  XNOR U9827 ( .A(\w3[6][88] ), .B(\w3[6][95] ), .Z(n7236) );
  XOR U9828 ( .A(\w3[6][78] ), .B(\w3[6][86] ), .Z(n7281) );
  XOR U9829 ( .A(n7236), .B(n7281), .Z(n7326) );
  XOR U9830 ( .A(\w3[6][94] ), .B(n7326), .Z(n7234) );
  XNOR U9831 ( .A(n7235), .B(n7234), .Z(\w1[7][70] ) );
  XNOR U9832 ( .A(\w3[6][79] ), .B(\w3[6][87] ), .Z(n7329) );
  XNOR U9833 ( .A(n7329), .B(key[967]), .Z(n7238) );
  XOR U9834 ( .A(\w3[6][64] ), .B(n7236), .Z(n7237) );
  XNOR U9835 ( .A(n7238), .B(n7237), .Z(\w1[7][71] ) );
  IV U9836 ( .A(\w3[6][65] ), .Z(n7298) );
  XOR U9837 ( .A(\w3[6][74] ), .B(key[969]), .Z(n7240) );
  XNOR U9838 ( .A(n7293), .B(\w3[6][66] ), .Z(n7239) );
  XNOR U9839 ( .A(n7240), .B(n7239), .Z(n7241) );
  XNOR U9840 ( .A(n7298), .B(n7241), .Z(\w1[7][73] ) );
  XOR U9841 ( .A(\w3[6][75] ), .B(key[970]), .Z(n7243) );
  IV U9842 ( .A(\w3[6][67] ), .Z(n7314) );
  XOR U9843 ( .A(\w3[6][82] ), .B(n7314), .Z(n7242) );
  XNOR U9844 ( .A(n7243), .B(n7242), .Z(n7244) );
  XNOR U9845 ( .A(n7244), .B(n7275), .Z(\w1[7][74] ) );
  IV U9846 ( .A(\w3[6][72] ), .Z(n7250) );
  XNOR U9847 ( .A(n7250), .B(n7245), .Z(n7246) );
  XOR U9848 ( .A(\w3[6][76] ), .B(n7246), .Z(n7276) );
  XNOR U9849 ( .A(n7276), .B(key[971]), .Z(n7249) );
  XNOR U9850 ( .A(\w3[6][83] ), .B(n7247), .Z(n7248) );
  XNOR U9851 ( .A(n7249), .B(n7248), .Z(\w1[7][75] ) );
  XOR U9852 ( .A(\w3[6][68] ), .B(\w3[6][77] ), .Z(n7252) );
  XOR U9853 ( .A(n7250), .B(\w3[6][92] ), .Z(n7251) );
  XOR U9854 ( .A(n7252), .B(n7251), .Z(n7277) );
  XNOR U9855 ( .A(n7277), .B(key[972]), .Z(n7255) );
  XNOR U9856 ( .A(\w3[6][84] ), .B(n7253), .Z(n7254) );
  XNOR U9857 ( .A(n7255), .B(n7254), .Z(\w1[7][76] ) );
  XNOR U9858 ( .A(\w3[6][93] ), .B(\w3[6][69] ), .Z(n7280) );
  XNOR U9859 ( .A(n7280), .B(key[973]), .Z(n7257) );
  XNOR U9860 ( .A(\w3[6][70] ), .B(\w3[6][78] ), .Z(n7256) );
  XNOR U9861 ( .A(n7257), .B(n7256), .Z(n7258) );
  XOR U9862 ( .A(\w3[6][85] ), .B(n7258), .Z(\w1[7][77] ) );
  XOR U9863 ( .A(\w3[6][72] ), .B(\w3[6][79] ), .Z(n7289) );
  XOR U9864 ( .A(n7259), .B(n7289), .Z(n7285) );
  XNOR U9865 ( .A(n7285), .B(key[974]), .Z(n7262) );
  XNOR U9866 ( .A(\w3[6][86] ), .B(n7260), .Z(n7261) );
  XNOR U9867 ( .A(n7262), .B(n7261), .Z(\w1[7][78] ) );
  XOR U9868 ( .A(\w3[6][95] ), .B(\w3[6][71] ), .Z(n7288) );
  XOR U9869 ( .A(n7288), .B(key[975]), .Z(n7264) );
  XNOR U9870 ( .A(\w3[6][72] ), .B(\w3[6][64] ), .Z(n7292) );
  XOR U9871 ( .A(\w3[6][87] ), .B(n7292), .Z(n7263) );
  XNOR U9872 ( .A(n7264), .B(n7263), .Z(\w1[7][79] ) );
  XNOR U9873 ( .A(n7265), .B(key[903]), .Z(n7268) );
  XOR U9874 ( .A(\w3[6][0] ), .B(n7266), .Z(n7267) );
  XNOR U9875 ( .A(n7268), .B(n7267), .Z(\w1[7][7] ) );
  XNOR U9876 ( .A(\w3[6][73] ), .B(\w3[6][81] ), .Z(n7297) );
  XNOR U9877 ( .A(n7297), .B(key[976]), .Z(n7270) );
  XOR U9878 ( .A(\w3[6][88] ), .B(n7292), .Z(n7269) );
  XNOR U9879 ( .A(n7270), .B(n7269), .Z(\w1[7][80] ) );
  XNOR U9880 ( .A(n7308), .B(key[977]), .Z(n7273) );
  XNOR U9881 ( .A(n7271), .B(\w3[6][73] ), .Z(n7272) );
  XNOR U9882 ( .A(n7273), .B(n7272), .Z(\w1[7][81] ) );
  IV U9883 ( .A(\w3[6][80] ), .Z(n7294) );
  XOR U9884 ( .A(n7294), .B(\w3[6][84] ), .Z(n7312) );
  XNOR U9885 ( .A(n7317), .B(key[980]), .Z(n7279) );
  XOR U9886 ( .A(\w3[6][76] ), .B(n7277), .Z(n7278) );
  XNOR U9887 ( .A(n7279), .B(n7278), .Z(\w1[7][84] ) );
  XNOR U9888 ( .A(n7280), .B(key[981]), .Z(n7284) );
  XOR U9889 ( .A(n7282), .B(n7281), .Z(n7283) );
  XNOR U9890 ( .A(n7284), .B(n7283), .Z(\w1[7][85] ) );
  XOR U9891 ( .A(n7294), .B(\w3[6][87] ), .Z(n7325) );
  XNOR U9892 ( .A(n7325), .B(key[982]), .Z(n7287) );
  XOR U9893 ( .A(\w3[6][78] ), .B(n7285), .Z(n7286) );
  XNOR U9894 ( .A(n7287), .B(n7286), .Z(\w1[7][86] ) );
  XOR U9895 ( .A(n7288), .B(key[983]), .Z(n7291) );
  XNOR U9896 ( .A(\w3[6][80] ), .B(n7289), .Z(n7290) );
  XNOR U9897 ( .A(n7291), .B(n7290), .Z(\w1[7][87] ) );
  XNOR U9898 ( .A(n7292), .B(key[984]), .Z(n7296) );
  XOR U9899 ( .A(n7294), .B(n7293), .Z(n7295) );
  XNOR U9900 ( .A(n7296), .B(n7295), .Z(\w1[7][88] ) );
  XNOR U9901 ( .A(n7297), .B(key[985]), .Z(n7300) );
  XOR U9902 ( .A(n7298), .B(\w3[6][82] ), .Z(n7299) );
  XNOR U9903 ( .A(n7300), .B(n7299), .Z(n7301) );
  XOR U9904 ( .A(\w3[6][90] ), .B(n7301), .Z(\w1[7][89] ) );
  XNOR U9905 ( .A(n7302), .B(key[904]), .Z(n7304) );
  XNOR U9906 ( .A(\w3[6][1] ), .B(\w3[6][0] ), .Z(n7303) );
  XNOR U9907 ( .A(n7304), .B(n7303), .Z(n7306) );
  XNOR U9908 ( .A(n7306), .B(n7305), .Z(\w1[7][8] ) );
  XNOR U9909 ( .A(n7307), .B(key[986]), .Z(n7310) );
  XOR U9910 ( .A(n7308), .B(\w3[6][91] ), .Z(n7309) );
  XNOR U9911 ( .A(n7310), .B(n7309), .Z(n7311) );
  XOR U9912 ( .A(\w3[6][66] ), .B(n7311), .Z(\w1[7][90] ) );
  XNOR U9913 ( .A(n7312), .B(key[987]), .Z(n7316) );
  XOR U9914 ( .A(n7314), .B(n7313), .Z(n7315) );
  XNOR U9915 ( .A(n7316), .B(n7315), .Z(\w1[7][91] ) );
  XNOR U9916 ( .A(n7317), .B(key[988]), .Z(n7320) );
  XOR U9917 ( .A(\w3[6][68] ), .B(n7318), .Z(n7319) );
  XNOR U9918 ( .A(n7320), .B(n7319), .Z(\w1[7][92] ) );
  XOR U9919 ( .A(\w3[6][86] ), .B(key[989]), .Z(n7323) );
  XOR U9920 ( .A(n7321), .B(\w3[6][94] ), .Z(n7322) );
  XNOR U9921 ( .A(n7323), .B(n7322), .Z(n7324) );
  XOR U9922 ( .A(\w3[6][69] ), .B(n7324), .Z(\w1[7][93] ) );
  XNOR U9923 ( .A(n7325), .B(key[990]), .Z(n7328) );
  XOR U9924 ( .A(\w3[6][70] ), .B(n7326), .Z(n7327) );
  XNOR U9925 ( .A(n7328), .B(n7327), .Z(\w1[7][94] ) );
  XNOR U9926 ( .A(n7329), .B(key[991]), .Z(n7332) );
  XOR U9927 ( .A(n7330), .B(\w3[6][71] ), .Z(n7331) );
  XNOR U9928 ( .A(n7332), .B(n7331), .Z(\w1[7][95] ) );
  XOR U9929 ( .A(\w3[6][104] ), .B(key[992]), .Z(n7336) );
  XOR U9930 ( .A(n7334), .B(n7333), .Z(n7335) );
  XNOR U9931 ( .A(n7336), .B(n7335), .Z(\w1[7][96] ) );
  XNOR U9932 ( .A(n7337), .B(key[993]), .Z(n7340) );
  XOR U9933 ( .A(\w3[6][121] ), .B(n7338), .Z(n7339) );
  XNOR U9934 ( .A(n7340), .B(n7339), .Z(\w1[7][97] ) );
  XNOR U9935 ( .A(n7341), .B(key[994]), .Z(n7344) );
  XOR U9936 ( .A(\w3[6][122] ), .B(n7342), .Z(n7343) );
  XNOR U9937 ( .A(n7344), .B(n7343), .Z(\w1[7][98] ) );
  XOR U9938 ( .A(n7345), .B(key[995]), .Z(n7348) );
  XOR U9939 ( .A(n7346), .B(\w3[6][123] ), .Z(n7347) );
  XNOR U9940 ( .A(n7348), .B(n7347), .Z(\w1[7][99] ) );
  XOR U9941 ( .A(\w3[6][10] ), .B(key[905]), .Z(n7350) );
  XNOR U9942 ( .A(\w3[6][2] ), .B(\w3[6][17] ), .Z(n7349) );
  XNOR U9943 ( .A(n7350), .B(n7349), .Z(n7351) );
  XNOR U9944 ( .A(n7352), .B(n7351), .Z(\w1[7][9] ) );
  XNOR U9945 ( .A(\w3[7][25] ), .B(\w3[7][1] ), .Z(n7778) );
  IV U9946 ( .A(\w3[7][16] ), .Z(n7480) );
  XOR U9947 ( .A(\w3[7][24] ), .B(n7480), .Z(n7730) );
  XNOR U9948 ( .A(\w3[7][8] ), .B(key[1024]), .Z(n7353) );
  XNOR U9949 ( .A(n7730), .B(n7353), .Z(n7354) );
  XOR U9950 ( .A(n7778), .B(n7354), .Z(\w1[8][0] ) );
  XOR U9951 ( .A(\w3[7][96] ), .B(\w3[7][101] ), .Z(n7377) );
  XOR U9952 ( .A(\w3[7][116] ), .B(\w3[7][125] ), .Z(n7356) );
  IV U9953 ( .A(\w3[7][120] ), .Z(n7429) );
  XOR U9954 ( .A(n7429), .B(\w3[7][108] ), .Z(n7355) );
  XOR U9955 ( .A(n7356), .B(n7355), .Z(n7435) );
  XOR U9956 ( .A(n7435), .B(key[1124]), .Z(n7357) );
  XOR U9957 ( .A(n7377), .B(n7357), .Z(n7358) );
  XNOR U9958 ( .A(\w3[7][124] ), .B(n7358), .Z(\w1[8][100] ) );
  XNOR U9959 ( .A(\w3[7][102] ), .B(\w3[7][126] ), .Z(n7386) );
  XNOR U9960 ( .A(n7386), .B(key[1125]), .Z(n7360) );
  XNOR U9961 ( .A(\w3[7][109] ), .B(\w3[7][117] ), .Z(n7438) );
  XOR U9962 ( .A(\w3[7][125] ), .B(n7438), .Z(n7359) );
  XNOR U9963 ( .A(n7360), .B(n7359), .Z(\w1[8][101] ) );
  XOR U9964 ( .A(\w3[7][96] ), .B(\w3[7][103] ), .Z(n7387) );
  XOR U9965 ( .A(n7387), .B(key[1126]), .Z(n7362) );
  XOR U9966 ( .A(n7429), .B(\w3[7][127] ), .Z(n7363) );
  XOR U9967 ( .A(\w3[7][110] ), .B(\w3[7][118] ), .Z(n7405) );
  XOR U9968 ( .A(n7363), .B(n7405), .Z(n7443) );
  XOR U9969 ( .A(\w3[7][126] ), .B(n7443), .Z(n7361) );
  XNOR U9970 ( .A(n7362), .B(n7361), .Z(\w1[8][102] ) );
  XNOR U9971 ( .A(\w3[7][111] ), .B(\w3[7][119] ), .Z(n7446) );
  XNOR U9972 ( .A(n7446), .B(key[1127]), .Z(n7365) );
  XOR U9973 ( .A(\w3[7][96] ), .B(n7363), .Z(n7364) );
  XNOR U9974 ( .A(n7365), .B(n7364), .Z(\w1[8][103] ) );
  IV U9975 ( .A(\w3[7][97] ), .Z(n7425) );
  IV U9976 ( .A(\w3[7][112] ), .Z(n7421) );
  XOR U9977 ( .A(\w3[7][120] ), .B(n7421), .Z(n7759) );
  XOR U9978 ( .A(\w3[7][106] ), .B(\w3[7][98] ), .Z(n7367) );
  XNOR U9979 ( .A(\w3[7][97] ), .B(\w3[7][121] ), .Z(n7758) );
  XOR U9980 ( .A(n7758), .B(key[1129]), .Z(n7366) );
  XNOR U9981 ( .A(n7367), .B(n7366), .Z(n7368) );
  XOR U9982 ( .A(\w3[7][113] ), .B(n7368), .Z(\w1[8][105] ) );
  XOR U9983 ( .A(\w3[7][107] ), .B(\w3[7][114] ), .Z(n7370) );
  XOR U9984 ( .A(\w3[7][98] ), .B(\w3[7][122] ), .Z(n7763) );
  XNOR U9985 ( .A(n7763), .B(key[1130]), .Z(n7369) );
  XNOR U9986 ( .A(n7370), .B(n7369), .Z(n7371) );
  XOR U9987 ( .A(\w3[7][99] ), .B(n7371), .Z(\w1[8][106] ) );
  IV U9988 ( .A(\w3[7][123] ), .Z(n7771) );
  XOR U9989 ( .A(\w3[7][99] ), .B(n7771), .Z(n7767) );
  XOR U9990 ( .A(\w3[7][108] ), .B(n7767), .Z(n7372) );
  XOR U9991 ( .A(\w3[7][104] ), .B(n7372), .Z(n7398) );
  XNOR U9992 ( .A(n7398), .B(key[1131]), .Z(n7374) );
  IV U9993 ( .A(\w3[7][100] ), .Z(n7434) );
  XOR U9994 ( .A(\w3[7][96] ), .B(n7434), .Z(n7772) );
  XOR U9995 ( .A(\w3[7][115] ), .B(n7772), .Z(n7373) );
  XNOR U9996 ( .A(n7374), .B(n7373), .Z(\w1[8][107] ) );
  XOR U9997 ( .A(\w3[7][100] ), .B(\w3[7][104] ), .Z(n7376) );
  XNOR U9998 ( .A(\w3[7][124] ), .B(\w3[7][109] ), .Z(n7375) );
  XOR U9999 ( .A(n7376), .B(n7375), .Z(n7401) );
  XNOR U10000 ( .A(n7401), .B(key[1132]), .Z(n7379) );
  XNOR U10001 ( .A(\w3[7][116] ), .B(n7377), .Z(n7378) );
  XNOR U10002 ( .A(n7379), .B(n7378), .Z(\w1[8][108] ) );
  XNOR U10003 ( .A(\w3[7][125] ), .B(\w3[7][101] ), .Z(n7404) );
  XNOR U10004 ( .A(n7404), .B(key[1133]), .Z(n7381) );
  XNOR U10005 ( .A(\w3[7][102] ), .B(\w3[7][110] ), .Z(n7380) );
  XNOR U10006 ( .A(n7381), .B(n7380), .Z(n7382) );
  XOR U10007 ( .A(\w3[7][117] ), .B(n7382), .Z(\w1[8][109] ) );
  IV U10008 ( .A(\w3[7][18] ), .Z(n7485) );
  XNOR U10009 ( .A(\w3[7][11] ), .B(n7485), .Z(n7384) );
  XNOR U10010 ( .A(\w3[7][2] ), .B(\w3[7][26] ), .Z(n7467) );
  XOR U10011 ( .A(n7467), .B(key[1034]), .Z(n7383) );
  XNOR U10012 ( .A(n7384), .B(n7383), .Z(n7385) );
  XOR U10013 ( .A(\w3[7][3] ), .B(n7385), .Z(\w1[8][10] ) );
  XOR U10014 ( .A(\w3[7][111] ), .B(\w3[7][104] ), .Z(n7412) );
  XOR U10015 ( .A(n7386), .B(n7412), .Z(n7408) );
  XNOR U10016 ( .A(n7408), .B(key[1134]), .Z(n7389) );
  XNOR U10017 ( .A(\w3[7][118] ), .B(n7387), .Z(n7388) );
  XNOR U10018 ( .A(n7389), .B(n7388), .Z(\w1[8][110] ) );
  XOR U10019 ( .A(\w3[7][127] ), .B(\w3[7][103] ), .Z(n7411) );
  XOR U10020 ( .A(n7411), .B(key[1135]), .Z(n7391) );
  XNOR U10021 ( .A(\w3[7][96] ), .B(\w3[7][104] ), .Z(n7417) );
  XOR U10022 ( .A(\w3[7][119] ), .B(n7417), .Z(n7390) );
  XNOR U10023 ( .A(n7391), .B(n7390), .Z(\w1[8][111] ) );
  XNOR U10024 ( .A(\w3[7][105] ), .B(\w3[7][113] ), .Z(n7762) );
  XNOR U10025 ( .A(n7762), .B(key[1136]), .Z(n7393) );
  XNOR U10026 ( .A(n7429), .B(n7417), .Z(n7392) );
  XNOR U10027 ( .A(n7393), .B(n7392), .Z(\w1[8][112] ) );
  XNOR U10028 ( .A(\w3[7][106] ), .B(\w3[7][114] ), .Z(n7766) );
  XNOR U10029 ( .A(n7766), .B(key[1137]), .Z(n7395) );
  XOR U10030 ( .A(\w3[7][105] ), .B(n7758), .Z(n7394) );
  XNOR U10031 ( .A(n7395), .B(n7394), .Z(\w1[8][113] ) );
  XNOR U10032 ( .A(\w3[7][107] ), .B(\w3[7][115] ), .Z(n7431) );
  XNOR U10033 ( .A(n7431), .B(key[1138]), .Z(n7397) );
  XNOR U10034 ( .A(\w3[7][106] ), .B(n7763), .Z(n7396) );
  XNOR U10035 ( .A(n7397), .B(n7396), .Z(\w1[8][114] ) );
  XOR U10036 ( .A(\w3[7][116] ), .B(n7421), .Z(n7432) );
  XNOR U10037 ( .A(n7432), .B(key[1139]), .Z(n7400) );
  XOR U10038 ( .A(\w3[7][107] ), .B(n7398), .Z(n7399) );
  XNOR U10039 ( .A(n7400), .B(n7399), .Z(\w1[8][115] ) );
  XOR U10040 ( .A(\w3[7][117] ), .B(n7421), .Z(n7433) );
  XNOR U10041 ( .A(n7433), .B(key[1140]), .Z(n7403) );
  XOR U10042 ( .A(\w3[7][108] ), .B(n7401), .Z(n7402) );
  XNOR U10043 ( .A(n7403), .B(n7402), .Z(\w1[8][116] ) );
  XNOR U10044 ( .A(n7404), .B(key[1141]), .Z(n7407) );
  XNOR U10045 ( .A(\w3[7][109] ), .B(n7405), .Z(n7406) );
  XNOR U10046 ( .A(n7407), .B(n7406), .Z(\w1[8][117] ) );
  XOR U10047 ( .A(\w3[7][119] ), .B(n7421), .Z(n7442) );
  XNOR U10048 ( .A(n7442), .B(key[1142]), .Z(n7410) );
  XOR U10049 ( .A(\w3[7][110] ), .B(n7408), .Z(n7409) );
  XNOR U10050 ( .A(n7410), .B(n7409), .Z(\w1[8][118] ) );
  XOR U10051 ( .A(n7411), .B(key[1143]), .Z(n7414) );
  XNOR U10052 ( .A(\w3[7][112] ), .B(n7412), .Z(n7413) );
  XNOR U10053 ( .A(n7414), .B(n7413), .Z(\w1[8][119] ) );
  XNOR U10054 ( .A(\w3[7][3] ), .B(\w3[7][27] ), .Z(n7506) );
  XNOR U10055 ( .A(n7466), .B(key[1035]), .Z(n7416) );
  XNOR U10056 ( .A(\w3[7][0] ), .B(\w3[7][4] ), .Z(n7538) );
  XOR U10057 ( .A(\w3[7][19] ), .B(n7538), .Z(n7415) );
  XNOR U10058 ( .A(n7416), .B(n7415), .Z(\w1[8][11] ) );
  XNOR U10059 ( .A(n7417), .B(key[1144]), .Z(n7419) );
  XNOR U10060 ( .A(\w3[7][113] ), .B(\w3[7][121] ), .Z(n7418) );
  XNOR U10061 ( .A(n7419), .B(n7418), .Z(n7420) );
  XNOR U10062 ( .A(n7421), .B(n7420), .Z(\w1[8][120] ) );
  XNOR U10063 ( .A(n7762), .B(key[1145]), .Z(n7423) );
  XNOR U10064 ( .A(\w3[7][122] ), .B(\w3[7][114] ), .Z(n7422) );
  XNOR U10065 ( .A(n7423), .B(n7422), .Z(n7424) );
  XNOR U10066 ( .A(n7425), .B(n7424), .Z(\w1[8][121] ) );
  XNOR U10067 ( .A(n7766), .B(key[1146]), .Z(n7427) );
  XNOR U10068 ( .A(\w3[7][115] ), .B(\w3[7][123] ), .Z(n7426) );
  XNOR U10069 ( .A(n7427), .B(n7426), .Z(n7428) );
  XOR U10070 ( .A(\w3[7][98] ), .B(n7428), .Z(\w1[8][122] ) );
  XOR U10071 ( .A(\w3[7][124] ), .B(n7429), .Z(n7430) );
  XOR U10072 ( .A(n7431), .B(n7430), .Z(n7770) );
  XNOR U10073 ( .A(n7433), .B(key[1148]), .Z(n7437) );
  XNOR U10074 ( .A(n7435), .B(n7434), .Z(n7436) );
  XNOR U10075 ( .A(n7437), .B(n7436), .Z(\w1[8][124] ) );
  XOR U10076 ( .A(\w3[7][118] ), .B(key[1149]), .Z(n7440) );
  XOR U10077 ( .A(n7438), .B(\w3[7][126] ), .Z(n7439) );
  XNOR U10078 ( .A(n7440), .B(n7439), .Z(n7441) );
  XOR U10079 ( .A(\w3[7][101] ), .B(n7441), .Z(\w1[8][125] ) );
  XNOR U10080 ( .A(n7442), .B(key[1150]), .Z(n7445) );
  XOR U10081 ( .A(\w3[7][102] ), .B(n7443), .Z(n7444) );
  XNOR U10082 ( .A(n7445), .B(n7444), .Z(\w1[8][126] ) );
  XNOR U10083 ( .A(n7759), .B(key[1151]), .Z(n7448) );
  XOR U10084 ( .A(\w3[7][103] ), .B(n7446), .Z(n7447) );
  XNOR U10085 ( .A(n7448), .B(n7447), .Z(\w1[8][127] ) );
  XOR U10086 ( .A(\w3[7][13] ), .B(\w3[7][28] ), .Z(n7450) );
  XNOR U10087 ( .A(\w3[7][8] ), .B(\w3[7][4] ), .Z(n7449) );
  XOR U10088 ( .A(n7450), .B(n7449), .Z(n7470) );
  XNOR U10089 ( .A(n7470), .B(key[1036]), .Z(n7452) );
  XNOR U10090 ( .A(\w3[7][0] ), .B(\w3[7][5] ), .Z(n7576) );
  XOR U10091 ( .A(\w3[7][20] ), .B(n7576), .Z(n7451) );
  XNOR U10092 ( .A(n7452), .B(n7451), .Z(\w1[8][12] ) );
  IV U10093 ( .A(\w3[7][6] ), .Z(n7512) );
  XNOR U10094 ( .A(\w3[7][14] ), .B(n7512), .Z(n7454) );
  XNOR U10095 ( .A(\w3[7][5] ), .B(\w3[7][29] ), .Z(n7473) );
  XOR U10096 ( .A(n7473), .B(key[1037]), .Z(n7453) );
  XNOR U10097 ( .A(n7454), .B(n7453), .Z(n7455) );
  XOR U10098 ( .A(\w3[7][21] ), .B(n7455), .Z(\w1[8][13] ) );
  IV U10099 ( .A(\w3[7][30] ), .Z(n7655) );
  XOR U10100 ( .A(\w3[7][6] ), .B(n7655), .Z(n7620) );
  XOR U10101 ( .A(\w3[7][8] ), .B(\w3[7][15] ), .Z(n7476) );
  XNOR U10102 ( .A(n7620), .B(n7476), .Z(n7474) );
  XOR U10103 ( .A(n7474), .B(key[1038]), .Z(n7457) );
  XNOR U10104 ( .A(\w3[7][0] ), .B(\w3[7][7] ), .Z(n7656) );
  XOR U10105 ( .A(\w3[7][22] ), .B(n7656), .Z(n7456) );
  XNOR U10106 ( .A(n7457), .B(n7456), .Z(\w1[8][14] ) );
  XNOR U10107 ( .A(\w3[7][7] ), .B(\w3[7][31] ), .Z(n7475) );
  XNOR U10108 ( .A(n7475), .B(key[1039]), .Z(n7459) );
  XOR U10109 ( .A(\w3[7][8] ), .B(\w3[7][0] ), .Z(n7479) );
  XNOR U10110 ( .A(\w3[7][23] ), .B(n7479), .Z(n7458) );
  XNOR U10111 ( .A(n7459), .B(n7458), .Z(\w1[8][15] ) );
  XNOR U10112 ( .A(\w3[7][17] ), .B(\w3[7][9] ), .Z(n7481) );
  XNOR U10113 ( .A(n7481), .B(key[1040]), .Z(n7461) );
  XNOR U10114 ( .A(\w3[7][24] ), .B(n7479), .Z(n7460) );
  XNOR U10115 ( .A(n7461), .B(n7460), .Z(\w1[8][16] ) );
  XNOR U10116 ( .A(\w3[7][18] ), .B(\w3[7][10] ), .Z(n7505) );
  XNOR U10117 ( .A(n7505), .B(key[1041]), .Z(n7463) );
  IV U10118 ( .A(\w3[7][9] ), .Z(n7727) );
  XNOR U10119 ( .A(n7778), .B(n7727), .Z(n7462) );
  XNOR U10120 ( .A(n7463), .B(n7462), .Z(\w1[8][17] ) );
  IV U10121 ( .A(\w3[7][19] ), .Z(n7486) );
  XOR U10122 ( .A(\w3[7][11] ), .B(n7486), .Z(n7491) );
  XNOR U10123 ( .A(n7491), .B(key[1042]), .Z(n7465) );
  XOR U10124 ( .A(n7467), .B(\w3[7][10] ), .Z(n7464) );
  XNOR U10125 ( .A(n7465), .B(n7464), .Z(\w1[8][18] ) );
  XOR U10126 ( .A(n7480), .B(\w3[7][20] ), .Z(n7492) );
  XNOR U10127 ( .A(n7481), .B(key[1025]), .Z(n7469) );
  XOR U10128 ( .A(\w3[7][25] ), .B(n7467), .Z(n7468) );
  XNOR U10129 ( .A(n7469), .B(n7468), .Z(\w1[8][1] ) );
  IV U10130 ( .A(\w3[7][21] ), .Z(n7500) );
  XOR U10131 ( .A(\w3[7][16] ), .B(n7500), .Z(n7497) );
  XNOR U10132 ( .A(n7497), .B(key[1044]), .Z(n7472) );
  XOR U10133 ( .A(\w3[7][12] ), .B(n7470), .Z(n7471) );
  XNOR U10134 ( .A(n7472), .B(n7471), .Z(\w1[8][20] ) );
  IV U10135 ( .A(\w3[7][22] ), .Z(n7501) );
  XOR U10136 ( .A(\w3[7][14] ), .B(n7501), .Z(n7510) );
  XOR U10137 ( .A(n7480), .B(\w3[7][23] ), .Z(n7511) );
  XNOR U10138 ( .A(n7475), .B(key[1047]), .Z(n7478) );
  XNOR U10139 ( .A(\w3[7][16] ), .B(n7476), .Z(n7477) );
  XNOR U10140 ( .A(n7478), .B(n7477), .Z(\w1[8][23] ) );
  XNOR U10141 ( .A(n7481), .B(key[1049]), .Z(n7483) );
  XNOR U10142 ( .A(\w3[7][1] ), .B(\w3[7][26] ), .Z(n7482) );
  XNOR U10143 ( .A(n7483), .B(n7482), .Z(n7484) );
  XNOR U10144 ( .A(n7485), .B(n7484), .Z(\w1[8][25] ) );
  XNOR U10145 ( .A(n7505), .B(key[1050]), .Z(n7488) );
  XOR U10146 ( .A(\w3[7][2] ), .B(n7486), .Z(n7487) );
  XNOR U10147 ( .A(n7488), .B(n7487), .Z(n7489) );
  XOR U10148 ( .A(\w3[7][27] ), .B(n7489), .Z(\w1[8][26] ) );
  IV U10149 ( .A(\w3[7][24] ), .Z(n7509) );
  XOR U10150 ( .A(n7509), .B(\w3[7][28] ), .Z(n7490) );
  XOR U10151 ( .A(n7491), .B(n7490), .Z(n7537) );
  XOR U10152 ( .A(n7537), .B(key[1051]), .Z(n7494) );
  XOR U10153 ( .A(\w3[7][3] ), .B(n7492), .Z(n7493) );
  XNOR U10154 ( .A(n7494), .B(n7493), .Z(\w1[8][27] ) );
  XOR U10155 ( .A(\w3[7][20] ), .B(\w3[7][29] ), .Z(n7496) );
  XOR U10156 ( .A(n7509), .B(\w3[7][12] ), .Z(n7495) );
  XOR U10157 ( .A(n7496), .B(n7495), .Z(n7575) );
  XNOR U10158 ( .A(n7575), .B(key[1052]), .Z(n7499) );
  XOR U10159 ( .A(\w3[7][4] ), .B(n7497), .Z(n7498) );
  XNOR U10160 ( .A(n7499), .B(n7498), .Z(\w1[8][28] ) );
  XOR U10161 ( .A(\w3[7][13] ), .B(n7500), .Z(n7619) );
  XNOR U10162 ( .A(n7619), .B(key[1053]), .Z(n7503) );
  XNOR U10163 ( .A(n7501), .B(n7655), .Z(n7502) );
  XNOR U10164 ( .A(n7503), .B(n7502), .Z(n7504) );
  XOR U10165 ( .A(\w3[7][5] ), .B(n7504), .Z(\w1[8][29] ) );
  XNOR U10166 ( .A(n7505), .B(key[1026]), .Z(n7508) );
  XOR U10167 ( .A(\w3[7][26] ), .B(n7506), .Z(n7507) );
  XNOR U10168 ( .A(n7508), .B(n7507), .Z(\w1[8][2] ) );
  XOR U10169 ( .A(n7509), .B(\w3[7][31] ), .Z(n7691) );
  XNOR U10170 ( .A(n7510), .B(n7691), .Z(n7654) );
  XNOR U10171 ( .A(n7654), .B(key[1054]), .Z(n7514) );
  XNOR U10172 ( .A(n7512), .B(n7511), .Z(n7513) );
  XNOR U10173 ( .A(n7514), .B(n7513), .Z(\w1[8][30] ) );
  XNOR U10174 ( .A(\w3[7][15] ), .B(\w3[7][23] ), .Z(n7690) );
  XNOR U10175 ( .A(n7690), .B(key[1055]), .Z(n7516) );
  XOR U10176 ( .A(n7730), .B(\w3[7][7] ), .Z(n7515) );
  XNOR U10177 ( .A(n7516), .B(n7515), .Z(\w1[8][31] ) );
  XNOR U10178 ( .A(\w3[7][48] ), .B(\w3[7][56] ), .Z(n7636) );
  XOR U10179 ( .A(\w3[7][33] ), .B(\w3[7][57] ), .Z(n7572) );
  XNOR U10180 ( .A(\w3[7][40] ), .B(key[1056]), .Z(n7517) );
  XOR U10181 ( .A(n7572), .B(n7517), .Z(n7518) );
  XOR U10182 ( .A(n7636), .B(n7518), .Z(\w1[8][32] ) );
  XOR U10183 ( .A(\w3[7][49] ), .B(\w3[7][41] ), .Z(n7569) );
  XOR U10184 ( .A(n7569), .B(key[1057]), .Z(n7520) );
  XNOR U10185 ( .A(\w3[7][34] ), .B(\w3[7][58] ), .Z(n7580) );
  XOR U10186 ( .A(\w3[7][57] ), .B(n7580), .Z(n7519) );
  XNOR U10187 ( .A(n7520), .B(n7519), .Z(\w1[8][33] ) );
  XNOR U10188 ( .A(n7549), .B(key[1058]), .Z(n7522) );
  XNOR U10189 ( .A(\w3[7][50] ), .B(\w3[7][42] ), .Z(n7610) );
  XOR U10190 ( .A(\w3[7][58] ), .B(n7610), .Z(n7521) );
  XNOR U10191 ( .A(n7522), .B(n7521), .Z(\w1[8][34] ) );
  XOR U10192 ( .A(\w3[7][36] ), .B(\w3[7][32] ), .Z(n7551) );
  XOR U10193 ( .A(n7551), .B(key[1059]), .Z(n7525) );
  IV U10194 ( .A(\w3[7][51] ), .Z(n7609) );
  XOR U10195 ( .A(\w3[7][43] ), .B(n7609), .Z(n7579) );
  XOR U10196 ( .A(\w3[7][56] ), .B(n7579), .Z(n7523) );
  XNOR U10197 ( .A(\w3[7][60] ), .B(n7523), .Z(n7615) );
  XNOR U10198 ( .A(\w3[7][59] ), .B(n7615), .Z(n7524) );
  XNOR U10199 ( .A(n7525), .B(n7524), .Z(\w1[8][35] ) );
  XOR U10200 ( .A(\w3[7][32] ), .B(\w3[7][37] ), .Z(n7557) );
  XOR U10201 ( .A(\w3[7][52] ), .B(\w3[7][61] ), .Z(n7527) );
  XNOR U10202 ( .A(\w3[7][56] ), .B(\w3[7][44] ), .Z(n7526) );
  XOR U10203 ( .A(n7527), .B(n7526), .Z(n7624) );
  XOR U10204 ( .A(n7624), .B(key[1060]), .Z(n7528) );
  XOR U10205 ( .A(n7557), .B(n7528), .Z(n7529) );
  XNOR U10206 ( .A(\w3[7][60] ), .B(n7529), .Z(\w1[8][36] ) );
  XNOR U10207 ( .A(\w3[7][38] ), .B(\w3[7][62] ), .Z(n7563) );
  XNOR U10208 ( .A(n7563), .B(key[1061]), .Z(n7531) );
  IV U10209 ( .A(\w3[7][45] ), .Z(n7589) );
  XOR U10210 ( .A(\w3[7][53] ), .B(n7589), .Z(n7627) );
  XOR U10211 ( .A(\w3[7][61] ), .B(n7627), .Z(n7530) );
  XNOR U10212 ( .A(n7531), .B(n7530), .Z(\w1[8][37] ) );
  XOR U10213 ( .A(\w3[7][32] ), .B(\w3[7][39] ), .Z(n7564) );
  XOR U10214 ( .A(n7564), .B(key[1062]), .Z(n7533) );
  XNOR U10215 ( .A(\w3[7][56] ), .B(\w3[7][63] ), .Z(n7534) );
  XOR U10216 ( .A(\w3[7][46] ), .B(\w3[7][54] ), .Z(n7588) );
  XOR U10217 ( .A(n7534), .B(n7588), .Z(n7632) );
  XOR U10218 ( .A(\w3[7][62] ), .B(n7632), .Z(n7532) );
  XNOR U10219 ( .A(n7533), .B(n7532), .Z(\w1[8][38] ) );
  XNOR U10220 ( .A(\w3[7][55] ), .B(\w3[7][47] ), .Z(n7635) );
  XNOR U10221 ( .A(n7635), .B(key[1063]), .Z(n7536) );
  XOR U10222 ( .A(\w3[7][32] ), .B(n7534), .Z(n7535) );
  XNOR U10223 ( .A(n7536), .B(n7535), .Z(\w1[8][39] ) );
  XOR U10224 ( .A(n7537), .B(key[1027]), .Z(n7540) );
  XOR U10225 ( .A(n7538), .B(\w3[7][27] ), .Z(n7539) );
  XNOR U10226 ( .A(n7540), .B(n7539), .Z(\w1[8][3] ) );
  XNOR U10227 ( .A(\w3[7][33] ), .B(\w3[7][41] ), .Z(n7604) );
  XNOR U10228 ( .A(n7604), .B(key[1064]), .Z(n7542) );
  XOR U10229 ( .A(n7636), .B(\w3[7][32] ), .Z(n7541) );
  XNOR U10230 ( .A(n7542), .B(n7541), .Z(\w1[8][40] ) );
  XOR U10231 ( .A(\w3[7][42] ), .B(key[1065]), .Z(n7544) );
  IV U10232 ( .A(\w3[7][49] ), .Z(n7605) );
  XOR U10233 ( .A(\w3[7][34] ), .B(n7605), .Z(n7543) );
  XNOR U10234 ( .A(n7544), .B(n7543), .Z(n7545) );
  XOR U10235 ( .A(n7545), .B(n7572), .Z(\w1[8][41] ) );
  XOR U10236 ( .A(\w3[7][43] ), .B(key[1066]), .Z(n7547) );
  IV U10237 ( .A(\w3[7][35] ), .Z(n7616) );
  XOR U10238 ( .A(\w3[7][50] ), .B(n7616), .Z(n7546) );
  XNOR U10239 ( .A(n7547), .B(n7546), .Z(n7548) );
  XNOR U10240 ( .A(n7580), .B(n7548), .Z(\w1[8][42] ) );
  IV U10241 ( .A(\w3[7][40] ), .Z(n7554) );
  XNOR U10242 ( .A(n7554), .B(n7549), .Z(n7550) );
  XOR U10243 ( .A(\w3[7][44] ), .B(n7550), .Z(n7583) );
  XNOR U10244 ( .A(n7583), .B(key[1067]), .Z(n7553) );
  XNOR U10245 ( .A(\w3[7][51] ), .B(n7551), .Z(n7552) );
  XNOR U10246 ( .A(n7553), .B(n7552), .Z(\w1[8][43] ) );
  XOR U10247 ( .A(\w3[7][36] ), .B(\w3[7][45] ), .Z(n7556) );
  XOR U10248 ( .A(n7554), .B(\w3[7][60] ), .Z(n7555) );
  XOR U10249 ( .A(n7556), .B(n7555), .Z(n7584) );
  XNOR U10250 ( .A(n7584), .B(key[1068]), .Z(n7559) );
  XNOR U10251 ( .A(\w3[7][52] ), .B(n7557), .Z(n7558) );
  XNOR U10252 ( .A(n7559), .B(n7558), .Z(\w1[8][44] ) );
  XNOR U10253 ( .A(\w3[7][61] ), .B(\w3[7][37] ), .Z(n7587) );
  XNOR U10254 ( .A(n7587), .B(key[1069]), .Z(n7561) );
  XNOR U10255 ( .A(\w3[7][38] ), .B(\w3[7][46] ), .Z(n7560) );
  XNOR U10256 ( .A(n7561), .B(n7560), .Z(n7562) );
  XOR U10257 ( .A(\w3[7][53] ), .B(n7562), .Z(\w1[8][45] ) );
  XOR U10258 ( .A(\w3[7][40] ), .B(\w3[7][47] ), .Z(n7596) );
  XOR U10259 ( .A(n7563), .B(n7596), .Z(n7592) );
  XNOR U10260 ( .A(n7592), .B(key[1070]), .Z(n7566) );
  XNOR U10261 ( .A(\w3[7][54] ), .B(n7564), .Z(n7565) );
  XNOR U10262 ( .A(n7566), .B(n7565), .Z(\w1[8][46] ) );
  XOR U10263 ( .A(\w3[7][63] ), .B(\w3[7][39] ), .Z(n7595) );
  XOR U10264 ( .A(n7595), .B(key[1071]), .Z(n7568) );
  XNOR U10265 ( .A(\w3[7][40] ), .B(\w3[7][32] ), .Z(n7599) );
  XOR U10266 ( .A(\w3[7][55] ), .B(n7599), .Z(n7567) );
  XNOR U10267 ( .A(n7568), .B(n7567), .Z(\w1[8][47] ) );
  XNOR U10268 ( .A(n7599), .B(key[1072]), .Z(n7571) );
  XNOR U10269 ( .A(\w3[7][56] ), .B(n7569), .Z(n7570) );
  XNOR U10270 ( .A(n7571), .B(n7570), .Z(\w1[8][48] ) );
  XNOR U10271 ( .A(n7610), .B(key[1073]), .Z(n7574) );
  XNOR U10272 ( .A(n7572), .B(\w3[7][41] ), .Z(n7573) );
  XNOR U10273 ( .A(n7574), .B(n7573), .Z(\w1[8][49] ) );
  XNOR U10274 ( .A(n7575), .B(key[1028]), .Z(n7578) );
  XOR U10275 ( .A(n7576), .B(\w3[7][28] ), .Z(n7577) );
  XNOR U10276 ( .A(n7578), .B(n7577), .Z(\w1[8][4] ) );
  XNOR U10277 ( .A(n7579), .B(key[1074]), .Z(n7582) );
  XOR U10278 ( .A(n7580), .B(\w3[7][42] ), .Z(n7581) );
  XNOR U10279 ( .A(n7582), .B(n7581), .Z(\w1[8][50] ) );
  IV U10280 ( .A(\w3[7][48] ), .Z(n7600) );
  XOR U10281 ( .A(n7600), .B(\w3[7][52] ), .Z(n7614) );
  XNOR U10282 ( .A(n7623), .B(key[1076]), .Z(n7586) );
  XOR U10283 ( .A(\w3[7][44] ), .B(n7584), .Z(n7585) );
  XNOR U10284 ( .A(n7586), .B(n7585), .Z(\w1[8][52] ) );
  XNOR U10285 ( .A(n7587), .B(key[1077]), .Z(n7591) );
  XOR U10286 ( .A(n7589), .B(n7588), .Z(n7590) );
  XNOR U10287 ( .A(n7591), .B(n7590), .Z(\w1[8][53] ) );
  XOR U10288 ( .A(n7600), .B(\w3[7][55] ), .Z(n7631) );
  XNOR U10289 ( .A(n7631), .B(key[1078]), .Z(n7594) );
  XOR U10290 ( .A(\w3[7][46] ), .B(n7592), .Z(n7593) );
  XNOR U10291 ( .A(n7594), .B(n7593), .Z(\w1[8][54] ) );
  XOR U10292 ( .A(n7595), .B(key[1079]), .Z(n7598) );
  XNOR U10293 ( .A(\w3[7][48] ), .B(n7596), .Z(n7597) );
  XNOR U10294 ( .A(n7598), .B(n7597), .Z(\w1[8][55] ) );
  XNOR U10295 ( .A(n7599), .B(key[1080]), .Z(n7602) );
  XOR U10296 ( .A(n7600), .B(\w3[7][49] ), .Z(n7601) );
  XNOR U10297 ( .A(n7602), .B(n7601), .Z(n7603) );
  XOR U10298 ( .A(\w3[7][57] ), .B(n7603), .Z(\w1[8][56] ) );
  XNOR U10299 ( .A(n7604), .B(key[1081]), .Z(n7607) );
  XOR U10300 ( .A(n7605), .B(\w3[7][50] ), .Z(n7606) );
  XNOR U10301 ( .A(n7607), .B(n7606), .Z(n7608) );
  XOR U10302 ( .A(\w3[7][58] ), .B(n7608), .Z(\w1[8][57] ) );
  XNOR U10303 ( .A(n7609), .B(key[1082]), .Z(n7612) );
  XOR U10304 ( .A(n7610), .B(\w3[7][59] ), .Z(n7611) );
  XNOR U10305 ( .A(n7612), .B(n7611), .Z(n7613) );
  XOR U10306 ( .A(\w3[7][34] ), .B(n7613), .Z(\w1[8][58] ) );
  XNOR U10307 ( .A(n7614), .B(key[1083]), .Z(n7618) );
  XOR U10308 ( .A(n7616), .B(n7615), .Z(n7617) );
  XNOR U10309 ( .A(n7618), .B(n7617), .Z(\w1[8][59] ) );
  XNOR U10310 ( .A(n7619), .B(key[1029]), .Z(n7622) );
  XOR U10311 ( .A(\w3[7][29] ), .B(n7620), .Z(n7621) );
  XNOR U10312 ( .A(n7622), .B(n7621), .Z(\w1[8][5] ) );
  XNOR U10313 ( .A(n7623), .B(key[1084]), .Z(n7626) );
  XOR U10314 ( .A(\w3[7][36] ), .B(n7624), .Z(n7625) );
  XNOR U10315 ( .A(n7626), .B(n7625), .Z(\w1[8][60] ) );
  XOR U10316 ( .A(\w3[7][54] ), .B(key[1085]), .Z(n7629) );
  XOR U10317 ( .A(n7627), .B(\w3[7][62] ), .Z(n7628) );
  XNOR U10318 ( .A(n7629), .B(n7628), .Z(n7630) );
  XOR U10319 ( .A(\w3[7][37] ), .B(n7630), .Z(\w1[8][61] ) );
  XNOR U10320 ( .A(n7631), .B(key[1086]), .Z(n7634) );
  XOR U10321 ( .A(\w3[7][38] ), .B(n7632), .Z(n7633) );
  XNOR U10322 ( .A(n7634), .B(n7633), .Z(\w1[8][62] ) );
  XNOR U10323 ( .A(n7635), .B(key[1087]), .Z(n7638) );
  XOR U10324 ( .A(n7636), .B(\w3[7][39] ), .Z(n7637) );
  XNOR U10325 ( .A(n7638), .B(n7637), .Z(\w1[8][63] ) );
  XOR U10326 ( .A(\w3[7][65] ), .B(\w3[7][89] ), .Z(n7696) );
  XOR U10327 ( .A(n7696), .B(key[1088]), .Z(n7640) );
  XNOR U10328 ( .A(\w3[7][80] ), .B(\w3[7][88] ), .Z(n7755) );
  XOR U10329 ( .A(n7755), .B(\w3[7][72] ), .Z(n7639) );
  XNOR U10330 ( .A(n7640), .B(n7639), .Z(\w1[8][64] ) );
  XNOR U10331 ( .A(\w3[7][66] ), .B(\w3[7][90] ), .Z(n7700) );
  XOR U10332 ( .A(\w3[7][89] ), .B(\w3[7][81] ), .Z(n7718) );
  XNOR U10333 ( .A(n7718), .B(key[1089]), .Z(n7641) );
  XNOR U10334 ( .A(n7700), .B(n7641), .Z(n7642) );
  XNOR U10335 ( .A(\w3[7][73] ), .B(n7642), .Z(\w1[8][65] ) );
  XNOR U10336 ( .A(n7670), .B(key[1090]), .Z(n7644) );
  XNOR U10337 ( .A(\w3[7][82] ), .B(\w3[7][74] ), .Z(n7733) );
  XOR U10338 ( .A(\w3[7][90] ), .B(n7733), .Z(n7643) );
  XNOR U10339 ( .A(n7644), .B(n7643), .Z(\w1[8][66] ) );
  XOR U10340 ( .A(\w3[7][68] ), .B(\w3[7][64] ), .Z(n7672) );
  XOR U10341 ( .A(n7672), .B(key[1091]), .Z(n7647) );
  IV U10342 ( .A(\w3[7][83] ), .Z(n7732) );
  XOR U10343 ( .A(\w3[7][75] ), .B(n7732), .Z(n7699) );
  XOR U10344 ( .A(\w3[7][88] ), .B(n7699), .Z(n7645) );
  XNOR U10345 ( .A(\w3[7][92] ), .B(n7645), .Z(n7738) );
  XNOR U10346 ( .A(\w3[7][91] ), .B(n7738), .Z(n7646) );
  XNOR U10347 ( .A(n7647), .B(n7646), .Z(\w1[8][67] ) );
  XOR U10348 ( .A(\w3[7][64] ), .B(\w3[7][69] ), .Z(n7678) );
  XOR U10349 ( .A(\w3[7][84] ), .B(\w3[7][93] ), .Z(n7649) );
  XNOR U10350 ( .A(\w3[7][88] ), .B(\w3[7][76] ), .Z(n7648) );
  XOR U10351 ( .A(n7649), .B(n7648), .Z(n7743) );
  XOR U10352 ( .A(n7743), .B(key[1092]), .Z(n7650) );
  XOR U10353 ( .A(n7678), .B(n7650), .Z(n7651) );
  XNOR U10354 ( .A(\w3[7][92] ), .B(n7651), .Z(\w1[8][68] ) );
  XNOR U10355 ( .A(\w3[7][70] ), .B(\w3[7][94] ), .Z(n7684) );
  XNOR U10356 ( .A(n7684), .B(key[1093]), .Z(n7653) );
  IV U10357 ( .A(\w3[7][77] ), .Z(n7707) );
  XOR U10358 ( .A(\w3[7][85] ), .B(n7707), .Z(n7746) );
  XOR U10359 ( .A(\w3[7][93] ), .B(n7746), .Z(n7652) );
  XNOR U10360 ( .A(n7653), .B(n7652), .Z(\w1[8][69] ) );
  XNOR U10361 ( .A(n7654), .B(key[1030]), .Z(n7658) );
  XNOR U10362 ( .A(n7656), .B(n7655), .Z(n7657) );
  XNOR U10363 ( .A(n7658), .B(n7657), .Z(\w1[8][6] ) );
  XOR U10364 ( .A(\w3[7][64] ), .B(\w3[7][71] ), .Z(n7685) );
  XOR U10365 ( .A(n7685), .B(key[1094]), .Z(n7660) );
  XNOR U10366 ( .A(\w3[7][88] ), .B(\w3[7][95] ), .Z(n7661) );
  XOR U10367 ( .A(\w3[7][78] ), .B(\w3[7][86] ), .Z(n7706) );
  XOR U10368 ( .A(n7661), .B(n7706), .Z(n7751) );
  XOR U10369 ( .A(\w3[7][94] ), .B(n7751), .Z(n7659) );
  XNOR U10370 ( .A(n7660), .B(n7659), .Z(\w1[8][70] ) );
  XNOR U10371 ( .A(\w3[7][79] ), .B(\w3[7][87] ), .Z(n7754) );
  XNOR U10372 ( .A(n7754), .B(key[1095]), .Z(n7663) );
  XOR U10373 ( .A(\w3[7][64] ), .B(n7661), .Z(n7662) );
  XNOR U10374 ( .A(n7663), .B(n7662), .Z(\w1[8][71] ) );
  IV U10375 ( .A(\w3[7][65] ), .Z(n7723) );
  XOR U10376 ( .A(\w3[7][74] ), .B(key[1097]), .Z(n7665) );
  XNOR U10377 ( .A(n7718), .B(\w3[7][66] ), .Z(n7664) );
  XNOR U10378 ( .A(n7665), .B(n7664), .Z(n7666) );
  XNOR U10379 ( .A(n7723), .B(n7666), .Z(\w1[8][73] ) );
  XOR U10380 ( .A(\w3[7][75] ), .B(key[1098]), .Z(n7668) );
  IV U10381 ( .A(\w3[7][67] ), .Z(n7739) );
  XOR U10382 ( .A(\w3[7][82] ), .B(n7739), .Z(n7667) );
  XNOR U10383 ( .A(n7668), .B(n7667), .Z(n7669) );
  XNOR U10384 ( .A(n7669), .B(n7700), .Z(\w1[8][74] ) );
  IV U10385 ( .A(\w3[7][72] ), .Z(n7675) );
  XNOR U10386 ( .A(n7675), .B(n7670), .Z(n7671) );
  XOR U10387 ( .A(\w3[7][76] ), .B(n7671), .Z(n7701) );
  XNOR U10388 ( .A(n7701), .B(key[1099]), .Z(n7674) );
  XNOR U10389 ( .A(\w3[7][83] ), .B(n7672), .Z(n7673) );
  XNOR U10390 ( .A(n7674), .B(n7673), .Z(\w1[8][75] ) );
  XOR U10391 ( .A(\w3[7][68] ), .B(\w3[7][77] ), .Z(n7677) );
  XOR U10392 ( .A(n7675), .B(\w3[7][92] ), .Z(n7676) );
  XOR U10393 ( .A(n7677), .B(n7676), .Z(n7702) );
  XNOR U10394 ( .A(n7702), .B(key[1100]), .Z(n7680) );
  XNOR U10395 ( .A(\w3[7][84] ), .B(n7678), .Z(n7679) );
  XNOR U10396 ( .A(n7680), .B(n7679), .Z(\w1[8][76] ) );
  XNOR U10397 ( .A(\w3[7][93] ), .B(\w3[7][69] ), .Z(n7705) );
  XNOR U10398 ( .A(n7705), .B(key[1101]), .Z(n7682) );
  XNOR U10399 ( .A(\w3[7][70] ), .B(\w3[7][78] ), .Z(n7681) );
  XNOR U10400 ( .A(n7682), .B(n7681), .Z(n7683) );
  XOR U10401 ( .A(\w3[7][85] ), .B(n7683), .Z(\w1[8][77] ) );
  XOR U10402 ( .A(\w3[7][72] ), .B(\w3[7][79] ), .Z(n7714) );
  XOR U10403 ( .A(n7684), .B(n7714), .Z(n7710) );
  XNOR U10404 ( .A(n7710), .B(key[1102]), .Z(n7687) );
  XNOR U10405 ( .A(\w3[7][86] ), .B(n7685), .Z(n7686) );
  XNOR U10406 ( .A(n7687), .B(n7686), .Z(\w1[8][78] ) );
  XOR U10407 ( .A(\w3[7][95] ), .B(\w3[7][71] ), .Z(n7713) );
  XOR U10408 ( .A(n7713), .B(key[1103]), .Z(n7689) );
  XNOR U10409 ( .A(\w3[7][72] ), .B(\w3[7][64] ), .Z(n7717) );
  XOR U10410 ( .A(\w3[7][87] ), .B(n7717), .Z(n7688) );
  XNOR U10411 ( .A(n7689), .B(n7688), .Z(\w1[8][79] ) );
  XNOR U10412 ( .A(n7690), .B(key[1031]), .Z(n7693) );
  XOR U10413 ( .A(\w3[7][0] ), .B(n7691), .Z(n7692) );
  XNOR U10414 ( .A(n7693), .B(n7692), .Z(\w1[8][7] ) );
  XNOR U10415 ( .A(\w3[7][73] ), .B(\w3[7][81] ), .Z(n7722) );
  XNOR U10416 ( .A(n7722), .B(key[1104]), .Z(n7695) );
  XOR U10417 ( .A(\w3[7][88] ), .B(n7717), .Z(n7694) );
  XNOR U10418 ( .A(n7695), .B(n7694), .Z(\w1[8][80] ) );
  XNOR U10419 ( .A(n7733), .B(key[1105]), .Z(n7698) );
  XNOR U10420 ( .A(n7696), .B(\w3[7][73] ), .Z(n7697) );
  XNOR U10421 ( .A(n7698), .B(n7697), .Z(\w1[8][81] ) );
  IV U10422 ( .A(\w3[7][80] ), .Z(n7719) );
  XOR U10423 ( .A(n7719), .B(\w3[7][84] ), .Z(n7737) );
  XNOR U10424 ( .A(n7742), .B(key[1108]), .Z(n7704) );
  XOR U10425 ( .A(\w3[7][76] ), .B(n7702), .Z(n7703) );
  XNOR U10426 ( .A(n7704), .B(n7703), .Z(\w1[8][84] ) );
  XNOR U10427 ( .A(n7705), .B(key[1109]), .Z(n7709) );
  XOR U10428 ( .A(n7707), .B(n7706), .Z(n7708) );
  XNOR U10429 ( .A(n7709), .B(n7708), .Z(\w1[8][85] ) );
  XOR U10430 ( .A(n7719), .B(\w3[7][87] ), .Z(n7750) );
  XNOR U10431 ( .A(n7750), .B(key[1110]), .Z(n7712) );
  XOR U10432 ( .A(\w3[7][78] ), .B(n7710), .Z(n7711) );
  XNOR U10433 ( .A(n7712), .B(n7711), .Z(\w1[8][86] ) );
  XOR U10434 ( .A(n7713), .B(key[1111]), .Z(n7716) );
  XNOR U10435 ( .A(\w3[7][80] ), .B(n7714), .Z(n7715) );
  XNOR U10436 ( .A(n7716), .B(n7715), .Z(\w1[8][87] ) );
  XNOR U10437 ( .A(n7717), .B(key[1112]), .Z(n7721) );
  XOR U10438 ( .A(n7719), .B(n7718), .Z(n7720) );
  XNOR U10439 ( .A(n7721), .B(n7720), .Z(\w1[8][88] ) );
  XNOR U10440 ( .A(n7722), .B(key[1113]), .Z(n7725) );
  XOR U10441 ( .A(n7723), .B(\w3[7][82] ), .Z(n7724) );
  XNOR U10442 ( .A(n7725), .B(n7724), .Z(n7726) );
  XOR U10443 ( .A(\w3[7][90] ), .B(n7726), .Z(\w1[8][89] ) );
  XNOR U10444 ( .A(n7727), .B(key[1032]), .Z(n7729) );
  XNOR U10445 ( .A(\w3[7][1] ), .B(\w3[7][0] ), .Z(n7728) );
  XNOR U10446 ( .A(n7729), .B(n7728), .Z(n7731) );
  XNOR U10447 ( .A(n7731), .B(n7730), .Z(\w1[8][8] ) );
  XNOR U10448 ( .A(n7732), .B(key[1114]), .Z(n7735) );
  XOR U10449 ( .A(n7733), .B(\w3[7][91] ), .Z(n7734) );
  XNOR U10450 ( .A(n7735), .B(n7734), .Z(n7736) );
  XOR U10451 ( .A(\w3[7][66] ), .B(n7736), .Z(\w1[8][90] ) );
  XNOR U10452 ( .A(n7737), .B(key[1115]), .Z(n7741) );
  XOR U10453 ( .A(n7739), .B(n7738), .Z(n7740) );
  XNOR U10454 ( .A(n7741), .B(n7740), .Z(\w1[8][91] ) );
  XNOR U10455 ( .A(n7742), .B(key[1116]), .Z(n7745) );
  XOR U10456 ( .A(\w3[7][68] ), .B(n7743), .Z(n7744) );
  XNOR U10457 ( .A(n7745), .B(n7744), .Z(\w1[8][92] ) );
  XOR U10458 ( .A(\w3[7][86] ), .B(key[1117]), .Z(n7748) );
  XOR U10459 ( .A(n7746), .B(\w3[7][94] ), .Z(n7747) );
  XNOR U10460 ( .A(n7748), .B(n7747), .Z(n7749) );
  XOR U10461 ( .A(\w3[7][69] ), .B(n7749), .Z(\w1[8][93] ) );
  XNOR U10462 ( .A(n7750), .B(key[1118]), .Z(n7753) );
  XOR U10463 ( .A(\w3[7][70] ), .B(n7751), .Z(n7752) );
  XNOR U10464 ( .A(n7753), .B(n7752), .Z(\w1[8][94] ) );
  XNOR U10465 ( .A(n7754), .B(key[1119]), .Z(n7757) );
  XOR U10466 ( .A(n7755), .B(\w3[7][71] ), .Z(n7756) );
  XNOR U10467 ( .A(n7757), .B(n7756), .Z(\w1[8][95] ) );
  XOR U10468 ( .A(\w3[7][104] ), .B(key[1120]), .Z(n7761) );
  XNOR U10469 ( .A(n7759), .B(n7758), .Z(n7760) );
  XNOR U10470 ( .A(n7761), .B(n7760), .Z(\w1[8][96] ) );
  XNOR U10471 ( .A(n7762), .B(key[1121]), .Z(n7765) );
  XNOR U10472 ( .A(\w3[7][121] ), .B(n7763), .Z(n7764) );
  XNOR U10473 ( .A(n7765), .B(n7764), .Z(\w1[8][97] ) );
  XNOR U10474 ( .A(n7766), .B(key[1122]), .Z(n7769) );
  XOR U10475 ( .A(\w3[7][122] ), .B(n7767), .Z(n7768) );
  XNOR U10476 ( .A(n7769), .B(n7768), .Z(\w1[8][98] ) );
  XOR U10477 ( .A(n7770), .B(key[1123]), .Z(n7774) );
  XNOR U10478 ( .A(n7772), .B(n7771), .Z(n7773) );
  XNOR U10479 ( .A(n7774), .B(n7773), .Z(\w1[8][99] ) );
  XOR U10480 ( .A(\w3[7][10] ), .B(key[1033]), .Z(n7776) );
  XNOR U10481 ( .A(\w3[7][2] ), .B(\w3[7][17] ), .Z(n7775) );
  XNOR U10482 ( .A(n7776), .B(n7775), .Z(n7777) );
  XNOR U10483 ( .A(n7778), .B(n7777), .Z(\w1[8][9] ) );
  XNOR U10484 ( .A(\w3[8][25] ), .B(\w3[8][1] ), .Z(n8202) );
  IV U10485 ( .A(\w3[8][16] ), .Z(n7906) );
  XOR U10486 ( .A(\w3[8][24] ), .B(n7906), .Z(n8153) );
  XNOR U10487 ( .A(\w3[8][8] ), .B(key[1152]), .Z(n7779) );
  XNOR U10488 ( .A(n8153), .B(n7779), .Z(n7780) );
  XOR U10489 ( .A(n8202), .B(n7780), .Z(\w1[9][0] ) );
  XOR U10490 ( .A(\w3[8][96] ), .B(\w3[8][101] ), .Z(n7806) );
  XOR U10491 ( .A(\w3[8][116] ), .B(\w3[8][125] ), .Z(n7782) );
  IV U10492 ( .A(\w3[8][120] ), .Z(n7853) );
  XOR U10493 ( .A(n7853), .B(\w3[8][108] ), .Z(n7781) );
  XOR U10494 ( .A(n7782), .B(n7781), .Z(n7861) );
  XOR U10495 ( .A(n7861), .B(key[1252]), .Z(n7783) );
  XOR U10496 ( .A(n7806), .B(n7783), .Z(n7784) );
  XNOR U10497 ( .A(\w3[8][124] ), .B(n7784), .Z(\w1[9][100] ) );
  XNOR U10498 ( .A(\w3[8][102] ), .B(\w3[8][126] ), .Z(n7815) );
  XNOR U10499 ( .A(n7815), .B(key[1253]), .Z(n7786) );
  XNOR U10500 ( .A(\w3[8][109] ), .B(\w3[8][117] ), .Z(n7867) );
  XOR U10501 ( .A(\w3[8][125] ), .B(n7867), .Z(n7785) );
  XNOR U10502 ( .A(n7786), .B(n7785), .Z(\w1[9][101] ) );
  XOR U10503 ( .A(\w3[8][96] ), .B(\w3[8][103] ), .Z(n7816) );
  XOR U10504 ( .A(n7816), .B(key[1254]), .Z(n7788) );
  XOR U10505 ( .A(n7853), .B(\w3[8][127] ), .Z(n7789) );
  XOR U10506 ( .A(\w3[8][110] ), .B(\w3[8][118] ), .Z(n7832) );
  XOR U10507 ( .A(n7789), .B(n7832), .Z(n7869) );
  XOR U10508 ( .A(\w3[8][126] ), .B(n7869), .Z(n7787) );
  XNOR U10509 ( .A(n7788), .B(n7787), .Z(\w1[9][102] ) );
  XNOR U10510 ( .A(\w3[8][111] ), .B(\w3[8][119] ), .Z(n7872) );
  XNOR U10511 ( .A(n7872), .B(key[1255]), .Z(n7791) );
  XOR U10512 ( .A(\w3[8][96] ), .B(n7789), .Z(n7790) );
  XNOR U10513 ( .A(n7791), .B(n7790), .Z(\w1[9][103] ) );
  XOR U10514 ( .A(key[1256]), .B(\w3[8][105] ), .Z(n7793) );
  XNOR U10515 ( .A(\w3[8][96] ), .B(\w3[8][97] ), .Z(n7792) );
  XNOR U10516 ( .A(n7793), .B(n7792), .Z(n7794) );
  IV U10517 ( .A(\w3[8][112] ), .Z(n7848) );
  XOR U10518 ( .A(\w3[8][120] ), .B(n7848), .Z(n8183) );
  XNOR U10519 ( .A(n7794), .B(n8183), .Z(\w1[9][104] ) );
  XOR U10520 ( .A(\w3[8][106] ), .B(\w3[8][113] ), .Z(n7796) );
  XNOR U10521 ( .A(\w3[8][97] ), .B(\w3[8][121] ), .Z(n8182) );
  XOR U10522 ( .A(n8182), .B(key[1257]), .Z(n7795) );
  XNOR U10523 ( .A(n7796), .B(n7795), .Z(n7797) );
  XOR U10524 ( .A(\w3[8][98] ), .B(n7797), .Z(\w1[9][105] ) );
  IV U10525 ( .A(\w3[8][99] ), .Z(n7857) );
  XNOR U10526 ( .A(\w3[8][107] ), .B(n7857), .Z(n7799) );
  XOR U10527 ( .A(\w3[8][98] ), .B(\w3[8][122] ), .Z(n8187) );
  XNOR U10528 ( .A(n8187), .B(key[1258]), .Z(n7798) );
  XNOR U10529 ( .A(n7799), .B(n7798), .Z(n7800) );
  XOR U10530 ( .A(\w3[8][114] ), .B(n7800), .Z(\w1[9][106] ) );
  IV U10531 ( .A(\w3[8][123] ), .Z(n8195) );
  XOR U10532 ( .A(\w3[8][99] ), .B(n8195), .Z(n8191) );
  XOR U10533 ( .A(\w3[8][108] ), .B(n8191), .Z(n7801) );
  XOR U10534 ( .A(\w3[8][104] ), .B(n7801), .Z(n7827) );
  XNOR U10535 ( .A(n7827), .B(key[1259]), .Z(n7803) );
  XNOR U10536 ( .A(\w3[8][96] ), .B(\w3[8][100] ), .Z(n8196) );
  XOR U10537 ( .A(\w3[8][115] ), .B(n8196), .Z(n7802) );
  XNOR U10538 ( .A(n7803), .B(n7802), .Z(\w1[9][107] ) );
  XOR U10539 ( .A(\w3[8][100] ), .B(\w3[8][104] ), .Z(n7805) );
  XNOR U10540 ( .A(\w3[8][124] ), .B(\w3[8][109] ), .Z(n7804) );
  XOR U10541 ( .A(n7805), .B(n7804), .Z(n7828) );
  XNOR U10542 ( .A(n7828), .B(key[1260]), .Z(n7808) );
  XNOR U10543 ( .A(\w3[8][116] ), .B(n7806), .Z(n7807) );
  XNOR U10544 ( .A(n7808), .B(n7807), .Z(\w1[9][108] ) );
  XNOR U10545 ( .A(\w3[8][125] ), .B(\w3[8][101] ), .Z(n7831) );
  XNOR U10546 ( .A(n7831), .B(key[1261]), .Z(n7810) );
  XNOR U10547 ( .A(\w3[8][102] ), .B(\w3[8][110] ), .Z(n7809) );
  XNOR U10548 ( .A(n7810), .B(n7809), .Z(n7811) );
  XOR U10549 ( .A(\w3[8][117] ), .B(n7811), .Z(\w1[9][109] ) );
  IV U10550 ( .A(\w3[8][18] ), .Z(n7911) );
  XNOR U10551 ( .A(\w3[8][11] ), .B(n7911), .Z(n7813) );
  XNOR U10552 ( .A(\w3[8][2] ), .B(\w3[8][26] ), .Z(n7893) );
  XOR U10553 ( .A(n7893), .B(key[1162]), .Z(n7812) );
  XNOR U10554 ( .A(n7813), .B(n7812), .Z(n7814) );
  XOR U10555 ( .A(\w3[8][3] ), .B(n7814), .Z(\w1[9][10] ) );
  XOR U10556 ( .A(\w3[8][111] ), .B(\w3[8][104] ), .Z(n7839) );
  XOR U10557 ( .A(n7815), .B(n7839), .Z(n7835) );
  XNOR U10558 ( .A(n7835), .B(key[1262]), .Z(n7818) );
  XNOR U10559 ( .A(\w3[8][118] ), .B(n7816), .Z(n7817) );
  XNOR U10560 ( .A(n7818), .B(n7817), .Z(\w1[9][110] ) );
  XOR U10561 ( .A(\w3[8][127] ), .B(\w3[8][103] ), .Z(n7838) );
  XOR U10562 ( .A(n7838), .B(key[1263]), .Z(n7820) );
  XNOR U10563 ( .A(\w3[8][96] ), .B(\w3[8][104] ), .Z(n7844) );
  XOR U10564 ( .A(\w3[8][119] ), .B(n7844), .Z(n7819) );
  XNOR U10565 ( .A(n7820), .B(n7819), .Z(\w1[9][111] ) );
  XNOR U10566 ( .A(\w3[8][105] ), .B(\w3[8][113] ), .Z(n8186) );
  XNOR U10567 ( .A(n8186), .B(key[1264]), .Z(n7822) );
  XNOR U10568 ( .A(n7853), .B(n7844), .Z(n7821) );
  XNOR U10569 ( .A(n7822), .B(n7821), .Z(\w1[9][112] ) );
  XNOR U10570 ( .A(\w3[8][106] ), .B(\w3[8][114] ), .Z(n7851) );
  XNOR U10571 ( .A(n7851), .B(key[1265]), .Z(n7824) );
  XOR U10572 ( .A(\w3[8][105] ), .B(n8182), .Z(n7823) );
  XNOR U10573 ( .A(n7824), .B(n7823), .Z(\w1[9][113] ) );
  IV U10574 ( .A(\w3[8][115] ), .Z(n7852) );
  XOR U10575 ( .A(\w3[8][107] ), .B(n7852), .Z(n7855) );
  XNOR U10576 ( .A(n7855), .B(key[1266]), .Z(n7826) );
  XNOR U10577 ( .A(\w3[8][106] ), .B(n8187), .Z(n7825) );
  XNOR U10578 ( .A(n7826), .B(n7825), .Z(\w1[9][114] ) );
  XOR U10579 ( .A(\w3[8][116] ), .B(n7848), .Z(n7856) );
  XOR U10580 ( .A(\w3[8][117] ), .B(n7848), .Z(n7860) );
  XNOR U10581 ( .A(n7860), .B(key[1268]), .Z(n7830) );
  XOR U10582 ( .A(\w3[8][108] ), .B(n7828), .Z(n7829) );
  XNOR U10583 ( .A(n7830), .B(n7829), .Z(\w1[9][116] ) );
  XNOR U10584 ( .A(n7831), .B(key[1269]), .Z(n7834) );
  XNOR U10585 ( .A(\w3[8][109] ), .B(n7832), .Z(n7833) );
  XNOR U10586 ( .A(n7834), .B(n7833), .Z(\w1[9][117] ) );
  XOR U10587 ( .A(\w3[8][119] ), .B(n7848), .Z(n7868) );
  XNOR U10588 ( .A(n7868), .B(key[1270]), .Z(n7837) );
  XOR U10589 ( .A(\w3[8][110] ), .B(n7835), .Z(n7836) );
  XNOR U10590 ( .A(n7837), .B(n7836), .Z(\w1[9][118] ) );
  XOR U10591 ( .A(n7838), .B(key[1271]), .Z(n7841) );
  XNOR U10592 ( .A(\w3[8][112] ), .B(n7839), .Z(n7840) );
  XNOR U10593 ( .A(n7841), .B(n7840), .Z(\w1[9][119] ) );
  XNOR U10594 ( .A(\w3[8][3] ), .B(\w3[8][27] ), .Z(n7932) );
  XNOR U10595 ( .A(n7892), .B(key[1163]), .Z(n7843) );
  XNOR U10596 ( .A(\w3[8][0] ), .B(\w3[8][4] ), .Z(n7961) );
  XOR U10597 ( .A(\w3[8][19] ), .B(n7961), .Z(n7842) );
  XNOR U10598 ( .A(n7843), .B(n7842), .Z(\w1[9][11] ) );
  XNOR U10599 ( .A(n7844), .B(key[1272]), .Z(n7846) );
  XNOR U10600 ( .A(\w3[8][121] ), .B(\w3[8][113] ), .Z(n7845) );
  XNOR U10601 ( .A(n7846), .B(n7845), .Z(n7847) );
  XNOR U10602 ( .A(n7848), .B(n7847), .Z(\w1[9][120] ) );
  XNOR U10603 ( .A(\w3[8][114] ), .B(\w3[8][122] ), .Z(n8190) );
  XNOR U10604 ( .A(n8190), .B(key[1273]), .Z(n7850) );
  XOR U10605 ( .A(\w3[8][97] ), .B(n8186), .Z(n7849) );
  XNOR U10606 ( .A(n7850), .B(n7849), .Z(\w1[9][121] ) );
  XOR U10607 ( .A(\w3[8][124] ), .B(n7853), .Z(n7854) );
  XOR U10608 ( .A(n7855), .B(n7854), .Z(n8194) );
  XOR U10609 ( .A(n8194), .B(key[1275]), .Z(n7859) );
  XNOR U10610 ( .A(n7857), .B(n7856), .Z(n7858) );
  XNOR U10611 ( .A(n7859), .B(n7858), .Z(\w1[9][123] ) );
  XNOR U10612 ( .A(n7860), .B(key[1276]), .Z(n7863) );
  XOR U10613 ( .A(n7861), .B(\w3[8][100] ), .Z(n7862) );
  XNOR U10614 ( .A(n7863), .B(n7862), .Z(\w1[9][124] ) );
  XOR U10615 ( .A(\w3[8][118] ), .B(key[1277]), .Z(n7865) );
  XNOR U10616 ( .A(\w3[8][101] ), .B(\w3[8][126] ), .Z(n7864) );
  XNOR U10617 ( .A(n7865), .B(n7864), .Z(n7866) );
  XNOR U10618 ( .A(n7867), .B(n7866), .Z(\w1[9][125] ) );
  XNOR U10619 ( .A(n7868), .B(key[1278]), .Z(n7871) );
  XOR U10620 ( .A(\w3[8][102] ), .B(n7869), .Z(n7870) );
  XNOR U10621 ( .A(n7871), .B(n7870), .Z(\w1[9][126] ) );
  XNOR U10622 ( .A(n8183), .B(key[1279]), .Z(n7874) );
  XOR U10623 ( .A(\w3[8][103] ), .B(n7872), .Z(n7873) );
  XNOR U10624 ( .A(n7874), .B(n7873), .Z(\w1[9][127] ) );
  XOR U10625 ( .A(\w3[8][13] ), .B(\w3[8][28] ), .Z(n7876) );
  XNOR U10626 ( .A(\w3[8][8] ), .B(\w3[8][4] ), .Z(n7875) );
  XOR U10627 ( .A(n7876), .B(n7875), .Z(n7896) );
  XNOR U10628 ( .A(n7896), .B(key[1164]), .Z(n7878) );
  XNOR U10629 ( .A(\w3[8][0] ), .B(\w3[8][5] ), .Z(n7996) );
  XOR U10630 ( .A(\w3[8][20] ), .B(n7996), .Z(n7877) );
  XNOR U10631 ( .A(n7878), .B(n7877), .Z(\w1[9][12] ) );
  IV U10632 ( .A(\w3[8][21] ), .Z(n7926) );
  XNOR U10633 ( .A(\w3[8][14] ), .B(n7926), .Z(n7880) );
  XNOR U10634 ( .A(\w3[8][5] ), .B(\w3[8][29] ), .Z(n7899) );
  XOR U10635 ( .A(n7899), .B(key[1165]), .Z(n7879) );
  XNOR U10636 ( .A(n7880), .B(n7879), .Z(n7881) );
  XOR U10637 ( .A(\w3[8][6] ), .B(n7881), .Z(\w1[9][13] ) );
  IV U10638 ( .A(\w3[8][30] ), .Z(n8074) );
  XOR U10639 ( .A(\w3[8][6] ), .B(n8074), .Z(n8039) );
  XOR U10640 ( .A(\w3[8][8] ), .B(\w3[8][15] ), .Z(n7902) );
  XNOR U10641 ( .A(n8039), .B(n7902), .Z(n7900) );
  XOR U10642 ( .A(n7900), .B(key[1166]), .Z(n7883) );
  XNOR U10643 ( .A(\w3[8][0] ), .B(\w3[8][7] ), .Z(n8075) );
  XOR U10644 ( .A(\w3[8][22] ), .B(n8075), .Z(n7882) );
  XNOR U10645 ( .A(n7883), .B(n7882), .Z(\w1[9][14] ) );
  XNOR U10646 ( .A(\w3[8][7] ), .B(\w3[8][31] ), .Z(n7901) );
  XNOR U10647 ( .A(n7901), .B(key[1167]), .Z(n7885) );
  XOR U10648 ( .A(\w3[8][8] ), .B(\w3[8][0] ), .Z(n7905) );
  XNOR U10649 ( .A(\w3[8][23] ), .B(n7905), .Z(n7884) );
  XNOR U10650 ( .A(n7885), .B(n7884), .Z(\w1[9][15] ) );
  XNOR U10651 ( .A(\w3[8][17] ), .B(\w3[8][9] ), .Z(n7907) );
  XNOR U10652 ( .A(n7907), .B(key[1168]), .Z(n7887) );
  XNOR U10653 ( .A(\w3[8][24] ), .B(n7905), .Z(n7886) );
  XNOR U10654 ( .A(n7887), .B(n7886), .Z(\w1[9][16] ) );
  XNOR U10655 ( .A(\w3[8][18] ), .B(\w3[8][10] ), .Z(n7931) );
  XNOR U10656 ( .A(n7931), .B(key[1169]), .Z(n7889) );
  IV U10657 ( .A(\w3[8][9] ), .Z(n8150) );
  XNOR U10658 ( .A(n8202), .B(n8150), .Z(n7888) );
  XNOR U10659 ( .A(n7889), .B(n7888), .Z(\w1[9][17] ) );
  IV U10660 ( .A(\w3[8][19] ), .Z(n7912) );
  XOR U10661 ( .A(\w3[8][11] ), .B(n7912), .Z(n7917) );
  XNOR U10662 ( .A(n7917), .B(key[1170]), .Z(n7891) );
  XOR U10663 ( .A(n7893), .B(\w3[8][10] ), .Z(n7890) );
  XNOR U10664 ( .A(n7891), .B(n7890), .Z(\w1[9][18] ) );
  XOR U10665 ( .A(n7906), .B(\w3[8][20] ), .Z(n7918) );
  XNOR U10666 ( .A(n7907), .B(key[1153]), .Z(n7895) );
  XOR U10667 ( .A(\w3[8][25] ), .B(n7893), .Z(n7894) );
  XNOR U10668 ( .A(n7895), .B(n7894), .Z(\w1[9][1] ) );
  XOR U10669 ( .A(\w3[8][16] ), .B(n7926), .Z(n7923) );
  XNOR U10670 ( .A(n7923), .B(key[1172]), .Z(n7898) );
  XOR U10671 ( .A(\w3[8][12] ), .B(n7896), .Z(n7897) );
  XNOR U10672 ( .A(n7898), .B(n7897), .Z(\w1[9][20] ) );
  IV U10673 ( .A(\w3[8][22] ), .Z(n7927) );
  XOR U10674 ( .A(\w3[8][14] ), .B(n7927), .Z(n7936) );
  XOR U10675 ( .A(n7906), .B(\w3[8][23] ), .Z(n7937) );
  XNOR U10676 ( .A(n7901), .B(key[1175]), .Z(n7904) );
  XNOR U10677 ( .A(\w3[8][16] ), .B(n7902), .Z(n7903) );
  XNOR U10678 ( .A(n7904), .B(n7903), .Z(\w1[9][23] ) );
  XNOR U10679 ( .A(n7907), .B(key[1177]), .Z(n7909) );
  XNOR U10680 ( .A(\w3[8][1] ), .B(\w3[8][26] ), .Z(n7908) );
  XNOR U10681 ( .A(n7909), .B(n7908), .Z(n7910) );
  XNOR U10682 ( .A(n7911), .B(n7910), .Z(\w1[9][25] ) );
  XNOR U10683 ( .A(n7931), .B(key[1178]), .Z(n7914) );
  XOR U10684 ( .A(\w3[8][2] ), .B(n7912), .Z(n7913) );
  XNOR U10685 ( .A(n7914), .B(n7913), .Z(n7915) );
  XOR U10686 ( .A(\w3[8][27] ), .B(n7915), .Z(\w1[9][26] ) );
  IV U10687 ( .A(\w3[8][24] ), .Z(n7935) );
  XOR U10688 ( .A(n7935), .B(\w3[8][28] ), .Z(n7916) );
  XOR U10689 ( .A(n7917), .B(n7916), .Z(n7960) );
  XOR U10690 ( .A(n7960), .B(key[1179]), .Z(n7920) );
  XOR U10691 ( .A(\w3[8][3] ), .B(n7918), .Z(n7919) );
  XNOR U10692 ( .A(n7920), .B(n7919), .Z(\w1[9][27] ) );
  XOR U10693 ( .A(\w3[8][20] ), .B(\w3[8][29] ), .Z(n7922) );
  XOR U10694 ( .A(n7935), .B(\w3[8][12] ), .Z(n7921) );
  XOR U10695 ( .A(n7922), .B(n7921), .Z(n7995) );
  XNOR U10696 ( .A(n7995), .B(key[1180]), .Z(n7925) );
  XOR U10697 ( .A(\w3[8][4] ), .B(n7923), .Z(n7924) );
  XNOR U10698 ( .A(n7925), .B(n7924), .Z(\w1[9][28] ) );
  XOR U10699 ( .A(\w3[8][13] ), .B(n7926), .Z(n8038) );
  XNOR U10700 ( .A(n8038), .B(key[1181]), .Z(n7929) );
  XNOR U10701 ( .A(n7927), .B(n8074), .Z(n7928) );
  XNOR U10702 ( .A(n7929), .B(n7928), .Z(n7930) );
  XOR U10703 ( .A(\w3[8][5] ), .B(n7930), .Z(\w1[9][29] ) );
  XNOR U10704 ( .A(n7931), .B(key[1154]), .Z(n7934) );
  XOR U10705 ( .A(\w3[8][26] ), .B(n7932), .Z(n7933) );
  XNOR U10706 ( .A(n7934), .B(n7933), .Z(\w1[9][2] ) );
  XOR U10707 ( .A(n7935), .B(\w3[8][31] ), .Z(n8113) );
  XNOR U10708 ( .A(n7936), .B(n8113), .Z(n8073) );
  XNOR U10709 ( .A(\w3[8][15] ), .B(\w3[8][23] ), .Z(n8112) );
  XNOR U10710 ( .A(n8112), .B(key[1183]), .Z(n7939) );
  XOR U10711 ( .A(n8153), .B(\w3[8][7] ), .Z(n7938) );
  XNOR U10712 ( .A(n7939), .B(n7938), .Z(\w1[9][31] ) );
  XNOR U10713 ( .A(\w3[8][48] ), .B(\w3[8][56] ), .Z(n8055) );
  XNOR U10714 ( .A(\w3[8][33] ), .B(\w3[8][57] ), .Z(n7992) );
  XNOR U10715 ( .A(\w3[8][40] ), .B(key[1184]), .Z(n7940) );
  XNOR U10716 ( .A(n7992), .B(n7940), .Z(n7941) );
  XOR U10717 ( .A(n8055), .B(n7941), .Z(\w1[9][32] ) );
  IV U10718 ( .A(\w3[8][34] ), .Z(n8032) );
  IV U10719 ( .A(\w3[8][58] ), .Z(n8001) );
  XOR U10720 ( .A(n8032), .B(n8001), .Z(n7969) );
  XOR U10721 ( .A(n7969), .B(key[1185]), .Z(n7943) );
  XNOR U10722 ( .A(\w3[8][41] ), .B(\w3[8][49] ), .Z(n8025) );
  XOR U10723 ( .A(\w3[8][57] ), .B(n8025), .Z(n7942) );
  XNOR U10724 ( .A(n7943), .B(n7942), .Z(\w1[9][33] ) );
  XNOR U10725 ( .A(n7970), .B(key[1186]), .Z(n7945) );
  XNOR U10726 ( .A(\w3[8][50] ), .B(\w3[8][42] ), .Z(n8028) );
  XOR U10727 ( .A(\w3[8][58] ), .B(n8028), .Z(n7944) );
  XNOR U10728 ( .A(n7945), .B(n7944), .Z(\w1[9][34] ) );
  XOR U10729 ( .A(\w3[8][36] ), .B(\w3[8][32] ), .Z(n7972) );
  XOR U10730 ( .A(n7972), .B(key[1187]), .Z(n7948) );
  IV U10731 ( .A(\w3[8][51] ), .Z(n8027) );
  XOR U10732 ( .A(\w3[8][43] ), .B(n8027), .Z(n8000) );
  XOR U10733 ( .A(\w3[8][56] ), .B(n8000), .Z(n7946) );
  XNOR U10734 ( .A(\w3[8][60] ), .B(n7946), .Z(n8034) );
  XNOR U10735 ( .A(\w3[8][59] ), .B(n8034), .Z(n7947) );
  XNOR U10736 ( .A(n7948), .B(n7947), .Z(\w1[9][35] ) );
  XOR U10737 ( .A(\w3[8][32] ), .B(\w3[8][37] ), .Z(n7978) );
  XOR U10738 ( .A(\w3[8][52] ), .B(\w3[8][61] ), .Z(n7950) );
  XNOR U10739 ( .A(\w3[8][56] ), .B(\w3[8][44] ), .Z(n7949) );
  XOR U10740 ( .A(n7950), .B(n7949), .Z(n8043) );
  XOR U10741 ( .A(n8043), .B(key[1188]), .Z(n7951) );
  XOR U10742 ( .A(n7978), .B(n7951), .Z(n7952) );
  XNOR U10743 ( .A(\w3[8][60] ), .B(n7952), .Z(\w1[9][36] ) );
  XNOR U10744 ( .A(\w3[8][38] ), .B(\w3[8][62] ), .Z(n7984) );
  XNOR U10745 ( .A(n7984), .B(key[1189]), .Z(n7954) );
  IV U10746 ( .A(\w3[8][45] ), .Z(n8010) );
  XOR U10747 ( .A(\w3[8][53] ), .B(n8010), .Z(n8049) );
  XOR U10748 ( .A(\w3[8][61] ), .B(n8049), .Z(n7953) );
  XNOR U10749 ( .A(n7954), .B(n7953), .Z(\w1[9][37] ) );
  XOR U10750 ( .A(\w3[8][32] ), .B(\w3[8][39] ), .Z(n7985) );
  XOR U10751 ( .A(n7985), .B(key[1190]), .Z(n7956) );
  XNOR U10752 ( .A(\w3[8][56] ), .B(\w3[8][63] ), .Z(n7957) );
  XOR U10753 ( .A(\w3[8][46] ), .B(\w3[8][54] ), .Z(n8009) );
  XOR U10754 ( .A(n7957), .B(n8009), .Z(n8051) );
  XOR U10755 ( .A(\w3[8][62] ), .B(n8051), .Z(n7955) );
  XNOR U10756 ( .A(n7956), .B(n7955), .Z(\w1[9][38] ) );
  XNOR U10757 ( .A(\w3[8][55] ), .B(\w3[8][47] ), .Z(n8054) );
  XNOR U10758 ( .A(n8054), .B(key[1191]), .Z(n7959) );
  XOR U10759 ( .A(\w3[8][32] ), .B(n7957), .Z(n7958) );
  XNOR U10760 ( .A(n7959), .B(n7958), .Z(\w1[9][39] ) );
  XOR U10761 ( .A(n7960), .B(key[1155]), .Z(n7963) );
  XOR U10762 ( .A(n7961), .B(\w3[8][27] ), .Z(n7962) );
  XNOR U10763 ( .A(n7963), .B(n7962), .Z(\w1[9][3] ) );
  IV U10764 ( .A(\w3[8][33] ), .Z(n8026) );
  XOR U10765 ( .A(\w3[8][34] ), .B(\w3[8][42] ), .Z(n7999) );
  XOR U10766 ( .A(n7999), .B(key[1193]), .Z(n7965) );
  XOR U10767 ( .A(n7992), .B(\w3[8][49] ), .Z(n7964) );
  XNOR U10768 ( .A(n7965), .B(n7964), .Z(\w1[9][41] ) );
  XOR U10769 ( .A(\w3[8][43] ), .B(key[1194]), .Z(n7967) );
  IV U10770 ( .A(\w3[8][35] ), .Z(n8035) );
  XOR U10771 ( .A(\w3[8][50] ), .B(n8035), .Z(n7966) );
  XNOR U10772 ( .A(n7967), .B(n7966), .Z(n7968) );
  XOR U10773 ( .A(n7969), .B(n7968), .Z(\w1[9][42] ) );
  IV U10774 ( .A(\w3[8][40] ), .Z(n7975) );
  XNOR U10775 ( .A(n7975), .B(n7970), .Z(n7971) );
  XOR U10776 ( .A(\w3[8][44] ), .B(n7971), .Z(n8004) );
  XNOR U10777 ( .A(n8004), .B(key[1195]), .Z(n7974) );
  XNOR U10778 ( .A(\w3[8][51] ), .B(n7972), .Z(n7973) );
  XNOR U10779 ( .A(n7974), .B(n7973), .Z(\w1[9][43] ) );
  XOR U10780 ( .A(\w3[8][36] ), .B(\w3[8][45] ), .Z(n7977) );
  XOR U10781 ( .A(n7975), .B(\w3[8][60] ), .Z(n7976) );
  XOR U10782 ( .A(n7977), .B(n7976), .Z(n8005) );
  XNOR U10783 ( .A(n8005), .B(key[1196]), .Z(n7980) );
  XNOR U10784 ( .A(\w3[8][52] ), .B(n7978), .Z(n7979) );
  XNOR U10785 ( .A(n7980), .B(n7979), .Z(\w1[9][44] ) );
  XNOR U10786 ( .A(\w3[8][61] ), .B(\w3[8][37] ), .Z(n8008) );
  XNOR U10787 ( .A(n8008), .B(key[1197]), .Z(n7982) );
  XNOR U10788 ( .A(\w3[8][38] ), .B(\w3[8][46] ), .Z(n7981) );
  XNOR U10789 ( .A(n7982), .B(n7981), .Z(n7983) );
  XOR U10790 ( .A(\w3[8][53] ), .B(n7983), .Z(\w1[9][45] ) );
  XOR U10791 ( .A(\w3[8][40] ), .B(\w3[8][47] ), .Z(n8017) );
  XOR U10792 ( .A(n7984), .B(n8017), .Z(n8013) );
  XNOR U10793 ( .A(n8013), .B(key[1198]), .Z(n7987) );
  XNOR U10794 ( .A(\w3[8][54] ), .B(n7985), .Z(n7986) );
  XNOR U10795 ( .A(n7987), .B(n7986), .Z(\w1[9][46] ) );
  XOR U10796 ( .A(\w3[8][63] ), .B(\w3[8][39] ), .Z(n8016) );
  XOR U10797 ( .A(n8016), .B(key[1199]), .Z(n7989) );
  XNOR U10798 ( .A(\w3[8][40] ), .B(\w3[8][32] ), .Z(n8020) );
  XOR U10799 ( .A(\w3[8][55] ), .B(n8020), .Z(n7988) );
  XNOR U10800 ( .A(n7989), .B(n7988), .Z(\w1[9][47] ) );
  XNOR U10801 ( .A(n8020), .B(key[1200]), .Z(n7991) );
  XOR U10802 ( .A(\w3[8][56] ), .B(n8025), .Z(n7990) );
  XNOR U10803 ( .A(n7991), .B(n7990), .Z(\w1[9][48] ) );
  XNOR U10804 ( .A(n8028), .B(key[1201]), .Z(n7994) );
  XOR U10805 ( .A(n7992), .B(\w3[8][41] ), .Z(n7993) );
  XNOR U10806 ( .A(n7994), .B(n7993), .Z(\w1[9][49] ) );
  XNOR U10807 ( .A(n7995), .B(key[1156]), .Z(n7998) );
  XOR U10808 ( .A(n7996), .B(\w3[8][28] ), .Z(n7997) );
  XNOR U10809 ( .A(n7998), .B(n7997), .Z(\w1[9][4] ) );
  XOR U10810 ( .A(n7999), .B(key[1202]), .Z(n8003) );
  XNOR U10811 ( .A(n8001), .B(n8000), .Z(n8002) );
  XNOR U10812 ( .A(n8003), .B(n8002), .Z(\w1[9][50] ) );
  IV U10813 ( .A(\w3[8][48] ), .Z(n8021) );
  XOR U10814 ( .A(n8021), .B(\w3[8][52] ), .Z(n8033) );
  XNOR U10815 ( .A(n8042), .B(key[1204]), .Z(n8007) );
  XOR U10816 ( .A(\w3[8][44] ), .B(n8005), .Z(n8006) );
  XNOR U10817 ( .A(n8007), .B(n8006), .Z(\w1[9][52] ) );
  XNOR U10818 ( .A(n8008), .B(key[1205]), .Z(n8012) );
  XOR U10819 ( .A(n8010), .B(n8009), .Z(n8011) );
  XNOR U10820 ( .A(n8012), .B(n8011), .Z(\w1[9][53] ) );
  XOR U10821 ( .A(n8021), .B(\w3[8][55] ), .Z(n8050) );
  XNOR U10822 ( .A(n8050), .B(key[1206]), .Z(n8015) );
  XOR U10823 ( .A(\w3[8][46] ), .B(n8013), .Z(n8014) );
  XNOR U10824 ( .A(n8015), .B(n8014), .Z(\w1[9][54] ) );
  XOR U10825 ( .A(n8016), .B(key[1207]), .Z(n8019) );
  XNOR U10826 ( .A(\w3[8][48] ), .B(n8017), .Z(n8018) );
  XNOR U10827 ( .A(n8019), .B(n8018), .Z(\w1[9][55] ) );
  XNOR U10828 ( .A(n8020), .B(key[1208]), .Z(n8023) );
  XOR U10829 ( .A(n8021), .B(\w3[8][49] ), .Z(n8022) );
  XNOR U10830 ( .A(n8023), .B(n8022), .Z(n8024) );
  XOR U10831 ( .A(\w3[8][57] ), .B(n8024), .Z(\w1[9][56] ) );
  XNOR U10832 ( .A(n8027), .B(key[1210]), .Z(n8030) );
  XOR U10833 ( .A(n8028), .B(\w3[8][59] ), .Z(n8029) );
  XNOR U10834 ( .A(n8030), .B(n8029), .Z(n8031) );
  XNOR U10835 ( .A(n8032), .B(n8031), .Z(\w1[9][58] ) );
  XNOR U10836 ( .A(n8033), .B(key[1211]), .Z(n8037) );
  XOR U10837 ( .A(n8035), .B(n8034), .Z(n8036) );
  XNOR U10838 ( .A(n8037), .B(n8036), .Z(\w1[9][59] ) );
  XNOR U10839 ( .A(n8038), .B(key[1157]), .Z(n8041) );
  XOR U10840 ( .A(\w3[8][29] ), .B(n8039), .Z(n8040) );
  XNOR U10841 ( .A(n8041), .B(n8040), .Z(\w1[9][5] ) );
  XNOR U10842 ( .A(n8042), .B(key[1212]), .Z(n8045) );
  XOR U10843 ( .A(\w3[8][36] ), .B(n8043), .Z(n8044) );
  XNOR U10844 ( .A(n8045), .B(n8044), .Z(\w1[9][60] ) );
  XOR U10845 ( .A(\w3[8][54] ), .B(key[1213]), .Z(n8047) );
  XNOR U10846 ( .A(\w3[8][37] ), .B(\w3[8][62] ), .Z(n8046) );
  XNOR U10847 ( .A(n8047), .B(n8046), .Z(n8048) );
  XNOR U10848 ( .A(n8049), .B(n8048), .Z(\w1[9][61] ) );
  XNOR U10849 ( .A(n8050), .B(key[1214]), .Z(n8053) );
  XOR U10850 ( .A(\w3[8][38] ), .B(n8051), .Z(n8052) );
  XNOR U10851 ( .A(n8053), .B(n8052), .Z(\w1[9][62] ) );
  XNOR U10852 ( .A(n8054), .B(key[1215]), .Z(n8057) );
  XOR U10853 ( .A(n8055), .B(\w3[8][39] ), .Z(n8056) );
  XNOR U10854 ( .A(n8057), .B(n8056), .Z(\w1[9][63] ) );
  IV U10855 ( .A(\w3[8][65] ), .Z(n8149) );
  IV U10856 ( .A(\w3[8][89] ), .Z(n8147) );
  XOR U10857 ( .A(n8149), .B(n8147), .Z(n8085) );
  XOR U10858 ( .A(n8085), .B(key[1216]), .Z(n8059) );
  XNOR U10859 ( .A(\w3[8][80] ), .B(\w3[8][88] ), .Z(n8179) );
  XOR U10860 ( .A(n8179), .B(\w3[8][72] ), .Z(n8058) );
  XNOR U10861 ( .A(n8059), .B(n8058), .Z(\w1[9][64] ) );
  IV U10862 ( .A(\w3[8][66] ), .Z(n8160) );
  IV U10863 ( .A(\w3[8][90] ), .Z(n8123) );
  XOR U10864 ( .A(n8160), .B(n8123), .Z(n8091) );
  XOR U10865 ( .A(n8091), .B(key[1217]), .Z(n8061) );
  XNOR U10866 ( .A(\w3[8][73] ), .B(\w3[8][81] ), .Z(n8148) );
  XOR U10867 ( .A(\w3[8][89] ), .B(n8148), .Z(n8060) );
  XNOR U10868 ( .A(n8061), .B(n8060), .Z(\w1[9][65] ) );
  XNOR U10869 ( .A(n8092), .B(key[1218]), .Z(n8063) );
  XNOR U10870 ( .A(\w3[8][82] ), .B(\w3[8][74] ), .Z(n8156) );
  XOR U10871 ( .A(\w3[8][90] ), .B(n8156), .Z(n8062) );
  XNOR U10872 ( .A(n8063), .B(n8062), .Z(\w1[9][66] ) );
  XOR U10873 ( .A(\w3[8][68] ), .B(\w3[8][64] ), .Z(n8094) );
  XOR U10874 ( .A(n8094), .B(key[1219]), .Z(n8066) );
  IV U10875 ( .A(\w3[8][83] ), .Z(n8155) );
  XOR U10876 ( .A(\w3[8][75] ), .B(n8155), .Z(n8122) );
  XOR U10877 ( .A(\w3[8][88] ), .B(n8122), .Z(n8064) );
  XNOR U10878 ( .A(\w3[8][92] ), .B(n8064), .Z(n8162) );
  XNOR U10879 ( .A(\w3[8][91] ), .B(n8162), .Z(n8065) );
  XNOR U10880 ( .A(n8066), .B(n8065), .Z(\w1[9][67] ) );
  XOR U10881 ( .A(\w3[8][64] ), .B(\w3[8][69] ), .Z(n8100) );
  XOR U10882 ( .A(\w3[8][84] ), .B(\w3[8][93] ), .Z(n8068) );
  XNOR U10883 ( .A(\w3[8][88] ), .B(\w3[8][76] ), .Z(n8067) );
  XOR U10884 ( .A(n8068), .B(n8067), .Z(n8167) );
  XOR U10885 ( .A(n8167), .B(key[1220]), .Z(n8069) );
  XOR U10886 ( .A(n8100), .B(n8069), .Z(n8070) );
  XNOR U10887 ( .A(\w3[8][92] ), .B(n8070), .Z(\w1[9][68] ) );
  XNOR U10888 ( .A(\w3[8][70] ), .B(\w3[8][94] ), .Z(n8106) );
  XNOR U10889 ( .A(n8106), .B(key[1221]), .Z(n8072) );
  IV U10890 ( .A(\w3[8][77] ), .Z(n8132) );
  XOR U10891 ( .A(\w3[8][85] ), .B(n8132), .Z(n8173) );
  XOR U10892 ( .A(\w3[8][93] ), .B(n8173), .Z(n8071) );
  XNOR U10893 ( .A(n8072), .B(n8071), .Z(\w1[9][69] ) );
  XNOR U10894 ( .A(n8073), .B(key[1158]), .Z(n8077) );
  XNOR U10895 ( .A(n8075), .B(n8074), .Z(n8076) );
  XNOR U10896 ( .A(n8077), .B(n8076), .Z(\w1[9][6] ) );
  XOR U10897 ( .A(\w3[8][64] ), .B(\w3[8][71] ), .Z(n8107) );
  XOR U10898 ( .A(n8107), .B(key[1222]), .Z(n8079) );
  XNOR U10899 ( .A(\w3[8][88] ), .B(\w3[8][95] ), .Z(n8080) );
  XOR U10900 ( .A(\w3[8][78] ), .B(\w3[8][86] ), .Z(n8131) );
  XOR U10901 ( .A(n8080), .B(n8131), .Z(n8175) );
  XOR U10902 ( .A(\w3[8][94] ), .B(n8175), .Z(n8078) );
  XNOR U10903 ( .A(n8079), .B(n8078), .Z(\w1[9][70] ) );
  XNOR U10904 ( .A(\w3[8][79] ), .B(\w3[8][87] ), .Z(n8178) );
  XNOR U10905 ( .A(n8178), .B(key[1223]), .Z(n8082) );
  XOR U10906 ( .A(\w3[8][64] ), .B(n8080), .Z(n8081) );
  XNOR U10907 ( .A(n8082), .B(n8081), .Z(\w1[9][71] ) );
  XOR U10908 ( .A(\w3[8][65] ), .B(\w3[8][73] ), .Z(n8118) );
  XOR U10909 ( .A(n8118), .B(key[1224]), .Z(n8084) );
  XOR U10910 ( .A(n8179), .B(\w3[8][64] ), .Z(n8083) );
  XNOR U10911 ( .A(n8084), .B(n8083), .Z(\w1[9][72] ) );
  XOR U10912 ( .A(\w3[8][66] ), .B(\w3[8][74] ), .Z(n8121) );
  XOR U10913 ( .A(n8121), .B(key[1225]), .Z(n8087) );
  XNOR U10914 ( .A(n8085), .B(\w3[8][81] ), .Z(n8086) );
  XNOR U10915 ( .A(n8087), .B(n8086), .Z(\w1[9][73] ) );
  XOR U10916 ( .A(\w3[8][75] ), .B(key[1226]), .Z(n8089) );
  IV U10917 ( .A(\w3[8][67] ), .Z(n8163) );
  XOR U10918 ( .A(\w3[8][82] ), .B(n8163), .Z(n8088) );
  XNOR U10919 ( .A(n8089), .B(n8088), .Z(n8090) );
  XOR U10920 ( .A(n8091), .B(n8090), .Z(\w1[9][74] ) );
  IV U10921 ( .A(\w3[8][72] ), .Z(n8097) );
  XNOR U10922 ( .A(n8097), .B(n8092), .Z(n8093) );
  XOR U10923 ( .A(\w3[8][76] ), .B(n8093), .Z(n8126) );
  XNOR U10924 ( .A(n8126), .B(key[1227]), .Z(n8096) );
  XNOR U10925 ( .A(\w3[8][83] ), .B(n8094), .Z(n8095) );
  XNOR U10926 ( .A(n8096), .B(n8095), .Z(\w1[9][75] ) );
  XOR U10927 ( .A(\w3[8][68] ), .B(\w3[8][77] ), .Z(n8099) );
  XOR U10928 ( .A(n8097), .B(\w3[8][92] ), .Z(n8098) );
  XOR U10929 ( .A(n8099), .B(n8098), .Z(n8127) );
  XNOR U10930 ( .A(n8127), .B(key[1228]), .Z(n8102) );
  XNOR U10931 ( .A(\w3[8][84] ), .B(n8100), .Z(n8101) );
  XNOR U10932 ( .A(n8102), .B(n8101), .Z(\w1[9][76] ) );
  XNOR U10933 ( .A(\w3[8][93] ), .B(\w3[8][69] ), .Z(n8130) );
  XNOR U10934 ( .A(n8130), .B(key[1229]), .Z(n8104) );
  XNOR U10935 ( .A(\w3[8][70] ), .B(\w3[8][78] ), .Z(n8103) );
  XNOR U10936 ( .A(n8104), .B(n8103), .Z(n8105) );
  XOR U10937 ( .A(\w3[8][85] ), .B(n8105), .Z(\w1[9][77] ) );
  XOR U10938 ( .A(\w3[8][72] ), .B(\w3[8][79] ), .Z(n8139) );
  XOR U10939 ( .A(n8106), .B(n8139), .Z(n8135) );
  XNOR U10940 ( .A(n8135), .B(key[1230]), .Z(n8109) );
  XNOR U10941 ( .A(\w3[8][86] ), .B(n8107), .Z(n8108) );
  XNOR U10942 ( .A(n8109), .B(n8108), .Z(\w1[9][78] ) );
  XOR U10943 ( .A(\w3[8][95] ), .B(\w3[8][71] ), .Z(n8138) );
  XOR U10944 ( .A(n8138), .B(key[1231]), .Z(n8111) );
  XNOR U10945 ( .A(\w3[8][72] ), .B(\w3[8][64] ), .Z(n8142) );
  XOR U10946 ( .A(\w3[8][87] ), .B(n8142), .Z(n8110) );
  XNOR U10947 ( .A(n8111), .B(n8110), .Z(\w1[9][79] ) );
  XNOR U10948 ( .A(n8112), .B(key[1159]), .Z(n8115) );
  XOR U10949 ( .A(\w3[8][0] ), .B(n8113), .Z(n8114) );
  XNOR U10950 ( .A(n8115), .B(n8114), .Z(\w1[9][7] ) );
  XNOR U10951 ( .A(n8142), .B(key[1232]), .Z(n8117) );
  XOR U10952 ( .A(\w3[8][88] ), .B(n8148), .Z(n8116) );
  XNOR U10953 ( .A(n8117), .B(n8116), .Z(\w1[9][80] ) );
  XOR U10954 ( .A(n8118), .B(key[1233]), .Z(n8120) );
  XOR U10955 ( .A(\w3[8][89] ), .B(n8156), .Z(n8119) );
  XNOR U10956 ( .A(n8120), .B(n8119), .Z(\w1[9][81] ) );
  XOR U10957 ( .A(n8121), .B(key[1234]), .Z(n8125) );
  XNOR U10958 ( .A(n8123), .B(n8122), .Z(n8124) );
  XNOR U10959 ( .A(n8125), .B(n8124), .Z(\w1[9][82] ) );
  IV U10960 ( .A(\w3[8][80] ), .Z(n8143) );
  XOR U10961 ( .A(n8143), .B(\w3[8][84] ), .Z(n8161) );
  XNOR U10962 ( .A(n8166), .B(key[1236]), .Z(n8129) );
  XOR U10963 ( .A(\w3[8][76] ), .B(n8127), .Z(n8128) );
  XNOR U10964 ( .A(n8129), .B(n8128), .Z(\w1[9][84] ) );
  XNOR U10965 ( .A(n8130), .B(key[1237]), .Z(n8134) );
  XOR U10966 ( .A(n8132), .B(n8131), .Z(n8133) );
  XNOR U10967 ( .A(n8134), .B(n8133), .Z(\w1[9][85] ) );
  XOR U10968 ( .A(n8143), .B(\w3[8][87] ), .Z(n8174) );
  XNOR U10969 ( .A(n8174), .B(key[1238]), .Z(n8137) );
  XOR U10970 ( .A(\w3[8][78] ), .B(n8135), .Z(n8136) );
  XNOR U10971 ( .A(n8137), .B(n8136), .Z(\w1[9][86] ) );
  XOR U10972 ( .A(n8138), .B(key[1239]), .Z(n8141) );
  XNOR U10973 ( .A(\w3[8][80] ), .B(n8139), .Z(n8140) );
  XNOR U10974 ( .A(n8141), .B(n8140), .Z(\w1[9][87] ) );
  XNOR U10975 ( .A(n8142), .B(key[1240]), .Z(n8145) );
  XOR U10976 ( .A(n8143), .B(\w3[8][81] ), .Z(n8144) );
  XNOR U10977 ( .A(n8145), .B(n8144), .Z(n8146) );
  XNOR U10978 ( .A(n8147), .B(n8146), .Z(\w1[9][88] ) );
  XNOR U10979 ( .A(n8150), .B(key[1160]), .Z(n8152) );
  XNOR U10980 ( .A(\w3[8][1] ), .B(\w3[8][0] ), .Z(n8151) );
  XNOR U10981 ( .A(n8152), .B(n8151), .Z(n8154) );
  XNOR U10982 ( .A(n8154), .B(n8153), .Z(\w1[9][8] ) );
  XNOR U10983 ( .A(n8155), .B(key[1242]), .Z(n8158) );
  XOR U10984 ( .A(n8156), .B(\w3[8][91] ), .Z(n8157) );
  XNOR U10985 ( .A(n8158), .B(n8157), .Z(n8159) );
  XNOR U10986 ( .A(n8160), .B(n8159), .Z(\w1[9][90] ) );
  XNOR U10987 ( .A(n8161), .B(key[1243]), .Z(n8165) );
  XOR U10988 ( .A(n8163), .B(n8162), .Z(n8164) );
  XNOR U10989 ( .A(n8165), .B(n8164), .Z(\w1[9][91] ) );
  XNOR U10990 ( .A(n8166), .B(key[1244]), .Z(n8169) );
  XOR U10991 ( .A(\w3[8][68] ), .B(n8167), .Z(n8168) );
  XNOR U10992 ( .A(n8169), .B(n8168), .Z(\w1[9][92] ) );
  XOR U10993 ( .A(\w3[8][86] ), .B(key[1245]), .Z(n8171) );
  XNOR U10994 ( .A(\w3[8][69] ), .B(\w3[8][94] ), .Z(n8170) );
  XNOR U10995 ( .A(n8171), .B(n8170), .Z(n8172) );
  XNOR U10996 ( .A(n8173), .B(n8172), .Z(\w1[9][93] ) );
  XNOR U10997 ( .A(n8174), .B(key[1246]), .Z(n8177) );
  XOR U10998 ( .A(\w3[8][70] ), .B(n8175), .Z(n8176) );
  XNOR U10999 ( .A(n8177), .B(n8176), .Z(\w1[9][94] ) );
  XNOR U11000 ( .A(n8178), .B(key[1247]), .Z(n8181) );
  XOR U11001 ( .A(n8179), .B(\w3[8][71] ), .Z(n8180) );
  XNOR U11002 ( .A(n8181), .B(n8180), .Z(\w1[9][95] ) );
  XOR U11003 ( .A(\w3[8][104] ), .B(key[1248]), .Z(n8185) );
  XNOR U11004 ( .A(n8183), .B(n8182), .Z(n8184) );
  XNOR U11005 ( .A(n8185), .B(n8184), .Z(\w1[9][96] ) );
  XNOR U11006 ( .A(n8186), .B(key[1249]), .Z(n8189) );
  XNOR U11007 ( .A(\w3[8][121] ), .B(n8187), .Z(n8188) );
  XNOR U11008 ( .A(n8189), .B(n8188), .Z(\w1[9][97] ) );
  XNOR U11009 ( .A(n8190), .B(key[1250]), .Z(n8193) );
  XOR U11010 ( .A(\w3[8][106] ), .B(n8191), .Z(n8192) );
  XNOR U11011 ( .A(n8193), .B(n8192), .Z(\w1[9][98] ) );
  XOR U11012 ( .A(n8194), .B(key[1251]), .Z(n8198) );
  XNOR U11013 ( .A(n8196), .B(n8195), .Z(n8197) );
  XNOR U11014 ( .A(n8198), .B(n8197), .Z(\w1[9][99] ) );
  XOR U11015 ( .A(\w3[8][10] ), .B(key[1161]), .Z(n8200) );
  XNOR U11016 ( .A(\w3[8][2] ), .B(\w3[8][17] ), .Z(n8199) );
  XNOR U11017 ( .A(n8200), .B(n8199), .Z(n8201) );
  XNOR U11018 ( .A(n8202), .B(n8201), .Z(\w1[9][9] ) );
endmodule

